magic
tech sky130A
magscale 1 2
timestamp 1655456512
<< pwell >>
rect 550695 586819 551333 586993
rect 571706 586850 572344 587024
rect 544594 572605 544768 573243
rect 525144 567939 525782 568113
rect 513830 562201 514004 562839
rect 505307 559956 505481 560594
rect 531100 552647 531274 553285
rect 544604 552356 544778 552994
rect 522369 549878 522543 550516
rect 513810 541759 513984 542397
rect 505417 539368 505591 540006
rect 544609 532130 544783 532768
rect 531055 531402 531229 532040
rect 522418 529101 522592 529739
rect 355859 521649 356033 522287
rect 513807 521788 513981 522426
rect 424083 519146 424721 519320
rect 444096 519205 444734 519379
rect 464279 519288 464917 519462
rect 484611 519249 485249 519423
rect 504085 519256 504723 519430
rect 537514 519401 538152 519575
rect 534412 508338 534586 508976
rect 515106 507471 515280 508109
rect 508800 505911 508974 506549
rect 355824 501740 355998 502378
rect 502246 499864 502420 500502
rect 521250 497785 521424 498423
rect 564206 497618 564844 497792
rect 527534 495539 527708 496177
rect 550534 491594 550708 492232
rect 373694 490060 373868 490698
rect 383346 490058 383520 490696
rect 387983 490139 388157 490777
rect 392886 490153 393060 490791
rect 534422 487938 534596 488576
rect 515069 487270 515243 487908
rect 508812 485860 508986 486498
rect 355886 481796 356060 482434
rect 384062 479678 384700 479852
rect 399517 479703 400155 479877
rect 419759 479643 420397 479817
rect 439997 479672 440635 479846
rect 460297 479684 460935 479858
rect 480479 479662 481117 479836
rect 522885 479711 523523 479885
rect 500435 479364 501073 479538
rect 545778 479368 546416 479542
rect 346850 477856 347024 478494
rect 379027 475577 379665 475751
rect 399517 475610 400155 475784
rect 419759 475550 420397 475724
rect 439997 475579 440635 475753
rect 460297 475591 460935 475765
rect 480479 475569 481117 475743
rect 500467 475587 501105 475761
rect 522917 475240 523555 475414
rect 545831 475276 546469 475450
rect 387992 469175 388166 469813
rect 392884 469175 393058 469813
rect 508844 468627 509018 469265
rect 515101 467217 515275 467855
rect 534454 466549 534628 467187
rect 355894 461776 356068 462414
rect 527389 458988 527563 459626
rect 550228 459117 550402 459755
rect 346864 456602 347038 457240
rect 521282 456702 521456 457340
rect 240779 455301 240953 455939
rect 251501 455279 251675 455917
rect 502278 454623 502452 455261
rect 564140 453363 564778 453537
rect 387953 448155 388127 448793
rect 392874 448223 393048 448861
rect 508832 448576 509006 449214
rect 515138 447016 515312 447654
rect 534444 446149 534618 446787
rect 355868 441783 356042 442421
rect 346836 435994 347010 436632
rect 240699 433784 240873 434422
rect 251484 433498 251658 434136
rect 387982 427112 388156 427750
rect 392906 427131 393080 427769
rect 252934 425835 253572 426009
rect 272880 425900 273518 426074
rect 293161 425934 293799 426108
rect 313310 425924 313948 426098
rect 335365 425909 336003 426083
rect 355355 425905 355993 426079
rect 375318 425999 375956 426173
rect 355873 421829 356047 422467
rect 258288 420337 258926 420511
rect 278422 420370 279060 420544
rect 299099 420376 299737 420550
rect 319427 420328 320065 420502
rect 353585 420337 354223 420511
rect 373928 420407 374566 420581
rect 324622 416564 324796 417202
rect 336632 416489 336806 417127
rect 346780 415360 346954 415998
rect 568022 408736 568660 408910
rect 549621 406734 549795 407372
rect 355862 401794 356036 402432
rect 324620 395774 324794 396412
rect 336657 395836 336831 396474
rect 346808 394682 346982 395320
rect 549638 387690 549812 388328
rect 347422 386472 348060 386646
rect 367438 386501 368076 386675
rect 387250 386491 387888 386665
rect 407509 386489 408147 386663
rect 427785 386544 428423 386718
rect 447944 386524 448582 386698
rect 467946 386519 468584 386693
rect 488064 386503 488702 386677
rect 508194 386526 508832 386700
rect 528303 386540 528941 386714
rect 355842 381730 356016 382368
rect 333053 380505 333691 380679
rect 357632 380513 358270 380687
rect 387079 380471 387717 380645
rect 407657 380502 408295 380676
rect 427631 380477 428269 380651
rect 447877 380481 448515 380655
rect 467861 380548 468499 380722
rect 488276 380473 488914 380647
rect 507959 380545 508597 380719
rect 528329 380479 528967 380653
rect 549446 378880 549620 379518
rect 346794 373400 346968 374038
rect 549407 363694 549581 364332
rect 355899 361747 356073 362385
rect 568178 362353 568816 362527
rect 346794 352550 346968 353188
rect 355899 341744 356073 342382
rect 346878 331954 347052 332592
rect 355823 321742 355997 322380
rect 346850 310086 347024 310724
rect 355861 301721 356035 302359
rect 370652 295792 371290 295966
rect 390661 295809 391299 295983
rect 410667 295780 411305 295954
rect 430663 295856 431301 296030
rect 450680 295823 451318 295997
rect 470682 295848 471320 296022
rect 490677 295881 491315 296055
rect 510670 295837 511308 296011
rect 530655 295881 531293 296055
rect 549415 292979 549589 293617
rect 346808 288428 346982 289066
rect 551273 273774 551911 273948
rect 571736 273734 572374 273908
rect 346766 263648 346940 264286
rect 346850 242274 347024 242912
rect 346878 222398 347052 223036
rect 346822 200570 346996 201208
rect 346836 179536 347010 180174
rect 346794 158148 346968 158786
rect 346738 136802 346912 137440
rect 346794 115668 346968 116306
rect 346822 95058 346996 95696
rect 346808 74376 346982 75014
rect 346878 50796 347052 51434
rect 47966 48854 48604 49028
rect 69260 48914 69898 49088
rect 90626 48840 91264 49014
rect 111686 48884 112324 49058
rect 133008 48928 133646 49102
rect 154566 48898 155204 49072
rect 175772 48870 176410 49044
rect 197154 48928 197792 49102
rect 219048 48840 219686 49014
rect 240034 48810 240672 48984
rect 260536 48870 261174 49044
rect 281348 48972 281986 49146
rect 302538 48766 303176 48940
rect 324086 48802 324724 48976
rect 34446 42542 34620 43180
rect 34446 20444 34620 21082
rect 6524 3530 7162 3704
rect 27716 3590 28354 3764
<< viali >>
rect 550871 586751 550937 586861
rect 551243 586741 551309 586851
rect 571882 586782 571948 586892
rect 572254 586772 572320 586882
rect 544736 573153 544846 573219
rect 544726 572781 544836 572847
rect 525320 567871 525386 567981
rect 525692 567861 525758 567971
rect 513762 562597 513872 562663
rect 513752 562225 513862 562291
rect 505449 560504 505559 560570
rect 505439 560132 505549 560198
rect 531032 553043 531142 553109
rect 544746 552904 544856 552970
rect 531022 552671 531132 552737
rect 544736 552532 544846 552598
rect 522511 550426 522621 550492
rect 522501 550054 522611 550120
rect 513742 542155 513852 542221
rect 513732 541783 513842 541849
rect 505559 539916 505669 539982
rect 505549 539544 505659 539610
rect 544751 532678 544861 532744
rect 544741 532306 544851 532372
rect 530987 531798 531097 531864
rect 530977 531426 531087 531492
rect 522560 529649 522670 529715
rect 522550 529277 522660 529343
rect 513739 522184 513849 522250
rect 355991 522045 356101 522111
rect 513729 521812 513839 521878
rect 356001 521673 356111 521739
rect 537690 519333 537756 519443
rect 424259 519078 424325 519188
rect 424631 519068 424697 519178
rect 444272 519137 444338 519247
rect 444644 519127 444710 519237
rect 464455 519220 464521 519330
rect 538062 519323 538128 519433
rect 464827 519210 464893 519320
rect 484787 519181 484853 519291
rect 485159 519171 485225 519281
rect 504261 519188 504327 519298
rect 504633 519178 504699 519288
rect 534334 508886 534444 508952
rect 534344 508514 534454 508580
rect 515038 507867 515148 507933
rect 515028 507495 515138 507561
rect 508942 506459 509052 506525
rect 508932 506087 509042 506153
rect 355956 502136 356066 502202
rect 355966 501764 356076 501830
rect 502178 500260 502288 500326
rect 502168 499888 502278 499954
rect 521392 498333 521502 498399
rect 521382 497961 521492 498027
rect 564230 497760 564296 497870
rect 564602 497750 564668 497860
rect 527466 495935 527576 496001
rect 527456 495563 527566 495629
rect 550466 491990 550576 492056
rect 550456 491618 550566 491684
rect 387905 490687 388015 490753
rect 392808 490701 392918 490767
rect 373616 490608 373726 490674
rect 383268 490606 383378 490672
rect 387915 490315 388025 490381
rect 392818 490329 392928 490395
rect 373626 490236 373736 490302
rect 383278 490234 383388 490300
rect 534344 488486 534454 488552
rect 534354 488114 534464 488180
rect 515001 487666 515111 487732
rect 514991 487294 515101 487360
rect 508954 486408 509064 486474
rect 508944 486036 509054 486102
rect 356018 482192 356128 482258
rect 356028 481820 356138 481886
rect 384086 479600 384152 479710
rect 384458 479610 384524 479720
rect 399541 479625 399607 479735
rect 399913 479635 399979 479745
rect 419783 479565 419849 479675
rect 420155 479575 420221 479685
rect 440021 479594 440087 479704
rect 440393 479604 440459 479714
rect 460321 479606 460387 479716
rect 460693 479616 460759 479726
rect 480503 479584 480569 479694
rect 480875 479594 480941 479704
rect 522909 479633 522975 479743
rect 523281 479643 523347 479753
rect 500459 479506 500525 479616
rect 500831 479496 500897 479606
rect 545802 479510 545868 479620
rect 546174 479500 546240 479610
rect 346982 478252 347092 478318
rect 346992 477880 347102 477946
rect 379051 475499 379117 475609
rect 379423 475509 379489 475619
rect 399541 475532 399607 475642
rect 399913 475542 399979 475652
rect 419783 475472 419849 475582
rect 420155 475482 420221 475592
rect 440021 475501 440087 475611
rect 440393 475511 440459 475621
rect 460321 475513 460387 475623
rect 460693 475523 460759 475633
rect 480503 475491 480569 475601
rect 480875 475501 480941 475611
rect 500491 475509 500557 475619
rect 500863 475519 500929 475629
rect 522941 475382 523007 475492
rect 523313 475372 523379 475482
rect 545855 475418 545921 475528
rect 546227 475408 546293 475518
rect 387914 469723 388024 469789
rect 392806 469723 392916 469789
rect 387924 469351 388034 469417
rect 392816 469351 392926 469417
rect 508976 469023 509086 469089
rect 508986 468651 509096 468717
rect 515023 467765 515133 467831
rect 515033 467393 515143 467459
rect 534386 466945 534496 467011
rect 534376 466573 534486 466639
rect 356026 462172 356136 462238
rect 356036 461800 356146 461866
rect 550370 459665 550480 459731
rect 527531 459536 527641 459602
rect 550360 459293 550470 459359
rect 527521 459164 527631 459230
rect 521414 457098 521524 457164
rect 346996 456998 347106 457064
rect 521424 456726 521534 456792
rect 347006 456626 347116 456692
rect 240701 455849 240811 455915
rect 251423 455827 251533 455893
rect 240711 455477 240821 455543
rect 251433 455455 251543 455521
rect 502200 455171 502310 455237
rect 502210 454799 502320 454865
rect 564164 453285 564230 453395
rect 564536 453295 564602 453405
rect 508964 448972 509074 449038
rect 392796 448771 392906 448837
rect 387875 448703 387985 448769
rect 508974 448600 509084 448666
rect 392806 448399 392916 448465
rect 387885 448331 387995 448397
rect 515060 447564 515170 447630
rect 515070 447192 515180 447258
rect 534376 446545 534486 446611
rect 534366 446173 534476 446239
rect 356000 442179 356110 442245
rect 356010 441807 356120 441873
rect 346968 436390 347078 436456
rect 346978 436018 347088 436084
rect 240621 434332 240731 434398
rect 251406 434046 251516 434112
rect 240631 433960 240741 434026
rect 251416 433674 251526 433740
rect 387904 427660 388014 427726
rect 392828 427679 392938 427745
rect 387914 427288 388024 427354
rect 392838 427307 392948 427373
rect 252958 425977 253024 426087
rect 253330 425967 253396 426077
rect 272904 426042 272970 426152
rect 273276 426032 273342 426142
rect 293185 426076 293251 426186
rect 293557 426066 293623 426176
rect 313334 426066 313400 426176
rect 313706 426056 313772 426166
rect 335541 426041 335607 426151
rect 335913 426051 335979 426161
rect 355531 426037 355597 426147
rect 355903 426047 355969 426157
rect 375494 426131 375560 426241
rect 375866 426141 375932 426251
rect 356005 422225 356115 422291
rect 356015 421853 356125 421919
rect 258312 420479 258378 420589
rect 258684 420469 258750 420579
rect 278446 420512 278512 420622
rect 278818 420502 278884 420612
rect 299123 420518 299189 420628
rect 299495 420508 299561 420618
rect 319451 420470 319517 420580
rect 319823 420460 319889 420570
rect 353761 420469 353827 420579
rect 354133 420479 354199 420589
rect 374104 420539 374170 420649
rect 374476 420549 374542 420659
rect 324544 417112 324654 417178
rect 336554 417037 336664 417103
rect 324554 416740 324664 416806
rect 336564 416665 336674 416731
rect 346912 415756 347022 415822
rect 346922 415384 347032 415450
rect 568046 408878 568112 408988
rect 568418 408868 568484 408978
rect 549553 407130 549663 407196
rect 549543 406758 549653 406824
rect 355994 402190 356104 402256
rect 356004 401818 356114 401884
rect 324542 396322 324652 396388
rect 336579 396384 336689 396450
rect 324552 395950 324662 396016
rect 336589 396012 336699 396078
rect 346940 395078 347050 395144
rect 346950 394706 347060 394772
rect 549570 388086 549680 388152
rect 549560 387714 549670 387780
rect 347446 386614 347512 386724
rect 347818 386604 347884 386714
rect 367462 386643 367528 386753
rect 367834 386633 367900 386743
rect 387274 386633 387340 386743
rect 387646 386623 387712 386733
rect 407533 386631 407599 386741
rect 407905 386621 407971 386731
rect 427809 386686 427875 386796
rect 428181 386676 428247 386786
rect 447968 386666 448034 386776
rect 448340 386656 448406 386766
rect 467970 386661 468036 386771
rect 468342 386651 468408 386761
rect 488088 386645 488154 386755
rect 488460 386635 488526 386745
rect 508218 386668 508284 386778
rect 508590 386658 508656 386768
rect 528327 386682 528393 386792
rect 528699 386672 528765 386782
rect 355974 382126 356084 382192
rect 355984 381754 356094 381820
rect 333077 380647 333143 380757
rect 333449 380637 333515 380747
rect 357656 380655 357722 380765
rect 358028 380645 358094 380755
rect 387103 380613 387169 380723
rect 387475 380603 387541 380713
rect 407681 380644 407747 380754
rect 408053 380634 408119 380744
rect 427655 380619 427721 380729
rect 428027 380609 428093 380719
rect 447901 380623 447967 380733
rect 448273 380613 448339 380723
rect 467885 380690 467951 380800
rect 468257 380680 468323 380790
rect 488300 380615 488366 380725
rect 488672 380605 488738 380715
rect 507983 380687 508049 380797
rect 508355 380677 508421 380787
rect 528353 380621 528419 380731
rect 528725 380611 528791 380721
rect 549368 379428 549478 379494
rect 549378 379056 549488 379122
rect 346926 373796 347036 373862
rect 346936 373424 347046 373490
rect 549329 364242 549439 364308
rect 549339 363870 549449 363936
rect 568202 362495 568268 362605
rect 568574 362485 568640 362595
rect 356031 362143 356141 362209
rect 356041 361771 356151 361837
rect 346926 352946 347036 353012
rect 346936 352574 347046 352640
rect 356031 342140 356141 342206
rect 356041 341768 356151 341834
rect 347010 332350 347120 332416
rect 347020 331978 347130 332044
rect 355955 322138 356065 322204
rect 355965 321766 356075 321832
rect 346982 310482 347092 310548
rect 346992 310110 347102 310176
rect 355993 302117 356103 302183
rect 356003 301745 356113 301811
rect 370828 295924 370894 296034
rect 371200 295934 371266 296044
rect 390837 295941 390903 296051
rect 391209 295951 391275 296061
rect 410843 295912 410909 296022
rect 411215 295922 411281 296032
rect 430839 295988 430905 296098
rect 431211 295998 431277 296108
rect 450856 295955 450922 296065
rect 451228 295965 451294 296075
rect 470858 295980 470924 296090
rect 471230 295990 471296 296100
rect 490853 296013 490919 296123
rect 491225 296023 491291 296133
rect 510846 295969 510912 296079
rect 511218 295979 511284 296089
rect 530831 296013 530897 296123
rect 531203 296023 531269 296133
rect 549547 293375 549657 293441
rect 549557 293003 549667 293069
rect 346940 288824 347050 288890
rect 346950 288452 347060 288518
rect 551449 273906 551515 274016
rect 551821 273916 551887 274026
rect 571912 273866 571978 273976
rect 572284 273876 572350 273986
rect 346898 264044 347008 264110
rect 346908 263672 347018 263738
rect 346982 242670 347092 242736
rect 346992 242298 347102 242364
rect 347010 222794 347120 222860
rect 347020 222422 347130 222488
rect 346954 200966 347064 201032
rect 346964 200594 347074 200660
rect 346968 179932 347078 179998
rect 346978 179560 347088 179626
rect 346926 158544 347036 158610
rect 346936 158172 347046 158238
rect 346870 137198 346980 137264
rect 346880 136826 346990 136892
rect 346926 116064 347036 116130
rect 346936 115692 347046 115758
rect 346954 95454 347064 95520
rect 346964 95082 347074 95148
rect 346940 74772 347050 74838
rect 346950 74400 347060 74466
rect 347010 51192 347120 51258
rect 347020 50820 347130 50886
rect 47990 48776 48056 48886
rect 48362 48786 48428 48896
rect 69284 48836 69350 48946
rect 69656 48846 69722 48956
rect 90650 48762 90716 48872
rect 91022 48772 91088 48882
rect 111710 48806 111776 48916
rect 112082 48816 112148 48926
rect 133032 48850 133098 48960
rect 133404 48860 133470 48970
rect 154590 48820 154656 48930
rect 154962 48830 155028 48940
rect 175796 48792 175862 48902
rect 176168 48802 176234 48912
rect 197178 48850 197244 48960
rect 197550 48860 197616 48970
rect 219072 48762 219138 48872
rect 219444 48772 219510 48882
rect 240058 48732 240124 48842
rect 240430 48742 240496 48852
rect 260560 48792 260626 48902
rect 260932 48802 260998 48912
rect 281372 48894 281438 49004
rect 281744 48904 281810 49014
rect 302562 48688 302628 48798
rect 302934 48698 303000 48808
rect 324110 48724 324176 48834
rect 324482 48734 324548 48844
rect 34578 42938 34688 43004
rect 34588 42566 34698 42632
rect 34578 20840 34688 20906
rect 34588 20468 34698 20534
rect 6548 3452 6614 3562
rect 6920 3462 6986 3572
rect 27740 3512 27806 3622
rect 28112 3522 28178 3632
<< metal1 >>
rect 537809 587971 572320 588573
rect 537809 579323 538411 587971
rect 550705 587051 551307 587971
rect 571718 587062 572320 587971
rect 571876 586892 571954 586904
rect 550865 586861 550943 586873
rect 550861 586751 550871 586861
rect 550937 586751 550947 586861
rect 551237 586851 551315 586863
rect 550865 586739 550943 586751
rect 551233 586741 551243 586851
rect 551309 586741 551319 586851
rect 571872 586782 571882 586892
rect 571948 586782 571958 586892
rect 572248 586882 572326 586894
rect 571876 586770 571954 586782
rect 572244 586772 572254 586882
rect 572320 586772 572330 586882
rect 572248 586760 572326 586772
rect 551237 586729 551315 586741
rect 550709 585241 551311 586439
rect 571723 585241 572325 586467
rect 547170 584639 572326 585241
rect 537803 578721 537809 579323
rect 538411 578721 538417 579323
rect 525158 573235 538424 573237
rect 525158 572635 544549 573235
rect 544736 573225 544846 573229
rect 544724 573219 544858 573225
rect 547170 573221 547772 584639
rect 544724 573153 544736 573219
rect 544846 573153 544858 573219
rect 544724 573147 544858 573153
rect 544736 573143 544846 573147
rect 544726 572853 544836 572857
rect 544714 572847 544848 572853
rect 544714 572781 544726 572847
rect 544836 572781 544848 572847
rect 544714 572775 544848 572781
rect 544726 572771 544836 572775
rect 525158 568164 525760 572635
rect 537822 572633 544549 572635
rect 525314 567981 525392 567993
rect 525310 567871 525320 567981
rect 525386 567871 525396 567981
rect 525686 567971 525764 567983
rect 525314 567859 525392 567871
rect 525682 567861 525692 567971
rect 525758 567861 525768 567971
rect 525686 567849 525764 567861
rect 525158 564049 525760 567606
rect 525158 563447 527213 564049
rect 509388 562231 513451 562833
rect 513762 562669 513872 562673
rect 513750 562663 513884 562669
rect 513750 562597 513762 562663
rect 513872 562597 513884 562663
rect 513750 562591 513884 562597
rect 513762 562587 513872 562591
rect 513752 562297 513862 562301
rect 513740 562291 513874 562297
rect 509388 560581 509990 562231
rect 513740 562225 513752 562291
rect 513862 562225 513874 562291
rect 514051 562238 518526 562840
rect 513740 562219 513874 562225
rect 513752 562215 513862 562219
rect 502344 559977 505253 560579
rect 505449 560576 505559 560580
rect 505437 560570 505571 560576
rect 505437 560504 505449 560570
rect 505559 560504 505571 560570
rect 505437 560498 505571 560504
rect 505449 560494 505559 560498
rect 505439 560204 505549 560208
rect 505427 560198 505561 560204
rect 505427 560132 505439 560198
rect 505549 560132 505561 560198
rect 505427 560126 505561 560132
rect 505439 560122 505549 560126
rect 505821 559979 509990 560581
rect 502344 540003 502946 559977
rect 509388 556160 509990 559979
rect 509388 554242 509408 556160
rect 509938 554242 509990 556160
rect 509388 542389 509990 554242
rect 517924 550499 518526 562238
rect 526606 556182 527208 563447
rect 526598 554236 526608 556182
rect 527208 554236 527218 556182
rect 526606 553273 527208 554236
rect 537822 553293 538424 572633
rect 545105 572619 547772 573221
rect 526606 552671 530737 553273
rect 531032 553115 531142 553119
rect 531020 553109 531154 553115
rect 531020 553043 531032 553109
rect 531142 553043 531154 553109
rect 531020 553037 531154 553043
rect 531032 553033 531142 553037
rect 531317 552987 538424 553293
rect 547170 556178 547772 572619
rect 547170 554212 547182 556178
rect 547758 554212 547772 556178
rect 531022 552743 531132 552747
rect 531010 552737 531144 552743
rect 531010 552671 531022 552737
rect 531132 552671 531144 552737
rect 531317 552691 544585 552987
rect 544746 552976 544856 552980
rect 544734 552970 544868 552976
rect 544734 552904 544746 552970
rect 544856 552904 544868 552970
rect 547170 552961 547772 554212
rect 544734 552898 544868 552904
rect 544746 552894 544856 552898
rect 517924 549897 522315 550499
rect 522511 550498 522621 550502
rect 522499 550492 522633 550498
rect 522499 550426 522511 550492
rect 522621 550426 522633 550492
rect 526606 550485 527208 552671
rect 531010 552665 531144 552671
rect 531022 552661 531132 552665
rect 522499 550420 522633 550426
rect 522511 550416 522621 550420
rect 522501 550126 522611 550130
rect 522489 550120 522623 550126
rect 522489 550054 522501 550120
rect 522611 550054 522623 550120
rect 522489 550048 522623 550054
rect 522501 550044 522611 550048
rect 517924 542393 518526 549897
rect 522891 549883 527208 550485
rect 509388 541787 513463 542389
rect 513742 542227 513852 542231
rect 513730 542221 513864 542227
rect 513730 542155 513742 542221
rect 513852 542155 513864 542221
rect 513730 542149 513864 542155
rect 513742 542145 513852 542149
rect 513732 541855 513842 541859
rect 513720 541849 513854 541855
rect 500443 539631 501045 539637
rect 502344 539631 505375 540003
rect 505559 539988 505669 539992
rect 505547 539982 505681 539988
rect 505547 539916 505559 539982
rect 505669 539916 505681 539982
rect 509388 539973 509990 541787
rect 513720 541783 513732 541849
rect 513842 541783 513854 541849
rect 514029 541791 518526 542393
rect 513720 541777 513854 541783
rect 513732 541773 513842 541777
rect 517924 540212 518526 541791
rect 505547 539910 505681 539916
rect 505559 539906 505669 539910
rect 464231 538845 464237 539447
rect 464839 538845 464845 539447
rect 484622 538955 484628 539557
rect 485230 538955 485236 539557
rect 501045 539401 505375 539631
rect 505549 539616 505659 539620
rect 505537 539610 505671 539616
rect 505537 539544 505549 539610
rect 505659 539544 505671 539610
rect 505537 539538 505671 539544
rect 505549 539534 505659 539538
rect 501045 539029 502946 539401
rect 505967 539371 509990 539973
rect 500443 539023 501045 539029
rect 353946 522265 354488 522268
rect 353946 521723 355823 522265
rect 357540 522237 358082 522238
rect 355991 522117 356101 522121
rect 355979 522111 356113 522117
rect 355979 522045 355991 522111
rect 356101 522045 356113 522111
rect 355979 522039 356113 522045
rect 355991 522035 356101 522039
rect 356001 521745 356111 521749
rect 355989 521739 356123 521745
rect 353946 502339 354488 521723
rect 355989 521673 356001 521739
rect 356111 521673 356123 521739
rect 356391 521695 358082 522237
rect 355989 521667 356123 521673
rect 356001 521663 356111 521667
rect 357540 502339 358082 521695
rect 464237 521667 464839 538845
rect 484628 521667 485230 538955
rect 509388 522407 509990 539371
rect 517864 538396 517874 540212
rect 518574 538396 518584 540212
rect 517924 529729 518526 538396
rect 526606 532039 527208 549883
rect 537822 552385 544585 552691
rect 544736 552604 544846 552608
rect 544724 552598 544858 552604
rect 544724 552532 544736 552598
rect 544846 552532 544858 552598
rect 544724 552526 544858 552532
rect 544736 552522 544846 552526
rect 537822 540294 538424 552385
rect 545149 552359 547772 552961
rect 537822 538328 537834 540294
rect 538410 538328 538424 540294
rect 537822 532741 538424 538328
rect 547170 532778 547772 552359
rect 544751 532750 544861 532754
rect 544739 532744 544873 532750
rect 537822 532139 544573 532741
rect 544739 532678 544751 532744
rect 544861 532678 544873 532744
rect 544739 532672 544873 532678
rect 544751 532668 544861 532672
rect 544741 532378 544851 532382
rect 544729 532372 544863 532378
rect 544729 532306 544741 532372
rect 544851 532306 544863 532372
rect 544729 532300 544863 532306
rect 544741 532296 544851 532300
rect 545161 532176 547772 532778
rect 537822 532043 538424 532139
rect 526606 531437 530679 532039
rect 530987 531870 531097 531874
rect 530975 531864 531109 531870
rect 530975 531798 530987 531864
rect 531097 531798 531109 531864
rect 530975 531792 531109 531798
rect 530987 531788 531097 531792
rect 530977 531498 531087 531502
rect 530965 531492 531099 531498
rect 526606 529737 527208 531437
rect 530965 531426 530977 531492
rect 531087 531426 531099 531492
rect 531271 531441 538424 532043
rect 530965 531420 531099 531426
rect 530977 531416 531087 531420
rect 517924 529127 522371 529729
rect 522560 529721 522670 529725
rect 522548 529715 522682 529721
rect 522548 529649 522560 529715
rect 522670 529649 522682 529715
rect 522548 529643 522682 529649
rect 522560 529639 522670 529643
rect 522550 529349 522660 529353
rect 522538 529343 522672 529349
rect 522538 529277 522550 529343
rect 522660 529277 522672 529343
rect 522538 529271 522672 529277
rect 522550 529267 522660 529271
rect 522947 529136 527208 529737
rect 522947 529135 526442 529136
rect 517924 522414 518526 529127
rect 509388 521805 513445 522407
rect 513739 522256 513849 522260
rect 513727 522250 513861 522256
rect 513727 522184 513739 522250
rect 513849 522184 513861 522250
rect 513727 522178 513861 522184
rect 513739 522174 513849 522178
rect 513729 521884 513839 521888
rect 513717 521878 513851 521884
rect 513717 521812 513729 521878
rect 513839 521812 513851 521878
rect 514031 521812 518526 522414
rect 513717 521806 513851 521812
rect 513729 521802 513839 521806
rect 424093 521065 504698 521667
rect 424093 519369 424695 521065
rect 444108 519417 444710 521065
rect 464290 519486 464892 521065
rect 484628 519458 485230 521065
rect 504096 519478 504698 521065
rect 464449 519330 464527 519342
rect 444266 519247 444344 519259
rect 424253 519188 424331 519200
rect 424249 519078 424259 519188
rect 424325 519078 424335 519188
rect 424625 519178 424703 519190
rect 424253 519066 424331 519078
rect 424621 519068 424631 519178
rect 424697 519068 424707 519178
rect 444262 519137 444272 519247
rect 444338 519137 444348 519247
rect 444638 519237 444716 519249
rect 444266 519125 444344 519137
rect 444634 519127 444644 519237
rect 444710 519127 444720 519237
rect 464445 519220 464455 519330
rect 464521 519220 464531 519330
rect 464821 519320 464899 519332
rect 464449 519208 464527 519220
rect 464817 519210 464827 519320
rect 464893 519210 464903 519320
rect 484781 519291 484859 519303
rect 504255 519298 504333 519310
rect 464821 519198 464899 519210
rect 484777 519181 484787 519291
rect 484853 519181 484863 519291
rect 485153 519281 485231 519293
rect 484781 519169 484859 519181
rect 485149 519171 485159 519281
rect 485225 519171 485235 519281
rect 504251 519188 504261 519298
rect 504327 519188 504337 519298
rect 504627 519288 504705 519300
rect 504255 519176 504333 519188
rect 504623 519178 504633 519288
rect 504699 519178 504709 519288
rect 485153 519159 485231 519171
rect 504627 519166 504705 519178
rect 444638 519115 444716 519127
rect 424625 519056 424703 519068
rect 424103 516881 424705 518769
rect 444108 516881 444710 518839
rect 464290 516881 464892 518926
rect 484628 516881 485230 518888
rect 504098 516881 504700 518874
rect 526606 517499 527208 529136
rect 537822 524181 538424 531441
rect 537530 523347 538424 524181
rect 537530 519612 538132 523347
rect 537684 519443 537762 519455
rect 537680 519333 537690 519443
rect 537756 519333 537766 519443
rect 538056 519433 538134 519445
rect 537684 519321 537762 519333
rect 538052 519323 538062 519433
rect 538128 519323 538138 519433
rect 538056 519311 538134 519323
rect 537541 517499 538143 519023
rect 526606 516897 538143 517499
rect 424093 516279 504700 516881
rect 353946 501797 355817 502339
rect 355956 502208 356066 502212
rect 355944 502202 356078 502208
rect 355944 502136 355956 502202
rect 356066 502136 356078 502202
rect 355944 502130 356078 502136
rect 355956 502126 356066 502130
rect 355966 501836 356076 501840
rect 355954 501830 356088 501836
rect 353946 482379 354488 501797
rect 355954 501764 355966 501830
rect 356076 501764 356088 501830
rect 356313 501797 358082 502339
rect 355954 501758 356088 501764
rect 355966 501754 356076 501758
rect 357540 485147 358082 501797
rect 374598 491783 384731 492325
rect 373616 490680 373726 490684
rect 373604 490674 373738 490680
rect 371709 490630 372251 490641
rect 371709 490088 373320 490630
rect 373604 490608 373616 490674
rect 373726 490608 373738 490674
rect 374609 490642 375151 491783
rect 383268 490678 383378 490682
rect 373604 490602 373738 490608
rect 373616 490598 373726 490602
rect 373626 490308 373736 490312
rect 373614 490302 373748 490308
rect 373614 490236 373626 490302
rect 373736 490236 373748 490302
rect 373614 490230 373748 490236
rect 373626 490226 373736 490230
rect 373894 490100 375151 490642
rect 383256 490672 383390 490678
rect 381671 490094 382966 490636
rect 383256 490606 383268 490672
rect 383378 490606 383390 490672
rect 384189 490660 384731 491783
rect 392808 490773 392918 490777
rect 392796 490767 392930 490773
rect 387905 490759 388015 490763
rect 387893 490753 388027 490759
rect 383256 490600 383390 490606
rect 383268 490596 383378 490600
rect 383278 490306 383388 490310
rect 383266 490300 383400 490306
rect 383266 490234 383278 490300
rect 383388 490234 383400 490300
rect 383266 490228 383400 490234
rect 383278 490224 383388 490228
rect 383564 490118 384731 490660
rect 386579 490189 387595 490731
rect 387893 490687 387905 490753
rect 388015 490687 388027 490753
rect 387893 490681 388027 490687
rect 387905 490677 388015 490681
rect 387915 490387 388025 490391
rect 387903 490381 388037 490387
rect 387903 490315 387915 490381
rect 388025 490315 388037 490381
rect 387903 490309 388037 490315
rect 387915 490305 388025 490309
rect 388195 490216 389225 490758
rect 371709 488181 372251 490088
rect 381671 488181 382213 490094
rect 371709 487639 382213 488181
rect 375489 485289 376031 485295
rect 360443 485147 360985 485153
rect 357540 484605 360443 485147
rect 357540 482381 358082 484605
rect 360443 484599 360985 484605
rect 386579 485219 387121 490189
rect 353946 481837 355843 482379
rect 356018 482264 356128 482268
rect 356006 482258 356140 482264
rect 356006 482192 356018 482258
rect 356128 482192 356140 482258
rect 356006 482186 356140 482192
rect 356018 482182 356128 482186
rect 356028 481892 356138 481896
rect 356016 481886 356150 481892
rect 345480 477897 346807 478439
rect 346982 478324 347092 478328
rect 346970 478318 347104 478324
rect 346970 478252 346982 478318
rect 347092 478252 347104 478318
rect 346970 478246 347104 478252
rect 346982 478242 347092 478246
rect 346992 477952 347102 477956
rect 346980 477946 347114 477952
rect 345480 457185 346022 477897
rect 346980 477880 346992 477946
rect 347102 477880 347114 477946
rect 347379 477899 348785 478441
rect 346980 477874 347114 477880
rect 346992 477870 347102 477874
rect 348243 457187 348785 477899
rect 353946 472981 354488 481837
rect 356016 481820 356028 481886
rect 356138 481820 356150 481886
rect 356415 481839 358082 482381
rect 356016 481814 356150 481820
rect 356028 481810 356138 481814
rect 352775 472439 352781 472981
rect 353323 472439 354488 472981
rect 345480 456643 346821 457185
rect 346996 457070 347106 457074
rect 346984 457064 347118 457070
rect 346984 456998 346996 457064
rect 347106 456998 347118 457064
rect 346984 456992 347118 456998
rect 346996 456988 347106 456992
rect 347006 456698 347116 456702
rect 346994 456692 347128 456698
rect 240701 455921 240811 455925
rect 238866 455377 240432 455918
rect 240689 455915 240823 455921
rect 240689 455849 240701 455915
rect 240811 455849 240823 455915
rect 251423 455899 251533 455903
rect 240689 455843 240823 455849
rect 240701 455839 240811 455843
rect 240711 455549 240821 455553
rect 240699 455543 240833 455549
rect 240699 455477 240711 455543
rect 240821 455477 240833 455543
rect 240699 455471 240833 455477
rect 240711 455467 240821 455471
rect 238866 434363 239407 455377
rect 240974 455353 242560 455894
rect 251411 455893 251545 455899
rect 240621 434404 240731 434408
rect 240609 434398 240743 434404
rect 238866 433822 240338 434363
rect 240609 434332 240621 434398
rect 240731 434332 240743 434398
rect 242019 434361 242560 455353
rect 240609 434326 240743 434332
rect 240621 434322 240731 434326
rect 240631 434032 240741 434036
rect 240619 434026 240753 434032
rect 240619 433960 240631 434026
rect 240741 433960 240753 434026
rect 240619 433954 240753 433960
rect 240631 433950 240741 433954
rect 238866 430259 239407 433822
rect 240912 433820 242560 434361
rect 249243 455318 251115 455860
rect 251411 455827 251423 455893
rect 251533 455827 251545 455893
rect 251411 455821 251545 455827
rect 251423 455817 251533 455821
rect 251433 455527 251543 455531
rect 251421 455521 251555 455527
rect 251421 455455 251433 455521
rect 251543 455455 251555 455521
rect 251421 455449 251555 455455
rect 251433 455445 251543 455449
rect 251703 455347 255815 455889
rect 249243 434082 249785 455318
rect 251406 434118 251516 434122
rect 251394 434112 251528 434118
rect 238860 429718 238866 430259
rect 239407 429718 239413 430259
rect 242019 415901 242560 433820
rect 249236 433540 251133 434082
rect 251394 434046 251406 434112
rect 251516 434046 251528 434112
rect 255273 434088 255815 455347
rect 251394 434040 251528 434046
rect 251406 434036 251516 434040
rect 251416 433746 251526 433750
rect 251404 433740 251538 433746
rect 251404 433674 251416 433740
rect 251526 433674 251538 433740
rect 251404 433668 251538 433674
rect 251416 433664 251526 433668
rect 251689 433546 255815 434088
rect 249236 433424 249777 433540
rect 249235 430379 249777 433424
rect 249229 429837 249235 430379
rect 249777 429837 249783 430379
rect 252980 430363 253522 430369
rect 252980 426336 253522 429821
rect 252952 426087 253030 426099
rect 252948 425977 252958 426087
rect 253024 425977 253034 426087
rect 253324 426077 253402 426089
rect 252952 425965 253030 425977
rect 253320 425967 253330 426077
rect 253396 425967 253406 426077
rect 253324 425955 253402 425967
rect 252972 415912 253512 425832
rect 252966 415372 252972 415912
rect 253512 415372 253518 415912
rect 255273 415727 255815 433546
rect 345480 436577 346022 456643
rect 346994 456626 347006 456692
rect 347116 456626 347128 456692
rect 347393 456645 348785 457187
rect 346994 456620 347128 456626
rect 347006 456616 347116 456620
rect 348243 436579 348785 456645
rect 353946 462365 354488 472439
rect 357540 462375 358082 481839
rect 375489 474787 376031 484747
rect 386095 485213 387121 485219
rect 386637 484671 387121 485213
rect 386095 484665 387121 484671
rect 380557 481753 381099 481779
rect 380557 481211 384638 481753
rect 380557 476939 381099 481211
rect 384096 479890 384638 481211
rect 384080 479710 384158 479722
rect 384452 479720 384530 479732
rect 384076 479600 384086 479710
rect 384152 479600 384162 479710
rect 384448 479610 384458 479720
rect 384524 479610 384534 479720
rect 384080 479588 384158 479600
rect 384452 479598 384530 479610
rect 384100 478639 384642 479320
rect 386579 478639 387121 484665
rect 384100 478097 387121 478639
rect 379046 476397 381099 476939
rect 379046 475789 379588 476397
rect 379045 475609 379123 475621
rect 379417 475619 379495 475631
rect 379041 475499 379051 475609
rect 379117 475499 379127 475609
rect 379413 475509 379423 475619
rect 379489 475509 379499 475619
rect 379045 475487 379123 475499
rect 379417 475497 379495 475509
rect 379068 474787 379610 475204
rect 375489 474245 379610 474787
rect 380557 473159 381099 476397
rect 380551 472617 380557 473159
rect 381099 472617 381105 473159
rect 386579 469780 387121 478097
rect 388683 473083 389225 490216
rect 391257 490198 392525 490740
rect 392796 490701 392808 490767
rect 392918 490701 392930 490767
rect 392796 490695 392930 490701
rect 392808 490691 392918 490695
rect 392818 490401 392928 490405
rect 392806 490395 392940 490401
rect 392806 490329 392818 490395
rect 392928 490329 392940 490395
rect 392806 490323 392940 490329
rect 392818 490319 392928 490323
rect 393081 490198 394227 490740
rect 390329 485211 390871 485217
rect 391257 485211 391799 490198
rect 390871 484669 391801 485211
rect 390329 484663 390871 484669
rect 389491 473083 390033 473089
rect 388683 472541 389491 473083
rect 387914 469795 388024 469799
rect 387902 469789 388036 469795
rect 386579 469238 387613 469780
rect 387902 469723 387914 469789
rect 388024 469723 388036 469789
rect 388683 469774 389225 472541
rect 389491 472535 390033 472541
rect 388300 469773 389225 469774
rect 387902 469717 388036 469723
rect 387914 469713 388024 469717
rect 387924 469423 388034 469427
rect 387912 469417 388046 469423
rect 387912 469351 387924 469417
rect 388034 469351 388046 469417
rect 387912 469345 388046 469351
rect 387924 469341 388034 469345
rect 388223 469231 389225 469773
rect 391259 469780 391801 484669
rect 393685 473157 394227 490198
rect 458519 485307 459121 485313
rect 434805 485229 435407 485235
rect 428641 485221 429183 485227
rect 400223 485181 400765 485187
rect 398067 484639 400223 485181
rect 398067 478677 398609 484639
rect 400223 484633 400765 484639
rect 417907 484679 428641 485221
rect 399570 480859 402357 481401
rect 399570 479920 400112 480859
rect 399535 479735 399613 479747
rect 399907 479745 399985 479757
rect 399531 479625 399541 479735
rect 399607 479625 399617 479735
rect 399903 479635 399913 479745
rect 399979 479635 399989 479745
rect 399535 479613 399613 479625
rect 399907 479623 399985 479635
rect 399570 478677 400112 479335
rect 398067 478135 400112 478677
rect 398067 474879 398609 478135
rect 401815 477111 402357 480859
rect 399570 476569 402357 477111
rect 399570 475838 400112 476569
rect 399535 475642 399613 475654
rect 399907 475652 399985 475664
rect 399531 475532 399541 475642
rect 399607 475532 399617 475642
rect 399903 475542 399913 475652
rect 399979 475542 399989 475652
rect 399535 475520 399613 475532
rect 399907 475530 399985 475542
rect 399565 474879 400107 475263
rect 398067 474337 400107 474879
rect 394697 473157 395239 473163
rect 393685 472615 394697 473157
rect 392806 469795 392916 469799
rect 392794 469789 392928 469795
rect 391259 469238 392499 469780
rect 392794 469723 392806 469789
rect 392916 469723 392928 469789
rect 393685 469788 394227 472615
rect 394697 472609 395239 472615
rect 400591 473109 401133 473115
rect 401815 473109 402357 476569
rect 417907 478783 418449 484679
rect 428641 484673 429183 484679
rect 419800 480645 422521 481187
rect 419800 479855 420342 480645
rect 419777 479675 419855 479687
rect 420149 479685 420227 479697
rect 419773 479565 419783 479675
rect 419849 479565 419859 479675
rect 420145 479575 420155 479685
rect 420221 479575 420231 479685
rect 419777 479553 419855 479565
rect 420149 479563 420227 479575
rect 419800 478783 420342 479286
rect 417907 478744 420342 478783
rect 417907 478241 420341 478744
rect 417907 474607 418449 478241
rect 421979 476759 422521 480645
rect 419799 476217 422521 476759
rect 419804 475780 420346 476217
rect 419777 475582 419855 475594
rect 420149 475592 420227 475604
rect 419773 475472 419783 475582
rect 419849 475472 419859 475582
rect 420145 475482 420155 475592
rect 420221 475482 420231 475592
rect 419777 475460 419855 475472
rect 420149 475470 420227 475482
rect 419804 474607 420346 475183
rect 417907 474065 420346 474607
rect 401133 472567 402357 473109
rect 421979 473109 422521 476217
rect 434805 478725 435407 484627
rect 440018 480579 443838 481181
rect 440018 479898 440620 480579
rect 440015 479704 440093 479716
rect 440387 479714 440465 479726
rect 440011 479594 440021 479704
rect 440087 479594 440097 479704
rect 440383 479604 440393 479714
rect 440459 479604 440469 479714
rect 440015 479582 440093 479594
rect 440387 479592 440465 479604
rect 440004 478725 440606 479306
rect 434805 478123 440606 478725
rect 434805 474565 435407 478123
rect 443236 476825 443838 480579
rect 440022 476223 443838 476825
rect 440022 475806 440624 476223
rect 440015 475611 440093 475623
rect 440387 475621 440465 475633
rect 440011 475501 440021 475611
rect 440087 475501 440097 475611
rect 440383 475511 440393 475621
rect 440459 475511 440469 475621
rect 440015 475489 440093 475501
rect 440387 475499 440465 475511
rect 440016 475109 440618 475198
rect 440015 474608 440618 475109
rect 440015 474565 440617 474608
rect 434805 473963 440617 474565
rect 428295 473109 428837 473115
rect 421979 472567 428295 473109
rect 400591 472561 401133 472567
rect 428295 472561 428837 472567
rect 443236 473047 443838 476223
rect 458519 478859 459121 484705
rect 464290 485157 464892 516279
rect 484628 485195 485230 516279
rect 534334 508958 534444 508962
rect 531125 508352 534028 508954
rect 534322 508952 534456 508958
rect 534322 508886 534334 508952
rect 534444 508886 534456 508952
rect 534322 508880 534456 508886
rect 534334 508876 534444 508880
rect 534344 508586 534454 508590
rect 534332 508580 534466 508586
rect 534332 508514 534344 508580
rect 534454 508514 534466 508580
rect 534332 508508 534466 508514
rect 534344 508504 534454 508508
rect 534619 508357 537545 508959
rect 511844 507491 514721 508093
rect 515038 507939 515148 507943
rect 515026 507933 515160 507939
rect 515026 507867 515038 507933
rect 515148 507867 515160 507933
rect 515026 507861 515160 507867
rect 515038 507857 515148 507861
rect 515028 507567 515138 507571
rect 515016 507561 515150 507567
rect 515016 507495 515028 507561
rect 515138 507495 515150 507561
rect 515325 507499 518395 508101
rect 511844 506543 512446 507491
rect 515016 507489 515150 507495
rect 515028 507485 515138 507489
rect 508942 506531 509052 506535
rect 508930 506525 509064 506531
rect 505369 505921 508757 506523
rect 508930 506459 508942 506525
rect 509052 506459 509064 506525
rect 508930 506453 509064 506459
rect 508942 506449 509052 506453
rect 508932 506159 509042 506163
rect 508920 506153 509054 506159
rect 508920 506087 508932 506153
rect 509042 506087 509054 506153
rect 508920 506081 509054 506087
rect 508932 506077 509042 506081
rect 509343 505941 512446 506543
rect 498503 499886 501872 500488
rect 505369 500461 505971 505921
rect 502178 500332 502288 500336
rect 502166 500326 502300 500332
rect 502166 500260 502178 500326
rect 502288 500260 502300 500326
rect 502166 500254 502300 500260
rect 502178 500250 502288 500254
rect 502168 499960 502278 499964
rect 502156 499954 502290 499960
rect 502156 499888 502168 499954
rect 502278 499888 502290 499954
rect 464290 484549 464892 484555
rect 475009 485127 475611 485133
rect 484622 484593 484628 485195
rect 485230 484593 485236 485195
rect 498503 485111 499105 499886
rect 502156 499882 502290 499888
rect 502168 499878 502278 499882
rect 502461 499859 505971 500461
rect 505369 488623 505971 499859
rect 505369 488021 507297 488623
rect 506695 486479 507297 488021
rect 511844 487883 512446 505941
rect 517793 498409 518395 507499
rect 531125 501411 531727 508352
rect 531125 500803 531727 500809
rect 517793 497807 521195 498409
rect 521392 498405 521502 498409
rect 521380 498399 521514 498405
rect 521380 498333 521392 498399
rect 521502 498333 521514 498399
rect 521380 498327 521514 498333
rect 521392 498323 521502 498327
rect 521382 498033 521492 498037
rect 521370 498027 521504 498033
rect 521370 497961 521382 498027
rect 521492 497961 521504 498027
rect 521370 497955 521504 497961
rect 521382 497951 521492 497955
rect 521777 497833 524892 498435
rect 517793 492219 518395 497807
rect 524290 496161 524892 497833
rect 524290 495559 527149 496161
rect 536943 496160 537545 508357
rect 564212 499797 568479 500427
rect 564212 498164 564842 499797
rect 564224 497870 564302 497882
rect 564220 497760 564230 497870
rect 564296 497760 564306 497870
rect 564596 497860 564674 497872
rect 564224 497748 564302 497760
rect 564592 497750 564602 497860
rect 564668 497750 564678 497860
rect 564596 497738 564674 497750
rect 527466 496007 527576 496011
rect 527454 496001 527588 496007
rect 527454 495935 527466 496001
rect 527576 495935 527588 496001
rect 527454 495929 527588 495935
rect 527466 495925 527576 495929
rect 527456 495635 527566 495639
rect 527444 495629 527578 495635
rect 527444 495563 527456 495629
rect 527566 495563 527578 495629
rect 517793 491617 522606 492219
rect 511844 487281 514699 487883
rect 517793 487881 518395 491617
rect 515001 487738 515111 487742
rect 514989 487732 515123 487738
rect 514989 487666 515001 487732
rect 515111 487666 515123 487732
rect 514989 487660 515123 487666
rect 515001 487656 515111 487660
rect 514991 487366 515101 487370
rect 514979 487360 515113 487366
rect 514979 487294 514991 487360
rect 515101 487294 515113 487360
rect 514979 487288 515113 487294
rect 514991 487284 515101 487288
rect 511844 486485 512446 487281
rect 515279 487279 518395 487881
rect 508954 486480 509064 486484
rect 506695 485877 508767 486479
rect 508942 486474 509076 486480
rect 508942 486408 508954 486474
rect 509064 486408 509076 486474
rect 508942 486402 509076 486408
rect 508954 486398 509064 486402
rect 508944 486108 509054 486112
rect 508932 486102 509066 486108
rect 508932 486036 508944 486102
rect 509054 486036 509066 486102
rect 508932 486030 509066 486036
rect 508944 486026 509054 486030
rect 509343 485883 512446 486485
rect 504627 485165 505229 485171
rect 460316 481435 462687 481439
rect 460316 480837 462737 481435
rect 460316 479914 460918 480837
rect 460315 479716 460393 479728
rect 460687 479726 460765 479738
rect 460311 479606 460321 479716
rect 460387 479606 460397 479716
rect 460683 479616 460693 479726
rect 460759 479616 460769 479726
rect 460315 479594 460393 479606
rect 460687 479604 460765 479616
rect 460312 478859 460914 479312
rect 458519 478257 460914 478859
rect 458519 474797 459121 478257
rect 462135 476931 462737 480837
rect 460318 476329 462737 476931
rect 460318 475810 460920 476329
rect 460315 475623 460393 475635
rect 460687 475633 460765 475645
rect 460311 475513 460321 475623
rect 460387 475513 460397 475623
rect 460683 475523 460693 475633
rect 460759 475523 460769 475633
rect 460315 475501 460393 475513
rect 460687 475511 460765 475523
rect 460300 474797 460902 475210
rect 458519 474195 460909 474797
rect 462135 473059 462737 476329
rect 475009 478753 475611 484525
rect 498497 484509 498503 485111
rect 499105 484509 499111 485111
rect 504627 481579 505229 484563
rect 480491 480473 485899 481075
rect 480506 479876 481108 480473
rect 480497 479694 480575 479706
rect 480869 479704 480947 479716
rect 480493 479584 480503 479694
rect 480569 479584 480579 479694
rect 480865 479594 480875 479704
rect 480941 479594 480951 479704
rect 480497 479572 480575 479584
rect 480869 479582 480947 479594
rect 480496 478753 481098 479284
rect 475009 478151 481098 478753
rect 475009 474789 475611 478151
rect 485297 476891 485899 480473
rect 500456 480977 505229 481579
rect 500456 479924 501058 480977
rect 500453 479616 500531 479628
rect 500449 479506 500459 479616
rect 500525 479506 500535 479616
rect 500825 479606 500903 479618
rect 500453 479494 500531 479506
rect 500821 479496 500831 479606
rect 500897 479496 500907 479606
rect 500825 479484 500903 479496
rect 500458 477887 501060 479334
rect 500458 477866 501086 477887
rect 480500 476289 485899 476891
rect 480500 475794 481102 476289
rect 480497 475601 480575 475613
rect 480869 475611 480947 475623
rect 480493 475491 480503 475601
rect 480569 475491 480579 475601
rect 480865 475501 480875 475611
rect 480941 475501 480951 475611
rect 480497 475479 480575 475491
rect 480869 475489 480947 475501
rect 480490 474789 481092 475184
rect 475009 474187 481092 474789
rect 445483 473047 446085 473053
rect 443236 472445 445483 473047
rect 485297 473103 485899 476289
rect 497352 477238 501086 477866
rect 497352 473194 497980 477238
rect 500458 477211 501086 477238
rect 500484 475794 501086 477211
rect 500485 475619 500563 475631
rect 500857 475629 500935 475641
rect 500481 475509 500491 475619
rect 500557 475509 500567 475619
rect 500853 475519 500863 475629
rect 500929 475519 500939 475629
rect 500485 475497 500563 475509
rect 500857 475507 500935 475519
rect 500479 474485 501081 475205
rect 504627 474485 505229 480977
rect 500479 473883 505229 474485
rect 497352 472560 497980 472566
rect 503860 472998 504488 473004
rect 506695 473001 507297 485877
rect 511844 485215 512446 485883
rect 511838 484613 511844 485215
rect 512446 484613 512452 485215
rect 518207 484585 518213 485215
rect 518843 484585 518849 485215
rect 518213 478003 518843 484585
rect 522004 480973 522606 491617
rect 524290 485159 524892 495559
rect 527444 495557 527578 495563
rect 527746 495558 537545 496160
rect 527456 495553 527566 495557
rect 531125 491757 531727 491763
rect 531125 488547 531727 491155
rect 534344 488558 534454 488562
rect 536943 488561 537545 495558
rect 534332 488552 534466 488558
rect 531125 487945 534041 488547
rect 534332 488486 534344 488552
rect 534454 488486 534466 488552
rect 534332 488480 534466 488486
rect 534344 488476 534454 488480
rect 534354 488186 534464 488190
rect 534342 488180 534476 488186
rect 534342 488114 534354 488180
rect 534464 488114 534476 488180
rect 534342 488108 534476 488114
rect 534354 488104 534464 488108
rect 534641 487959 537545 488561
rect 530389 485173 530991 485179
rect 531125 485173 531727 487945
rect 531891 485221 532521 485227
rect 524284 484557 524290 485159
rect 524892 484557 524898 485159
rect 530991 484591 531891 485173
rect 530991 484571 532521 484591
rect 530389 484565 530991 484571
rect 524525 480973 525127 480976
rect 522004 480371 525127 480973
rect 522004 480355 522606 480371
rect 522900 479928 523502 480371
rect 522903 479743 522981 479755
rect 523275 479753 523353 479765
rect 522899 479633 522909 479743
rect 522975 479633 522985 479743
rect 523271 479643 523281 479753
rect 523347 479643 523357 479753
rect 522903 479621 522981 479633
rect 523275 479631 523353 479643
rect 522906 478107 523508 479328
rect 522906 478003 523536 478107
rect 518213 477373 523536 478003
rect 522906 477211 523536 477373
rect 522934 475800 523536 477211
rect 522935 475492 523013 475504
rect 522931 475382 522941 475492
rect 523007 475382 523017 475492
rect 523307 475482 523385 475494
rect 522935 475370 523013 475382
rect 523303 475372 523313 475482
rect 523379 475372 523389 475482
rect 523307 475360 523385 475372
rect 522944 473097 523546 475226
rect 524525 473097 525127 480371
rect 485297 472495 485899 472501
rect 462135 472451 462737 472457
rect 445483 472439 446085 472445
rect 392794 469717 392928 469723
rect 392806 469713 392916 469717
rect 392816 469423 392926 469427
rect 392804 469417 392938 469423
rect 392804 469351 392816 469417
rect 392926 469351 392938 469417
rect 392804 469345 392938 469351
rect 392816 469341 392926 469345
rect 393105 469246 394227 469788
rect 393685 469243 394227 469246
rect 506689 472399 506695 473001
rect 507297 472399 507303 473001
rect 518229 472485 518235 473087
rect 518837 472485 518843 473087
rect 522934 472495 522944 473097
rect 525127 472495 525137 473097
rect 353946 461823 355831 462365
rect 356026 462244 356136 462248
rect 356014 462238 356148 462244
rect 356014 462172 356026 462238
rect 356136 462172 356148 462238
rect 356014 462166 356148 462172
rect 356026 462162 356136 462166
rect 356036 461872 356146 461876
rect 356024 461866 356158 461872
rect 353946 442359 354488 461823
rect 356024 461800 356036 461866
rect 356146 461800 356158 461866
rect 356461 461833 358082 462375
rect 356024 461794 356158 461800
rect 356036 461790 356146 461794
rect 357540 442375 358082 461833
rect 503860 455262 504488 472370
rect 506695 469236 507297 472399
rect 506695 468634 508803 469236
rect 508976 469095 509086 469099
rect 508964 469089 509098 469095
rect 508964 469023 508976 469089
rect 509086 469023 509098 469089
rect 508964 469017 509098 469023
rect 508976 469013 509086 469017
rect 508986 468723 509096 468727
rect 508974 468717 509108 468723
rect 508974 468651 508986 468717
rect 509096 468651 509108 468717
rect 508974 468645 509108 468651
rect 508986 468641 509096 468645
rect 509394 468640 510884 469242
rect 497210 454616 501886 455244
rect 502200 455243 502310 455247
rect 502188 455237 502322 455243
rect 502188 455171 502200 455237
rect 502310 455171 502322 455237
rect 502188 455165 502322 455171
rect 502200 455161 502310 455165
rect 502210 454871 502320 454875
rect 502198 454865 502332 454871
rect 502198 454799 502210 454865
rect 502320 454799 502332 454865
rect 502198 454793 502332 454799
rect 502210 454789 502320 454793
rect 502480 454634 504488 455262
rect 510283 468398 510884 468640
rect 392796 448843 392906 448847
rect 392784 448837 392918 448843
rect 387875 448775 387985 448779
rect 387863 448769 387997 448775
rect 353946 441817 355831 442359
rect 356000 442251 356110 442255
rect 355988 442245 356122 442251
rect 355988 442179 356000 442245
rect 356110 442179 356122 442245
rect 355988 442173 356122 442179
rect 356000 442169 356110 442173
rect 356010 441879 356120 441883
rect 355998 441873 356132 441879
rect 353946 441787 354488 441817
rect 355998 441807 356010 441873
rect 356120 441807 356132 441873
rect 356407 441833 358082 442375
rect 355998 441801 356132 441807
rect 356010 441797 356120 441801
rect 345480 436035 346793 436577
rect 346968 436462 347078 436466
rect 346956 436456 347090 436462
rect 346956 436390 346968 436456
rect 347078 436390 347090 436456
rect 346956 436384 347090 436390
rect 346968 436380 347078 436384
rect 346978 436090 347088 436094
rect 346966 436084 347100 436090
rect 258332 429822 258338 430362
rect 258878 429822 258884 430362
rect 272940 430299 273482 430305
rect 258338 420854 258878 429822
rect 278444 429801 278450 430343
rect 278992 429801 278998 430343
rect 293208 429813 293214 430355
rect 293756 429813 293762 430355
rect 272940 426398 273482 429757
rect 272898 426152 272976 426164
rect 272894 426042 272904 426152
rect 272970 426042 272980 426152
rect 273270 426142 273348 426154
rect 272898 426030 272976 426042
rect 273266 426032 273276 426142
rect 273342 426032 273352 426142
rect 273270 426020 273348 426032
rect 258306 420589 258384 420601
rect 258302 420479 258312 420589
rect 258378 420479 258388 420589
rect 258678 420579 258756 420591
rect 258306 420467 258384 420479
rect 258674 420469 258684 420579
rect 258750 420469 258760 420579
rect 258678 420457 258756 420469
rect 242019 415354 242560 415360
rect 258336 415876 258876 420318
rect 258336 415330 258876 415336
rect 272932 415809 273474 425855
rect 278450 420897 278992 429801
rect 293214 426463 293756 429813
rect 299156 429713 299162 430255
rect 299704 429713 299710 430255
rect 313348 430191 313890 430197
rect 293179 426186 293257 426198
rect 293175 426076 293185 426186
rect 293251 426076 293261 426186
rect 293551 426176 293629 426188
rect 293179 426064 293257 426076
rect 293547 426066 293557 426176
rect 293623 426066 293633 426176
rect 293551 426054 293629 426066
rect 278440 420622 278518 420634
rect 278436 420512 278446 420622
rect 278512 420512 278522 420622
rect 278812 420612 278890 420624
rect 278440 420500 278518 420512
rect 278808 420502 278818 420612
rect 278884 420502 278894 420612
rect 278812 420490 278890 420502
rect 278450 415815 278992 420339
rect 293214 415789 293756 425895
rect 299162 420901 299704 429713
rect 313348 426453 313890 429649
rect 319470 429615 319476 430157
rect 320018 429615 320024 430157
rect 322079 429673 322085 430215
rect 322627 429673 322633 430215
rect 335388 429711 335394 430253
rect 335936 429711 335942 430253
rect 313328 426176 313406 426188
rect 313324 426066 313334 426176
rect 313400 426066 313410 426176
rect 313700 426166 313778 426178
rect 313328 426054 313406 426066
rect 313696 426056 313706 426166
rect 313772 426056 313782 426166
rect 313700 426044 313778 426056
rect 299117 420628 299195 420640
rect 299113 420518 299123 420628
rect 299189 420518 299199 420628
rect 299489 420618 299567 420630
rect 299117 420506 299195 420518
rect 299485 420508 299495 420618
rect 299561 420508 299571 420618
rect 299489 420496 299567 420508
rect 299136 415813 299678 420375
rect 313354 415871 313896 425907
rect 319476 420847 320018 429615
rect 319445 420580 319523 420592
rect 319441 420470 319451 420580
rect 319517 420470 319527 420580
rect 319817 420570 319895 420582
rect 319445 420458 319523 420470
rect 319813 420460 319823 420570
rect 319889 420460 319899 420570
rect 319817 420448 319895 420460
rect 319466 415947 320008 420323
rect 322085 417138 322627 429673
rect 335394 426431 335936 429711
rect 335535 426151 335613 426163
rect 335907 426161 335985 426173
rect 335531 426041 335541 426151
rect 335607 426041 335617 426151
rect 335903 426051 335913 426161
rect 335979 426051 335989 426161
rect 335535 426029 335613 426041
rect 335907 426039 335985 426051
rect 335404 423817 335946 425862
rect 328033 423275 335946 423817
rect 324544 417184 324654 417188
rect 324532 417178 324666 417184
rect 322085 416596 324256 417138
rect 324532 417112 324544 417178
rect 324654 417112 324666 417178
rect 328033 417166 328575 423275
rect 332869 420847 333411 420853
rect 324532 417106 324666 417112
rect 324544 417102 324654 417106
rect 324554 416812 324664 416816
rect 324542 416806 324676 416812
rect 324542 416740 324554 416806
rect 324664 416740 324676 416806
rect 324542 416734 324676 416740
rect 324554 416730 324664 416734
rect 324836 416624 328701 417166
rect 278450 415267 278992 415273
rect 272932 415261 273474 415267
rect 293208 415247 293214 415789
rect 293756 415247 293762 415789
rect 313348 415329 313354 415871
rect 313896 415329 313902 415871
rect 319460 415405 319466 415947
rect 320008 415405 320014 415947
rect 328159 415901 328701 416624
rect 332869 417080 333411 420305
rect 336554 417109 336664 417113
rect 336542 417103 336676 417109
rect 332869 416538 336266 417080
rect 336542 417037 336554 417103
rect 336664 417037 336676 417103
rect 336542 417031 336676 417037
rect 336554 417027 336664 417031
rect 336564 416737 336674 416741
rect 336552 416731 336686 416737
rect 336552 416665 336564 416731
rect 336674 416665 336686 416731
rect 336552 416659 336686 416665
rect 336564 416655 336674 416659
rect 336844 416546 340417 417088
rect 328153 415359 328159 415901
rect 328701 415359 328707 415901
rect 339875 415863 340417 416546
rect 345480 416210 346022 436035
rect 346966 436018 346978 436084
rect 347088 436018 347100 436084
rect 347365 436037 348785 436579
rect 346966 436012 347100 436018
rect 346978 436008 347088 436012
rect 348243 430698 348785 436037
rect 348084 429382 348094 430698
rect 348522 429382 348785 430698
rect 357540 430443 358082 441833
rect 385933 448206 387583 448748
rect 387863 448703 387875 448769
rect 387985 448703 387997 448769
rect 387863 448697 387997 448703
rect 387875 448693 387985 448697
rect 387885 448403 387995 448407
rect 387873 448397 388007 448403
rect 387873 448331 387885 448397
rect 387995 448331 388007 448397
rect 387873 448325 388007 448331
rect 387885 448321 387995 448325
rect 388181 448215 389159 448757
rect 360001 430443 360543 430445
rect 362171 430443 362713 430449
rect 357540 430439 362171 430443
rect 339869 415321 339875 415863
rect 340417 415321 340423 415863
rect 299136 415265 299678 415271
rect 255273 415179 255815 415185
rect 345480 414894 345550 416210
rect 345978 415943 346022 416210
rect 348243 415945 348785 429382
rect 353636 430275 354787 430291
rect 353636 430269 354899 430275
rect 353636 429749 354357 430269
rect 353636 420851 354178 429749
rect 354899 429727 355932 430269
rect 354357 429721 354899 429727
rect 355390 426447 355932 429727
rect 357540 429897 360001 430439
rect 360543 429901 362171 430439
rect 385933 430287 386475 448206
rect 375352 430195 375894 430201
rect 355525 426147 355603 426159
rect 355897 426157 355975 426169
rect 355521 426037 355531 426147
rect 355597 426037 355607 426147
rect 355893 426047 355903 426157
rect 355969 426047 355979 426157
rect 355525 426025 355603 426037
rect 355897 426035 355975 426047
rect 355390 424503 355932 425869
rect 355065 423961 355932 424503
rect 355065 422435 355607 423961
rect 355065 421893 355887 422435
rect 357540 422409 358082 429897
rect 360001 429891 360543 429897
rect 362171 429895 362713 429901
rect 373944 429649 373950 430191
rect 374492 429649 374498 430191
rect 385927 429745 385933 430287
rect 386475 429745 386481 430287
rect 356005 422297 356115 422301
rect 355993 422291 356127 422297
rect 355993 422225 356005 422291
rect 356115 422225 356127 422291
rect 355993 422219 356127 422225
rect 356005 422215 356115 422219
rect 356015 421925 356125 421929
rect 356003 421919 356137 421925
rect 353755 420579 353833 420591
rect 354127 420589 354205 420601
rect 353751 420469 353761 420579
rect 353827 420469 353837 420579
rect 354123 420479 354133 420589
rect 354199 420479 354209 420589
rect 353755 420457 353833 420469
rect 354127 420467 354205 420479
rect 345978 415401 346737 415943
rect 346912 415828 347022 415832
rect 346900 415822 347034 415828
rect 346900 415756 346912 415822
rect 347022 415756 347034 415822
rect 346900 415750 347034 415756
rect 346912 415746 347022 415750
rect 346922 415456 347032 415460
rect 346910 415450 347044 415456
rect 345978 414894 346022 415401
rect 346910 415384 346922 415450
rect 347032 415384 347044 415450
rect 347309 415403 348785 415945
rect 353626 415781 354168 420293
rect 346910 415378 347044 415384
rect 346922 415374 347032 415378
rect 336579 396456 336689 396460
rect 336567 396450 336701 396456
rect 324542 396394 324652 396398
rect 324530 396388 324664 396394
rect 322895 395804 324257 396346
rect 324530 396322 324542 396388
rect 324652 396322 324664 396388
rect 324530 396316 324664 396322
rect 324542 396312 324652 396316
rect 324552 396022 324662 396026
rect 324540 396016 324674 396022
rect 324540 395950 324552 396016
rect 324662 395950 324674 396016
rect 324540 395944 324674 395950
rect 324552 395940 324662 395944
rect 322895 391347 323437 395804
rect 324813 395802 326307 396344
rect 322889 390805 322895 391347
rect 323437 390805 323443 391347
rect 325765 376095 326307 395802
rect 334879 395900 336291 396442
rect 336567 396384 336579 396450
rect 336689 396384 336701 396450
rect 336567 396378 336701 396384
rect 336579 396374 336689 396378
rect 336589 396084 336699 396088
rect 336577 396078 336711 396084
rect 336577 396012 336589 396078
rect 336699 396012 336711 396078
rect 336577 396006 336711 396012
rect 336589 396002 336699 396006
rect 336863 395900 337875 396442
rect 333086 390825 333092 391367
rect 333634 390825 333640 391367
rect 334879 391309 335421 395900
rect 333092 381059 333634 390825
rect 334873 390767 334879 391309
rect 335421 390767 335427 391309
rect 333071 380757 333149 380769
rect 333067 380647 333077 380757
rect 333143 380647 333153 380757
rect 333443 380747 333521 380759
rect 333071 380635 333149 380647
rect 333439 380637 333449 380747
rect 333515 380637 333525 380747
rect 333443 380625 333521 380637
rect 333090 376209 333632 380469
rect 325759 375553 325765 376095
rect 326307 375553 326313 376095
rect 333090 375661 333632 375667
rect 337333 376115 337875 395900
rect 345480 395265 346022 414894
rect 348243 395267 348785 415403
rect 353573 415775 354168 415781
rect 355065 415775 355607 421893
rect 356003 421853 356015 421919
rect 356125 421853 356137 421919
rect 356403 421867 358082 422409
rect 356003 421847 356137 421853
rect 356015 421843 356125 421847
rect 373950 420915 374492 429649
rect 375352 426531 375894 429653
rect 385933 427718 386475 429745
rect 387904 427732 388014 427736
rect 387892 427726 388026 427732
rect 385933 427176 387605 427718
rect 387892 427660 387904 427726
rect 388014 427660 388026 427726
rect 388617 427706 389159 448215
rect 391205 448275 392489 448817
rect 392784 448771 392796 448837
rect 392906 448771 392918 448837
rect 392784 448765 392918 448771
rect 392796 448761 392906 448765
rect 392806 448471 392916 448475
rect 392794 448465 392928 448471
rect 392794 448399 392806 448465
rect 392916 448399 392928 448465
rect 392794 448393 392928 448399
rect 392806 448389 392916 448393
rect 391205 430371 391747 448275
rect 393089 448262 394207 448804
rect 391199 429829 391205 430371
rect 391747 429829 391753 430371
rect 387892 427654 388026 427660
rect 387904 427650 388014 427654
rect 387914 427360 388024 427364
rect 387902 427354 388036 427360
rect 387902 427288 387914 427354
rect 388024 427288 388036 427354
rect 387902 427282 388036 427288
rect 387914 427278 388024 427282
rect 388129 427164 389159 427706
rect 391205 427714 391747 429829
rect 392828 427751 392938 427755
rect 392816 427745 392950 427751
rect 391205 427172 392540 427714
rect 392816 427679 392828 427745
rect 392938 427679 392950 427745
rect 393665 427718 394207 448262
rect 497210 430398 497838 454616
rect 503867 449198 504469 454634
rect 510283 449200 510885 468398
rect 515023 467837 515133 467841
rect 503867 448596 508774 449198
rect 508964 449044 509074 449048
rect 508952 449038 509086 449044
rect 508952 448972 508964 449038
rect 509074 448972 509086 449038
rect 508952 448966 509086 448972
rect 508964 448962 509074 448966
rect 508974 448672 509084 448676
rect 508962 448666 509096 448672
rect 508962 448600 508974 448666
rect 509084 448600 509096 448666
rect 508962 448594 509096 448600
rect 509384 448598 510885 449200
rect 508974 448590 509084 448594
rect 497210 429764 497838 429770
rect 510283 430285 510885 448598
rect 513067 467230 514710 467832
rect 515011 467831 515145 467837
rect 515011 467765 515023 467831
rect 515133 467765 515145 467831
rect 518235 467830 518837 472485
rect 515011 467759 515145 467765
rect 515023 467755 515133 467759
rect 515033 467465 515143 467469
rect 515021 467459 515155 467465
rect 515021 467393 515033 467459
rect 515143 467393 515155 467459
rect 515021 467387 515155 467393
rect 515033 467383 515143 467387
rect 513067 447647 513669 467230
rect 515313 467228 518837 467830
rect 518235 457319 518837 467228
rect 523715 459620 524345 472495
rect 531891 467186 532521 484571
rect 536943 473163 537545 487959
rect 545784 492230 549875 492231
rect 545784 491601 550146 492230
rect 550466 492062 550576 492066
rect 550454 492056 550588 492062
rect 550454 491990 550466 492056
rect 550576 491990 550588 492056
rect 550454 491984 550588 491990
rect 550466 491980 550576 491984
rect 550456 491690 550566 491694
rect 550444 491684 550578 491690
rect 550444 491618 550456 491684
rect 550566 491618 550578 491684
rect 550444 491612 550578 491618
rect 550456 491608 550566 491612
rect 550736 491602 553793 492232
rect 545784 485127 546414 491601
rect 549516 491600 550146 491601
rect 545778 484497 545784 485127
rect 546414 484497 546420 485127
rect 542602 482075 543232 482083
rect 545784 482075 546414 484497
rect 542602 481445 546414 482075
rect 542602 477185 543232 481445
rect 545784 479912 546414 481445
rect 545796 479620 545874 479632
rect 545792 479510 545802 479620
rect 545868 479510 545878 479620
rect 546168 479610 546246 479622
rect 545796 479498 545874 479510
rect 546164 479500 546174 479610
rect 546240 479500 546250 479610
rect 546168 479488 546246 479500
rect 545774 478829 546404 479312
rect 545774 478199 548783 478829
rect 542602 476555 546463 477185
rect 545833 475831 546463 476555
rect 545849 475528 545927 475540
rect 545845 475418 545855 475528
rect 545921 475418 545931 475528
rect 546221 475518 546299 475530
rect 545849 475406 545927 475418
rect 546217 475408 546227 475518
rect 546293 475408 546303 475518
rect 546221 475396 546299 475408
rect 545838 474731 546468 475228
rect 548153 474731 548783 478199
rect 545838 474101 548783 474731
rect 548153 473207 548783 474101
rect 536937 472561 536943 473163
rect 537545 472561 537551 473163
rect 537951 472511 537957 473141
rect 538587 472511 538593 473141
rect 548147 472577 548153 473207
rect 548783 472577 548789 473207
rect 553163 473131 553793 491602
rect 531891 466556 534080 467186
rect 537957 467184 538587 472511
rect 553157 472501 553163 473131
rect 553793 472501 553799 473131
rect 562803 473059 563433 473065
rect 564214 473059 564844 497566
rect 567849 485171 568479 499797
rect 567843 484541 567849 485171
rect 568479 484541 568485 485171
rect 534386 467017 534496 467021
rect 534374 467011 534508 467017
rect 534374 466945 534386 467011
rect 534496 466945 534508 467011
rect 534374 466939 534508 466945
rect 534386 466935 534496 466939
rect 534376 466645 534486 466649
rect 534364 466639 534498 466645
rect 534364 466573 534376 466639
rect 534486 466573 534498 466639
rect 534364 466567 534498 466573
rect 534376 466563 534486 466567
rect 534672 466554 538587 467184
rect 523715 458990 527356 459620
rect 527531 459608 527641 459612
rect 527519 459602 527653 459608
rect 527519 459536 527531 459602
rect 527641 459536 527653 459602
rect 527519 459530 527653 459536
rect 527531 459526 527641 459530
rect 527521 459236 527631 459240
rect 527509 459230 527643 459236
rect 527509 459164 527521 459230
rect 527631 459164 527643 459230
rect 527509 459158 527643 459164
rect 527521 459154 527631 459158
rect 527900 458994 529589 459624
rect 518235 456717 521291 457319
rect 521414 457170 521524 457174
rect 521402 457164 521536 457170
rect 521402 457098 521414 457164
rect 521524 457098 521536 457164
rect 521402 457092 521536 457098
rect 521414 457088 521524 457092
rect 521424 456798 521534 456802
rect 521412 456792 521546 456798
rect 521412 456726 521424 456792
rect 521534 456726 521546 456792
rect 521412 456720 521546 456726
rect 521830 456722 522913 457324
rect 513067 447045 514771 447647
rect 518235 447640 518837 456717
rect 521424 456716 521534 456720
rect 515060 447636 515170 447640
rect 515048 447630 515182 447636
rect 515048 447564 515060 447630
rect 515170 447564 515182 447630
rect 515048 447558 515182 447564
rect 515060 447554 515170 447558
rect 515070 447264 515180 447268
rect 515058 447258 515192 447264
rect 515058 447192 515070 447258
rect 515180 447192 515192 447258
rect 515058 447186 515192 447192
rect 515070 447182 515180 447186
rect 513067 430335 513669 447045
rect 515336 447038 518837 447640
rect 522311 430301 522913 456722
rect 528959 446776 529589 458994
rect 537957 446795 538587 466554
rect 553163 459752 553793 472501
rect 563433 472429 564844 473059
rect 562803 472423 563433 472429
rect 528959 446146 534082 446776
rect 534376 446617 534486 446621
rect 534364 446611 534498 446617
rect 534364 446545 534376 446611
rect 534486 446545 534498 446611
rect 534364 446539 534498 446545
rect 534376 446535 534486 446539
rect 534366 446245 534476 446249
rect 534354 446239 534488 446245
rect 534354 446173 534366 446239
rect 534476 446173 534488 446239
rect 534354 446167 534488 446173
rect 534366 446163 534476 446167
rect 534663 446165 538587 446795
rect 545783 459122 550190 459752
rect 550370 459737 550480 459741
rect 550358 459731 550492 459737
rect 550358 459665 550370 459731
rect 550480 459665 550492 459731
rect 550358 459659 550492 459665
rect 550370 459655 550480 459659
rect 550360 459365 550470 459369
rect 550348 459359 550482 459365
rect 550348 459293 550360 459359
rect 550470 459293 550482 459359
rect 550348 459287 550482 459293
rect 550360 459283 550470 459287
rect 550778 459122 553793 459752
rect 564146 471173 564844 472429
rect 528959 430329 529589 446146
rect 545783 430403 546413 459122
rect 564146 453575 564776 471173
rect 564158 453395 564236 453407
rect 564530 453405 564608 453417
rect 564154 453285 564164 453395
rect 564230 453285 564240 453395
rect 564526 453295 564536 453405
rect 564602 453295 564612 453405
rect 564158 453273 564236 453285
rect 564530 453283 564608 453295
rect 513067 429727 513669 429733
rect 522305 429699 522311 430301
rect 522913 429699 522919 430301
rect 528953 429699 528959 430329
rect 529589 429699 529595 430329
rect 545777 429773 545783 430403
rect 546413 429773 546419 430403
rect 562801 430329 563431 430335
rect 564148 430329 564778 452976
rect 563431 429699 564778 430329
rect 510283 429677 510885 429683
rect 528959 429675 529589 429699
rect 562801 429693 563431 429699
rect 392816 427673 392950 427679
rect 392828 427669 392938 427673
rect 392838 427379 392948 427383
rect 392826 427373 392960 427379
rect 392826 427307 392838 427373
rect 392948 427307 392960 427373
rect 392826 427301 392960 427307
rect 392838 427297 392948 427301
rect 393124 427176 394207 427718
rect 375488 426241 375566 426253
rect 375860 426251 375938 426263
rect 375484 426131 375494 426241
rect 375560 426131 375570 426241
rect 375856 426141 375866 426251
rect 375932 426141 375942 426251
rect 375488 426119 375566 426131
rect 375860 426129 375938 426141
rect 374098 420649 374176 420661
rect 374470 420659 374548 420671
rect 374094 420539 374104 420649
rect 374170 420539 374180 420649
rect 374466 420549 374476 420659
rect 374542 420549 374552 420659
rect 374098 420527 374176 420539
rect 374470 420537 374548 420549
rect 373944 415845 374486 420379
rect 354115 415233 355607 415775
rect 373938 415303 373944 415845
rect 374486 415303 374492 415845
rect 375340 415649 375882 425961
rect 388617 415849 389159 427164
rect 393665 415927 394207 427176
rect 353573 415227 354419 415233
rect 353877 402378 354419 415227
rect 375334 415107 375340 415649
rect 375882 415107 375888 415649
rect 388611 415307 388617 415849
rect 389159 415307 389165 415849
rect 393665 415379 394207 415385
rect 568059 410195 571789 410757
rect 568059 409942 568621 410195
rect 568052 409380 568621 409942
rect 568059 409253 568621 409380
rect 568040 408988 568118 409000
rect 568036 408878 568046 408988
rect 568112 408878 568122 408988
rect 568412 408978 568490 408990
rect 568040 408866 568118 408878
rect 568408 408868 568418 408978
rect 568484 408868 568494 408978
rect 568412 408856 568490 408868
rect 546403 407353 546965 407431
rect 546403 406791 549239 407353
rect 552361 407335 552923 407359
rect 549553 407202 549663 407206
rect 549541 407196 549675 407202
rect 549541 407130 549553 407196
rect 549663 407130 549675 407196
rect 549541 407124 549675 407130
rect 549553 407120 549663 407124
rect 549543 406830 549653 406834
rect 549531 406824 549665 406830
rect 356805 402394 358232 402405
rect 353877 401836 355803 402378
rect 355994 402262 356104 402266
rect 355982 402256 356116 402262
rect 355982 402190 355994 402256
rect 356104 402190 356116 402256
rect 355982 402184 356116 402190
rect 355994 402180 356104 402184
rect 356004 401890 356114 401894
rect 355992 401884 356126 401890
rect 355992 401818 356004 401884
rect 356114 401818 356126 401884
rect 356422 401863 358232 402394
rect 356422 401852 356964 401863
rect 355992 401812 356126 401818
rect 356004 401808 356114 401812
rect 345477 394723 346765 395265
rect 346940 395150 347050 395154
rect 346928 395144 347062 395150
rect 346928 395078 346940 395144
rect 347050 395078 347062 395144
rect 346928 395072 347062 395078
rect 346940 395068 347050 395072
rect 346950 394778 347060 394782
rect 346938 394772 347072 394778
rect 346938 394706 346950 394772
rect 347060 394706 347072 394772
rect 347337 394725 348785 395267
rect 346938 394700 347072 394706
rect 346950 394696 347060 394700
rect 357690 391157 358232 401863
rect 428501 391297 429043 391303
rect 353565 390939 354107 390945
rect 347476 390397 353565 390939
rect 357684 390615 357690 391157
rect 358232 390615 358238 391157
rect 367478 390651 367484 391193
rect 368026 390651 368032 391193
rect 347476 387029 348018 390397
rect 353565 390391 354107 390397
rect 347440 386724 347518 386736
rect 347436 386614 347446 386724
rect 347512 386614 347522 386724
rect 347812 386714 347890 386726
rect 347440 386602 347518 386614
rect 347808 386604 347818 386714
rect 347884 386604 347894 386714
rect 347812 386592 347890 386604
rect 347468 382360 348010 386427
rect 347468 381818 355792 382360
rect 357690 382359 358232 390615
rect 367484 387063 368026 390651
rect 385263 390627 385269 391169
rect 385811 390627 385817 391169
rect 400431 390647 400437 391189
rect 400979 390647 400985 391189
rect 425687 390755 428501 391297
rect 546403 391241 546965 406791
rect 549531 406758 549543 406824
rect 549653 406758 549665 406824
rect 549821 406773 552923 407335
rect 549531 406752 549665 406758
rect 549543 406748 549653 406752
rect 385269 388729 385811 390627
rect 385269 388187 387838 388729
rect 367456 386753 367534 386765
rect 367452 386643 367462 386753
rect 367528 386643 367538 386753
rect 367828 386743 367906 386755
rect 367456 386631 367534 386643
rect 367824 386633 367834 386743
rect 367900 386633 367910 386743
rect 367828 386621 367906 386633
rect 355974 382198 356084 382202
rect 355962 382192 356096 382198
rect 355962 382126 355974 382192
rect 356084 382126 356096 382192
rect 355962 382120 356096 382126
rect 355974 382116 356084 382120
rect 355984 381826 356094 381830
rect 355972 381820 356106 381826
rect 347468 376199 348010 381818
rect 355972 381754 355984 381820
rect 356094 381754 356106 381820
rect 356347 381817 358232 382359
rect 355972 381748 356106 381754
rect 355984 381744 356094 381748
rect 357690 381073 358232 381817
rect 357650 380765 357728 380777
rect 357646 380655 357656 380765
rect 357722 380655 357732 380765
rect 358022 380755 358100 380767
rect 357650 380643 357728 380655
rect 358018 380645 358028 380755
rect 358094 380645 358104 380755
rect 358022 380633 358100 380645
rect 352320 376199 352330 376280
rect 337333 375567 337875 375573
rect 345681 376089 346223 376095
rect 347468 375657 352330 376199
rect 352307 375655 352330 375657
rect 352320 375608 352330 375655
rect 353838 376197 353848 376280
rect 353838 375655 354583 376197
rect 357684 376101 358226 380451
rect 353838 375608 353848 375655
rect 345681 373983 346223 375547
rect 345681 373441 346751 373983
rect 346926 373868 347036 373872
rect 346914 373862 347048 373868
rect 346914 373796 346926 373862
rect 347036 373796 347048 373862
rect 346914 373790 347048 373796
rect 346926 373786 347036 373790
rect 346936 373496 347046 373500
rect 346924 373490 347058 373496
rect 345681 353133 346223 373441
rect 346924 373424 346936 373490
rect 347046 373424 347058 373490
rect 347323 373443 348671 373985
rect 346924 373418 347058 373424
rect 346936 373414 347046 373418
rect 348129 353135 348671 373443
rect 345681 352591 346751 353133
rect 346926 353018 347036 353022
rect 346914 353012 347048 353018
rect 346914 352946 346926 353012
rect 347036 352946 347048 353012
rect 346914 352940 347048 352946
rect 346926 352936 347036 352940
rect 346936 352646 347046 352650
rect 346924 352640 347058 352646
rect 345681 332537 346223 352591
rect 346924 352574 346936 352640
rect 347046 352574 347058 352640
rect 347323 352593 348671 353135
rect 346924 352568 347058 352574
rect 346936 352564 347046 352568
rect 348129 332539 348671 352593
rect 345681 331995 346835 332537
rect 347010 332422 347120 332426
rect 346998 332416 347132 332422
rect 346998 332350 347010 332416
rect 347120 332350 347132 332416
rect 346998 332344 347132 332350
rect 347010 332340 347120 332344
rect 347020 332050 347130 332054
rect 347008 332044 347142 332050
rect 345681 310669 346223 331995
rect 347008 331978 347020 332044
rect 347130 331978 347142 332044
rect 347407 331997 348671 332539
rect 347008 331972 347142 331978
rect 347020 331968 347130 331972
rect 348129 310671 348671 331997
rect 345681 310127 346807 310669
rect 346982 310554 347092 310558
rect 346970 310548 347104 310554
rect 346970 310482 346982 310548
rect 347092 310482 347104 310548
rect 346970 310476 347104 310482
rect 346982 310472 347092 310476
rect 346992 310182 347102 310186
rect 346980 310176 347114 310182
rect 345681 289011 346223 310127
rect 346980 310110 346992 310176
rect 347102 310110 347114 310176
rect 347379 310129 348671 310671
rect 346980 310104 347114 310110
rect 346992 310100 347102 310104
rect 348129 307618 348671 310129
rect 348014 305644 348024 307618
rect 348476 305644 348671 307618
rect 348129 289013 348671 305644
rect 345681 288469 346765 289011
rect 346940 288896 347050 288900
rect 346928 288890 347062 288896
rect 346928 288824 346940 288890
rect 347050 288824 347062 288890
rect 346928 288818 347062 288824
rect 346940 288814 347050 288818
rect 346950 288524 347060 288528
rect 346938 288518 347072 288524
rect 345681 287588 346223 288469
rect 346938 288452 346950 288518
rect 347060 288452 347072 288518
rect 347337 288471 348671 289013
rect 346938 288446 347072 288452
rect 346950 288442 347060 288446
rect 345681 285614 345710 287588
rect 346162 285614 346223 287588
rect 345681 264231 346223 285614
rect 348129 264233 348671 288471
rect 354041 362352 354583 375655
rect 357678 375559 357684 376101
rect 358226 375559 358232 376101
rect 367484 376051 368026 386463
rect 385269 382711 385811 388187
rect 387296 387041 387838 388187
rect 400437 388487 400979 390647
rect 425687 388569 426229 390755
rect 428501 390749 429043 390755
rect 446389 390507 446395 391049
rect 446937 390507 446943 391049
rect 470021 390513 470027 391055
rect 470569 390513 470575 391055
rect 490263 390563 490269 391105
rect 490811 390563 490817 391105
rect 400437 387945 408104 388487
rect 387268 386743 387346 386755
rect 387264 386633 387274 386743
rect 387340 386633 387350 386743
rect 387640 386733 387718 386745
rect 387268 386621 387346 386633
rect 387636 386623 387646 386733
rect 387712 386623 387722 386733
rect 387640 386611 387718 386623
rect 387295 386054 387837 386451
rect 387295 385691 387838 386054
rect 387295 385149 389101 385691
rect 385269 382169 387659 382711
rect 387117 381778 387659 382169
rect 387112 381236 387659 381778
rect 387117 381015 387659 381236
rect 387097 380723 387175 380735
rect 387093 380613 387103 380723
rect 387169 380613 387179 380723
rect 387469 380713 387547 380725
rect 387097 380601 387175 380613
rect 387465 380603 387475 380713
rect 387541 380603 387551 380713
rect 387469 380591 387547 380603
rect 387112 379667 387654 380429
rect 388559 379667 389101 385149
rect 406151 382205 406693 387945
rect 407562 387049 408104 387945
rect 425687 388027 428360 388569
rect 407527 386741 407605 386753
rect 407523 386631 407533 386741
rect 407599 386631 407609 386741
rect 407899 386731 407977 386743
rect 407527 386619 407605 386631
rect 407895 386621 407905 386731
rect 407971 386621 407981 386731
rect 407899 386609 407977 386621
rect 407564 385635 408106 386457
rect 407564 385093 409803 385635
rect 406151 381746 408237 382205
rect 406151 381663 408250 381746
rect 407695 381204 408250 381663
rect 407695 381061 408237 381204
rect 407675 380754 407753 380766
rect 407671 380644 407681 380754
rect 407747 380644 407757 380754
rect 408047 380744 408125 380756
rect 407675 380632 407753 380644
rect 408043 380634 408053 380744
rect 408119 380634 408129 380744
rect 408047 380622 408125 380634
rect 387112 379125 389101 379667
rect 407710 379613 408252 380473
rect 409261 379613 409803 385093
rect 425687 382259 426229 388027
rect 427818 387071 428360 388027
rect 446395 388537 446937 390507
rect 446395 387995 448520 388537
rect 470027 388131 470569 390513
rect 490269 388471 490811 390563
rect 510717 390533 510723 391075
rect 511265 390533 511271 391075
rect 530379 390605 530385 391147
rect 530927 390605 530933 391147
rect 546397 390679 546403 391241
rect 546965 390679 546971 391241
rect 510723 388541 511265 390533
rect 427803 386796 427881 386808
rect 427799 386686 427809 386796
rect 427875 386686 427885 386796
rect 428175 386786 428253 386798
rect 427803 386674 427881 386686
rect 428171 386676 428181 386786
rect 428247 386676 428257 386786
rect 428175 386664 428253 386676
rect 427825 386250 428367 386489
rect 427824 385999 428367 386250
rect 427824 385708 429691 385999
rect 427825 385457 429691 385708
rect 425687 382258 427630 382259
rect 425687 381717 428218 382258
rect 427676 381039 428218 381717
rect 427649 380729 427727 380741
rect 427645 380619 427655 380729
rect 427721 380619 427731 380729
rect 428021 380719 428099 380731
rect 427649 380607 427727 380619
rect 428017 380609 428027 380719
rect 428093 380609 428103 380719
rect 428021 380597 428099 380609
rect 427676 379680 428218 380421
rect 429149 379680 429691 385457
rect 446395 382191 446937 387995
rect 447978 387043 448520 387995
rect 467998 387589 470569 388131
rect 467998 387079 468540 387589
rect 447962 386776 448040 386788
rect 447958 386666 447968 386776
rect 448034 386666 448044 386776
rect 448334 386766 448412 386778
rect 467964 386771 468042 386783
rect 447962 386654 448040 386666
rect 448330 386656 448340 386766
rect 448406 386656 448416 386766
rect 467960 386661 467970 386771
rect 468036 386661 468046 386771
rect 468336 386761 468414 386773
rect 448334 386644 448412 386656
rect 467964 386649 468042 386661
rect 468332 386651 468342 386761
rect 468408 386651 468418 386761
rect 468336 386639 468414 386651
rect 447978 385789 448520 386501
rect 468001 386184 468543 386489
rect 467996 386123 468543 386184
rect 447978 385247 450417 385789
rect 446395 381649 448473 382191
rect 447930 381220 448473 381649
rect 447931 381033 448473 381220
rect 447895 380733 447973 380745
rect 447891 380623 447901 380733
rect 447967 380623 447977 380733
rect 448267 380723 448345 380735
rect 447895 380611 447973 380623
rect 448263 380613 448273 380723
rect 448339 380613 448349 380723
rect 448267 380601 448345 380613
rect 447932 379823 448474 380435
rect 449875 379823 450417 385247
rect 367478 375509 367484 376051
rect 368026 375509 368032 376051
rect 388559 375919 389101 379125
rect 400425 379071 409805 379613
rect 427676 379138 429691 379680
rect 400425 376101 400967 379071
rect 388553 375377 388559 375919
rect 389101 375377 389107 375919
rect 400419 375559 400425 376101
rect 400967 375559 400973 376101
rect 429149 376007 429691 379138
rect 446411 379281 450417 379823
rect 466549 385581 468543 386123
rect 466549 380069 467091 385581
rect 470027 382451 470569 387589
rect 488130 387929 490811 388471
rect 488130 387037 488672 387929
rect 488082 386755 488160 386767
rect 488078 386645 488088 386755
rect 488154 386645 488164 386755
rect 488454 386745 488532 386757
rect 488082 386633 488160 386645
rect 488450 386635 488460 386745
rect 488526 386635 488536 386745
rect 488454 386623 488532 386635
rect 488117 386276 488659 386465
rect 488116 385827 488659 386276
rect 467909 381909 470569 382451
rect 485509 385285 488659 385827
rect 467909 381746 468451 381909
rect 467902 381204 468451 381746
rect 467909 381085 468451 381204
rect 467879 380800 467957 380812
rect 467875 380690 467885 380800
rect 467951 380690 467961 380800
rect 468251 380790 468329 380802
rect 467879 380678 467957 380690
rect 468247 380680 468257 380790
rect 468323 380680 468333 380790
rect 468251 380668 468329 380680
rect 467900 380069 468442 380531
rect 466549 379527 468442 380069
rect 485509 380052 486051 385285
rect 490269 382483 490811 387929
rect 508262 387999 511265 388541
rect 530385 388103 530927 390605
rect 508262 387086 508804 387999
rect 508212 386778 508290 386790
rect 508208 386668 508218 386778
rect 508284 386668 508294 386778
rect 508584 386768 508662 386780
rect 508212 386656 508290 386668
rect 508580 386658 508590 386768
rect 508656 386658 508666 386768
rect 508584 386646 508662 386658
rect 508238 386017 508780 386486
rect 488330 381941 490811 382483
rect 505733 385475 508780 386017
rect 488330 381043 488872 381941
rect 488294 380725 488372 380737
rect 488290 380615 488300 380725
rect 488366 380615 488376 380725
rect 488666 380715 488744 380727
rect 488294 380603 488372 380615
rect 488662 380605 488672 380715
rect 488738 380605 488748 380715
rect 488666 380593 488744 380605
rect 488322 380052 488864 380427
rect 446411 376065 446953 379281
rect 429143 375465 429149 376007
rect 429691 375465 429697 376007
rect 446405 375523 446411 376065
rect 446953 375523 446959 376065
rect 466549 376049 467091 379527
rect 485509 379510 488864 380052
rect 505733 380053 506275 385475
rect 510723 382593 511265 387999
rect 528360 387561 530927 388103
rect 528360 387092 528902 387561
rect 528321 386792 528399 386804
rect 528317 386682 528327 386792
rect 528393 386682 528403 386792
rect 528693 386782 528771 386794
rect 528321 386670 528399 386682
rect 528689 386672 528699 386782
rect 528765 386672 528775 386782
rect 528693 386660 528771 386672
rect 528336 385693 528878 386514
rect 527028 385692 528878 385693
rect 526297 385151 528878 385692
rect 508018 382051 511265 382593
rect 508018 381098 508560 382051
rect 507977 380797 508055 380809
rect 507973 380687 507983 380797
rect 508049 380687 508059 380797
rect 508349 380787 508427 380799
rect 507977 380675 508055 380687
rect 508345 380677 508355 380787
rect 508421 380677 508431 380787
rect 508349 380665 508427 380677
rect 507994 380053 508536 380520
rect 505733 379511 508536 380053
rect 526305 379745 526847 385151
rect 530385 382097 530927 387561
rect 528388 381555 530927 382097
rect 546403 388288 546965 390679
rect 552361 388300 552923 406773
rect 568048 406629 568610 408690
rect 546403 387726 549272 388288
rect 549570 388158 549680 388162
rect 549558 388152 549692 388158
rect 549558 388086 549570 388152
rect 549680 388086 549692 388152
rect 549558 388080 549692 388086
rect 549570 388076 549680 388080
rect 549560 387786 549670 387790
rect 549548 387780 549682 387786
rect 528388 381026 528930 381555
rect 528347 380731 528425 380743
rect 528343 380621 528353 380731
rect 528419 380621 528429 380731
rect 528719 380721 528797 380733
rect 528347 380609 528425 380621
rect 528715 380611 528725 380721
rect 528791 380611 528801 380721
rect 528719 380599 528797 380611
rect 528364 379745 528906 380448
rect 466543 375507 466549 376049
rect 467091 375507 467097 376049
rect 485509 376005 486051 379510
rect 485503 375463 485509 376005
rect 486051 375463 486057 376005
rect 505733 375989 506275 379511
rect 526305 379203 528906 379745
rect 546403 379464 546965 387726
rect 549548 387714 549560 387780
rect 549670 387714 549682 387780
rect 549850 387738 552923 388300
rect 549548 387708 549682 387714
rect 549560 387704 549670 387708
rect 549368 379500 549478 379504
rect 549356 379494 549490 379500
rect 526305 376169 526847 379203
rect 546403 378904 549080 379464
rect 549356 379428 549368 379494
rect 549478 379428 549490 379494
rect 552361 379480 552923 387738
rect 549356 379422 549490 379428
rect 549368 379418 549478 379422
rect 549378 379128 549488 379132
rect 549366 379122 549500 379128
rect 549366 379056 549378 379122
rect 549488 379056 549500 379122
rect 549366 379050 549500 379056
rect 549378 379046 549488 379050
rect 549664 378918 552923 379480
rect 505727 375447 505733 375989
rect 506275 375447 506281 375989
rect 526299 375627 526305 376169
rect 526847 375627 526853 376169
rect 546403 364265 546965 378904
rect 548520 378902 549062 378904
rect 552361 376047 552923 378918
rect 564047 406067 568610 406629
rect 562709 376121 563271 376127
rect 564047 376121 564609 406067
rect 571227 391205 571789 410195
rect 571221 390643 571227 391205
rect 571789 390643 571795 391205
rect 552355 375485 552361 376047
rect 552923 375485 552929 376047
rect 563271 375559 564609 376121
rect 562709 375553 563271 375559
rect 549329 364314 549439 364318
rect 549317 364308 549451 364314
rect 546403 363703 549029 364265
rect 549317 364242 549329 364308
rect 549439 364242 549451 364308
rect 552361 364305 552923 375485
rect 549317 364236 549451 364242
rect 549329 364232 549439 364236
rect 549339 363942 549449 363946
rect 549327 363936 549461 363942
rect 549327 363870 549339 363936
rect 549449 363870 549461 363936
rect 549327 363864 549461 363870
rect 549339 363860 549449 363864
rect 549637 363743 552923 364305
rect 354041 361810 355861 362352
rect 356446 362319 358483 362350
rect 356031 362215 356141 362219
rect 356019 362209 356153 362215
rect 356019 362143 356031 362209
rect 356141 362143 356153 362209
rect 356019 362137 356153 362143
rect 356031 362133 356141 362137
rect 356041 361843 356151 361847
rect 356029 361837 356163 361843
rect 354041 342326 354583 361810
rect 356029 361771 356041 361837
rect 356151 361771 356163 361837
rect 356446 361808 358487 362319
rect 356029 361765 356163 361771
rect 356041 361761 356151 361765
rect 354041 341784 355861 342326
rect 357945 342324 358487 361808
rect 564047 360213 564609 375559
rect 571227 365957 571789 390643
rect 568218 365395 571789 365957
rect 568218 362912 568780 365395
rect 568196 362605 568274 362617
rect 568192 362495 568202 362605
rect 568268 362495 568278 362605
rect 568568 362595 568646 362607
rect 568196 362483 568274 362495
rect 568564 362485 568574 362595
rect 568640 362485 568650 362595
rect 568568 362473 568646 362485
rect 568226 362069 568788 362302
rect 568226 361740 568793 362069
rect 568231 360213 568793 361740
rect 564047 359651 568793 360213
rect 356031 342212 356141 342216
rect 356019 342206 356153 342212
rect 356019 342140 356031 342206
rect 356141 342140 356153 342206
rect 356019 342134 356153 342140
rect 356031 342130 356141 342134
rect 356041 341840 356151 341844
rect 356029 341834 356163 341840
rect 354041 322328 354583 341784
rect 356029 341768 356041 341834
rect 356151 341768 356163 341834
rect 356438 341782 358487 342324
rect 356029 341762 356163 341768
rect 356041 341758 356151 341762
rect 354041 321786 355773 322328
rect 357945 322326 358487 341782
rect 355955 322210 356065 322214
rect 355943 322204 356077 322210
rect 355943 322138 355955 322204
rect 356065 322138 356077 322204
rect 355943 322132 356077 322138
rect 355955 322128 356065 322132
rect 355965 321838 356075 321842
rect 355953 321832 356087 321838
rect 354041 302314 354583 321786
rect 355953 321766 355965 321832
rect 356075 321766 356087 321832
rect 356372 321784 358487 322326
rect 355953 321760 356087 321766
rect 355965 321756 356075 321760
rect 357945 306779 358487 321784
rect 390700 306940 391249 306946
rect 354041 301772 355807 302314
rect 357945 302312 358487 306237
rect 355993 302189 356103 302193
rect 355981 302183 356115 302189
rect 355981 302117 355993 302183
rect 356103 302117 356115 302183
rect 355981 302111 356115 302117
rect 355993 302107 356103 302111
rect 356003 301817 356113 301821
rect 355991 301811 356125 301817
rect 354041 286813 354583 301772
rect 355991 301745 356003 301811
rect 356113 301745 356125 301811
rect 356406 301770 358487 302312
rect 370688 306812 371237 306818
rect 355991 301739 356125 301745
rect 356003 301735 356113 301739
rect 370688 296332 371237 306263
rect 390700 296362 391249 306391
rect 400264 306898 400813 306904
rect 400813 306349 411265 306898
rect 445440 306860 445989 306866
rect 400264 306343 400813 306349
rect 410716 296330 411265 306349
rect 430714 306662 431263 306668
rect 445989 306311 451273 306860
rect 445440 306305 445989 306311
rect 430714 296408 431263 306113
rect 450724 296374 451273 306311
rect 470712 306231 470718 306780
rect 471267 306231 471273 306780
rect 490708 306455 490714 307004
rect 491263 306455 491269 307004
rect 470718 296392 471267 306231
rect 490714 296426 491263 306455
rect 510694 306347 510700 306896
rect 511249 306347 511255 306896
rect 569358 306806 569927 306812
rect 510700 296377 511249 306347
rect 530680 306193 530686 306742
rect 531235 306193 531241 306742
rect 530686 296421 531235 306193
rect 552161 306173 552167 306730
rect 552724 306173 552730 306730
rect 569927 306237 572331 306806
rect 569358 306231 569927 306237
rect 490847 296123 490925 296135
rect 491219 296133 491297 296145
rect 430833 296098 430911 296110
rect 431205 296108 431283 296120
rect 370822 296034 370900 296046
rect 371194 296044 371272 296056
rect 390831 296051 390909 296063
rect 391203 296061 391281 296073
rect 370818 295924 370828 296034
rect 370894 295924 370904 296034
rect 371190 295934 371200 296044
rect 371266 295934 371276 296044
rect 390827 295941 390837 296051
rect 390903 295941 390913 296051
rect 391199 295951 391209 296061
rect 391275 295951 391285 296061
rect 410837 296022 410915 296034
rect 411209 296032 411287 296044
rect 370822 295912 370900 295924
rect 371194 295922 371272 295934
rect 390831 295929 390909 295941
rect 391203 295939 391281 295951
rect 410833 295912 410843 296022
rect 410909 295912 410919 296022
rect 411205 295922 411215 296032
rect 411281 295922 411291 296032
rect 430829 295988 430839 296098
rect 430905 295988 430915 296098
rect 431201 295998 431211 296108
rect 431277 295998 431287 296108
rect 470852 296090 470930 296102
rect 471224 296100 471302 296112
rect 450850 296065 450928 296077
rect 451222 296075 451300 296087
rect 430833 295976 430911 295988
rect 431205 295986 431283 295998
rect 450846 295955 450856 296065
rect 450922 295955 450932 296065
rect 451218 295965 451228 296075
rect 451294 295965 451304 296075
rect 470848 295980 470858 296090
rect 470924 295980 470934 296090
rect 471220 295990 471230 296100
rect 471296 295990 471306 296100
rect 490843 296013 490853 296123
rect 490919 296013 490929 296123
rect 491215 296023 491225 296133
rect 491291 296023 491301 296133
rect 530825 296123 530903 296135
rect 531197 296133 531275 296145
rect 510840 296079 510918 296091
rect 511212 296089 511290 296101
rect 490847 296001 490925 296013
rect 491219 296011 491297 296023
rect 470852 295968 470930 295980
rect 471224 295978 471302 295990
rect 510836 295969 510846 296079
rect 510912 295969 510922 296079
rect 511208 295979 511218 296089
rect 511284 295979 511294 296089
rect 530821 296013 530831 296123
rect 530897 296013 530907 296123
rect 531193 296023 531203 296133
rect 531269 296023 531279 296133
rect 530825 296001 530903 296013
rect 531197 296011 531275 296023
rect 450850 295943 450928 295955
rect 451222 295953 451300 295965
rect 510840 295957 510918 295969
rect 511212 295967 511290 295979
rect 410837 295900 410915 295912
rect 411209 295910 411287 295922
rect 354035 286271 354041 286813
rect 354583 286271 354589 286813
rect 370688 286607 371237 295745
rect 390700 286691 391249 295784
rect 370682 286058 370688 286607
rect 371237 286058 371243 286607
rect 400180 286903 400729 286909
rect 410716 286903 411265 295752
rect 400729 286354 411265 286903
rect 430714 286809 431263 295830
rect 450724 292777 451273 295796
rect 400180 286348 400729 286354
rect 445452 292228 451273 292777
rect 445452 287021 446001 292228
rect 470718 286753 471267 295814
rect 490714 286883 491263 295848
rect 445452 286466 446001 286472
rect 430714 286254 431263 286260
rect 470712 286204 470718 286753
rect 471267 286204 471273 286753
rect 490708 286334 490714 286883
rect 491263 286334 491269 286883
rect 510700 286819 511249 295808
rect 510694 286270 510700 286819
rect 511249 286270 511255 286819
rect 530686 286807 531235 295848
rect 552167 293595 552724 306173
rect 546320 293036 549377 293593
rect 549547 293447 549657 293451
rect 549535 293441 549669 293447
rect 549535 293375 549547 293441
rect 549657 293375 549669 293441
rect 549535 293369 549669 293375
rect 549547 293365 549657 293369
rect 549557 293075 549667 293079
rect 549545 293069 549679 293075
rect 546320 286983 546877 293036
rect 549545 293003 549557 293069
rect 549667 293003 549679 293069
rect 549958 293038 552724 293595
rect 549545 292997 549679 293003
rect 549557 292993 549667 292997
rect 530680 286258 530686 286807
rect 531235 286258 531241 286807
rect 546314 286426 546320 286983
rect 546877 286426 546883 286983
rect 390700 286136 391249 286142
rect 546320 272119 546877 286426
rect 552167 275741 552724 293038
rect 551280 275184 552724 275741
rect 568318 286882 568887 286888
rect 551298 274881 551865 275184
rect 551296 274324 551865 274881
rect 551298 274314 551865 274324
rect 551443 274016 551521 274028
rect 551815 274026 551893 274038
rect 551439 273906 551449 274016
rect 551515 273906 551525 274016
rect 551811 273916 551821 274026
rect 551887 273916 551897 274026
rect 551443 273894 551521 273906
rect 551815 273904 551893 273916
rect 551307 273729 551871 273736
rect 551302 273172 551871 273729
rect 551307 272119 551871 273172
rect 568318 272935 568887 286313
rect 571762 274274 572331 306237
rect 571906 273976 571984 273988
rect 572278 273986 572356 273998
rect 571902 273866 571912 273976
rect 571978 273866 571988 273976
rect 572274 273876 572284 273986
rect 572350 273876 572360 273986
rect 571906 273854 571984 273866
rect 572278 273864 572356 273876
rect 571762 272935 572331 273696
rect 568318 272366 572331 272935
rect 546320 271562 551871 272119
rect 551307 271528 551871 271562
rect 345681 263689 346723 264231
rect 346898 264116 347008 264120
rect 346886 264110 347020 264116
rect 346886 264044 346898 264110
rect 347008 264044 347020 264110
rect 346886 264038 347020 264044
rect 346898 264034 347008 264038
rect 346908 263744 347018 263748
rect 346896 263738 347030 263744
rect 345681 242857 346223 263689
rect 346896 263672 346908 263738
rect 347018 263672 347030 263738
rect 347295 263691 348671 264233
rect 346896 263666 347030 263672
rect 346908 263662 347018 263666
rect 348129 242859 348671 263691
rect 345681 242315 346807 242857
rect 346982 242742 347092 242746
rect 346970 242736 347104 242742
rect 346970 242670 346982 242736
rect 347092 242670 347104 242736
rect 346970 242664 347104 242670
rect 346982 242660 347092 242664
rect 346992 242370 347102 242374
rect 346980 242364 347114 242370
rect 345681 222981 346223 242315
rect 346980 242298 346992 242364
rect 347102 242298 347114 242364
rect 347379 242317 348671 242859
rect 346980 242292 347114 242298
rect 346992 242288 347102 242292
rect 348129 222983 348671 242317
rect 345681 222439 346835 222981
rect 347010 222866 347120 222870
rect 346998 222860 347132 222866
rect 346998 222794 347010 222860
rect 347120 222794 347132 222860
rect 346998 222788 347132 222794
rect 347010 222784 347120 222788
rect 347020 222494 347130 222498
rect 347008 222488 347142 222494
rect 345681 201153 346223 222439
rect 347008 222422 347020 222488
rect 347130 222422 347142 222488
rect 347407 222441 348671 222983
rect 347008 222416 347142 222422
rect 347020 222412 347130 222416
rect 348129 213096 348671 222441
rect 347972 208088 347982 213096
rect 348448 208088 348671 213096
rect 348129 201155 348671 208088
rect 345681 200611 346779 201153
rect 346954 201038 347064 201042
rect 346942 201032 347076 201038
rect 346942 200966 346954 201032
rect 347064 200966 347076 201032
rect 346942 200960 347076 200966
rect 346954 200956 347064 200960
rect 346964 200666 347074 200670
rect 346952 200660 347086 200666
rect 345681 180119 346223 200611
rect 346952 200594 346964 200660
rect 347074 200594 347086 200660
rect 347351 200613 348671 201155
rect 346952 200588 347086 200594
rect 346964 200584 347074 200588
rect 348129 180121 348671 200613
rect 345681 179577 346793 180119
rect 346968 180004 347078 180008
rect 346956 179998 347090 180004
rect 346956 179932 346968 179998
rect 347078 179932 347090 179998
rect 346956 179926 347090 179932
rect 346968 179922 347078 179926
rect 346978 179632 347088 179636
rect 346966 179626 347100 179632
rect 345681 177826 346223 179577
rect 346966 179560 346978 179626
rect 347088 179560 347100 179626
rect 347365 179579 348671 180121
rect 346966 179554 347100 179560
rect 346978 179550 347088 179554
rect 345681 172818 345722 177826
rect 346188 172818 346223 177826
rect 345681 167836 346223 172818
rect 345681 162828 345698 167836
rect 346164 162828 346223 167836
rect 345681 158731 346223 162828
rect 348129 158733 348671 179579
rect 345681 158189 346751 158731
rect 346926 158616 347036 158620
rect 346914 158610 347048 158616
rect 346914 158544 346926 158610
rect 347036 158544 347048 158610
rect 346914 158538 347048 158544
rect 346926 158534 347036 158538
rect 346936 158244 347046 158248
rect 346924 158238 347058 158244
rect 345681 137385 346223 158189
rect 346924 158172 346936 158238
rect 347046 158172 347058 158238
rect 347323 158191 348671 158733
rect 346924 158166 347058 158172
rect 346936 158162 347046 158166
rect 348129 137387 348671 158191
rect 334821 136843 334827 137385
rect 335369 136843 346695 137385
rect 347267 137369 348671 137387
rect 346870 137270 346980 137274
rect 346858 137264 346992 137270
rect 346858 137198 346870 137264
rect 346980 137198 346992 137264
rect 346858 137192 346992 137198
rect 346870 137188 346980 137192
rect 346880 136898 346990 136902
rect 346868 136892 347002 136898
rect 345681 116251 346223 136843
rect 346868 136826 346880 136892
rect 346990 136826 347002 136892
rect 347267 136845 358795 137369
rect 346868 136820 347002 136826
rect 348129 136827 358795 136845
rect 359337 136827 359343 137369
rect 346880 136816 346990 136820
rect 348129 116253 348671 136827
rect 345681 115709 346751 116251
rect 346926 116136 347036 116140
rect 346914 116130 347048 116136
rect 346914 116064 346926 116130
rect 347036 116064 347048 116130
rect 346914 116058 347048 116064
rect 346926 116054 347036 116058
rect 346936 115764 347046 115768
rect 346924 115758 347058 115764
rect 345681 95641 346223 115709
rect 346924 115692 346936 115758
rect 347046 115692 347058 115758
rect 347323 115711 348671 116253
rect 346924 115686 347058 115692
rect 346936 115682 347046 115686
rect 348129 95643 348671 115711
rect 345681 95639 346779 95641
rect 334793 95097 334799 95639
rect 335341 95099 346779 95639
rect 347351 95639 348671 95643
rect 346954 95526 347064 95530
rect 346942 95520 347076 95526
rect 346942 95454 346954 95520
rect 347064 95454 347076 95520
rect 346942 95448 347076 95454
rect 346954 95444 347064 95448
rect 346964 95154 347074 95158
rect 346952 95148 347086 95154
rect 335341 95097 346223 95099
rect 345681 74959 346223 95097
rect 346952 95082 346964 95148
rect 347074 95082 347086 95148
rect 347351 95101 359143 95639
rect 346952 95076 347086 95082
rect 348129 95097 359143 95101
rect 359685 95097 359691 95639
rect 346964 95072 347074 95076
rect 348129 74961 348671 95097
rect 345681 74417 346765 74959
rect 346940 74844 347050 74848
rect 346928 74838 347062 74844
rect 346928 74772 346940 74838
rect 347050 74772 347062 74838
rect 346928 74766 347062 74772
rect 346940 74762 347050 74766
rect 346950 74472 347060 74476
rect 346938 74466 347072 74472
rect 90274 58752 90284 60006
rect 91538 58752 91548 60006
rect 240075 59381 240617 59387
rect 133049 59371 133591 59377
rect 111727 59361 112269 59367
rect 39905 52861 40867 52867
rect 90667 52861 91209 58752
rect 30825 51899 39905 52861
rect 40867 51899 91209 52861
rect 30833 43125 31375 51899
rect 39905 51893 40867 51899
rect 48007 49071 48549 51899
rect 69301 49131 69843 51899
rect 90667 49057 91209 51899
rect 111727 49101 112269 58819
rect 133049 49145 133591 58829
rect 154607 59327 155149 59333
rect 154607 49115 155149 58785
rect 175813 59327 176355 59333
rect 219089 59305 219631 59311
rect 175813 49087 176355 58785
rect 197195 59283 197737 59289
rect 197195 49145 197737 58741
rect 219089 49057 219631 58763
rect 240075 49027 240617 58839
rect 260571 58837 260577 59379
rect 261119 58837 261125 59379
rect 260577 49087 261119 58837
rect 281383 58593 281389 59135
rect 281931 58593 281937 59135
rect 302573 58961 302579 59503
rect 303121 58961 303127 59503
rect 324121 58961 324127 59503
rect 324669 58961 324675 59503
rect 281389 49189 281931 58593
rect 281366 49004 281444 49016
rect 281738 49014 281816 49026
rect 69278 48946 69356 48958
rect 69650 48956 69728 48968
rect 133026 48960 133104 48972
rect 133398 48970 133476 48982
rect 47984 48886 48062 48898
rect 48356 48896 48434 48908
rect 47980 48776 47990 48886
rect 48056 48776 48066 48886
rect 48352 48786 48362 48896
rect 48428 48786 48438 48896
rect 69274 48836 69284 48946
rect 69350 48836 69360 48946
rect 69646 48846 69656 48956
rect 69722 48846 69732 48956
rect 111704 48916 111782 48928
rect 112076 48926 112154 48938
rect 90644 48872 90722 48884
rect 91016 48882 91094 48894
rect 69278 48824 69356 48836
rect 69650 48834 69728 48846
rect 47984 48764 48062 48776
rect 48356 48774 48434 48786
rect 90640 48762 90650 48872
rect 90716 48762 90726 48872
rect 91012 48772 91022 48882
rect 91088 48772 91098 48882
rect 111700 48806 111710 48916
rect 111776 48806 111786 48916
rect 112072 48816 112082 48926
rect 112148 48816 112158 48926
rect 133022 48850 133032 48960
rect 133098 48850 133108 48960
rect 133394 48860 133404 48970
rect 133470 48860 133480 48970
rect 197172 48960 197250 48972
rect 197544 48970 197622 48982
rect 154584 48930 154662 48942
rect 154956 48940 155034 48952
rect 133026 48838 133104 48850
rect 133398 48848 133476 48860
rect 154580 48820 154590 48930
rect 154656 48820 154666 48930
rect 154952 48830 154962 48940
rect 155028 48830 155038 48940
rect 175790 48902 175868 48914
rect 176162 48912 176240 48924
rect 111704 48794 111782 48806
rect 112076 48804 112154 48816
rect 154584 48808 154662 48820
rect 154956 48818 155034 48830
rect 175786 48792 175796 48902
rect 175862 48792 175872 48902
rect 176158 48802 176168 48912
rect 176234 48802 176244 48912
rect 197168 48850 197178 48960
rect 197244 48850 197254 48960
rect 197540 48860 197550 48970
rect 197616 48860 197626 48970
rect 260554 48902 260632 48914
rect 260926 48912 261004 48924
rect 219066 48872 219144 48884
rect 219438 48882 219516 48894
rect 197172 48838 197250 48850
rect 197544 48848 197622 48860
rect 175790 48780 175868 48792
rect 176162 48790 176240 48802
rect 90644 48750 90722 48762
rect 91016 48760 91094 48772
rect 219062 48762 219072 48872
rect 219138 48762 219148 48872
rect 219434 48772 219444 48882
rect 219510 48772 219520 48882
rect 240052 48842 240130 48854
rect 240424 48852 240502 48864
rect 219066 48750 219144 48762
rect 219438 48760 219516 48772
rect 240048 48732 240058 48842
rect 240124 48732 240134 48842
rect 240420 48742 240430 48852
rect 240496 48742 240506 48852
rect 260550 48792 260560 48902
rect 260626 48792 260636 48902
rect 260922 48802 260932 48912
rect 260998 48802 261008 48912
rect 281362 48894 281372 49004
rect 281438 48894 281448 49004
rect 281734 48904 281744 49014
rect 281810 48904 281820 49014
rect 302579 48983 303121 58961
rect 324127 49019 324669 58961
rect 334723 54525 335265 54531
rect 345681 54525 346223 74417
rect 346938 74400 346950 74466
rect 347060 74400 347072 74466
rect 347337 74419 348671 74961
rect 346938 74394 347072 74400
rect 346950 74390 347060 74394
rect 335265 53983 346223 54525
rect 334723 53977 335265 53983
rect 345681 51379 346223 53983
rect 348129 54525 348671 74419
rect 348129 53983 358805 54525
rect 359347 53983 359353 54525
rect 348129 51381 348671 53983
rect 345681 50837 346835 51379
rect 347010 51264 347120 51268
rect 346998 51258 347132 51264
rect 346998 51192 347010 51258
rect 347120 51192 347132 51258
rect 346998 51186 347132 51192
rect 347010 51182 347120 51186
rect 347020 50892 347130 50896
rect 347008 50886 347142 50892
rect 345681 50815 346223 50837
rect 347008 50820 347020 50886
rect 347130 50820 347142 50886
rect 347407 50839 348671 51381
rect 347008 50814 347142 50820
rect 347020 50810 347130 50814
rect 281366 48882 281444 48894
rect 281738 48892 281816 48904
rect 324104 48834 324182 48846
rect 324476 48844 324554 48856
rect 260554 48780 260632 48792
rect 260926 48790 261004 48802
rect 302556 48798 302634 48810
rect 302928 48808 303006 48820
rect 240052 48720 240130 48732
rect 240424 48730 240502 48742
rect 302552 48688 302562 48798
rect 302628 48688 302638 48798
rect 302924 48698 302934 48808
rect 303000 48698 303010 48808
rect 324100 48724 324110 48834
rect 324176 48724 324186 48834
rect 324472 48734 324482 48844
rect 324548 48734 324558 48844
rect 324104 48712 324182 48724
rect 324476 48722 324554 48734
rect 302556 48676 302634 48688
rect 302928 48686 303006 48698
rect 30833 42583 34403 43125
rect 34578 43010 34688 43014
rect 34566 43004 34700 43010
rect 34566 42938 34578 43004
rect 34688 42938 34700 43004
rect 34566 42932 34700 42938
rect 34578 42928 34688 42932
rect 34588 42638 34698 42642
rect 34576 42632 34710 42638
rect 30833 21027 31375 42583
rect 34576 42566 34588 42632
rect 34698 42566 34710 42632
rect 34975 42585 41467 43127
rect 34576 42560 34710 42566
rect 34588 42556 34698 42560
rect 40925 39258 41467 42585
rect 39640 36270 39650 39258
rect 42762 36270 42772 39258
rect 48009 37907 48551 48499
rect 69303 38013 69845 48559
rect 69303 37465 69845 37471
rect 90669 37695 91211 48485
rect 48009 37359 48551 37365
rect 111729 37747 112271 48529
rect 133051 37667 133593 48573
rect 154609 37835 155151 48543
rect 111729 37199 112271 37205
rect 90669 37147 91211 37153
rect 133045 37125 133051 37667
rect 133593 37125 133599 37667
rect 154609 37287 155151 37293
rect 175815 37835 176357 48515
rect 197197 37933 197739 48573
rect 197197 37385 197739 37391
rect 219091 37883 219633 48485
rect 240077 37781 240619 48455
rect 219091 37335 219633 37341
rect 175815 37287 176357 37293
rect 240071 37239 240077 37781
rect 240619 37239 240625 37781
rect 260579 37719 261121 48515
rect 281391 37815 281933 48617
rect 302581 37919 303123 48411
rect 260573 37177 260579 37719
rect 261121 37177 261127 37719
rect 281385 37273 281391 37815
rect 281933 37273 281939 37815
rect 302575 37377 302581 37919
rect 303123 37377 303129 37919
rect 324129 37867 324671 48447
rect 324123 37325 324129 37867
rect 324671 37325 324677 37867
rect 40925 21029 41467 36270
rect 30833 20485 34403 21027
rect 34578 20912 34688 20916
rect 34566 20906 34700 20912
rect 34566 20840 34578 20906
rect 34688 20840 34700 20906
rect 34566 20834 34700 20840
rect 34578 20830 34688 20834
rect 34588 20540 34698 20544
rect 34576 20534 34710 20540
rect 30833 5865 31375 20485
rect 34576 20468 34588 20534
rect 34698 20468 34710 20534
rect 34975 20487 41467 21029
rect 34576 20462 34710 20468
rect 34588 20458 34698 20462
rect 6571 5861 31375 5865
rect 6565 5323 31375 5861
rect 6565 3747 7107 5323
rect 27757 3807 28299 5323
rect 27734 3622 27812 3634
rect 28106 3632 28184 3644
rect 6542 3562 6620 3574
rect 6914 3572 6992 3584
rect 6538 3452 6548 3562
rect 6614 3452 6624 3562
rect 6910 3462 6920 3572
rect 6986 3462 6996 3572
rect 27730 3512 27740 3622
rect 27806 3512 27816 3622
rect 28102 3522 28112 3632
rect 28178 3522 28188 3632
rect 27734 3500 27812 3512
rect 28106 3510 28184 3522
rect 6542 3440 6620 3452
rect 6914 3450 6992 3462
rect 6567 2205 7109 3175
rect 27759 2205 28301 3235
rect 40925 2205 41467 20487
rect 6567 1671 41467 2205
rect 6571 1663 41467 1671
<< via1 >>
rect 550871 586751 550937 586861
rect 551243 586741 551309 586851
rect 571882 586782 571948 586892
rect 572254 586772 572320 586882
rect 537809 578721 538411 579323
rect 544736 573153 544846 573219
rect 544726 572781 544836 572847
rect 525320 567871 525386 567981
rect 525692 567861 525758 567971
rect 513762 562597 513872 562663
rect 513752 562225 513862 562291
rect 505449 560504 505559 560570
rect 505439 560132 505549 560198
rect 509408 554242 509938 556160
rect 526608 554236 527208 556182
rect 531032 553043 531142 553109
rect 547182 554212 547758 556178
rect 531022 552671 531132 552737
rect 544746 552904 544856 552970
rect 522511 550426 522621 550492
rect 522501 550054 522611 550120
rect 513742 542155 513852 542221
rect 505559 539916 505669 539982
rect 513732 541783 513842 541849
rect 464237 538845 464839 539447
rect 484628 538955 485230 539557
rect 500443 539029 501045 539631
rect 505549 539544 505659 539610
rect 355991 522045 356101 522111
rect 356001 521673 356111 521739
rect 517874 538396 518574 540212
rect 544736 552532 544846 552598
rect 537834 538328 538410 540294
rect 544751 532678 544861 532744
rect 544741 532306 544851 532372
rect 530987 531798 531097 531864
rect 530977 531426 531087 531492
rect 522560 529649 522670 529715
rect 522550 529277 522660 529343
rect 513739 522184 513849 522250
rect 513729 521812 513839 521878
rect 424259 519078 424325 519188
rect 424631 519068 424697 519178
rect 444272 519137 444338 519247
rect 444644 519127 444710 519237
rect 464455 519220 464521 519330
rect 464827 519210 464893 519320
rect 484787 519181 484853 519291
rect 485159 519171 485225 519281
rect 504261 519188 504327 519298
rect 504633 519178 504699 519288
rect 537690 519333 537756 519443
rect 538062 519323 538128 519433
rect 355956 502136 356066 502202
rect 355966 501764 356076 501830
rect 373616 490608 373726 490674
rect 373626 490236 373736 490302
rect 383268 490606 383378 490672
rect 383278 490234 383388 490300
rect 387905 490687 388015 490753
rect 387915 490315 388025 490381
rect 360443 484605 360985 485147
rect 375489 484747 376031 485289
rect 356018 482192 356128 482258
rect 346982 478252 347092 478318
rect 346992 477880 347102 477946
rect 356028 481820 356138 481886
rect 352781 472439 353323 472981
rect 346996 456998 347106 457064
rect 240701 455849 240811 455915
rect 240711 455477 240821 455543
rect 240621 434332 240731 434398
rect 240631 433960 240741 434026
rect 251423 455827 251533 455893
rect 251433 455455 251543 455521
rect 238866 429718 239407 430259
rect 251406 434046 251516 434112
rect 251416 433674 251526 433740
rect 249235 429837 249777 430379
rect 252980 429821 253522 430363
rect 252958 425977 253024 426087
rect 253330 425967 253396 426077
rect 242019 415360 242560 415901
rect 252972 415372 253512 415912
rect 347006 456626 347116 456692
rect 386095 484671 386637 485213
rect 384086 479600 384152 479710
rect 384458 479610 384524 479720
rect 379051 475499 379117 475609
rect 379423 475509 379489 475619
rect 380557 472617 381099 473159
rect 392808 490701 392918 490767
rect 392818 490329 392928 490395
rect 390329 484669 390871 485211
rect 389491 472541 390033 473083
rect 387914 469723 388024 469789
rect 387924 469351 388034 469417
rect 400223 484639 400765 485181
rect 428641 484679 429183 485221
rect 399541 479625 399607 479735
rect 399913 479635 399979 479745
rect 399541 475532 399607 475642
rect 399913 475542 399979 475652
rect 394697 472615 395239 473157
rect 392806 469723 392916 469789
rect 434805 484627 435407 485229
rect 419783 479565 419849 479675
rect 420155 479575 420221 479685
rect 419783 475472 419849 475582
rect 420155 475482 420221 475592
rect 400591 472567 401133 473109
rect 458519 484705 459121 485307
rect 440021 479594 440087 479704
rect 440393 479604 440459 479714
rect 440021 475501 440087 475611
rect 440393 475511 440459 475621
rect 428295 472567 428837 473109
rect 534334 508886 534444 508952
rect 534344 508514 534454 508580
rect 515038 507867 515148 507933
rect 515028 507495 515138 507561
rect 508942 506459 509052 506525
rect 508932 506087 509042 506153
rect 502178 500260 502288 500326
rect 502168 499888 502278 499954
rect 464290 484555 464892 485157
rect 475009 484525 475611 485127
rect 484628 484593 485230 485195
rect 531125 500809 531727 501411
rect 521392 498333 521502 498399
rect 521382 497961 521492 498027
rect 564230 497760 564296 497870
rect 564602 497750 564668 497860
rect 527466 495935 527576 496001
rect 527456 495563 527566 495629
rect 515001 487666 515111 487732
rect 514991 487294 515101 487360
rect 508954 486408 509064 486474
rect 508944 486036 509054 486102
rect 460321 479606 460387 479716
rect 460693 479616 460759 479726
rect 460321 475513 460387 475623
rect 460693 475523 460759 475633
rect 498503 484509 499105 485111
rect 504627 484563 505229 485165
rect 480503 479584 480569 479694
rect 480875 479594 480941 479704
rect 500459 479506 500525 479616
rect 500831 479496 500897 479606
rect 480503 475491 480569 475601
rect 480875 475501 480941 475611
rect 445483 472445 446085 473047
rect 462135 472457 462737 473059
rect 485297 472501 485899 473103
rect 500491 475509 500557 475619
rect 500863 475519 500929 475629
rect 497352 472566 497980 473194
rect 511844 484613 512446 485215
rect 518213 484585 518843 485215
rect 531125 491155 531727 491757
rect 534344 488486 534454 488552
rect 534354 488114 534464 488180
rect 524290 484557 524892 485159
rect 530389 484571 530991 485173
rect 531891 484591 532521 485221
rect 522909 479633 522975 479743
rect 523281 479643 523347 479753
rect 522941 475382 523007 475492
rect 523313 475372 523379 475482
rect 392816 469351 392926 469417
rect 503860 472370 504488 472998
rect 506695 472399 507297 473001
rect 518235 472485 518837 473087
rect 522944 472495 525127 473097
rect 356026 462172 356136 462238
rect 356036 461800 356146 461866
rect 508976 469023 509086 469089
rect 508986 468651 509096 468717
rect 502200 455171 502310 455237
rect 502210 454799 502320 454865
rect 356000 442179 356110 442245
rect 356010 441807 356120 441873
rect 346968 436390 347078 436456
rect 258338 429822 258878 430362
rect 272940 429757 273482 430299
rect 278450 429801 278992 430343
rect 293214 429813 293756 430355
rect 272904 426042 272970 426152
rect 273276 426032 273342 426142
rect 258312 420479 258378 420589
rect 258684 420469 258750 420579
rect 255273 415185 255815 415727
rect 258336 415336 258876 415876
rect 299162 429713 299704 430255
rect 293185 426076 293251 426186
rect 293557 426066 293623 426176
rect 278446 420512 278512 420622
rect 278818 420502 278884 420612
rect 272932 415267 273474 415809
rect 278450 415273 278992 415815
rect 313348 429649 313890 430191
rect 319476 429615 320018 430157
rect 322085 429673 322627 430215
rect 335394 429711 335936 430253
rect 313334 426066 313400 426176
rect 313706 426056 313772 426166
rect 299123 420518 299189 420628
rect 299495 420508 299561 420618
rect 319451 420470 319517 420580
rect 319823 420460 319889 420570
rect 335541 426041 335607 426151
rect 335913 426051 335979 426161
rect 324544 417112 324654 417178
rect 332869 420305 333411 420847
rect 324554 416740 324664 416806
rect 293214 415247 293756 415789
rect 299136 415271 299678 415813
rect 313354 415329 313896 415871
rect 319466 415405 320008 415947
rect 336554 417037 336664 417103
rect 336564 416665 336674 416731
rect 328159 415359 328701 415901
rect 346978 436018 347088 436084
rect 348094 429382 348522 430698
rect 387875 448703 387985 448769
rect 387885 448331 387995 448397
rect 339875 415321 340417 415863
rect 345550 414894 345978 416210
rect 354357 429727 354899 430269
rect 360001 429897 360543 430439
rect 362171 429901 362713 430443
rect 355531 426037 355597 426147
rect 355903 426047 355969 426157
rect 373950 429649 374492 430191
rect 375352 429653 375894 430195
rect 385933 429745 386475 430287
rect 356005 422225 356115 422291
rect 353761 420469 353827 420579
rect 354133 420479 354199 420589
rect 346912 415756 347022 415822
rect 346922 415384 347032 415450
rect 324542 396322 324652 396388
rect 324552 395950 324662 396016
rect 322895 390805 323437 391347
rect 336579 396384 336689 396450
rect 336589 396012 336699 396078
rect 333092 390825 333634 391367
rect 334879 390767 335421 391309
rect 333077 380647 333143 380757
rect 333449 380637 333515 380747
rect 325765 375553 326307 376095
rect 333090 375667 333632 376209
rect 356015 421853 356125 421919
rect 387904 427660 388014 427726
rect 392796 448771 392906 448837
rect 392806 448399 392916 448465
rect 391205 429829 391747 430371
rect 387914 427288 388024 427354
rect 392828 427679 392938 427745
rect 508964 448972 509074 449038
rect 508974 448600 509084 448666
rect 497210 429770 497838 430398
rect 510283 429683 510885 430285
rect 515023 467765 515133 467831
rect 515033 467393 515143 467459
rect 550466 491990 550576 492056
rect 550456 491618 550566 491684
rect 545784 484497 546414 485127
rect 545802 479510 545868 479620
rect 546174 479500 546240 479610
rect 545855 475418 545921 475528
rect 546227 475408 546293 475518
rect 536943 472561 537545 473163
rect 537957 472511 538587 473141
rect 548153 472577 548783 473207
rect 553163 472501 553793 473131
rect 567849 484541 568479 485171
rect 534386 466945 534496 467011
rect 534376 466573 534486 466639
rect 527531 459536 527641 459602
rect 527521 459164 527631 459230
rect 521414 457098 521524 457164
rect 521424 456726 521534 456792
rect 515060 447564 515170 447630
rect 515070 447192 515180 447258
rect 513067 429733 513669 430335
rect 562803 472429 563433 473059
rect 534376 446545 534486 446611
rect 534366 446173 534476 446239
rect 550370 459665 550480 459731
rect 550360 459293 550470 459359
rect 564164 453285 564230 453395
rect 564536 453295 564602 453405
rect 522311 429699 522913 430301
rect 528959 429699 529589 430329
rect 545783 429773 546413 430403
rect 562801 429699 563431 430329
rect 392838 427307 392948 427373
rect 375494 426131 375560 426241
rect 375866 426141 375932 426251
rect 374104 420539 374170 420649
rect 374476 420549 374542 420659
rect 353573 415233 354115 415775
rect 373944 415303 374486 415845
rect 375340 415107 375882 415649
rect 388617 415307 389159 415849
rect 393665 415385 394207 415927
rect 568046 408878 568112 408988
rect 568418 408868 568484 408978
rect 549553 407130 549663 407196
rect 355994 402190 356104 402256
rect 356004 401818 356114 401884
rect 346940 395078 347050 395144
rect 346950 394706 347060 394772
rect 353565 390397 354107 390939
rect 357690 390615 358232 391157
rect 367484 390651 368026 391193
rect 347446 386614 347512 386724
rect 347818 386604 347884 386714
rect 337333 375573 337875 376115
rect 385269 390627 385811 391169
rect 400437 390647 400979 391189
rect 428501 390755 429043 391297
rect 549543 406758 549653 406824
rect 367462 386643 367528 386753
rect 367834 386633 367900 386743
rect 355974 382126 356084 382192
rect 355984 381754 356094 381820
rect 357656 380655 357722 380765
rect 358028 380645 358094 380755
rect 345681 375547 346223 376089
rect 352330 375608 353838 376280
rect 346926 373796 347036 373862
rect 346936 373424 347046 373490
rect 346926 352946 347036 353012
rect 346936 352574 347046 352640
rect 347010 332350 347120 332416
rect 347020 331978 347130 332044
rect 346982 310482 347092 310548
rect 346992 310110 347102 310176
rect 348024 305644 348476 307618
rect 346940 288824 347050 288890
rect 346950 288452 347060 288518
rect 345710 285614 346162 287588
rect 357684 375559 358226 376101
rect 446395 390507 446937 391049
rect 470027 390513 470569 391055
rect 490269 390563 490811 391105
rect 387274 386633 387340 386743
rect 387646 386623 387712 386733
rect 387103 380613 387169 380723
rect 387475 380603 387541 380713
rect 407533 386631 407599 386741
rect 407905 386621 407971 386731
rect 407681 380644 407747 380754
rect 408053 380634 408119 380744
rect 510723 390533 511265 391075
rect 530385 390605 530927 391147
rect 546403 390679 546965 391241
rect 427809 386686 427875 386796
rect 428181 386676 428247 386786
rect 427655 380619 427721 380729
rect 428027 380609 428093 380719
rect 447968 386666 448034 386776
rect 448340 386656 448406 386766
rect 467970 386661 468036 386771
rect 468342 386651 468408 386761
rect 447901 380623 447967 380733
rect 448273 380613 448339 380723
rect 367484 375509 368026 376051
rect 388559 375377 389101 375919
rect 400425 375559 400967 376101
rect 488088 386645 488154 386755
rect 488460 386635 488526 386745
rect 467885 380690 467951 380800
rect 468257 380680 468323 380790
rect 508218 386668 508284 386778
rect 508590 386658 508656 386768
rect 488300 380615 488366 380725
rect 488672 380605 488738 380715
rect 429149 375465 429691 376007
rect 446411 375523 446953 376065
rect 528327 386682 528393 386792
rect 528699 386672 528765 386782
rect 507983 380687 508049 380797
rect 508355 380677 508421 380787
rect 549570 388086 549680 388152
rect 528353 380621 528419 380731
rect 528725 380611 528791 380721
rect 466549 375507 467091 376049
rect 485509 375463 486051 376005
rect 549560 387714 549670 387780
rect 549368 379428 549478 379494
rect 549378 379056 549488 379122
rect 505733 375447 506275 375989
rect 526305 375627 526847 376169
rect 571227 390643 571789 391205
rect 552361 375485 552923 376047
rect 562709 375559 563271 376121
rect 549329 364242 549439 364308
rect 549339 363870 549449 363936
rect 356031 362143 356141 362209
rect 356041 361771 356151 361837
rect 568202 362495 568268 362605
rect 568574 362485 568640 362595
rect 356031 342140 356141 342206
rect 356041 341768 356151 341834
rect 355955 322138 356065 322204
rect 355965 321766 356075 321832
rect 357945 306237 358487 306779
rect 355993 302117 356103 302183
rect 356003 301745 356113 301811
rect 370688 306263 371237 306812
rect 390700 306391 391249 306940
rect 400264 306349 400813 306898
rect 430714 306113 431263 306662
rect 445440 306311 445989 306860
rect 470718 306231 471267 306780
rect 490714 306455 491263 307004
rect 510700 306347 511249 306896
rect 530686 306193 531235 306742
rect 552167 306173 552724 306730
rect 569358 306237 569927 306806
rect 370828 295924 370894 296034
rect 371200 295934 371266 296044
rect 390837 295941 390903 296051
rect 391209 295951 391275 296061
rect 410843 295912 410909 296022
rect 411215 295922 411281 296032
rect 430839 295988 430905 296098
rect 431211 295998 431277 296108
rect 450856 295955 450922 296065
rect 451228 295965 451294 296075
rect 470858 295980 470924 296090
rect 471230 295990 471296 296100
rect 490853 296013 490919 296123
rect 491225 296023 491291 296133
rect 510846 295969 510912 296079
rect 511218 295979 511284 296089
rect 530831 296013 530897 296123
rect 531203 296023 531269 296133
rect 354041 286271 354583 286813
rect 370688 286058 371237 286607
rect 390700 286142 391249 286691
rect 400180 286354 400729 286903
rect 430714 286260 431263 286809
rect 445452 286472 446001 287021
rect 470718 286204 471267 286753
rect 490714 286334 491263 286883
rect 510700 286270 511249 286819
rect 549547 293375 549657 293441
rect 549557 293003 549667 293069
rect 530686 286258 531235 286807
rect 546320 286426 546877 286983
rect 568318 286313 568887 286882
rect 551449 273906 551515 274016
rect 551821 273916 551887 274026
rect 571912 273866 571978 273976
rect 572284 273876 572350 273986
rect 346898 264044 347008 264110
rect 346908 263672 347018 263738
rect 346982 242670 347092 242736
rect 346992 242298 347102 242364
rect 347010 222794 347120 222860
rect 347020 222422 347130 222488
rect 347982 208088 348448 213096
rect 346954 200966 347064 201032
rect 346964 200594 347074 200660
rect 346968 179932 347078 179998
rect 346978 179560 347088 179626
rect 345722 172818 346188 177826
rect 345698 162828 346164 167836
rect 346926 158544 347036 158610
rect 346936 158172 347046 158238
rect 334827 136843 335369 137385
rect 346870 137198 346980 137264
rect 346880 136826 346990 136892
rect 358795 136827 359337 137369
rect 346926 116064 347036 116130
rect 346936 115692 347046 115758
rect 334799 95097 335341 95639
rect 346954 95454 347064 95520
rect 346964 95082 347074 95148
rect 359143 95097 359685 95639
rect 346940 74772 347050 74838
rect 90284 58752 91538 60006
rect 111727 58819 112269 59361
rect 39905 51899 40867 52861
rect 133049 58829 133591 59371
rect 154607 58785 155149 59327
rect 175813 58785 176355 59327
rect 197195 58741 197737 59283
rect 219089 58763 219631 59305
rect 240075 58839 240617 59381
rect 260577 58837 261119 59379
rect 281389 58593 281931 59135
rect 302579 58961 303121 59503
rect 324127 58961 324669 59503
rect 47990 48776 48056 48886
rect 48362 48786 48428 48896
rect 69284 48836 69350 48946
rect 69656 48846 69722 48956
rect 90650 48762 90716 48872
rect 91022 48772 91088 48882
rect 111710 48806 111776 48916
rect 112082 48816 112148 48926
rect 133032 48850 133098 48960
rect 133404 48860 133470 48970
rect 154590 48820 154656 48930
rect 154962 48830 155028 48940
rect 175796 48792 175862 48902
rect 176168 48802 176234 48912
rect 197178 48850 197244 48960
rect 197550 48860 197616 48970
rect 219072 48762 219138 48872
rect 219444 48772 219510 48882
rect 240058 48732 240124 48842
rect 240430 48742 240496 48852
rect 260560 48792 260626 48902
rect 260932 48802 260998 48912
rect 281372 48894 281438 49004
rect 281744 48904 281810 49014
rect 346950 74400 347060 74466
rect 334723 53983 335265 54525
rect 358805 53983 359347 54525
rect 347010 51192 347120 51258
rect 347020 50820 347130 50886
rect 302562 48688 302628 48798
rect 302934 48698 303000 48808
rect 324110 48724 324176 48834
rect 324482 48734 324548 48844
rect 34578 42938 34688 43004
rect 34588 42566 34698 42632
rect 39650 36270 42762 39258
rect 48009 37365 48551 37907
rect 69303 37471 69845 38013
rect 90669 37153 91211 37695
rect 111729 37205 112271 37747
rect 133051 37125 133593 37667
rect 154609 37293 155151 37835
rect 175815 37293 176357 37835
rect 197197 37391 197739 37933
rect 219091 37341 219633 37883
rect 240077 37239 240619 37781
rect 260579 37177 261121 37719
rect 281391 37273 281933 37815
rect 302581 37377 303123 37919
rect 324129 37325 324671 37867
rect 34578 20840 34688 20906
rect 34588 20468 34698 20534
rect 6548 3452 6614 3562
rect 6920 3462 6986 3572
rect 27740 3512 27806 3622
rect 28112 3522 28178 3632
<< metal2 >>
rect 571882 586892 571948 586902
rect 550871 586861 550937 586871
rect 550861 586751 550871 586861
rect 550937 586751 550947 586861
rect 551243 586851 551309 586861
rect 550871 586741 550937 586751
rect 551233 586741 551243 586851
rect 551309 586741 551319 586851
rect 571872 586782 571882 586892
rect 571948 586782 571958 586892
rect 572254 586882 572320 586892
rect 571882 586772 571948 586782
rect 572244 586772 572254 586882
rect 572320 586772 572330 586882
rect 572254 586762 572320 586772
rect 551243 586731 551309 586741
rect 537809 579323 538411 579329
rect 537800 578721 537809 579323
rect 538411 578721 538420 579323
rect 537809 578715 538411 578721
rect 544736 573219 544846 573229
rect 544726 573153 544736 573219
rect 544846 573153 544856 573219
rect 544736 573143 544846 573153
rect 544726 572847 544836 572857
rect 544716 572781 544726 572847
rect 544836 572781 544846 572847
rect 544726 572771 544836 572781
rect 525320 567981 525386 567991
rect 525310 567871 525320 567981
rect 525386 567871 525396 567981
rect 525692 567971 525758 567981
rect 525320 567861 525386 567871
rect 525682 567861 525692 567971
rect 525758 567861 525768 567971
rect 525692 567851 525758 567861
rect 513762 562663 513872 562673
rect 513752 562597 513762 562663
rect 513872 562597 513882 562663
rect 513762 562587 513872 562597
rect 513752 562291 513862 562301
rect 513742 562225 513752 562291
rect 513862 562225 513872 562291
rect 513752 562215 513862 562225
rect 505449 560570 505559 560580
rect 505439 560504 505449 560570
rect 505559 560504 505569 560570
rect 505449 560494 505559 560504
rect 505439 560198 505549 560208
rect 505429 560132 505439 560198
rect 505549 560132 505559 560198
rect 505439 560122 505549 560132
rect 526608 556182 527208 556192
rect 509408 556160 509938 556170
rect 509408 554232 509938 554242
rect 526608 554226 527208 554236
rect 547182 556178 547758 556188
rect 547182 554202 547758 554212
rect 531032 553109 531142 553119
rect 531022 553043 531032 553109
rect 531142 553043 531152 553109
rect 531032 553033 531142 553043
rect 544746 552970 544856 552980
rect 544736 552904 544746 552970
rect 544856 552904 544866 552970
rect 544746 552894 544856 552904
rect 531022 552737 531132 552747
rect 531012 552671 531022 552737
rect 531132 552671 531142 552737
rect 531022 552661 531132 552671
rect 544736 552598 544846 552608
rect 544726 552532 544736 552598
rect 544846 552532 544856 552598
rect 544736 552522 544846 552532
rect 522511 550492 522621 550502
rect 522501 550426 522511 550492
rect 522621 550426 522631 550492
rect 522511 550416 522621 550426
rect 522501 550120 522611 550130
rect 522491 550054 522501 550120
rect 522611 550054 522621 550120
rect 522501 550044 522611 550054
rect 513742 542221 513852 542231
rect 513732 542155 513742 542221
rect 513852 542155 513862 542221
rect 513742 542145 513852 542155
rect 513732 541849 513842 541859
rect 513722 541783 513732 541849
rect 513842 541783 513852 541849
rect 513732 541773 513842 541783
rect 537834 540294 538410 540304
rect 517874 540212 518574 540222
rect 505559 539982 505669 539992
rect 505549 539916 505559 539982
rect 505669 539916 505679 539982
rect 505559 539906 505669 539916
rect 500443 539631 501045 539640
rect 484628 539557 485230 539563
rect 464237 539447 464839 539453
rect 464228 538845 464237 539447
rect 464839 538845 464848 539447
rect 484619 538955 484628 539557
rect 485230 538955 485239 539557
rect 500437 539029 500443 539631
rect 501045 539029 501051 539631
rect 505549 539610 505659 539620
rect 505539 539544 505549 539610
rect 505659 539544 505669 539610
rect 505549 539534 505659 539544
rect 500443 539020 501045 539029
rect 484628 538949 485230 538955
rect 464237 538839 464839 538845
rect 517874 538386 518574 538396
rect 537834 538318 538410 538328
rect 373663 535258 373691 535458
rect 402367 535238 402395 535432
rect 544751 532744 544861 532754
rect 544741 532678 544751 532744
rect 544861 532678 544871 532744
rect 544751 532668 544861 532678
rect 544741 532372 544851 532382
rect 544731 532306 544741 532372
rect 544851 532306 544861 532372
rect 544741 532296 544851 532306
rect 530987 531864 531097 531874
rect 530977 531798 530987 531864
rect 531097 531798 531107 531864
rect 530987 531788 531097 531798
rect 530977 531492 531087 531502
rect 530967 531426 530977 531492
rect 531087 531426 531097 531492
rect 530977 531416 531087 531426
rect 522560 529715 522670 529725
rect 522550 529649 522560 529715
rect 522670 529649 522680 529715
rect 522560 529639 522670 529649
rect 522550 529343 522660 529353
rect 522540 529277 522550 529343
rect 522660 529277 522670 529343
rect 522550 529267 522660 529277
rect 355981 522045 355991 522111
rect 356101 522045 356111 522111
rect 355991 521673 356001 521739
rect 356111 521673 356121 521739
rect 372200 516868 372209 516928
rect 372269 516912 372278 516928
rect 373663 516912 373691 522678
rect 513739 522250 513849 522260
rect 513729 522184 513739 522250
rect 513849 522184 513859 522250
rect 513739 522174 513849 522184
rect 513729 521878 513839 521888
rect 513719 521812 513729 521878
rect 513839 521812 513849 521878
rect 513729 521802 513839 521812
rect 402367 519092 402395 520676
rect 537690 519443 537756 519453
rect 464455 519330 464521 519340
rect 537680 519333 537690 519443
rect 537756 519333 537766 519443
rect 538062 519433 538128 519443
rect 444272 519247 444338 519257
rect 424259 519188 424325 519198
rect 403600 519092 403609 519108
rect 402367 519064 403609 519092
rect 403600 519048 403609 519064
rect 403669 519092 403678 519108
rect 403669 519064 403709 519092
rect 424259 519068 424325 519078
rect 424631 519178 424697 519188
rect 444272 519127 444338 519137
rect 444644 519237 444710 519247
rect 464455 519210 464521 519220
rect 464827 519320 464893 519330
rect 537690 519323 537756 519333
rect 538052 519323 538062 519433
rect 538128 519323 538138 519433
rect 538062 519313 538128 519323
rect 464827 519200 464893 519210
rect 484787 519291 484853 519301
rect 504261 519298 504327 519308
rect 484787 519171 484853 519181
rect 485159 519281 485225 519291
rect 504261 519178 504327 519188
rect 504633 519288 504699 519298
rect 485159 519161 485225 519171
rect 504633 519168 504699 519178
rect 444644 519117 444710 519127
rect 403669 519048 403678 519064
rect 424631 519058 424697 519068
rect 372269 516884 373691 516912
rect 372269 516868 372278 516884
rect 534334 508952 534444 508962
rect 534324 508886 534334 508952
rect 534444 508886 534454 508952
rect 534334 508876 534444 508886
rect 534344 508580 534454 508590
rect 534334 508514 534344 508580
rect 534454 508514 534464 508580
rect 534344 508504 534454 508514
rect 373663 504711 373691 507736
rect 383231 504757 383259 507813
rect 373647 504702 373707 504711
rect 383206 504697 383215 504757
rect 383275 504697 383284 504757
rect 392799 504716 392827 507951
rect 515038 507933 515148 507943
rect 402367 507506 402395 507914
rect 515028 507867 515038 507933
rect 515148 507867 515158 507933
rect 515038 507857 515148 507867
rect 515028 507561 515138 507571
rect 515018 507495 515028 507561
rect 515138 507495 515148 507561
rect 515028 507485 515138 507495
rect 508942 506525 509052 506535
rect 508932 506459 508942 506525
rect 509052 506459 509062 506525
rect 508942 506449 509052 506459
rect 508932 506153 509042 506163
rect 508922 506087 508932 506153
rect 509042 506087 509052 506153
rect 508932 506077 509042 506087
rect 392774 504656 392783 504716
rect 392843 504656 392852 504716
rect 373647 504633 373707 504642
rect 355946 502136 355956 502202
rect 356066 502136 356076 502202
rect 355956 501764 355966 501830
rect 356076 501764 356086 501830
rect 531119 500809 531125 501411
rect 531727 500809 531733 501411
rect 502178 500326 502288 500336
rect 502168 500260 502178 500326
rect 502288 500260 502298 500326
rect 502178 500250 502288 500260
rect 502168 499954 502278 499964
rect 502158 499888 502168 499954
rect 502278 499888 502288 499954
rect 502168 499878 502278 499888
rect 521392 498399 521502 498409
rect 521382 498333 521392 498399
rect 521502 498333 521512 498399
rect 521392 498323 521502 498333
rect 521382 498027 521492 498037
rect 521372 497961 521382 498027
rect 521492 497961 521502 498027
rect 521382 497951 521492 497961
rect 527466 496001 527576 496011
rect 527456 495935 527466 496001
rect 527576 495935 527586 496001
rect 527466 495925 527576 495935
rect 527456 495629 527566 495639
rect 527446 495563 527456 495629
rect 527566 495563 527576 495629
rect 527456 495553 527566 495563
rect 531125 491757 531727 500809
rect 564230 497870 564296 497880
rect 564220 497760 564230 497870
rect 564296 497760 564306 497870
rect 564602 497860 564668 497870
rect 564230 497750 564296 497760
rect 564592 497750 564602 497860
rect 564668 497750 564678 497860
rect 564602 497740 564668 497750
rect 550466 492056 550576 492066
rect 550456 491990 550466 492056
rect 550576 491990 550586 492056
rect 550466 491980 550576 491990
rect 531119 491155 531125 491757
rect 531727 491155 531733 491757
rect 550456 491684 550566 491694
rect 550446 491618 550456 491684
rect 550566 491618 550576 491684
rect 550456 491608 550566 491618
rect 387895 490687 387905 490753
rect 388015 490687 388025 490753
rect 392798 490701 392808 490767
rect 392918 490701 392928 490767
rect 373606 490608 373616 490674
rect 373726 490608 373736 490674
rect 383258 490606 383268 490672
rect 383378 490606 383388 490672
rect 387905 490315 387915 490381
rect 388025 490315 388035 490381
rect 392808 490329 392818 490395
rect 392928 490329 392938 490395
rect 373616 490236 373626 490302
rect 373736 490236 373746 490302
rect 383268 490234 383278 490300
rect 383388 490234 383398 490300
rect 534344 488552 534454 488562
rect 534334 488486 534344 488552
rect 534454 488486 534464 488552
rect 534344 488476 534454 488486
rect 534354 488180 534464 488190
rect 534344 488114 534354 488180
rect 534464 488114 534474 488180
rect 534354 488104 534464 488114
rect 515001 487732 515111 487742
rect 514991 487666 515001 487732
rect 515111 487666 515121 487732
rect 515001 487656 515111 487666
rect 514991 487360 515101 487370
rect 514981 487294 514991 487360
rect 515101 487294 515111 487360
rect 514991 487284 515101 487294
rect 508954 486474 509064 486484
rect 508944 486408 508954 486474
rect 509064 486408 509074 486474
rect 508954 486398 509064 486408
rect 508944 486102 509054 486112
rect 508934 486036 508944 486102
rect 509054 486036 509064 486102
rect 508944 486026 509054 486036
rect 458519 485307 459121 485316
rect 375489 485289 376031 485298
rect 360443 485147 360985 485156
rect 360437 484605 360443 485147
rect 360985 484605 360991 485147
rect 375483 484747 375489 485289
rect 376031 484747 376037 485289
rect 386095 485213 386637 485222
rect 428641 485221 429183 485230
rect 434805 485229 435407 485238
rect 375489 484738 376031 484747
rect 386089 484671 386095 485213
rect 386637 484671 386643 485213
rect 390329 485211 390871 485220
rect 386095 484662 386637 484671
rect 390323 484669 390329 485211
rect 390871 484669 390877 485211
rect 400223 485181 400765 485190
rect 390329 484660 390871 484669
rect 400217 484639 400223 485181
rect 400765 484639 400771 485181
rect 428635 484679 428641 485221
rect 429183 484679 429189 485221
rect 428641 484670 429183 484679
rect 400223 484630 400765 484639
rect 434799 484627 434805 485229
rect 435407 484627 435413 485229
rect 458513 484705 458519 485307
rect 459121 484705 459127 485307
rect 531891 485221 532521 485230
rect 511844 485215 512446 485221
rect 518213 485215 518843 485221
rect 484628 485195 485230 485201
rect 464290 485157 464892 485166
rect 458519 484696 459121 484705
rect 434805 484618 435407 484627
rect 360443 484596 360985 484605
rect 464284 484555 464290 485157
rect 464892 484555 464898 485157
rect 475009 485127 475611 485136
rect 464290 484546 464892 484555
rect 475003 484525 475009 485127
rect 475611 484525 475617 485127
rect 484619 484593 484628 485195
rect 485230 484593 485239 485195
rect 504627 485165 505229 485174
rect 498503 485111 499105 485117
rect 484628 484587 485230 484593
rect 475009 484516 475611 484525
rect 498494 484509 498503 485111
rect 499105 484509 499114 485111
rect 504621 484563 504627 485165
rect 505229 484563 505235 485165
rect 511835 484613 511844 485215
rect 512446 484613 512455 485215
rect 511844 484607 512446 484613
rect 518204 484585 518213 485215
rect 518843 484585 518852 485215
rect 530389 485173 530991 485182
rect 524290 485159 524892 485165
rect 518213 484579 518843 484585
rect 504627 484554 505229 484563
rect 524281 484557 524290 485159
rect 524892 484557 524901 485159
rect 530383 484571 530389 485173
rect 530991 484571 530997 485173
rect 531885 484591 531891 485221
rect 532521 484591 532527 485221
rect 567849 485171 568479 485177
rect 545784 485127 546414 485133
rect 531891 484582 532521 484591
rect 530389 484562 530991 484571
rect 524290 484551 524892 484557
rect 498503 484503 499105 484509
rect 545775 484497 545784 485127
rect 546414 484497 546423 485127
rect 567840 484541 567849 485171
rect 568479 484541 568488 485171
rect 567849 484535 568479 484541
rect 545784 484491 546414 484497
rect 356008 482192 356018 482258
rect 356128 482192 356138 482258
rect 356018 481820 356028 481886
rect 356138 481820 356148 481886
rect 399913 479745 399979 479755
rect 523281 479753 523347 479763
rect 399541 479735 399607 479745
rect 384458 479720 384524 479730
rect 384086 479710 384152 479720
rect 522909 479743 522975 479753
rect 460693 479726 460759 479736
rect 440393 479714 440459 479724
rect 440021 479704 440087 479714
rect 420155 479685 420221 479695
rect 399913 479625 399979 479635
rect 419783 479675 419849 479685
rect 399541 479615 399607 479625
rect 384458 479600 384524 479610
rect 384086 479590 384152 479600
rect 440393 479594 440459 479604
rect 460321 479716 460387 479726
rect 480875 479704 480941 479714
rect 460693 479606 460759 479616
rect 480503 479694 480569 479704
rect 460321 479596 460387 479606
rect 440021 479584 440087 479594
rect 523281 479633 523347 479643
rect 480875 479584 480941 479594
rect 500459 479616 500525 479626
rect 522909 479623 522975 479633
rect 545802 479620 545868 479630
rect 420155 479565 420221 479575
rect 480503 479574 480569 479584
rect 419783 479555 419849 479565
rect 500459 479496 500525 479506
rect 500831 479606 500897 479616
rect 545792 479510 545802 479620
rect 545868 479510 545878 479620
rect 546174 479610 546240 479620
rect 545802 479500 545868 479510
rect 546164 479500 546174 479610
rect 546240 479500 546250 479610
rect 500831 479486 500897 479496
rect 546174 479490 546240 479500
rect 346972 478252 346982 478318
rect 347092 478252 347102 478318
rect 346982 477880 346992 477946
rect 347102 477880 347112 477946
rect 399913 475652 399979 475662
rect 399541 475642 399607 475652
rect 379423 475619 379489 475629
rect 379051 475609 379117 475619
rect 460693 475633 460759 475643
rect 440393 475621 440459 475631
rect 440021 475611 440087 475621
rect 420155 475592 420221 475602
rect 399913 475532 399979 475542
rect 419783 475582 419849 475592
rect 399541 475522 399607 475532
rect 379423 475499 379489 475509
rect 379051 475489 379117 475499
rect 440393 475501 440459 475511
rect 460321 475623 460387 475633
rect 500863 475629 500929 475639
rect 480875 475611 480941 475621
rect 460693 475513 460759 475523
rect 480503 475601 480569 475611
rect 460321 475503 460387 475513
rect 440021 475491 440087 475501
rect 480875 475491 480941 475501
rect 500491 475619 500557 475629
rect 545855 475528 545921 475538
rect 500863 475509 500929 475519
rect 500491 475499 500557 475509
rect 522941 475492 523007 475502
rect 420155 475472 420221 475482
rect 480503 475481 480569 475491
rect 419783 475462 419849 475472
rect 522941 475372 523007 475382
rect 523313 475482 523379 475492
rect 545845 475418 545855 475528
rect 545921 475418 545931 475528
rect 546227 475518 546293 475528
rect 545855 475408 545921 475418
rect 546217 475408 546227 475518
rect 546293 475408 546303 475518
rect 546227 475398 546293 475408
rect 523313 475362 523379 475372
rect 548153 473207 548783 473213
rect 497352 473194 497980 473203
rect 380557 473159 381099 473165
rect 352781 472981 353323 472987
rect 352772 472439 352781 472981
rect 353323 472439 353332 472981
rect 380548 472617 380557 473159
rect 381099 472617 381108 473159
rect 394697 473157 395239 473166
rect 389491 473083 390033 473092
rect 380557 472611 381099 472617
rect 389485 472541 389491 473083
rect 390033 472541 390039 473083
rect 394691 472615 394697 473157
rect 395239 472615 395245 473157
rect 400591 473109 401133 473118
rect 428295 473109 428837 473118
rect 394697 472606 395239 472615
rect 400585 472567 400591 473109
rect 401133 472567 401139 473109
rect 428289 472567 428295 473109
rect 428837 472567 428843 473109
rect 485297 473103 485899 473112
rect 462135 473059 462737 473068
rect 445483 473047 446085 473056
rect 400591 472558 401133 472567
rect 428295 472558 428837 472567
rect 389491 472532 390033 472541
rect 445477 472445 445483 473047
rect 446085 472445 446091 473047
rect 462129 472457 462135 473059
rect 462737 472457 462743 473059
rect 485291 472501 485297 473103
rect 485899 472501 485905 473103
rect 497346 472566 497352 473194
rect 497980 472566 497986 473194
rect 536943 473163 537545 473169
rect 522944 473097 525127 473107
rect 518235 473087 518837 473093
rect 503860 472998 504488 473007
rect 506695 473001 507297 473007
rect 497352 472557 497980 472566
rect 485297 472492 485899 472501
rect 462135 472448 462737 472457
rect 352781 472433 353323 472439
rect 445483 472436 446085 472445
rect 503854 472370 503860 472998
rect 504488 472370 504494 472998
rect 506686 472399 506695 473001
rect 507297 472399 507306 473001
rect 518226 472485 518235 473087
rect 518837 472485 518846 473087
rect 536934 472561 536943 473163
rect 537545 472561 537554 473163
rect 537957 473141 538587 473147
rect 536943 472555 537545 472561
rect 537948 472511 537957 473141
rect 538587 472511 538596 473141
rect 548144 472577 548153 473207
rect 548783 472577 548792 473207
rect 553163 473131 553793 473137
rect 548153 472571 548783 472577
rect 537957 472505 538587 472511
rect 553154 472501 553163 473131
rect 553793 472501 553802 473131
rect 562803 473059 563433 473068
rect 553163 472495 553793 472501
rect 522944 472485 525127 472495
rect 518235 472479 518837 472485
rect 562797 472429 562803 473059
rect 563433 472429 563439 473059
rect 562803 472420 563433 472429
rect 506695 472393 507297 472399
rect 503860 472361 504488 472370
rect 387904 469723 387914 469789
rect 388024 469723 388034 469789
rect 392796 469723 392806 469789
rect 392916 469723 392926 469789
rect 387914 469351 387924 469417
rect 388034 469351 388044 469417
rect 392806 469351 392816 469417
rect 392926 469351 392936 469417
rect 508976 469089 509086 469099
rect 508966 469023 508976 469089
rect 509086 469023 509096 469089
rect 508976 469013 509086 469023
rect 508986 468717 509096 468727
rect 508976 468651 508986 468717
rect 509096 468651 509106 468717
rect 508986 468641 509096 468651
rect 515023 467831 515133 467841
rect 515013 467765 515023 467831
rect 515133 467765 515143 467831
rect 515023 467755 515133 467765
rect 515033 467459 515143 467469
rect 515023 467393 515033 467459
rect 515143 467393 515153 467459
rect 515033 467383 515143 467393
rect 534386 467011 534496 467021
rect 534376 466945 534386 467011
rect 534496 466945 534506 467011
rect 534386 466935 534496 466945
rect 534376 466639 534486 466649
rect 534366 466573 534376 466639
rect 534486 466573 534496 466639
rect 534376 466563 534486 466573
rect 356016 462172 356026 462238
rect 356136 462172 356146 462238
rect 356026 461800 356036 461866
rect 356146 461800 356156 461866
rect 550370 459731 550480 459741
rect 550360 459665 550370 459731
rect 550480 459665 550490 459731
rect 550370 459655 550480 459665
rect 527531 459602 527641 459612
rect 527521 459536 527531 459602
rect 527641 459536 527651 459602
rect 527531 459526 527641 459536
rect 550360 459359 550470 459369
rect 550350 459293 550360 459359
rect 550470 459293 550480 459359
rect 550360 459283 550470 459293
rect 527521 459230 527631 459240
rect 527511 459164 527521 459230
rect 527631 459164 527641 459230
rect 527521 459154 527631 459164
rect 521414 457164 521524 457174
rect 521404 457098 521414 457164
rect 521524 457098 521534 457164
rect 521414 457088 521524 457098
rect 346986 456998 346996 457064
rect 347106 456998 347116 457064
rect 521424 456792 521534 456802
rect 521414 456726 521424 456792
rect 521534 456726 521544 456792
rect 521424 456716 521534 456726
rect 346996 456626 347006 456692
rect 347116 456626 347126 456692
rect 240691 455849 240701 455915
rect 240811 455849 240821 455915
rect 251413 455827 251423 455893
rect 251533 455827 251543 455893
rect 240701 455477 240711 455543
rect 240821 455477 240831 455543
rect 251423 455455 251433 455521
rect 251543 455455 251553 455521
rect 502200 455237 502310 455247
rect 502190 455171 502200 455237
rect 502310 455171 502320 455237
rect 502200 455161 502310 455171
rect 502210 454865 502320 454875
rect 502200 454799 502210 454865
rect 502320 454799 502330 454865
rect 502210 454789 502320 454799
rect 564536 453405 564602 453415
rect 564164 453395 564230 453405
rect 564154 453285 564164 453395
rect 564230 453285 564240 453395
rect 564526 453295 564536 453405
rect 564602 453295 564612 453405
rect 564536 453285 564602 453295
rect 564164 453275 564230 453285
rect 508964 449038 509074 449048
rect 508954 448972 508964 449038
rect 509074 448972 509084 449038
rect 508964 448962 509074 448972
rect 392786 448771 392796 448837
rect 392906 448771 392916 448837
rect 387865 448703 387875 448769
rect 387985 448703 387995 448769
rect 508974 448666 509084 448676
rect 508964 448600 508974 448666
rect 509084 448600 509094 448666
rect 508974 448590 509084 448600
rect 392796 448399 392806 448465
rect 392916 448399 392926 448465
rect 387875 448331 387885 448397
rect 387995 448331 388005 448397
rect 515060 447630 515170 447640
rect 515050 447564 515060 447630
rect 515170 447564 515180 447630
rect 515060 447554 515170 447564
rect 515070 447258 515180 447268
rect 515060 447192 515070 447258
rect 515180 447192 515190 447258
rect 515070 447182 515180 447192
rect 534376 446611 534486 446621
rect 534366 446545 534376 446611
rect 534486 446545 534496 446611
rect 534376 446535 534486 446545
rect 534366 446239 534476 446249
rect 534356 446173 534366 446239
rect 534476 446173 534486 446239
rect 534366 446163 534476 446173
rect 355990 442179 356000 442245
rect 356110 442179 356120 442245
rect 356000 441807 356010 441873
rect 356120 441807 356130 441873
rect 346958 436390 346968 436456
rect 347078 436390 347088 436456
rect 346968 436018 346978 436084
rect 347088 436018 347098 436084
rect 240611 434332 240621 434398
rect 240731 434332 240741 434398
rect 251396 434046 251406 434112
rect 251516 434046 251526 434112
rect 240621 433960 240631 434026
rect 240741 433960 240751 434026
rect 251406 433674 251416 433740
rect 251526 433674 251536 433740
rect 348094 430698 348522 430708
rect 249235 430379 249777 430385
rect 238866 430259 239407 430265
rect 238857 429718 238866 430259
rect 239407 429718 239416 430259
rect 249226 429837 249235 430379
rect 249777 429837 249786 430379
rect 252980 430363 253522 430372
rect 332869 430371 333411 430380
rect 249235 429831 249777 429837
rect 252974 429821 252980 430363
rect 253522 429821 253528 430363
rect 258338 430362 258878 430368
rect 258329 429822 258338 430362
rect 258878 429822 258887 430362
rect 293214 430355 293756 430361
rect 278450 430343 278992 430349
rect 272940 430299 273482 430308
rect 252980 429812 253522 429821
rect 258338 429816 258878 429822
rect 272934 429757 272940 430299
rect 273482 429757 273488 430299
rect 278441 429801 278450 430343
rect 278992 429801 279001 430343
rect 293205 429813 293214 430355
rect 293756 429813 293765 430355
rect 299162 430255 299704 430261
rect 293214 429807 293756 429813
rect 278450 429795 278992 429801
rect 272940 429748 273482 429757
rect 238866 429712 239407 429718
rect 299153 429713 299162 430255
rect 299704 429713 299713 430255
rect 322085 430215 322627 430221
rect 313348 430191 313890 430200
rect 299162 429707 299704 429713
rect 313342 429649 313348 430191
rect 313890 429649 313896 430191
rect 319476 430157 320018 430163
rect 313348 429640 313890 429649
rect 319467 429615 319476 430157
rect 320018 429615 320027 430157
rect 322076 429673 322085 430215
rect 322627 429673 322636 430215
rect 335394 430253 335936 430259
rect 322085 429667 322627 429673
rect 319476 429609 320018 429615
rect 293185 426186 293251 426196
rect 272904 426152 272970 426162
rect 252958 426087 253024 426097
rect 252958 425967 253024 425977
rect 253330 426077 253396 426087
rect 272904 426032 272970 426042
rect 273276 426142 273342 426152
rect 293185 426066 293251 426076
rect 293557 426176 293623 426186
rect 293557 426056 293623 426066
rect 313334 426176 313400 426186
rect 313334 426056 313400 426066
rect 313706 426166 313772 426176
rect 313706 426046 313772 426056
rect 273276 426022 273342 426032
rect 253330 425957 253396 425967
rect 332869 420847 333411 429829
rect 335385 429711 335394 430253
rect 335936 429711 335945 430253
rect 335394 429705 335936 429711
rect 360001 430439 360543 430448
rect 362171 430443 362713 430452
rect 354357 430269 354899 430278
rect 354351 429727 354357 430269
rect 354899 429727 354905 430269
rect 359995 429897 360001 430439
rect 360543 429897 360549 430439
rect 362165 429901 362171 430443
rect 362713 429901 362719 430443
rect 497210 430398 497838 430407
rect 545783 430403 546413 430409
rect 391205 430371 391747 430377
rect 385933 430287 386475 430293
rect 373950 430191 374492 430197
rect 375352 430195 375894 430204
rect 360001 429888 360543 429897
rect 362171 429892 362713 429901
rect 354357 429718 354899 429727
rect 373941 429649 373950 430191
rect 374492 429649 374501 430191
rect 375346 429653 375352 430195
rect 375894 429653 375900 430195
rect 385924 429745 385933 430287
rect 386475 429745 386484 430287
rect 391196 429829 391205 430371
rect 391747 429829 391756 430371
rect 391205 429823 391747 429829
rect 497204 429770 497210 430398
rect 497838 429770 497844 430398
rect 513067 430335 513669 430344
rect 510283 430285 510885 430294
rect 497210 429761 497838 429770
rect 385933 429739 386475 429745
rect 510277 429683 510283 430285
rect 510885 429683 510891 430285
rect 513061 429733 513067 430335
rect 513669 429733 513675 430335
rect 528959 430329 529589 430335
rect 522311 430301 522913 430307
rect 513067 429724 513669 429733
rect 522302 429699 522311 430301
rect 522913 429699 522922 430301
rect 528950 429699 528959 430329
rect 529589 429699 529598 430329
rect 545774 429773 545783 430403
rect 546413 429773 546422 430403
rect 562801 430329 563431 430338
rect 545783 429767 546413 429773
rect 562795 429699 562801 430329
rect 563431 429699 563437 430329
rect 522311 429693 522913 429699
rect 528959 429693 529589 429699
rect 562801 429690 563431 429699
rect 510283 429674 510885 429683
rect 373950 429643 374492 429649
rect 375352 429644 375894 429653
rect 348094 429372 348522 429382
rect 387894 427660 387904 427726
rect 388014 427660 388024 427726
rect 392818 427679 392828 427745
rect 392938 427679 392948 427745
rect 387904 427288 387914 427354
rect 388024 427288 388034 427354
rect 392828 427307 392838 427373
rect 392948 427307 392958 427373
rect 375866 426251 375932 426261
rect 375494 426241 375560 426251
rect 335913 426161 335979 426171
rect 335541 426151 335607 426161
rect 355903 426157 355969 426167
rect 335913 426041 335979 426051
rect 355531 426147 355597 426157
rect 335541 426031 335607 426041
rect 375866 426131 375932 426141
rect 375494 426121 375560 426131
rect 355903 426037 355969 426047
rect 355531 426027 355597 426037
rect 355995 422225 356005 422291
rect 356115 422225 356125 422291
rect 356005 421853 356015 421919
rect 356125 421853 356135 421919
rect 278446 420622 278512 420632
rect 299123 420628 299189 420638
rect 258312 420589 258378 420599
rect 258312 420469 258378 420479
rect 258684 420579 258750 420589
rect 278446 420502 278512 420512
rect 278818 420612 278884 420622
rect 299123 420508 299189 420518
rect 299495 420618 299561 420628
rect 278818 420492 278884 420502
rect 299495 420498 299561 420508
rect 319451 420580 319517 420590
rect 258684 420459 258750 420469
rect 319451 420460 319517 420470
rect 319823 420570 319889 420580
rect 319823 420450 319889 420460
rect 332863 420305 332869 420847
rect 333411 420305 333417 420847
rect 374476 420659 374542 420669
rect 374104 420649 374170 420659
rect 354133 420589 354199 420599
rect 353761 420579 353827 420589
rect 374476 420539 374542 420549
rect 374104 420529 374170 420539
rect 354133 420469 354199 420479
rect 353761 420459 353827 420469
rect 324544 417178 324654 417188
rect 324534 417112 324544 417178
rect 324654 417112 324664 417178
rect 324544 417102 324654 417112
rect 336554 417103 336664 417113
rect 336544 417037 336554 417103
rect 336664 417037 336674 417103
rect 336554 417027 336664 417037
rect 324544 416740 324554 416806
rect 324664 416740 324674 416806
rect 336554 416665 336564 416731
rect 336674 416665 336684 416731
rect 345550 416210 345978 416220
rect 319466 415947 320008 415953
rect 252972 415912 253512 415918
rect 242019 415901 242560 415910
rect 242013 415360 242019 415901
rect 242560 415360 242566 415901
rect 252963 415372 252972 415912
rect 253512 415372 253521 415912
rect 258336 415876 258876 415885
rect 255273 415727 255815 415736
rect 252972 415366 253512 415372
rect 242019 415351 242560 415360
rect 255267 415185 255273 415727
rect 255815 415185 255821 415727
rect 258330 415336 258336 415876
rect 258876 415336 258882 415876
rect 313354 415871 313896 415877
rect 272932 415809 273474 415818
rect 278450 415815 278992 415824
rect 258336 415327 258876 415336
rect 272926 415267 272932 415809
rect 273474 415267 273480 415809
rect 278444 415273 278450 415815
rect 278992 415273 278998 415815
rect 299136 415813 299678 415822
rect 293214 415789 293756 415795
rect 272932 415258 273474 415267
rect 278450 415264 278992 415273
rect 293205 415247 293214 415789
rect 293756 415247 293765 415789
rect 299130 415271 299136 415813
rect 299678 415271 299684 415813
rect 313345 415329 313354 415871
rect 313896 415329 313905 415871
rect 319457 415405 319466 415947
rect 320008 415405 320017 415947
rect 328159 415901 328701 415907
rect 319466 415399 320008 415405
rect 328150 415359 328159 415901
rect 328701 415359 328710 415901
rect 339875 415863 340417 415869
rect 328159 415353 328701 415359
rect 313354 415323 313896 415329
rect 339866 415321 339875 415863
rect 340417 415321 340426 415863
rect 339875 415315 340417 415321
rect 299136 415262 299678 415271
rect 293214 415241 293756 415247
rect 255273 415176 255815 415185
rect 393665 415927 394207 415936
rect 373944 415845 374486 415851
rect 388617 415849 389159 415855
rect 346902 415756 346912 415822
rect 347022 415756 347032 415822
rect 353573 415775 354115 415784
rect 346912 415384 346922 415450
rect 347032 415384 347042 415450
rect 353567 415233 353573 415775
rect 354115 415233 354121 415775
rect 373935 415303 373944 415845
rect 374486 415303 374495 415845
rect 375340 415649 375882 415655
rect 373944 415297 374486 415303
rect 353573 415224 354115 415233
rect 375331 415107 375340 415649
rect 375882 415107 375891 415649
rect 388608 415307 388617 415849
rect 389159 415307 389168 415849
rect 393659 415385 393665 415927
rect 394207 415385 394213 415927
rect 393665 415376 394207 415385
rect 388617 415301 389159 415307
rect 375340 415101 375882 415107
rect 345550 414884 345978 414894
rect 568046 408988 568112 408998
rect 568036 408878 568046 408988
rect 568112 408878 568122 408988
rect 568418 408978 568484 408988
rect 568046 408868 568112 408878
rect 568418 408858 568484 408868
rect 549543 407130 549553 407196
rect 549663 407130 549673 407196
rect 549543 406824 549653 406834
rect 549533 406758 549543 406824
rect 549653 406758 549663 406824
rect 549543 406748 549653 406758
rect 355984 402190 355994 402256
rect 356104 402190 356114 402256
rect 355994 401818 356004 401884
rect 356114 401818 356124 401884
rect 336579 396450 336689 396460
rect 324542 396388 324652 396398
rect 324532 396322 324542 396388
rect 324652 396322 324662 396388
rect 336569 396384 336579 396450
rect 336689 396384 336699 396450
rect 336579 396374 336689 396384
rect 324542 396312 324652 396322
rect 324542 395950 324552 396016
rect 324662 395950 324672 396016
rect 336579 396012 336589 396078
rect 336699 396012 336709 396078
rect 346930 395078 346940 395144
rect 347050 395078 347060 395144
rect 346940 394706 346950 394772
rect 347060 394706 347070 394772
rect 333092 391367 333634 391373
rect 322895 391347 323437 391353
rect 322886 390805 322895 391347
rect 323437 390805 323446 391347
rect 333083 390825 333092 391367
rect 333634 390825 333643 391367
rect 334879 391309 335421 391315
rect 333092 390819 333634 390825
rect 322895 390799 323437 390805
rect 334870 390767 334879 391309
rect 335421 390767 335430 391309
rect 428501 391297 429043 391306
rect 367484 391193 368026 391199
rect 357690 391157 358232 391163
rect 353565 390939 354107 390948
rect 334879 390761 335421 390767
rect 353559 390397 353565 390939
rect 354107 390397 354113 390939
rect 357681 390615 357690 391157
rect 358232 390615 358241 391157
rect 367475 390651 367484 391193
rect 368026 390651 368035 391193
rect 400437 391189 400979 391195
rect 385269 391169 385811 391175
rect 367484 390645 368026 390651
rect 385260 390627 385269 391169
rect 385811 390627 385820 391169
rect 400428 390647 400437 391189
rect 400979 390647 400988 391189
rect 428495 390755 428501 391297
rect 429043 390755 429049 391297
rect 546403 391241 546965 391247
rect 530385 391147 530927 391153
rect 490269 391105 490811 391111
rect 470027 391055 470569 391061
rect 446395 391049 446937 391055
rect 428501 390746 429043 390755
rect 400437 390641 400979 390647
rect 385269 390621 385811 390627
rect 357690 390609 358232 390615
rect 446386 390507 446395 391049
rect 446937 390507 446946 391049
rect 470018 390513 470027 391055
rect 470569 390513 470578 391055
rect 490260 390563 490269 391105
rect 490811 390563 490820 391105
rect 510723 391075 511265 391081
rect 490269 390557 490811 390563
rect 510714 390533 510723 391075
rect 511265 390533 511274 391075
rect 530376 390605 530385 391147
rect 530927 390605 530936 391147
rect 546394 390679 546403 391241
rect 546965 390679 546974 391241
rect 571227 391205 571789 391211
rect 546403 390673 546965 390679
rect 571218 390643 571227 391205
rect 571789 390643 571798 391205
rect 571227 390637 571789 390643
rect 530385 390599 530927 390605
rect 510723 390527 511265 390533
rect 470027 390507 470569 390513
rect 446395 390501 446937 390507
rect 353565 390388 354107 390397
rect 549560 388086 549570 388152
rect 549680 388086 549690 388152
rect 549560 387780 549670 387790
rect 549550 387714 549560 387780
rect 549670 387714 549680 387780
rect 549560 387704 549670 387714
rect 427809 386796 427875 386806
rect 367462 386753 367528 386763
rect 347446 386724 347512 386734
rect 347436 386614 347446 386724
rect 347512 386614 347522 386724
rect 347818 386714 347884 386724
rect 347446 386604 347512 386614
rect 367452 386643 367462 386753
rect 367528 386643 367538 386753
rect 367834 386743 367900 386753
rect 387274 386743 387340 386753
rect 367462 386633 367528 386643
rect 387264 386633 387274 386743
rect 387340 386633 387350 386743
rect 387646 386733 387712 386743
rect 407533 386741 407599 386751
rect 367834 386623 367900 386633
rect 387274 386623 387340 386633
rect 407523 386631 407533 386741
rect 407599 386631 407609 386741
rect 407905 386731 407971 386741
rect 387646 386613 387712 386623
rect 407533 386621 407599 386631
rect 427799 386686 427809 386796
rect 427875 386686 427885 386796
rect 428181 386786 428247 386796
rect 528327 386792 528393 386802
rect 427809 386676 427875 386686
rect 447968 386776 448034 386786
rect 428181 386666 428247 386676
rect 447958 386666 447968 386776
rect 448034 386666 448044 386776
rect 448340 386766 448406 386776
rect 467970 386771 468036 386781
rect 508218 386778 508284 386788
rect 447968 386656 448034 386666
rect 467960 386661 467970 386771
rect 468036 386661 468046 386771
rect 468342 386761 468408 386771
rect 448340 386646 448406 386656
rect 467970 386651 468036 386661
rect 488088 386755 488154 386765
rect 468342 386641 468408 386651
rect 488078 386645 488088 386755
rect 488154 386645 488164 386755
rect 488460 386745 488526 386755
rect 488088 386635 488154 386645
rect 508208 386668 508218 386778
rect 508284 386668 508294 386778
rect 508590 386768 508656 386778
rect 508218 386658 508284 386668
rect 528317 386682 528327 386792
rect 528393 386682 528403 386792
rect 528699 386782 528765 386792
rect 528327 386672 528393 386682
rect 528699 386662 528765 386672
rect 508590 386648 508656 386658
rect 488460 386625 488526 386635
rect 407905 386611 407971 386621
rect 347818 386594 347884 386604
rect 355964 382126 355974 382192
rect 356084 382126 356094 382192
rect 355974 381754 355984 381820
rect 356094 381754 356104 381820
rect 467885 380800 467951 380810
rect 333077 380757 333143 380767
rect 357656 380765 357722 380775
rect 333067 380647 333077 380757
rect 333143 380647 333153 380757
rect 333449 380747 333515 380757
rect 333077 380637 333143 380647
rect 357646 380655 357656 380765
rect 357722 380655 357732 380765
rect 358028 380755 358094 380765
rect 357656 380645 357722 380655
rect 407681 380754 407747 380764
rect 387103 380723 387169 380733
rect 333449 380627 333515 380637
rect 358028 380635 358094 380645
rect 387093 380613 387103 380723
rect 387169 380613 387179 380723
rect 387475 380713 387541 380723
rect 387103 380603 387169 380613
rect 407671 380644 407681 380754
rect 407747 380644 407757 380754
rect 408053 380744 408119 380754
rect 407681 380634 407747 380644
rect 427655 380729 427721 380739
rect 447901 380733 447967 380743
rect 408053 380624 408119 380634
rect 427645 380619 427655 380729
rect 427721 380619 427731 380729
rect 428027 380719 428093 380729
rect 427655 380609 427721 380619
rect 447891 380623 447901 380733
rect 447967 380623 447977 380733
rect 448273 380723 448339 380733
rect 447901 380613 447967 380623
rect 467875 380690 467885 380800
rect 467951 380690 467961 380800
rect 468257 380790 468323 380800
rect 507983 380797 508049 380807
rect 467885 380680 467951 380690
rect 488300 380725 488366 380735
rect 468257 380670 468323 380680
rect 488290 380615 488300 380725
rect 488366 380615 488376 380725
rect 488672 380715 488738 380725
rect 387475 380593 387541 380603
rect 428027 380599 428093 380609
rect 448273 380603 448339 380613
rect 488300 380605 488366 380615
rect 507973 380687 507983 380797
rect 508049 380687 508059 380797
rect 508355 380787 508421 380797
rect 507983 380677 508049 380687
rect 528353 380731 528419 380741
rect 508355 380667 508421 380677
rect 528343 380621 528353 380731
rect 528419 380621 528429 380731
rect 528725 380721 528791 380731
rect 528353 380611 528419 380621
rect 488672 380595 488738 380605
rect 528725 380601 528791 380611
rect 549368 379494 549478 379504
rect 549358 379428 549368 379494
rect 549478 379428 549488 379494
rect 549368 379418 549478 379428
rect 549378 379122 549488 379132
rect 549368 379056 549378 379122
rect 549488 379056 549498 379122
rect 549378 379046 549488 379056
rect 352330 376280 353838 376290
rect 333090 376209 333632 376218
rect 325765 376095 326307 376101
rect 325756 375553 325765 376095
rect 326307 375553 326316 376095
rect 333084 375667 333090 376209
rect 333632 375667 333638 376209
rect 337333 376115 337875 376124
rect 333090 375658 333632 375667
rect 337327 375573 337333 376115
rect 337875 375573 337881 376115
rect 345681 376089 346223 376098
rect 337333 375564 337875 375573
rect 325765 375547 326307 375553
rect 345675 375547 345681 376089
rect 346223 375547 346229 376089
rect 526305 376169 526847 376175
rect 357684 376101 358226 376107
rect 400425 376101 400967 376107
rect 352330 375598 353838 375608
rect 357675 375559 357684 376101
rect 358226 375559 358235 376101
rect 367484 376051 368026 376057
rect 357684 375553 358226 375559
rect 345681 375538 346223 375547
rect 367475 375509 367484 376051
rect 368026 375509 368035 376051
rect 388559 375919 389101 375925
rect 367484 375503 368026 375509
rect 388550 375377 388559 375919
rect 389101 375377 389110 375919
rect 400416 375559 400425 376101
rect 400967 375559 400976 376101
rect 446411 376065 446953 376071
rect 429149 376007 429691 376013
rect 400425 375553 400967 375559
rect 429140 375465 429149 376007
rect 429691 375465 429700 376007
rect 446402 375523 446411 376065
rect 446953 375523 446962 376065
rect 466549 376049 467091 376055
rect 446411 375517 446953 375523
rect 466540 375507 466549 376049
rect 467091 375507 467100 376049
rect 485509 376005 486051 376011
rect 466549 375501 467091 375507
rect 429149 375459 429691 375465
rect 485500 375463 485509 376005
rect 486051 375463 486060 376005
rect 505733 375989 506275 375995
rect 485509 375457 486051 375463
rect 505724 375447 505733 375989
rect 506275 375447 506284 375989
rect 526296 375627 526305 376169
rect 526847 375627 526856 376169
rect 562709 376121 563271 376130
rect 552361 376047 552923 376053
rect 526305 375621 526847 375627
rect 552352 375485 552361 376047
rect 552923 375485 552932 376047
rect 562703 375559 562709 376121
rect 563271 375559 563277 376121
rect 562709 375550 563271 375559
rect 552361 375479 552923 375485
rect 505733 375441 506275 375447
rect 388559 375371 389101 375377
rect 346916 373796 346926 373862
rect 347036 373796 347046 373862
rect 346926 373424 346936 373490
rect 347046 373424 347056 373490
rect 549329 364308 549439 364318
rect 549319 364242 549329 364308
rect 549439 364242 549449 364308
rect 549329 364232 549439 364242
rect 549339 363936 549449 363946
rect 549329 363870 549339 363936
rect 549449 363870 549459 363936
rect 549339 363860 549449 363870
rect 568202 362605 568268 362615
rect 568192 362495 568202 362605
rect 568268 362495 568278 362605
rect 568574 362595 568640 362605
rect 568202 362485 568268 362495
rect 568574 362475 568640 362485
rect 356021 362143 356031 362209
rect 356141 362143 356151 362209
rect 356031 361771 356041 361837
rect 356151 361771 356161 361837
rect 346916 352946 346926 353012
rect 347036 352946 347046 353012
rect 346926 352574 346936 352640
rect 347046 352574 347056 352640
rect 356021 342140 356031 342206
rect 356141 342140 356151 342206
rect 356031 341768 356041 341834
rect 356151 341768 356161 341834
rect 347000 332350 347010 332416
rect 347120 332350 347130 332416
rect 347010 331978 347020 332044
rect 347130 331978 347140 332044
rect 355945 322138 355955 322204
rect 356065 322138 356075 322204
rect 355955 321766 355965 321832
rect 356075 321766 356085 321832
rect 346972 310482 346982 310548
rect 347092 310482 347102 310548
rect 346982 310110 346992 310176
rect 347102 310110 347112 310176
rect 348024 307618 348476 307628
rect 490714 307004 491263 307010
rect 390700 306940 391249 306949
rect 370688 306812 371237 306821
rect 357945 306779 358487 306788
rect 357939 306237 357945 306779
rect 358487 306237 358493 306779
rect 370682 306263 370688 306812
rect 371237 306263 371243 306812
rect 390694 306391 390700 306940
rect 391249 306391 391255 306940
rect 400264 306898 400813 306907
rect 390700 306382 391249 306391
rect 400258 306349 400264 306898
rect 400813 306349 400819 306898
rect 445440 306860 445989 306869
rect 430714 306662 431263 306671
rect 400264 306340 400813 306349
rect 370688 306254 371237 306263
rect 357945 306228 358487 306237
rect 430708 306113 430714 306662
rect 431263 306113 431269 306662
rect 445434 306311 445440 306860
rect 445989 306311 445995 306860
rect 470718 306780 471267 306786
rect 445440 306302 445989 306311
rect 470709 306231 470718 306780
rect 471267 306231 471276 306780
rect 490705 306455 490714 307004
rect 491263 306455 491272 307004
rect 510700 306896 511249 306902
rect 490714 306449 491263 306455
rect 510691 306347 510700 306896
rect 511249 306347 511258 306896
rect 569358 306806 569927 306815
rect 530686 306742 531235 306748
rect 510700 306341 511249 306347
rect 470718 306225 471267 306231
rect 530677 306193 530686 306742
rect 531235 306193 531244 306742
rect 552167 306730 552724 306736
rect 530686 306187 531235 306193
rect 552158 306173 552167 306730
rect 552724 306173 552733 306730
rect 569352 306237 569358 306806
rect 569927 306237 569933 306806
rect 569358 306228 569927 306237
rect 552167 306167 552724 306173
rect 430714 306104 431263 306113
rect 348024 305634 348476 305644
rect 355983 302117 355993 302183
rect 356103 302117 356113 302183
rect 355993 301745 356003 301811
rect 356113 301745 356123 301811
rect 491225 296133 491291 296143
rect 531203 296133 531269 296143
rect 490853 296123 490919 296133
rect 431211 296108 431277 296118
rect 430839 296098 430905 296108
rect 391209 296061 391275 296071
rect 371200 296044 371266 296054
rect 370828 296034 370894 296044
rect 371200 295924 371266 295934
rect 390837 296051 390903 296061
rect 411215 296032 411281 296042
rect 391209 295941 391275 295951
rect 410843 296022 410909 296032
rect 390837 295931 390903 295941
rect 370828 295914 370894 295924
rect 471230 296100 471296 296110
rect 470858 296090 470924 296100
rect 451228 296075 451294 296085
rect 431211 295988 431277 295998
rect 450856 296065 450922 296075
rect 430839 295978 430905 295988
rect 530831 296123 530897 296133
rect 511218 296089 511284 296099
rect 491225 296013 491291 296023
rect 510846 296079 510912 296089
rect 490853 296003 490919 296013
rect 471230 295980 471296 295990
rect 470858 295970 470924 295980
rect 451228 295955 451294 295965
rect 531203 296013 531269 296023
rect 530831 296003 530897 296013
rect 511218 295969 511284 295979
rect 510846 295959 510912 295969
rect 450856 295945 450922 295955
rect 411215 295912 411281 295922
rect 410843 295902 410909 295912
rect 549547 293441 549657 293451
rect 549537 293375 549547 293441
rect 549657 293375 549667 293441
rect 549547 293365 549657 293375
rect 549557 293069 549667 293079
rect 549547 293003 549557 293069
rect 549667 293003 549677 293069
rect 549557 292993 549667 293003
rect 346930 288824 346940 288890
rect 347050 288824 347060 288890
rect 346940 288452 346950 288518
rect 347060 288452 347070 288518
rect 345710 287588 346162 287598
rect 445452 287021 446001 287030
rect 400180 286903 400729 286912
rect 354041 286813 354583 286819
rect 354032 286271 354041 286813
rect 354583 286271 354592 286813
rect 390700 286691 391249 286700
rect 370688 286607 371237 286613
rect 354041 286265 354583 286271
rect 370679 286058 370688 286607
rect 371237 286058 371246 286607
rect 390694 286142 390700 286691
rect 391249 286142 391255 286691
rect 400174 286354 400180 286903
rect 400729 286354 400735 286903
rect 430714 286809 431263 286818
rect 400180 286345 400729 286354
rect 430708 286260 430714 286809
rect 431263 286260 431269 286809
rect 445446 286472 445452 287021
rect 446001 286472 446007 287021
rect 546320 286983 546877 286989
rect 490714 286883 491263 286889
rect 470718 286753 471267 286759
rect 445452 286463 446001 286472
rect 430714 286251 431263 286260
rect 470709 286204 470718 286753
rect 471267 286204 471276 286753
rect 490705 286334 490714 286883
rect 491263 286334 491272 286883
rect 510700 286819 511249 286825
rect 490714 286328 491263 286334
rect 510691 286270 510700 286819
rect 511249 286270 511258 286819
rect 530686 286807 531235 286813
rect 510700 286264 511249 286270
rect 530677 286258 530686 286807
rect 531235 286258 531244 286807
rect 546311 286426 546320 286983
rect 546877 286426 546886 286983
rect 568318 286882 568887 286891
rect 546320 286420 546877 286426
rect 568312 286313 568318 286882
rect 568887 286313 568893 286882
rect 568318 286304 568887 286313
rect 530686 286252 531235 286258
rect 470718 286198 471267 286204
rect 390700 286133 391249 286142
rect 370688 286052 371237 286058
rect 345710 285604 346162 285614
rect 551821 274026 551887 274036
rect 551449 274016 551515 274026
rect 572284 273986 572350 273996
rect 551821 273906 551887 273916
rect 571912 273976 571978 273986
rect 551449 273896 551515 273906
rect 572284 273866 572350 273876
rect 571912 273856 571978 273866
rect 346888 264044 346898 264110
rect 347008 264044 347018 264110
rect 346898 263672 346908 263738
rect 347018 263672 347028 263738
rect 346972 242670 346982 242736
rect 347092 242670 347102 242736
rect 346982 242298 346992 242364
rect 347102 242298 347112 242364
rect 347000 222794 347010 222860
rect 347120 222794 347130 222860
rect 347010 222422 347020 222488
rect 347130 222422 347140 222488
rect 347982 213096 348448 213106
rect 347982 208078 348448 208088
rect 346944 200966 346954 201032
rect 347064 200966 347074 201032
rect 346954 200594 346964 200660
rect 347074 200594 347084 200660
rect 346958 179932 346968 179998
rect 347078 179932 347088 179998
rect 346968 179560 346978 179626
rect 347088 179560 347098 179626
rect 345722 177826 346188 177836
rect 345722 172808 346188 172818
rect 345698 167836 346164 167846
rect 345698 162818 346164 162828
rect 346916 158544 346926 158610
rect 347036 158544 347046 158610
rect 346926 158172 346936 158238
rect 347046 158172 347056 158238
rect 334827 137385 335369 137391
rect 334818 136843 334827 137385
rect 335369 136843 335378 137385
rect 358795 137369 359337 137375
rect 346860 137198 346870 137264
rect 346980 137198 346990 137264
rect 334827 136837 335369 136843
rect 346870 136826 346880 136892
rect 346990 136826 347000 136892
rect 358786 136827 358795 137369
rect 359337 136827 359346 137369
rect 358795 136821 359337 136827
rect 346916 116064 346926 116130
rect 347036 116064 347046 116130
rect 346926 115692 346936 115758
rect 347046 115692 347056 115758
rect 334799 95639 335341 95645
rect 359143 95639 359685 95645
rect 334790 95097 334799 95639
rect 335341 95097 335350 95639
rect 346944 95454 346954 95520
rect 347064 95454 347074 95520
rect 334799 95091 335341 95097
rect 346954 95082 346964 95148
rect 347074 95082 347084 95148
rect 359134 95097 359143 95639
rect 359685 95097 359694 95639
rect 359143 95091 359685 95097
rect 346930 74772 346940 74838
rect 347050 74772 347060 74838
rect 346940 74400 346950 74466
rect 347060 74400 347070 74466
rect 90284 60006 91538 60016
rect 302579 59503 303121 59509
rect 324127 59503 324669 59509
rect 240075 59381 240617 59390
rect 133049 59371 133591 59380
rect 111727 59361 112269 59370
rect 111721 58819 111727 59361
rect 112269 58819 112275 59361
rect 133043 58829 133049 59371
rect 133591 58829 133597 59371
rect 154607 59327 155149 59336
rect 175813 59327 176355 59336
rect 133049 58820 133591 58829
rect 111727 58810 112269 58819
rect 154601 58785 154607 59327
rect 155149 58785 155155 59327
rect 175807 58785 175813 59327
rect 176355 58785 176361 59327
rect 219089 59305 219631 59314
rect 197195 59283 197737 59292
rect 154607 58776 155149 58785
rect 175813 58776 176355 58785
rect 90284 58742 91538 58752
rect 197189 58741 197195 59283
rect 197737 58741 197743 59283
rect 219083 58763 219089 59305
rect 219631 58763 219637 59305
rect 240069 58839 240075 59381
rect 240617 58839 240623 59381
rect 260577 59379 261119 59385
rect 240075 58830 240617 58839
rect 260568 58837 260577 59379
rect 261119 58837 261128 59379
rect 281389 59135 281931 59141
rect 260577 58831 261119 58837
rect 219089 58754 219631 58763
rect 197195 58732 197737 58741
rect 281380 58593 281389 59135
rect 281931 58593 281940 59135
rect 302570 58961 302579 59503
rect 303121 58961 303130 59503
rect 324118 58961 324127 59503
rect 324669 58961 324678 59503
rect 302579 58955 303121 58961
rect 324127 58955 324669 58961
rect 281389 58587 281931 58593
rect 334723 54525 335265 54534
rect 358805 54525 359347 54531
rect 334717 53983 334723 54525
rect 335265 53983 335271 54525
rect 358796 53983 358805 54525
rect 359347 53983 359356 54525
rect 334723 53974 335265 53983
rect 358805 53977 359347 53983
rect 39905 52861 40867 52870
rect 39899 51899 39905 52861
rect 40867 51899 40873 52861
rect 39905 51890 40867 51899
rect 347000 51192 347010 51258
rect 347120 51192 347130 51258
rect 347010 50820 347020 50886
rect 347130 50820 347140 50886
rect 281744 49014 281810 49024
rect 281372 49004 281438 49014
rect 133404 48970 133470 48980
rect 197550 48970 197616 48980
rect 69656 48956 69722 48966
rect 69284 48946 69350 48956
rect 48362 48896 48428 48906
rect 47990 48886 48056 48896
rect 133032 48960 133098 48970
rect 112082 48926 112148 48936
rect 111710 48916 111776 48926
rect 91022 48882 91088 48892
rect 69656 48836 69722 48846
rect 90650 48872 90716 48882
rect 69284 48826 69350 48836
rect 48362 48776 48428 48786
rect 47990 48766 48056 48776
rect 197178 48960 197244 48970
rect 154962 48940 155028 48950
rect 133404 48850 133470 48860
rect 154590 48930 154656 48940
rect 133032 48840 133098 48850
rect 112082 48806 112148 48816
rect 176168 48912 176234 48922
rect 154962 48820 155028 48830
rect 175796 48902 175862 48912
rect 154590 48810 154656 48820
rect 111710 48796 111776 48806
rect 260932 48912 260998 48922
rect 260560 48902 260626 48912
rect 219444 48882 219510 48892
rect 197550 48850 197616 48860
rect 219072 48872 219138 48882
rect 197178 48840 197244 48850
rect 176168 48792 176234 48802
rect 175796 48782 175862 48792
rect 91022 48762 91088 48772
rect 240430 48852 240496 48862
rect 219444 48762 219510 48772
rect 240058 48842 240124 48852
rect 90650 48752 90716 48762
rect 219072 48752 219138 48762
rect 281744 48894 281810 48904
rect 281372 48884 281438 48894
rect 324482 48844 324548 48854
rect 324110 48834 324176 48844
rect 302934 48808 303000 48818
rect 260932 48792 260998 48802
rect 302562 48798 302628 48808
rect 260560 48782 260626 48792
rect 240430 48732 240496 48742
rect 240058 48722 240124 48732
rect 324482 48724 324548 48734
rect 324110 48714 324176 48724
rect 302934 48688 303000 48698
rect 302562 48678 302628 48688
rect 34568 42938 34578 43004
rect 34688 42938 34698 43004
rect 34578 42566 34588 42632
rect 34698 42566 34708 42632
rect 39650 39258 42762 39268
rect 69303 38013 69845 38022
rect 48009 37907 48551 37916
rect 48003 37365 48009 37907
rect 48551 37365 48557 37907
rect 69297 37471 69303 38013
rect 69845 37471 69851 38013
rect 197197 37933 197739 37942
rect 154609 37835 155151 37844
rect 175815 37835 176357 37844
rect 111729 37747 112271 37756
rect 90669 37695 91211 37704
rect 69303 37462 69845 37471
rect 48009 37356 48551 37365
rect 90663 37153 90669 37695
rect 91211 37153 91217 37695
rect 111723 37205 111729 37747
rect 112271 37205 112277 37747
rect 133051 37667 133593 37673
rect 111729 37196 112271 37205
rect 90669 37144 91211 37153
rect 133042 37125 133051 37667
rect 133593 37125 133602 37667
rect 154603 37293 154609 37835
rect 155151 37293 155157 37835
rect 175809 37293 175815 37835
rect 176357 37293 176363 37835
rect 197191 37391 197197 37933
rect 197739 37391 197745 37933
rect 302581 37919 303123 37925
rect 219091 37883 219633 37892
rect 197197 37382 197739 37391
rect 219085 37341 219091 37883
rect 219633 37341 219639 37883
rect 281391 37815 281933 37821
rect 240077 37781 240619 37787
rect 219091 37332 219633 37341
rect 154609 37284 155151 37293
rect 175815 37284 176357 37293
rect 240068 37239 240077 37781
rect 240619 37239 240628 37781
rect 260579 37719 261121 37725
rect 240077 37233 240619 37239
rect 260570 37177 260579 37719
rect 261121 37177 261130 37719
rect 281382 37273 281391 37815
rect 281933 37273 281942 37815
rect 302572 37377 302581 37919
rect 303123 37377 303132 37919
rect 324129 37867 324671 37873
rect 302581 37371 303123 37377
rect 324120 37325 324129 37867
rect 324671 37325 324680 37867
rect 324129 37319 324671 37325
rect 281391 37267 281933 37273
rect 260579 37171 261121 37177
rect 133051 37119 133593 37125
rect 39650 36260 42762 36270
rect 34568 20840 34578 20906
rect 34688 20840 34698 20906
rect 34578 20468 34588 20534
rect 34698 20468 34708 20534
rect 338567 8478 338576 8590
rect 338688 8478 338697 8590
rect 28112 3632 28178 3642
rect 27740 3622 27806 3632
rect 6920 3572 6986 3582
rect 6548 3562 6614 3572
rect 28112 3512 28178 3522
rect 27740 3502 27806 3512
rect 6920 3452 6986 3462
rect 6548 3442 6614 3452
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 494
rect 337394 -800 337506 480
rect 338576 -800 338688 8478
rect 356297 8088 356306 8200
rect 356418 8088 356427 8200
rect 342113 7742 342122 7854
rect 342234 7742 342243 7854
rect 339758 -800 339870 494
rect 340940 -800 341052 480
rect 342122 -800 342234 7742
rect 345659 7144 345668 7256
rect 345780 7144 345789 7256
rect 352751 7184 352760 7296
rect 352872 7184 352881 7296
rect 343304 -800 343416 494
rect 344486 -800 344598 480
rect 345668 -800 345780 7144
rect 349584 6628 349696 6637
rect 349214 6516 349584 6628
rect 346850 -800 346962 494
rect 348032 -800 348144 480
rect 349214 -800 349326 6516
rect 349584 6507 349696 6516
rect 350396 -800 350508 494
rect 351578 -800 351690 480
rect 352760 -800 352872 7184
rect 353942 -800 354054 494
rect 355124 -800 355236 480
rect 356306 -800 356418 8088
rect 476870 4020 476982 4029
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 3908
rect 480416 4020 480528 4029
rect 483953 3912 483962 4024
rect 484074 3912 484083 4024
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 3908
rect 481598 -800 481710 492
rect 482780 -800 482892 492
rect 483962 -800 484074 3912
rect 485144 -800 485256 492
rect 486326 -800 486438 492
rect 487508 -800 487620 480
rect 488690 -800 488802 492
rect 489872 -800 489984 492
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 550871 586751 550937 586861
rect 551243 586741 551309 586851
rect 571882 586782 571948 586892
rect 572254 586772 572320 586882
rect 537809 578721 538411 579323
rect 544736 573153 544846 573219
rect 544726 572781 544836 572847
rect 525320 567871 525386 567981
rect 525692 567861 525758 567971
rect 513762 562597 513872 562663
rect 513752 562225 513862 562291
rect 505449 560504 505559 560570
rect 505439 560132 505549 560198
rect 509408 554242 509938 556160
rect 526608 554236 527208 556182
rect 547182 554212 547758 556178
rect 531032 553043 531142 553109
rect 544746 552904 544856 552970
rect 531022 552671 531132 552737
rect 544736 552532 544846 552598
rect 522511 550426 522621 550492
rect 522501 550054 522611 550120
rect 513742 542155 513852 542221
rect 513732 541783 513842 541849
rect 505559 539916 505669 539982
rect 464237 538845 464839 539447
rect 484628 538955 485230 539557
rect 500443 539029 501045 539631
rect 505549 539544 505659 539610
rect 517874 538396 518574 540212
rect 537834 538328 538410 540294
rect 544751 532678 544861 532744
rect 544741 532306 544851 532372
rect 530987 531798 531097 531864
rect 530977 531426 531087 531492
rect 522560 529649 522670 529715
rect 522550 529277 522660 529343
rect 355991 522045 356101 522111
rect 356001 521673 356111 521739
rect 372209 516868 372269 516928
rect 513739 522184 513849 522250
rect 513729 521812 513839 521878
rect 537690 519333 537756 519443
rect 403609 519048 403669 519108
rect 424259 519078 424325 519188
rect 424631 519068 424697 519178
rect 444272 519137 444338 519247
rect 444644 519127 444710 519237
rect 464455 519220 464521 519330
rect 538062 519323 538128 519433
rect 464827 519210 464893 519320
rect 484787 519181 484853 519291
rect 485159 519171 485225 519281
rect 504261 519188 504327 519298
rect 504633 519178 504699 519288
rect 534334 508886 534444 508952
rect 534344 508514 534454 508580
rect 373647 504642 373707 504702
rect 383215 504697 383275 504757
rect 515038 507867 515148 507933
rect 515028 507495 515138 507561
rect 508942 506459 509052 506525
rect 508932 506087 509042 506153
rect 392783 504656 392843 504716
rect 355956 502136 356066 502202
rect 355966 501764 356076 501830
rect 502178 500260 502288 500326
rect 502168 499888 502278 499954
rect 521392 498333 521502 498399
rect 521382 497961 521492 498027
rect 527466 495935 527576 496001
rect 527456 495563 527566 495629
rect 564230 497760 564296 497870
rect 564602 497750 564668 497860
rect 550466 491990 550576 492056
rect 550456 491618 550566 491684
rect 387905 490687 388015 490753
rect 392808 490701 392918 490767
rect 373616 490608 373726 490674
rect 383268 490606 383378 490672
rect 387915 490315 388025 490381
rect 392818 490329 392928 490395
rect 373626 490236 373736 490302
rect 383278 490234 383388 490300
rect 534344 488486 534454 488552
rect 534354 488114 534464 488180
rect 515001 487666 515111 487732
rect 514991 487294 515101 487360
rect 508954 486408 509064 486474
rect 508944 486036 509054 486102
rect 360443 484605 360985 485147
rect 375489 484747 376031 485289
rect 386095 484671 386637 485213
rect 390329 484669 390871 485211
rect 400223 484639 400765 485181
rect 428641 484679 429183 485221
rect 434805 484627 435407 485229
rect 458519 484705 459121 485307
rect 464290 484555 464892 485157
rect 475009 484525 475611 485127
rect 484628 484593 485230 485195
rect 498503 484509 499105 485111
rect 504627 484563 505229 485165
rect 511844 484613 512446 485215
rect 518213 484585 518843 485215
rect 524290 484557 524892 485159
rect 530389 484571 530991 485173
rect 531891 484591 532521 485221
rect 545784 484497 546414 485127
rect 567849 484541 568479 485171
rect 356018 482192 356128 482258
rect 356028 481820 356138 481886
rect 384086 479600 384152 479710
rect 384458 479610 384524 479720
rect 399541 479625 399607 479735
rect 399913 479635 399979 479745
rect 419783 479565 419849 479675
rect 420155 479575 420221 479685
rect 440021 479594 440087 479704
rect 440393 479604 440459 479714
rect 460321 479606 460387 479716
rect 460693 479616 460759 479726
rect 480503 479584 480569 479694
rect 480875 479594 480941 479704
rect 522909 479633 522975 479743
rect 523281 479643 523347 479753
rect 500459 479506 500525 479616
rect 500831 479496 500897 479606
rect 545802 479510 545868 479620
rect 546174 479500 546240 479610
rect 346982 478252 347092 478318
rect 346992 477880 347102 477946
rect 379051 475499 379117 475609
rect 379423 475509 379489 475619
rect 399541 475532 399607 475642
rect 399913 475542 399979 475652
rect 419783 475472 419849 475582
rect 420155 475482 420221 475592
rect 440021 475501 440087 475611
rect 440393 475511 440459 475621
rect 460321 475513 460387 475623
rect 460693 475523 460759 475633
rect 480503 475491 480569 475601
rect 480875 475501 480941 475611
rect 500491 475509 500557 475619
rect 500863 475519 500929 475629
rect 522941 475382 523007 475492
rect 523313 475372 523379 475482
rect 545855 475418 545921 475528
rect 546227 475408 546293 475518
rect 352781 472439 353323 472981
rect 380557 472617 381099 473159
rect 389491 472541 390033 473083
rect 394697 472615 395239 473157
rect 400591 472567 401133 473109
rect 428295 472567 428837 473109
rect 445483 472445 446085 473047
rect 462135 472457 462737 473059
rect 485297 472501 485899 473103
rect 497352 472566 497980 473194
rect 503860 472370 504488 472998
rect 506695 472399 507297 473001
rect 518235 472485 518837 473087
rect 522944 472495 525127 473097
rect 536943 472561 537545 473163
rect 537957 472511 538587 473141
rect 548153 472577 548783 473207
rect 553163 472501 553793 473131
rect 562803 472429 563433 473059
rect 387914 469723 388024 469789
rect 392806 469723 392916 469789
rect 387924 469351 388034 469417
rect 392816 469351 392926 469417
rect 508976 469023 509086 469089
rect 508986 468651 509096 468717
rect 515023 467765 515133 467831
rect 515033 467393 515143 467459
rect 534386 466945 534496 467011
rect 534376 466573 534486 466639
rect 356026 462172 356136 462238
rect 356036 461800 356146 461866
rect 550370 459665 550480 459731
rect 527531 459536 527641 459602
rect 550360 459293 550470 459359
rect 527521 459164 527631 459230
rect 521414 457098 521524 457164
rect 346996 456998 347106 457064
rect 521424 456726 521534 456792
rect 347006 456626 347116 456692
rect 240701 455849 240811 455915
rect 251423 455827 251533 455893
rect 240711 455477 240821 455543
rect 251433 455455 251543 455521
rect 502200 455171 502310 455237
rect 502210 454799 502320 454865
rect 564164 453285 564230 453395
rect 564536 453295 564602 453405
rect 508964 448972 509074 449038
rect 392796 448771 392906 448837
rect 387875 448703 387985 448769
rect 508974 448600 509084 448666
rect 392806 448399 392916 448465
rect 387885 448331 387995 448397
rect 515060 447564 515170 447630
rect 515070 447192 515180 447258
rect 534376 446545 534486 446611
rect 534366 446173 534476 446239
rect 356000 442179 356110 442245
rect 356010 441807 356120 441873
rect 346968 436390 347078 436456
rect 346978 436018 347088 436084
rect 240621 434332 240731 434398
rect 251406 434046 251516 434112
rect 240631 433960 240741 434026
rect 251416 433674 251526 433740
rect 238866 429718 239407 430259
rect 249235 429837 249777 430379
rect 252980 429821 253522 430363
rect 258338 429822 258878 430362
rect 272940 429757 273482 430299
rect 278450 429801 278992 430343
rect 293214 429813 293756 430355
rect 299162 429713 299704 430255
rect 313348 429649 313890 430191
rect 319476 429615 320018 430157
rect 322085 429673 322627 430215
rect 332869 429829 333411 430371
rect 252958 425977 253024 426087
rect 253330 425967 253396 426077
rect 272904 426042 272970 426152
rect 273276 426032 273342 426142
rect 293185 426076 293251 426186
rect 293557 426066 293623 426176
rect 313334 426066 313400 426176
rect 313706 426056 313772 426166
rect 335394 429711 335936 430253
rect 348094 429382 348522 430698
rect 354357 429727 354899 430269
rect 360001 429897 360543 430439
rect 362171 429901 362713 430443
rect 373950 429649 374492 430191
rect 375352 429653 375894 430195
rect 385933 429745 386475 430287
rect 391205 429829 391747 430371
rect 497210 429770 497838 430398
rect 510283 429683 510885 430285
rect 513067 429733 513669 430335
rect 522311 429699 522913 430301
rect 528959 429699 529589 430329
rect 545783 429773 546413 430403
rect 562801 429699 563431 430329
rect 387904 427660 388014 427726
rect 392828 427679 392938 427745
rect 387914 427288 388024 427354
rect 392838 427307 392948 427373
rect 335541 426041 335607 426151
rect 335913 426051 335979 426161
rect 355531 426037 355597 426147
rect 355903 426047 355969 426157
rect 375494 426131 375560 426241
rect 375866 426141 375932 426251
rect 356005 422225 356115 422291
rect 356015 421853 356125 421919
rect 258312 420479 258378 420589
rect 258684 420469 258750 420579
rect 278446 420512 278512 420622
rect 278818 420502 278884 420612
rect 299123 420518 299189 420628
rect 299495 420508 299561 420618
rect 319451 420470 319517 420580
rect 319823 420460 319889 420570
rect 353761 420469 353827 420579
rect 354133 420479 354199 420589
rect 374104 420539 374170 420649
rect 374476 420549 374542 420659
rect 324544 417112 324654 417178
rect 336554 417037 336664 417103
rect 324554 416740 324664 416806
rect 336564 416665 336674 416731
rect 242019 415360 242560 415901
rect 252972 415372 253512 415912
rect 255273 415185 255815 415727
rect 258336 415336 258876 415876
rect 272932 415267 273474 415809
rect 278450 415273 278992 415815
rect 293214 415247 293756 415789
rect 299136 415271 299678 415813
rect 313354 415329 313896 415871
rect 319466 415405 320008 415947
rect 328159 415359 328701 415901
rect 339875 415321 340417 415863
rect 345550 414894 345978 416210
rect 346912 415756 347022 415822
rect 346922 415384 347032 415450
rect 353573 415233 354115 415775
rect 373944 415303 374486 415845
rect 375340 415107 375882 415649
rect 388617 415307 389159 415849
rect 393665 415385 394207 415927
rect 568046 408878 568112 408988
rect 568418 408868 568484 408978
rect 549553 407130 549663 407196
rect 549543 406758 549653 406824
rect 355994 402190 356104 402256
rect 356004 401818 356114 401884
rect 324542 396322 324652 396388
rect 336579 396384 336689 396450
rect 324552 395950 324662 396016
rect 336589 396012 336699 396078
rect 346940 395078 347050 395144
rect 346950 394706 347060 394772
rect 322895 390805 323437 391347
rect 333092 390825 333634 391367
rect 334879 390767 335421 391309
rect 353565 390397 354107 390939
rect 357690 390615 358232 391157
rect 367484 390651 368026 391193
rect 385269 390627 385811 391169
rect 400437 390647 400979 391189
rect 428501 390755 429043 391297
rect 446395 390507 446937 391049
rect 470027 390513 470569 391055
rect 490269 390563 490811 391105
rect 510723 390533 511265 391075
rect 530385 390605 530927 391147
rect 546403 390679 546965 391241
rect 571227 390643 571789 391205
rect 549570 388086 549680 388152
rect 549560 387714 549670 387780
rect 347446 386614 347512 386724
rect 347818 386604 347884 386714
rect 367462 386643 367528 386753
rect 367834 386633 367900 386743
rect 387274 386633 387340 386743
rect 387646 386623 387712 386733
rect 407533 386631 407599 386741
rect 407905 386621 407971 386731
rect 427809 386686 427875 386796
rect 428181 386676 428247 386786
rect 447968 386666 448034 386776
rect 448340 386656 448406 386766
rect 467970 386661 468036 386771
rect 468342 386651 468408 386761
rect 488088 386645 488154 386755
rect 488460 386635 488526 386745
rect 508218 386668 508284 386778
rect 508590 386658 508656 386768
rect 528327 386682 528393 386792
rect 528699 386672 528765 386782
rect 355974 382126 356084 382192
rect 355984 381754 356094 381820
rect 333077 380647 333143 380757
rect 333449 380637 333515 380747
rect 357656 380655 357722 380765
rect 358028 380645 358094 380755
rect 387103 380613 387169 380723
rect 387475 380603 387541 380713
rect 407681 380644 407747 380754
rect 408053 380634 408119 380744
rect 427655 380619 427721 380729
rect 428027 380609 428093 380719
rect 447901 380623 447967 380733
rect 448273 380613 448339 380723
rect 467885 380690 467951 380800
rect 468257 380680 468323 380790
rect 488300 380615 488366 380725
rect 488672 380605 488738 380715
rect 507983 380687 508049 380797
rect 508355 380677 508421 380787
rect 528353 380621 528419 380731
rect 528725 380611 528791 380721
rect 549368 379428 549478 379494
rect 549378 379056 549488 379122
rect 325765 375553 326307 376095
rect 333090 375667 333632 376209
rect 337333 375573 337875 376115
rect 345681 375547 346223 376089
rect 352330 375608 353838 376280
rect 357684 375559 358226 376101
rect 367484 375509 368026 376051
rect 388559 375377 389101 375919
rect 400425 375559 400967 376101
rect 429149 375465 429691 376007
rect 446411 375523 446953 376065
rect 466549 375507 467091 376049
rect 485509 375463 486051 376005
rect 505733 375447 506275 375989
rect 526305 375627 526847 376169
rect 552361 375485 552923 376047
rect 562709 375559 563271 376121
rect 346926 373796 347036 373862
rect 346936 373424 347046 373490
rect 549329 364242 549439 364308
rect 549339 363870 549449 363936
rect 568202 362495 568268 362605
rect 568574 362485 568640 362595
rect 356031 362143 356141 362209
rect 356041 361771 356151 361837
rect 346926 352946 347036 353012
rect 346936 352574 347046 352640
rect 356031 342140 356141 342206
rect 356041 341768 356151 341834
rect 347010 332350 347120 332416
rect 347020 331978 347130 332044
rect 355955 322138 356065 322204
rect 355965 321766 356075 321832
rect 346982 310482 347092 310548
rect 346992 310110 347102 310176
rect 348024 305644 348476 307618
rect 357945 306237 358487 306779
rect 370688 306263 371237 306812
rect 390700 306391 391249 306940
rect 400264 306349 400813 306898
rect 430714 306113 431263 306662
rect 445440 306311 445989 306860
rect 470718 306231 471267 306780
rect 490714 306455 491263 307004
rect 510700 306347 511249 306896
rect 530686 306193 531235 306742
rect 552167 306173 552724 306730
rect 569358 306237 569927 306806
rect 355993 302117 356103 302183
rect 356003 301745 356113 301811
rect 370828 295924 370894 296034
rect 371200 295934 371266 296044
rect 390837 295941 390903 296051
rect 391209 295951 391275 296061
rect 410843 295912 410909 296022
rect 411215 295922 411281 296032
rect 430839 295988 430905 296098
rect 431211 295998 431277 296108
rect 450856 295955 450922 296065
rect 451228 295965 451294 296075
rect 470858 295980 470924 296090
rect 471230 295990 471296 296100
rect 490853 296013 490919 296123
rect 491225 296023 491291 296133
rect 510846 295969 510912 296079
rect 511218 295979 511284 296089
rect 530831 296013 530897 296123
rect 531203 296023 531269 296133
rect 549547 293375 549657 293441
rect 549557 293003 549667 293069
rect 346940 288824 347050 288890
rect 346950 288452 347060 288518
rect 345710 285614 346162 287588
rect 354041 286271 354583 286813
rect 370688 286058 371237 286607
rect 390700 286142 391249 286691
rect 400180 286354 400729 286903
rect 430714 286260 431263 286809
rect 445452 286472 446001 287021
rect 470718 286204 471267 286753
rect 490714 286334 491263 286883
rect 510700 286270 511249 286819
rect 530686 286258 531235 286807
rect 546320 286426 546877 286983
rect 568318 286313 568887 286882
rect 551449 273906 551515 274016
rect 551821 273916 551887 274026
rect 571912 273866 571978 273976
rect 572284 273876 572350 273986
rect 346898 264044 347008 264110
rect 346908 263672 347018 263738
rect 346982 242670 347092 242736
rect 346992 242298 347102 242364
rect 347010 222794 347120 222860
rect 347020 222422 347130 222488
rect 347982 208088 348448 213096
rect 346954 200966 347064 201032
rect 346964 200594 347074 200660
rect 346968 179932 347078 179998
rect 346978 179560 347088 179626
rect 345722 172818 346188 177826
rect 345698 162828 346164 167836
rect 346926 158544 347036 158610
rect 346936 158172 347046 158238
rect 334827 136843 335369 137385
rect 346870 137198 346980 137264
rect 346880 136826 346990 136892
rect 358795 136827 359337 137369
rect 346926 116064 347036 116130
rect 346936 115692 347046 115758
rect 334799 95097 335341 95639
rect 346954 95454 347064 95520
rect 346964 95082 347074 95148
rect 359143 95097 359685 95639
rect 346940 74772 347050 74838
rect 346950 74400 347060 74466
rect 90284 58752 91538 60006
rect 111727 58819 112269 59361
rect 133049 58829 133591 59371
rect 154607 58785 155149 59327
rect 175813 58785 176355 59327
rect 197195 58741 197737 59283
rect 219089 58763 219631 59305
rect 240075 58839 240617 59381
rect 260577 58837 261119 59379
rect 281389 58593 281931 59135
rect 302579 58961 303121 59503
rect 324127 58961 324669 59503
rect 334723 53983 335265 54525
rect 358805 53983 359347 54525
rect 39905 51899 40867 52861
rect 347010 51192 347120 51258
rect 347020 50820 347130 50886
rect 47990 48776 48056 48886
rect 48362 48786 48428 48896
rect 69284 48836 69350 48946
rect 69656 48846 69722 48956
rect 90650 48762 90716 48872
rect 91022 48772 91088 48882
rect 111710 48806 111776 48916
rect 112082 48816 112148 48926
rect 133032 48850 133098 48960
rect 133404 48860 133470 48970
rect 154590 48820 154656 48930
rect 154962 48830 155028 48940
rect 175796 48792 175862 48902
rect 176168 48802 176234 48912
rect 197178 48850 197244 48960
rect 197550 48860 197616 48970
rect 219072 48762 219138 48872
rect 219444 48772 219510 48882
rect 240058 48732 240124 48842
rect 240430 48742 240496 48852
rect 260560 48792 260626 48902
rect 260932 48802 260998 48912
rect 281372 48894 281438 49004
rect 281744 48904 281810 49014
rect 302562 48688 302628 48798
rect 302934 48698 303000 48808
rect 324110 48724 324176 48834
rect 324482 48734 324548 48844
rect 34578 42938 34688 43004
rect 34588 42566 34698 42632
rect 39650 36270 42762 39258
rect 48009 37365 48551 37907
rect 69303 37471 69845 38013
rect 90669 37153 91211 37695
rect 111729 37205 112271 37747
rect 133051 37125 133593 37667
rect 154609 37293 155151 37835
rect 175815 37293 176357 37835
rect 197197 37391 197739 37933
rect 219091 37341 219633 37883
rect 240077 37239 240619 37781
rect 260579 37177 261121 37719
rect 281391 37273 281933 37815
rect 302581 37377 303123 37919
rect 324129 37325 324671 37867
rect 34578 20840 34688 20906
rect 34588 20468 34698 20534
rect 338576 8478 338688 8590
rect 6548 3452 6614 3562
rect 6920 3462 6986 3572
rect 27740 3512 27806 3622
rect 28112 3522 28178 3632
rect 356306 8088 356418 8200
rect 342122 7742 342234 7854
rect 345668 7144 345780 7256
rect 352760 7184 352872 7296
rect 349584 6516 349696 6628
rect 476870 3908 476982 4020
rect 480416 3908 480528 4020
rect 483962 3912 484074 4024
<< metal3 >>
rect 16194 702737 21194 704800
rect 15877 695646 21331 702737
rect 68194 702547 73194 704800
rect 120194 702701 125194 704800
rect 49727 695646 55181 695653
rect 15877 690192 55181 695646
rect 558 685242 41326 685356
rect -800 680242 41326 685242
rect 558 679902 41326 680242
rect 5371 648752 8383 648776
rect 805 648642 8383 648752
rect -800 643842 8383 648642
rect 805 643688 8383 643842
rect 13471 643688 13477 648776
rect 805 643686 5945 643688
rect 5371 638726 8391 638742
rect 805 638642 8391 638726
rect -800 633842 8391 638642
rect 805 633670 8391 633842
rect 13463 633670 13469 638742
rect 805 633660 5945 633670
rect 35872 617459 41326 679902
rect 49727 657865 55181 690192
rect 68098 673045 73321 702547
rect 119810 690196 125221 702701
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702955 418394 704800
rect 465394 703014 470394 704800
rect 413191 690689 418453 702955
rect 119810 684785 260348 690196
rect 68098 667822 227958 673045
rect 49727 652411 203813 657865
rect 198359 646060 203813 652411
rect 222735 646060 227958 667822
rect 254937 646060 260348 684785
rect 285478 685427 418453 690689
rect 465252 702300 470394 703014
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 703689 571594 704800
rect 285478 646060 290740 685427
rect 465252 675437 470365 702300
rect 566410 693330 571704 703689
rect 308691 670324 470365 675437
rect 501739 688036 571704 693330
rect 308691 646060 313804 670324
rect 501739 655869 507033 688036
rect 571542 682984 582953 683337
rect 571542 677984 584800 682984
rect 571542 677569 582953 677984
rect 571542 665727 577310 677569
rect 342062 650575 507033 655869
rect 530161 659959 577310 665727
rect 342062 646060 347356 650575
rect 199510 623965 200510 646060
rect 224356 628106 225356 646060
rect 257844 640529 258844 646060
rect 238371 639529 258844 640529
rect 224356 627106 232299 628106
rect 199510 622965 217854 623965
rect 35872 615141 171201 617459
rect 35872 614141 210863 615141
rect 35872 612005 171201 614141
rect 209863 588028 210863 614141
rect 216854 588501 217854 622965
rect 231299 588737 232299 627106
rect 238371 587555 239371 639529
rect 287552 633507 288552 646060
rect 248373 632507 288552 633507
rect 248373 588028 249373 632507
rect 310957 628466 311957 646060
rect 259248 627466 311957 628466
rect 259248 587083 260248 627466
rect 344265 622344 345265 646060
rect 267558 621344 345265 622344
rect 267558 587733 268558 621344
rect 530161 618189 535929 659959
rect 570812 639592 570818 644694
rect 575920 644684 580012 644694
rect 575920 644584 583353 644684
rect 575920 639784 584800 644584
rect 575920 639592 583353 639784
rect 578927 639578 583353 639592
rect 579387 634674 583813 634748
rect 570867 629638 570873 634674
rect 575909 634584 583813 634674
rect 575909 629784 584800 634584
rect 575909 629642 583813 629784
rect 575909 629638 580012 629642
rect 356710 616223 535929 618189
rect 276898 615223 535929 616223
rect 276898 587124 277898 615223
rect 356710 612421 535929 615223
rect 286354 602558 487607 603558
rect 488607 602558 488613 603558
rect 286354 587425 287354 602558
rect 288354 596090 482433 597090
rect 483433 596090 483439 597090
rect 288354 587536 289354 596090
rect 290346 589077 477776 590077
rect 478776 589077 478782 590077
rect 565585 589584 565697 589590
rect 565697 589472 584800 589584
rect 565585 589466 565697 589472
rect 290346 589012 291354 589077
rect 290346 586827 291346 589012
rect 577012 588290 584800 588402
rect 544391 587292 550550 587293
rect 544386 586294 544392 587292
rect 545390 586885 550550 587292
rect 551431 586924 571518 587293
rect 572580 586958 576060 587293
rect 577012 586958 577124 588290
rect 583473 587108 584800 587220
rect 551431 586892 571980 586924
rect 572580 586921 577124 586958
rect 545390 586861 550966 586885
rect 551431 586883 571882 586892
rect 545390 586751 550871 586861
rect 550937 586751 550966 586861
rect 545390 586721 550966 586751
rect 551225 586851 571882 586883
rect 551225 586741 551243 586851
rect 551309 586782 571882 586851
rect 571948 586782 571980 586892
rect 551309 586741 571980 586782
rect 551225 586740 571980 586741
rect 572211 586882 577124 586921
rect 572211 586772 572254 586882
rect 572320 586846 577124 586882
rect 572320 586772 576060 586846
rect 545390 586294 550550 586721
rect 551225 586716 571518 586740
rect 572211 586737 576060 586772
rect 544391 586293 550550 586294
rect 551431 586293 571518 586716
rect 572580 586293 576060 586737
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 537798 578716 537804 579328
rect 538406 579323 538416 579328
rect 538411 578721 538416 579323
rect 538406 578716 538416 578721
rect 544726 573219 544856 573224
rect 544726 573153 544736 573219
rect 544846 573153 544856 573219
rect 544726 573148 544856 573153
rect 544716 572847 544846 572852
rect 544716 572781 544726 572847
rect 544836 572781 544846 572847
rect 544716 572776 544846 572781
rect 522151 568442 525018 568443
rect 505085 568273 506083 568278
rect 505084 568272 513276 568273
rect 505084 567274 505085 568272
rect 506083 567274 513276 568272
rect 505084 567273 513276 567274
rect 514276 567273 514282 568273
rect 522146 567444 522152 568442
rect 523150 568017 525018 568442
rect 523150 567981 525424 568017
rect 525876 568005 530514 568443
rect 523150 567871 525320 567981
rect 525386 567871 525424 567981
rect 523150 567827 525424 567871
rect 525641 567971 530514 568005
rect 525641 567861 525692 567971
rect 525758 567861 530514 567971
rect 523150 567444 525018 567827
rect 525641 567815 530514 567861
rect 522151 567443 525018 567444
rect 525876 567443 530514 567815
rect 531514 567443 531520 568443
rect 505085 567268 506083 567273
rect -800 559442 1660 564242
rect 513752 562663 513882 562668
rect 513752 562597 513762 562663
rect 513872 562597 513882 562663
rect 513752 562592 513882 562597
rect 513742 562291 513872 562296
rect 513742 562225 513752 562291
rect 513862 562225 513872 562291
rect 513742 562220 513872 562225
rect 505439 560570 505569 560575
rect 505439 560504 505449 560570
rect 505559 560504 505569 560570
rect 505439 560499 505569 560504
rect 505429 560198 505559 560203
rect 505429 560132 505439 560198
rect 505549 560132 505559 560198
rect 505429 560127 505559 560132
rect 526598 556182 527218 556187
rect 509398 556160 509948 556165
rect 509398 554242 509408 556160
rect 509938 554242 509948 556160
rect -800 549442 1660 554242
rect 509398 554237 509948 554242
rect 526598 554236 526608 556182
rect 527208 554236 527218 556182
rect 526598 554231 527218 554236
rect 547172 556178 547768 556183
rect 547172 554212 547182 556178
rect 547758 554212 547768 556178
rect 547172 554207 547768 554212
rect 531022 553109 531152 553114
rect 531022 553043 531032 553109
rect 531142 553043 531152 553109
rect 531022 553038 531152 553043
rect 544736 552970 544866 552975
rect 544736 552904 544746 552970
rect 544856 552904 544866 552970
rect 544736 552899 544866 552904
rect 531012 552737 531142 552742
rect 531012 552671 531022 552737
rect 531132 552671 531142 552737
rect 531012 552666 531142 552671
rect 544726 552598 544856 552603
rect 544726 552532 544736 552598
rect 544846 552532 544856 552598
rect 544726 552527 544856 552532
rect 582340 550562 584800 555362
rect 522501 550492 522631 550497
rect 522501 550426 522511 550492
rect 522621 550426 522631 550492
rect 522501 550421 522631 550426
rect 522491 550120 522621 550125
rect 522491 550054 522501 550120
rect 522611 550054 522621 550120
rect 522491 550049 522621 550054
rect 118329 542857 123445 542862
rect 118328 542856 147895 542857
rect 118328 537740 118329 542856
rect 123445 537740 147895 542856
rect 513732 542221 513862 542226
rect 513732 542155 513742 542221
rect 513852 542155 513862 542221
rect 513732 542150 513862 542155
rect 513722 541849 513852 541854
rect 513722 541783 513732 541849
rect 513842 541783 513852 541849
rect 513722 541778 513852 541783
rect 582340 540562 584800 545362
rect 537824 540294 538420 540299
rect 517864 540212 518584 540217
rect 505549 539982 505679 539987
rect 505549 539916 505559 539982
rect 505669 539916 505679 539982
rect 505549 539911 505679 539916
rect 500438 539636 501050 539642
rect 484623 539557 484633 539562
rect 464232 539447 464242 539452
rect 464232 538845 464237 539447
rect 464232 538840 464242 538845
rect 464844 538840 464850 539452
rect 484623 538955 484628 539557
rect 484623 538950 484633 538955
rect 485235 538950 485241 539562
rect 505539 539610 505669 539615
rect 505539 539544 505549 539610
rect 505659 539544 505669 539610
rect 505539 539539 505669 539544
rect 500438 539029 500443 539034
rect 501045 539029 501050 539034
rect 500438 539024 501050 539029
rect 517864 538396 517874 540212
rect 518574 538396 518584 540212
rect 517864 538391 518584 538396
rect 537824 538328 537834 540294
rect 538410 538328 538420 540294
rect 565228 538344 565238 540236
rect 566160 538344 566170 540236
rect 537824 538323 538420 538328
rect 118328 537739 147895 537740
rect 118329 537734 123445 537739
rect 425730 535389 425794 535395
rect 402219 535327 425730 535387
rect 425730 535319 425794 535325
rect 423449 532949 423513 532955
rect 402264 532887 423449 532947
rect 423449 532879 423513 532885
rect 544741 532744 544871 532749
rect 544741 532678 544751 532744
rect 544861 532678 544871 532744
rect 544741 532673 544871 532678
rect 355561 532597 356561 532603
rect 338673 531597 355561 532597
rect 356561 531597 366475 532597
rect 544731 532372 544861 532377
rect 544731 532306 544741 532372
rect 544851 532306 544861 532372
rect 544731 532301 544861 532306
rect 530977 531864 531107 531869
rect 530977 531798 530987 531864
rect 531097 531798 531107 531864
rect 530977 531793 531107 531798
rect 355561 531591 356561 531597
rect 118329 526347 123445 526352
rect 118328 526346 148605 526347
rect 118328 521230 118329 526346
rect 123445 521230 148605 526346
rect 355986 522111 356106 522121
rect 355981 522045 355991 522111
rect 356101 522045 356111 522111
rect 355986 522035 356106 522045
rect 365475 522025 366475 531597
rect 530967 531492 531097 531497
rect 530967 531426 530977 531492
rect 531087 531426 531097 531492
rect 530967 531421 531097 531426
rect 421586 530387 421650 530393
rect 402219 530325 421586 530385
rect 421586 530317 421650 530323
rect 522550 529715 522680 529720
rect 522550 529649 522560 529715
rect 522670 529649 522680 529715
rect 522550 529644 522680 529649
rect 522540 529343 522670 529348
rect 522540 529277 522550 529343
rect 522660 529277 522670 529343
rect 522540 529272 522670 529277
rect 419511 527947 419575 527953
rect 402230 527885 419511 527945
rect 419511 527877 419575 527883
rect 417539 525383 417545 525385
rect 402078 525323 417545 525383
rect 417539 525321 417545 525323
rect 417609 525321 417615 525385
rect 415539 522943 415545 522945
rect 401983 522883 415545 522943
rect 415539 522881 415545 522883
rect 415609 522881 415615 522945
rect 513729 522250 513859 522255
rect 513729 522184 513739 522250
rect 513849 522184 513859 522250
rect 513729 522179 513859 522184
rect 365475 522007 368109 522025
rect 355996 521739 356116 521749
rect 355991 521673 356001 521739
rect 356111 521673 356121 521739
rect 355996 521663 356116 521673
rect 118328 521229 148605 521230
rect 365475 521479 372498 522007
rect 513719 521878 513849 521883
rect 513719 521812 513729 521878
rect 513839 521812 513849 521878
rect 513719 521807 513849 521812
rect 365475 521419 373965 521479
rect 118329 521224 123445 521229
rect 365475 521025 372498 521419
rect 367231 521007 372498 521025
rect 413516 520383 413580 520389
rect 401504 520321 413516 520381
rect 413516 520313 413580 520319
rect 522151 519803 523151 519809
rect 513276 519802 522151 519803
rect 505084 519692 506084 519698
rect 403846 519227 423959 519345
rect 424869 519273 443786 519692
rect 444987 519356 463996 519692
rect 465154 519565 484281 519692
rect 444987 519330 464547 519356
rect 465156 519350 484281 519565
rect 424869 519247 444364 519273
rect 444987 519267 464455 519330
rect 403846 519188 424355 519227
rect 424869 519214 444272 519247
rect 403604 519108 403674 519113
rect 403846 519108 424259 519188
rect 403604 519048 403609 519108
rect 403669 519078 424259 519108
rect 424325 519078 424355 519188
rect 403669 519048 424355 519078
rect 403604 519043 403674 519048
rect 403846 519034 424355 519048
rect 424592 519178 444272 519214
rect 424592 519068 424631 519178
rect 424697 519137 444272 519178
rect 444338 519137 444364 519247
rect 424697 519113 444364 519137
rect 444624 519237 464455 519267
rect 444624 519127 444644 519237
rect 444710 519220 464455 519237
rect 464521 519220 464547 519330
rect 444710 519196 464547 519220
rect 464807 519320 484281 519350
rect 464807 519210 464827 519320
rect 464893 519317 484281 519320
rect 485492 519324 503896 519692
rect 464893 519291 484879 519317
rect 485492 519311 504353 519324
rect 504960 519318 505084 519692
rect 464893 519210 484787 519291
rect 444710 519127 463996 519196
rect 464807 519190 484787 519210
rect 424697 519068 443786 519113
rect 444624 519107 463996 519127
rect 403846 518839 423959 519034
rect 424592 519021 443786 519068
rect 424869 518692 443786 519021
rect 444987 518692 463996 519107
rect 465154 519181 484787 519190
rect 484853 519181 484879 519291
rect 465154 519157 484879 519181
rect 485139 519298 504353 519311
rect 485139 519281 504261 519298
rect 485139 519171 485159 519281
rect 485225 519188 504261 519281
rect 504327 519188 504353 519298
rect 485225 519171 504353 519188
rect 485139 519164 504353 519171
rect 504613 519288 505084 519318
rect 504613 519178 504633 519288
rect 504699 519178 505084 519288
rect 465154 518692 484281 519157
rect 485139 519151 503896 519164
rect 504613 519158 505084 519178
rect 485492 518692 503896 519151
rect 504960 518692 505084 519158
rect 506084 518692 506218 519692
rect 513271 518804 513277 519802
rect 514275 518804 522151 519802
rect 513276 518803 522151 518804
rect 530514 519802 537373 519803
rect 530509 518804 530515 519802
rect 531513 519466 537373 519802
rect 538383 519792 542371 519803
rect 544391 519792 545391 519798
rect 531513 519443 537783 519466
rect 538383 519458 544391 519792
rect 531513 519333 537690 519443
rect 537756 519333 537783 519443
rect 531513 519304 537783 519333
rect 538037 519433 544391 519458
rect 538037 519323 538062 519433
rect 538128 519323 544391 519433
rect 531513 518804 537373 519304
rect 538037 519296 544391 519323
rect 530514 518803 537373 518804
rect 522151 518797 523151 518803
rect 538383 518792 544391 519296
rect 544391 518786 545391 518792
rect 505084 518686 506084 518692
rect 411487 517943 411551 517949
rect 402002 517881 411487 517941
rect 411487 517873 411551 517879
rect 365528 517349 366528 517355
rect 366528 516928 372498 517349
rect 366528 516868 372209 516928
rect 372269 516868 372498 516928
rect 366528 516349 372498 516868
rect 365528 516343 366528 516349
rect 409483 515381 409547 515387
rect 402220 515319 409483 515379
rect 409483 515311 409547 515317
rect 407542 512941 407606 512947
rect 402309 512879 407542 512939
rect 407542 512871 407606 512877
rect -800 511530 480 511642
rect 501674 510564 502674 510570
rect 508549 510564 509547 510569
rect -800 510348 480 510460
rect 405502 510379 405566 510385
rect 401843 510317 405502 510377
rect 405502 510309 405566 510315
rect 502674 510563 509548 510564
rect 502674 509565 508549 510563
rect 509547 509565 509548 510563
rect 502674 509564 509548 509565
rect 514542 510484 515542 510490
rect 501674 509558 502674 509564
rect 508549 509559 509547 509564
rect 515542 510483 522016 510484
rect 515542 509485 521017 510483
rect 522015 509485 522021 510483
rect 515542 509484 522016 509485
rect 514542 509478 515542 509484
rect 527084 509404 527090 510404
rect 528090 510403 534844 510404
rect 528090 509405 533845 510403
rect 534843 509405 534849 510403
rect 528090 509404 534844 509405
rect -800 509166 480 509278
rect 83456 509247 84454 509252
rect 13939 509246 84455 509247
rect 12230 508887 12340 508892
rect 13939 508887 83456 509246
rect 12229 508886 83456 508887
rect 12229 508776 12230 508886
rect 12340 508776 83456 508886
rect 12229 508775 83456 508776
rect 12230 508770 12340 508775
rect 13939 508248 83456 508775
rect 84454 508248 84455 509246
rect 534324 508952 534454 508957
rect 534324 508886 534334 508952
rect 534444 508886 534454 508952
rect 534324 508881 534454 508886
rect 534334 508580 534464 508585
rect 534334 508514 534344 508580
rect 534454 508514 534464 508580
rect 534334 508509 534464 508514
rect 13939 508247 84455 508248
rect 83456 508242 84454 508247
rect -800 507984 480 508096
rect 515028 507933 515158 507938
rect 515028 507867 515038 507933
rect 515148 507867 515158 507933
rect 515028 507862 515158 507867
rect 403541 507817 403605 507823
rect 118329 507811 123445 507816
rect 118328 507810 148401 507811
rect 12229 506914 12341 506920
rect -800 506802 12229 506914
rect 12229 506796 12341 506802
rect -800 505620 25370 505732
rect 25482 505620 25488 505732
rect 118328 502694 118329 507810
rect 123445 502694 148401 507810
rect 387908 507753 387914 507817
rect 387978 507815 387984 507817
rect 387978 507755 388477 507815
rect 402339 507755 403541 507815
rect 387978 507753 387984 507755
rect 403541 507747 403605 507753
rect 515018 507561 515148 507566
rect 515018 507495 515028 507561
rect 515138 507495 515148 507561
rect 515018 507490 515148 507495
rect 508932 506525 509062 506530
rect 508932 506459 508942 506525
rect 509052 506459 509062 506525
rect 508932 506454 509062 506459
rect 508922 506153 509052 506158
rect 508922 506087 508932 506153
rect 509042 506087 509052 506153
rect 508922 506082 509052 506087
rect 350839 504930 351065 504936
rect 340115 504704 350839 504930
rect 350839 504698 351065 504704
rect 373560 504707 373808 504793
rect 373560 504637 373642 504707
rect 373712 504637 373808 504707
rect 383174 504762 383339 504801
rect 383174 504757 383216 504762
rect 383174 504697 383215 504757
rect 383174 504692 383216 504697
rect 383280 504692 383339 504762
rect 383174 504647 383339 504692
rect 373560 504536 373808 504637
rect 387425 504447 388425 504968
rect 392669 504721 392960 504847
rect 392669 504716 392784 504721
rect 392669 504656 392783 504716
rect 392669 504651 392784 504656
rect 392848 504651 392960 504721
rect 392669 504545 392960 504651
rect 350185 502978 350411 502984
rect 340341 502752 350185 502978
rect 350185 502746 350411 502752
rect 118328 502693 148401 502694
rect 118329 502688 123445 502693
rect 355951 502202 356071 502212
rect 355946 502136 355956 502202
rect 356066 502136 356076 502202
rect 355951 502126 356071 502136
rect 355961 501830 356081 501840
rect 355956 501764 355966 501830
rect 356076 501764 356086 501830
rect 355961 501754 356081 501764
rect 502168 500326 502298 500331
rect 502168 500260 502178 500326
rect 502288 500260 502298 500326
rect 502168 500255 502298 500260
rect 559955 500162 560067 500168
rect 559949 500052 559955 500162
rect 560067 500050 584800 500162
rect 559955 500044 560067 500050
rect 502158 499954 502288 499959
rect 502158 499888 502168 499954
rect 502278 499888 502288 499954
rect 502158 499883 502288 499888
rect 583520 498868 584800 498980
rect 521382 498399 521512 498404
rect 521382 498333 521392 498399
rect 521502 498333 521512 498399
rect 521382 498328 521512 498333
rect 549985 498323 563892 498324
rect 521372 498027 521502 498032
rect 521372 497961 521382 498027
rect 521492 497961 521502 498027
rect 521372 497956 521502 497961
rect 549980 497325 549986 498323
rect 550984 497915 563892 498323
rect 550984 497870 564335 497915
rect 565132 497899 578145 498324
rect 550984 497760 564230 497870
rect 564296 497760 564335 497870
rect 550984 497724 564335 497760
rect 564566 497860 578145 497899
rect 564566 497750 564602 497860
rect 564668 497798 578145 497860
rect 564668 497750 584800 497798
rect 550984 497325 563892 497724
rect 564566 497708 584800 497750
rect 549985 497324 563892 497325
rect 565132 497686 584800 497708
rect 565132 497324 578145 497686
rect 339345 496736 349515 496962
rect 349741 496736 349747 496962
rect 583520 496504 584800 496616
rect 527456 496001 527586 496006
rect 527456 495935 527466 496001
rect 527576 495935 527586 496001
rect 527456 495930 527586 495935
rect 527446 495629 527576 495634
rect 527446 495563 527456 495629
rect 527566 495563 527576 495629
rect 527446 495558 527576 495563
rect 583520 495322 584800 495434
rect 348839 494918 349065 494924
rect 339771 494692 348839 494918
rect 348839 494686 349065 494692
rect 583520 494140 584800 494252
rect 550456 492056 550586 492061
rect 550456 491990 550466 492056
rect 550576 491990 550586 492056
rect 550456 491985 550586 491990
rect 550446 491684 550576 491689
rect 550446 491618 550456 491684
rect 550566 491618 550576 491684
rect 550446 491613 550576 491618
rect 392803 490767 392923 490777
rect 387900 490753 388020 490763
rect 387895 490687 387905 490753
rect 388015 490687 388025 490753
rect 392798 490701 392808 490767
rect 392918 490701 392928 490767
rect 392803 490691 392923 490701
rect 373611 490674 373731 490684
rect 373606 490608 373616 490674
rect 373726 490608 373736 490674
rect 383263 490672 383383 490682
rect 387900 490677 388020 490687
rect 373611 490598 373731 490608
rect 383258 490606 383268 490672
rect 383378 490606 383388 490672
rect 383263 490596 383383 490606
rect 392813 490395 392933 490405
rect 387910 490381 388030 490391
rect 387905 490315 387915 490381
rect 388025 490315 388035 490381
rect 392808 490329 392818 490395
rect 392928 490329 392938 490395
rect 392813 490319 392933 490329
rect 373621 490302 373741 490312
rect 373616 490236 373626 490302
rect 373736 490236 373746 490302
rect 383273 490300 383393 490310
rect 387910 490305 388030 490315
rect 373621 490226 373741 490236
rect 383268 490234 383278 490300
rect 383388 490234 383398 490300
rect 383273 490224 383393 490234
rect 534334 488552 534464 488557
rect 534334 488486 534344 488552
rect 534454 488486 534464 488552
rect 534334 488481 534464 488486
rect 534344 488180 534474 488185
rect 534344 488114 534354 488180
rect 534464 488114 534474 488180
rect 534344 488109 534474 488114
rect 514991 487732 515121 487737
rect 514991 487666 515001 487732
rect 515111 487666 515121 487732
rect 514991 487661 515121 487666
rect 514981 487360 515111 487365
rect 335518 486302 346574 487302
rect 347574 486302 347580 487302
rect 514981 487294 514991 487360
rect 515101 487294 515111 487360
rect 514981 487289 515111 487294
rect 508944 486474 509074 486479
rect 508944 486408 508954 486474
rect 509064 486408 509074 486474
rect 508944 486403 509074 486408
rect 508934 486102 509064 486107
rect 508934 486036 508944 486102
rect 509054 486036 509064 486102
rect 508934 486031 509064 486036
rect 458514 485312 459126 485318
rect 375484 485289 376036 485294
rect 375484 485284 375489 485289
rect 376031 485284 376036 485289
rect 360438 485152 360990 485158
rect 345009 484722 345235 484728
rect 340171 484496 345009 484722
rect 434800 485229 435412 485234
rect 375484 484736 376036 484742
rect 386090 485213 386642 485218
rect 386090 485208 386095 485213
rect 386637 485208 386642 485213
rect 386090 484660 386642 484666
rect 390324 485216 390876 485222
rect 428636 485221 429188 485226
rect 428636 485216 428641 485221
rect 429183 485216 429188 485221
rect 390324 484669 390329 484674
rect 390871 484669 390876 484674
rect 390324 484664 390876 484669
rect 400218 485186 400770 485192
rect 428636 484668 429188 484674
rect 434800 485224 434805 485229
rect 435407 485224 435412 485229
rect 400218 484639 400223 484644
rect 400765 484639 400770 484644
rect 400218 484634 400770 484639
rect 531886 485221 532526 485226
rect 458514 484705 458519 484710
rect 459121 484705 459126 484710
rect 458514 484700 459126 484705
rect 464285 485162 464897 485168
rect 434800 484616 435412 484622
rect 360438 484605 360443 484610
rect 360985 484605 360990 484610
rect 360438 484600 360990 484605
rect 464285 484555 464290 484560
rect 464892 484555 464897 484560
rect 464285 484550 464897 484555
rect 475004 485132 475616 485138
rect 484617 484588 484623 485200
rect 485225 485195 485235 485200
rect 485230 484593 485235 485195
rect 504622 485170 505234 485176
rect 485225 484588 485235 484593
rect 475004 484525 475009 484530
rect 475611 484525 475616 484530
rect 475004 484520 475616 484525
rect 498492 484504 498498 485116
rect 499100 485111 499110 485116
rect 499105 484509 499110 485111
rect 511833 484608 511839 485220
rect 512441 485215 512451 485220
rect 512446 484613 512451 485215
rect 512441 484608 512451 484613
rect 518202 484580 518208 485220
rect 518838 485215 518848 485220
rect 518843 484585 518848 485215
rect 531886 485216 531891 485221
rect 532521 485216 532526 485221
rect 530384 485178 530996 485184
rect 518838 484580 518848 484585
rect 524285 485159 524295 485164
rect 504622 484563 504627 484568
rect 505229 484563 505234 484568
rect 504622 484558 505234 484563
rect 524285 484557 524290 485159
rect 524285 484552 524295 484557
rect 524897 484552 524903 485164
rect 567844 485171 567854 485176
rect 531886 484580 532526 484586
rect 530384 484571 530389 484576
rect 530991 484571 530996 484576
rect 530384 484566 530996 484571
rect 499100 484504 499110 484509
rect 345009 484490 345235 484496
rect 545773 484492 545779 485132
rect 546409 485127 546419 485132
rect 546414 484497 546419 485127
rect 567844 484541 567849 485171
rect 567844 484536 567854 484541
rect 568484 484536 568490 485176
rect 546409 484492 546419 484497
rect 344281 482404 344507 482410
rect 340351 482178 344281 482404
rect 356013 482258 356133 482268
rect 356008 482192 356018 482258
rect 356128 482192 356138 482258
rect 356013 482182 356133 482192
rect 344281 482172 344507 482178
rect 356023 481886 356143 481896
rect 356018 481820 356028 481886
rect 356138 481820 356148 481886
rect 356023 481810 356143 481820
rect 501402 480113 502774 480116
rect 382734 480108 383958 480109
rect 382729 479110 382735 480108
rect 383733 479740 383958 480108
rect 384879 479765 399342 480109
rect 400445 479771 419546 480109
rect 384879 479746 399627 479765
rect 383733 479710 384172 479740
rect 383733 479600 384086 479710
rect 384152 479600 384172 479710
rect 383733 479580 384172 479600
rect 384432 479735 399627 479746
rect 384432 479720 399541 479735
rect 384432 479610 384458 479720
rect 384524 479625 399541 479720
rect 399607 479625 399627 479735
rect 384524 479610 399627 479625
rect 399887 479745 419546 479771
rect 399887 479635 399913 479745
rect 399979 479705 419546 479745
rect 420619 479734 439798 480109
rect 440819 479746 460112 480109
rect 461175 479752 480245 480109
rect 440819 479740 460407 479746
rect 420619 479711 440107 479734
rect 399979 479675 419869 479705
rect 399979 479635 419783 479675
rect 399887 479611 419783 479635
rect 384432 479605 399627 479610
rect 384432 479586 399342 479605
rect 383733 479110 383958 479580
rect 382734 479109 383958 479110
rect 384879 479109 399342 479586
rect 400445 479565 419783 479611
rect 419849 479565 419869 479675
rect 400445 479545 419869 479565
rect 420129 479704 440107 479711
rect 420129 479685 440021 479704
rect 420129 479575 420155 479685
rect 420221 479594 440021 479685
rect 440087 479594 440107 479704
rect 420221 479575 440107 479594
rect 440367 479716 460407 479740
rect 440367 479714 460321 479716
rect 440367 479604 440393 479714
rect 440459 479606 460321 479714
rect 460387 479606 460407 479716
rect 440459 479604 460407 479606
rect 440367 479586 460407 479604
rect 460667 479726 480245 479752
rect 481410 479730 500313 480109
rect 460667 479616 460693 479726
rect 460759 479724 480245 479726
rect 460759 479694 480589 479724
rect 460759 479616 480503 479694
rect 460667 479592 480503 479616
rect 440367 479580 460112 479586
rect 420129 479574 440107 479575
rect 420129 479551 439798 479574
rect 400445 479109 419546 479545
rect 420619 479109 439798 479551
rect 440819 479109 460112 479580
rect 461175 479584 480503 479592
rect 480569 479584 480589 479694
rect 461175 479564 480589 479584
rect 480849 479704 500313 479730
rect 480849 479594 480875 479704
rect 480941 479636 500313 479704
rect 480941 479616 500545 479636
rect 501402 479630 501675 480113
rect 480941 479594 500459 479616
rect 480849 479570 500459 479594
rect 461175 479109 480245 479564
rect 481410 479506 500459 479570
rect 500525 479506 500545 479616
rect 481410 479476 500545 479506
rect 500805 479606 501675 479630
rect 500805 479496 500831 479606
rect 500897 479496 501675 479606
rect 481410 479109 500313 479476
rect 500805 479470 501675 479496
rect 501402 479116 501675 479470
rect 501669 479115 501675 479116
rect 502673 479116 502774 480113
rect 502673 479115 502679 479116
rect 508542 479114 508548 480114
rect 509548 480113 515542 480114
rect 509548 479115 514543 480113
rect 515541 479115 515547 480113
rect 509548 479114 515542 479115
rect 521010 479114 521016 480114
rect 522016 479779 522636 480114
rect 523714 480113 528090 480114
rect 523714 479792 527091 480113
rect 522016 479743 523014 479779
rect 522016 479633 522909 479743
rect 522975 479633 523014 479743
rect 522016 479586 523014 479633
rect 523251 479753 527091 479792
rect 523251 479643 523281 479753
rect 523347 479643 527091 479753
rect 523251 479599 527091 479643
rect 522016 479114 522636 479586
rect 523714 479115 527091 479599
rect 528089 479115 528095 480113
rect 533838 479116 533844 480116
rect 534844 480109 536275 480116
rect 549985 480109 550985 480115
rect 534844 480108 545444 480109
rect 546779 480108 549985 480109
rect 534844 479663 545541 480108
rect 534844 479620 545919 479663
rect 546674 479644 549985 480108
rect 534844 479510 545802 479620
rect 545868 479510 545919 479620
rect 534844 479463 545919 479510
rect 546149 479610 549985 479644
rect 546149 479500 546174 479610
rect 546240 479500 549985 479610
rect 534844 479116 545541 479463
rect 546149 479459 549985 479500
rect 523714 479114 528090 479115
rect 535757 479109 545541 479116
rect 545195 479108 545541 479109
rect 546674 479109 549985 479459
rect 546674 479108 546922 479109
rect 549985 479103 550985 479109
rect 346977 478318 347097 478328
rect 346972 478252 346982 478318
rect 347092 478252 347102 478318
rect 346977 478242 347097 478252
rect 346987 477946 347107 477956
rect 346982 477880 346992 477946
rect 347102 477880 347112 477946
rect 346987 477870 347107 477880
rect 373156 476016 374154 476021
rect 373155 476015 378904 476016
rect 373155 475017 373156 476015
rect 374154 475639 378904 476015
rect 379826 475672 399342 476016
rect 400445 475678 419546 476016
rect 379826 475645 399627 475672
rect 379397 475642 399627 475645
rect 374154 475609 379137 475639
rect 374154 475499 379051 475609
rect 379117 475499 379137 475609
rect 374154 475479 379137 475499
rect 379397 475619 399541 475642
rect 379397 475509 379423 475619
rect 379489 475532 399541 475619
rect 399607 475532 399627 475642
rect 379489 475512 399627 475532
rect 399887 475652 419546 475678
rect 399887 475542 399913 475652
rect 399979 475612 419546 475652
rect 420619 475641 439798 476016
rect 440819 475653 460112 476016
rect 461175 475659 480245 476016
rect 440819 475647 460407 475653
rect 420619 475618 440107 475641
rect 399979 475582 419869 475612
rect 399979 475542 419783 475582
rect 399887 475518 419783 475542
rect 379489 475509 399342 475512
rect 379397 475485 399342 475509
rect 374154 475017 378904 475479
rect 373155 475016 378904 475017
rect 379826 475016 399342 475485
rect 400445 475472 419783 475518
rect 419849 475472 419869 475582
rect 400445 475452 419869 475472
rect 420129 475611 440107 475618
rect 420129 475592 440021 475611
rect 420129 475482 420155 475592
rect 420221 475501 440021 475592
rect 440087 475501 440107 475611
rect 420221 475482 440107 475501
rect 440367 475623 460407 475647
rect 440367 475621 460321 475623
rect 440367 475511 440393 475621
rect 440459 475513 460321 475621
rect 460387 475513 460407 475623
rect 440459 475511 460407 475513
rect 440367 475493 460407 475511
rect 460667 475633 480245 475659
rect 481410 475649 500345 476016
rect 501701 476009 501707 476010
rect 501434 475655 501707 476009
rect 481410 475637 500577 475649
rect 460667 475523 460693 475633
rect 460759 475631 480245 475633
rect 460759 475601 480589 475631
rect 460759 475523 480503 475601
rect 460667 475499 480503 475523
rect 440367 475487 460112 475493
rect 420129 475481 440107 475482
rect 420129 475458 439798 475481
rect 400445 475016 419546 475452
rect 420619 475016 439798 475458
rect 440819 475016 460112 475487
rect 461175 475491 480503 475499
rect 480569 475491 480589 475601
rect 461175 475471 480589 475491
rect 480849 475619 500577 475637
rect 480849 475611 500491 475619
rect 480849 475501 480875 475611
rect 480941 475509 500491 475611
rect 500557 475509 500577 475619
rect 480941 475501 500577 475509
rect 480849 475489 500577 475501
rect 500837 475629 501707 475655
rect 500837 475519 500863 475629
rect 500929 475519 501707 475629
rect 500837 475495 501707 475519
rect 480849 475477 500345 475489
rect 461175 475016 480245 475471
rect 481410 475016 500345 475477
rect 373156 475011 374154 475016
rect 501434 475012 501707 475495
rect 502705 476009 502711 476010
rect 502705 475012 502806 476009
rect 501434 475009 502806 475012
rect 508574 475011 508580 476011
rect 509580 476010 515574 476011
rect 509580 475012 514575 476010
rect 515573 475012 515579 476010
rect 509580 475011 515574 475012
rect 521042 475011 521048 476011
rect 522048 475539 522668 476011
rect 523746 476010 528122 476011
rect 522048 475492 523046 475539
rect 523746 475526 527123 476010
rect 522048 475382 522941 475492
rect 523007 475382 523046 475492
rect 522048 475346 523046 475382
rect 523283 475482 527123 475526
rect 523283 475372 523313 475482
rect 523379 475372 527123 475482
rect 522048 475011 522668 475346
rect 523283 475333 527123 475372
rect 523746 475012 527123 475333
rect 528121 475012 528127 476010
rect 536254 476009 545594 476016
rect 523746 475011 528122 475012
rect 533870 475009 533876 476009
rect 534876 475571 545594 476009
rect 534876 475528 545972 475571
rect 546727 475552 549890 476016
rect 534876 475418 545855 475528
rect 545921 475418 545972 475528
rect 534876 475371 545972 475418
rect 546202 475518 549890 475552
rect 546202 475408 546227 475518
rect 546293 475408 549890 475518
rect 534876 475016 545594 475371
rect 546202 475367 549890 475408
rect 546727 475016 549890 475367
rect 550890 475016 550896 476016
rect 534876 475009 536526 475016
rect 497347 473194 497985 473199
rect 497347 473189 497352 473194
rect 497980 473189 497985 473194
rect 380552 473159 380562 473164
rect 352770 472434 352776 472986
rect 353318 472981 353328 472986
rect 353323 472439 353328 472981
rect 380552 472617 380557 473159
rect 380552 472612 380562 472617
rect 381104 472612 381110 473164
rect 394692 473157 395244 473162
rect 394692 473152 394697 473157
rect 395239 473152 395244 473157
rect 389486 473083 390038 473088
rect 389486 473078 389491 473083
rect 390033 473078 390038 473083
rect 428290 473114 428842 473120
rect 394692 472604 395244 472610
rect 400586 473109 401138 473114
rect 400586 473104 400591 473109
rect 401133 473104 401138 473109
rect 485292 473103 485904 473108
rect 485292 473098 485297 473103
rect 485899 473098 485904 473103
rect 462130 473059 462742 473064
rect 428290 472567 428295 472572
rect 428837 472567 428842 472572
rect 428290 472562 428842 472567
rect 445478 473052 446090 473058
rect 400586 472556 401138 472562
rect 389486 472530 390038 472536
rect 445478 472445 445483 472450
rect 446085 472445 446090 472450
rect 462130 473054 462135 473059
rect 462737 473054 462742 473059
rect 536938 473163 536948 473168
rect 522934 473097 525137 473102
rect 497347 472555 497985 472561
rect 503855 472998 504493 473003
rect 503855 472993 503860 472998
rect 504488 472993 504493 472998
rect 485292 472490 485904 472496
rect 462130 472446 462742 472452
rect 445478 472440 446090 472445
rect 353318 472434 353328 472439
rect 506684 472394 506690 473006
rect 507292 473001 507302 473006
rect 507297 472399 507302 473001
rect 518224 472480 518230 473092
rect 518832 473087 518842 473092
rect 518837 472485 518842 473087
rect 522934 472495 522944 473097
rect 525127 472495 525137 473097
rect 536938 472561 536943 473163
rect 536938 472556 536948 472561
rect 537550 472556 537556 473168
rect 537952 473141 537962 473146
rect 537952 472511 537957 473141
rect 537952 472506 537962 472511
rect 538592 472506 538598 473146
rect 548142 472572 548148 473212
rect 548778 473207 548788 473212
rect 548783 472577 548788 473207
rect 548778 472572 548788 472577
rect 553158 473131 553168 473136
rect 553158 472501 553163 473131
rect 553158 472496 553168 472501
rect 553798 472496 553804 473136
rect 562798 473064 563438 473070
rect 522934 472490 525137 472495
rect 518832 472480 518842 472485
rect 562798 472429 562803 472434
rect 563433 472429 563438 472434
rect 562798 472424 563438 472429
rect 507292 472394 507302 472399
rect 503855 472359 504493 472365
rect 387909 469789 388029 469799
rect 392801 469789 392921 469799
rect 387904 469723 387914 469789
rect 388024 469723 388034 469789
rect 392796 469723 392806 469789
rect 392916 469723 392926 469789
rect 387909 469713 388029 469723
rect 392801 469713 392921 469723
rect 387919 469417 388039 469427
rect 392811 469417 392931 469427
rect 387914 469351 387924 469417
rect 388034 469351 388044 469417
rect 392806 469351 392816 469417
rect 392926 469351 392936 469417
rect 387919 469341 388039 469351
rect 392811 469341 392931 469351
rect 508966 469089 509096 469094
rect 508966 469023 508976 469089
rect 509086 469023 509096 469089
rect 508966 469018 509096 469023
rect 508976 468717 509106 468722
rect 508976 468651 508986 468717
rect 509096 468651 509106 468717
rect 508976 468646 509106 468651
rect -800 468308 480 468420
rect 515013 467831 515143 467836
rect 515013 467765 515023 467831
rect 515133 467765 515143 467831
rect 515013 467760 515143 467765
rect 515023 467459 515153 467464
rect 515023 467393 515033 467459
rect 515143 467393 515153 467459
rect 515023 467388 515153 467393
rect -800 467126 480 467238
rect 534376 467011 534506 467016
rect 534376 466945 534386 467011
rect 534496 466945 534506 467011
rect 534376 466940 534506 466945
rect 534366 466639 534496 466644
rect 534366 466573 534376 466639
rect 534486 466573 534496 466639
rect 534366 466568 534496 466573
rect -800 465944 480 466056
rect 78270 465202 79268 465207
rect 15018 465201 79269 465202
rect -800 464762 480 464874
rect 15018 464769 78270 465201
rect 13362 464768 78270 464769
rect 13357 464658 13363 464768
rect 13473 464658 78270 464768
rect 13362 464657 78270 464658
rect 15018 464203 78270 464657
rect 79268 464203 79269 465201
rect 15018 464202 79269 464203
rect 78270 464197 79268 464202
rect 13362 463692 13474 463698
rect -800 463580 13362 463692
rect 13362 463574 13474 463580
rect 25407 462510 25519 462516
rect -800 462398 25407 462510
rect 25407 462392 25519 462398
rect 356021 462238 356141 462248
rect 356016 462172 356026 462238
rect 356136 462172 356146 462238
rect 356021 462162 356141 462172
rect 356031 461866 356151 461876
rect 356026 461800 356036 461866
rect 356146 461800 356156 461866
rect 356031 461790 356151 461800
rect 550360 459731 550490 459736
rect 550360 459665 550370 459731
rect 550480 459665 550490 459731
rect 550360 459660 550490 459665
rect 527521 459602 527651 459607
rect 527521 459536 527531 459602
rect 527641 459536 527651 459602
rect 527521 459531 527651 459536
rect 240180 457761 241180 459480
rect 550350 459359 550480 459364
rect 550350 459293 550360 459359
rect 550470 459293 550480 459359
rect 550350 459288 550480 459293
rect 527511 459230 527641 459235
rect 240180 456755 241180 456761
rect 250981 457761 251981 459175
rect 527511 459164 527521 459230
rect 527631 459164 527641 459230
rect 527511 459159 527641 459164
rect 521404 457164 521534 457169
rect 521404 457098 521414 457164
rect 521524 457098 521534 457164
rect 521404 457093 521534 457098
rect 346991 457064 347111 457074
rect 346986 456998 346996 457064
rect 347106 456998 347116 457064
rect 346991 456988 347111 456998
rect 250981 456755 251981 456761
rect 521414 456792 521544 456797
rect 521414 456726 521424 456792
rect 521534 456726 521544 456792
rect 521414 456721 521544 456726
rect 347001 456692 347121 456702
rect 346996 456626 347006 456692
rect 347116 456626 347126 456692
rect 347001 456616 347121 456626
rect 240696 455915 240816 455925
rect 240691 455849 240701 455915
rect 240811 455849 240821 455915
rect 251418 455893 251538 455903
rect 240696 455839 240816 455849
rect 251413 455827 251423 455893
rect 251533 455827 251543 455893
rect 251418 455817 251538 455827
rect 560008 455740 560120 455746
rect 560120 455628 584800 455740
rect 560008 455622 560120 455628
rect 240706 455543 240826 455553
rect 240701 455477 240711 455543
rect 240821 455477 240831 455543
rect 251428 455521 251548 455531
rect 240706 455467 240826 455477
rect 251423 455455 251433 455521
rect 251543 455455 251553 455521
rect 251428 455445 251548 455455
rect 502190 455237 502320 455242
rect 502190 455171 502200 455237
rect 502310 455171 502320 455237
rect 502190 455166 502320 455171
rect 502200 454865 502330 454870
rect 502200 454799 502210 454865
rect 502320 454799 502330 454865
rect 502200 454794 502330 454799
rect 583520 454446 584800 454558
rect 549890 453859 563921 453860
rect 549885 452861 549891 453859
rect 550889 453426 563921 453859
rect 565046 453433 578427 453860
rect 550889 453395 564260 453426
rect 550889 453285 564164 453395
rect 564230 453285 564260 453395
rect 550889 453253 564260 453285
rect 564499 453405 578427 453433
rect 564499 453295 564536 453405
rect 564602 453376 578427 453405
rect 564602 453295 584800 453376
rect 564499 453264 584800 453295
rect 564499 453260 578427 453264
rect 550889 452861 563921 453253
rect 549890 452860 563921 452861
rect 565046 452860 578427 453260
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 508954 449038 509084 449043
rect 508954 448972 508964 449038
rect 509074 448972 509084 449038
rect 508954 448967 509084 448972
rect 392791 448837 392911 448847
rect 387870 448769 387990 448779
rect 392786 448771 392796 448837
rect 392906 448771 392916 448837
rect 387865 448703 387875 448769
rect 387985 448703 387995 448769
rect 392791 448761 392911 448771
rect 387870 448693 387990 448703
rect 508964 448666 509094 448671
rect 508964 448600 508974 448666
rect 509084 448600 509094 448666
rect 508964 448595 509094 448600
rect 392801 448465 392921 448475
rect 387880 448397 388000 448407
rect 392796 448399 392806 448465
rect 392916 448399 392926 448465
rect 387875 448331 387885 448397
rect 387995 448331 388005 448397
rect 392801 448389 392921 448399
rect 387880 448321 388000 448331
rect 515050 447630 515180 447635
rect 515050 447564 515060 447630
rect 515170 447564 515180 447630
rect 515050 447559 515180 447564
rect 515060 447258 515190 447263
rect 515060 447192 515070 447258
rect 515180 447192 515190 447258
rect 515060 447187 515190 447192
rect 534366 446611 534496 446616
rect 534366 446545 534376 446611
rect 534486 446545 534496 446611
rect 534366 446540 534496 446545
rect 534356 446239 534486 446244
rect 534356 446173 534366 446239
rect 534476 446173 534486 446239
rect 534356 446168 534486 446173
rect 514574 445641 515574 445647
rect 501706 445561 502706 445567
rect 508581 445561 509579 445566
rect 502706 445560 509580 445561
rect 502706 444562 508581 445560
rect 509579 444562 509580 445560
rect 515574 445640 522048 445641
rect 515574 444642 521049 445640
rect 522047 444642 522053 445640
rect 527116 444721 527122 445721
rect 528122 445720 534876 445721
rect 528122 444722 533877 445720
rect 534875 444722 534881 445720
rect 528122 444721 534876 444722
rect 515574 444641 522048 444642
rect 514574 444635 515574 444641
rect 502706 444561 509580 444562
rect 501706 444555 502706 444561
rect 508581 444556 509579 444561
rect 355995 442245 356115 442255
rect 355990 442179 356000 442245
rect 356110 442179 356120 442245
rect 355995 442169 356115 442179
rect 356005 441873 356125 441883
rect 356000 441807 356010 441873
rect 356120 441807 356130 441873
rect 356005 441797 356125 441807
rect 346963 436456 347083 436466
rect 346958 436390 346968 436456
rect 347078 436390 347088 436456
rect 346963 436380 347083 436390
rect 346973 436084 347093 436094
rect 346968 436018 346978 436084
rect 347088 436018 347098 436084
rect 346973 436008 347093 436018
rect 240616 434398 240736 434408
rect 240611 434332 240621 434398
rect 240731 434332 240741 434398
rect 240616 434322 240736 434332
rect 251401 434112 251521 434122
rect 251396 434046 251406 434112
rect 251516 434046 251526 434112
rect 251401 434036 251521 434046
rect 240626 434026 240746 434036
rect 240621 433960 240631 434026
rect 240741 433960 240751 434026
rect 240626 433950 240746 433960
rect 251411 433740 251531 433750
rect 251406 433674 251416 433740
rect 251526 433674 251536 433740
rect 251411 433664 251531 433674
rect 348084 430698 348532 430703
rect 238855 429713 238861 430264
rect 239402 430259 239412 430264
rect 239407 429718 239412 430259
rect 249224 429832 249230 430384
rect 249772 430379 249782 430384
rect 249777 429837 249782 430379
rect 332864 430376 333416 430382
rect 249772 429832 249782 429837
rect 252975 430368 253527 430374
rect 252975 429821 252980 429826
rect 253522 429821 253527 429826
rect 252975 429816 253527 429821
rect 258333 430362 258343 430367
rect 258333 429822 258338 430362
rect 258333 429817 258343 429822
rect 258883 429817 258889 430367
rect 293209 430355 293219 430360
rect 278445 430343 278455 430348
rect 272935 430299 273487 430304
rect 272935 430294 272940 430299
rect 273482 430294 273487 430299
rect 278445 429801 278450 430343
rect 278445 429796 278455 429801
rect 278997 429796 279003 430348
rect 293209 429813 293214 430355
rect 293209 429808 293219 429813
rect 293761 429808 293767 430360
rect 299157 430255 299167 430260
rect 272935 429746 273487 429752
rect 239402 429713 239412 429718
rect 299157 429713 299162 430255
rect 299157 429708 299167 429713
rect 299709 429708 299715 430260
rect 322080 430215 322090 430220
rect 313343 430196 313895 430202
rect 313343 429649 313348 429654
rect 313890 429649 313895 429654
rect 313343 429644 313895 429649
rect 319471 430157 319481 430162
rect 319471 429615 319476 430157
rect 319471 429610 319481 429615
rect 320023 429610 320029 430162
rect 322080 429673 322085 430215
rect 322080 429668 322090 429673
rect 322632 429668 322638 430220
rect 332864 429829 332869 429834
rect 333411 429829 333416 429834
rect 332864 429824 333416 429829
rect 335389 430253 335399 430258
rect 335389 429711 335394 430253
rect 335389 429706 335399 429711
rect 335941 429706 335947 430258
rect 348084 429382 348094 430698
rect 348522 429382 348532 430698
rect 359996 430444 360548 430450
rect 354352 430269 354904 430274
rect 354352 430264 354357 430269
rect 354899 430264 354904 430269
rect 359996 429897 360001 429902
rect 360543 429897 360548 429902
rect 359996 429892 360548 429897
rect 362166 430443 362718 430448
rect 362166 430438 362171 430443
rect 362713 430438 362718 430443
rect 497205 430403 497843 430409
rect 375347 430200 375899 430206
rect 362166 429890 362718 429896
rect 373945 430191 373955 430196
rect 354352 429716 354904 429722
rect 373945 429649 373950 430191
rect 373945 429644 373955 429649
rect 374497 429644 374503 430196
rect 385922 429740 385928 430292
rect 386470 430287 386480 430292
rect 386475 429745 386480 430287
rect 391194 429824 391200 430376
rect 391742 430371 391752 430376
rect 391747 429829 391752 430371
rect 391742 429824 391752 429829
rect 513062 430340 513674 430346
rect 497205 429770 497210 429775
rect 497838 429770 497843 429775
rect 497205 429765 497843 429770
rect 510278 430290 510890 430296
rect 386470 429740 386480 429745
rect 528954 430329 528964 430334
rect 513062 429733 513067 429738
rect 513669 429733 513674 429738
rect 513062 429728 513674 429733
rect 522300 429694 522306 430306
rect 522908 430301 522918 430306
rect 522913 429699 522918 430301
rect 522908 429694 522918 429699
rect 528954 429699 528959 430329
rect 528954 429694 528964 429699
rect 529594 429694 529600 430334
rect 545772 429768 545778 430408
rect 546408 430403 546418 430408
rect 546413 429773 546418 430403
rect 546408 429768 546418 429773
rect 562796 430329 563436 430334
rect 562796 430324 562801 430329
rect 563431 430324 563436 430329
rect 562796 429688 563436 429694
rect 510278 429683 510283 429688
rect 510885 429683 510890 429688
rect 510278 429678 510890 429683
rect 375347 429653 375352 429658
rect 375894 429653 375899 429658
rect 375347 429648 375899 429653
rect 348084 429377 348532 429382
rect 392823 427745 392943 427755
rect 387899 427726 388019 427736
rect 387894 427660 387904 427726
rect 388014 427660 388024 427726
rect 392818 427679 392828 427745
rect 392938 427679 392948 427745
rect 392823 427669 392943 427679
rect 387899 427650 388019 427660
rect 392833 427373 392953 427383
rect 387909 427354 388029 427364
rect 387904 427288 387914 427354
rect 388024 427288 388034 427354
rect 392828 427307 392838 427373
rect 392948 427307 392958 427373
rect 392833 427297 392953 427307
rect 387909 427278 388029 427288
rect 392312 426639 393310 426644
rect 243838 426633 252655 426639
rect 240180 426632 252655 426633
rect 240175 425634 240181 426632
rect 241179 426126 252655 426632
rect 253865 426191 272666 426639
rect 273694 426225 292901 426639
rect 253865 426152 273003 426191
rect 273694 426186 293284 426225
rect 294000 426215 313058 426639
rect 294000 426214 313433 426215
rect 273694 426180 293185 426186
rect 241179 426087 253057 426126
rect 253865 426115 272904 426152
rect 241179 425977 252958 426087
rect 253024 425977 253057 426087
rect 241179 425955 253057 425977
rect 253298 426077 272904 426115
rect 253298 425967 253330 426077
rect 253396 426042 272904 426077
rect 272970 426042 273003 426152
rect 253396 426020 273003 426042
rect 273244 426142 293185 426180
rect 273244 426032 273276 426142
rect 273342 426076 293185 426142
rect 293251 426076 293284 426186
rect 273342 426054 293284 426076
rect 293525 426176 313433 426214
rect 314235 426204 324048 426639
rect 293525 426066 293557 426176
rect 293623 426066 313334 426176
rect 313400 426066 313433 426176
rect 273342 426032 292901 426054
rect 293525 426044 313433 426066
rect 313674 426166 324048 426204
rect 313674 426056 313706 426166
rect 313772 426056 324048 426166
rect 293525 426043 313058 426044
rect 253396 425967 272666 426020
rect 273244 426009 292901 426032
rect 241179 425639 252655 425955
rect 253298 425944 272666 425967
rect 253865 425639 272666 425944
rect 273694 425639 292901 426009
rect 294000 425639 313058 426043
rect 313674 426033 324048 426056
rect 314235 425639 324048 426033
rect 325048 426189 335115 426639
rect 336297 426200 355101 426639
rect 325048 426151 335639 426189
rect 325048 426041 335541 426151
rect 335607 426041 335639 426151
rect 325048 426018 335639 426041
rect 335880 426185 355101 426200
rect 356268 426279 375002 426639
rect 376360 426638 393311 426639
rect 376360 426290 392312 426638
rect 356268 426241 375592 426279
rect 356268 426196 375494 426241
rect 335880 426161 355629 426185
rect 335880 426051 335913 426161
rect 335979 426147 355629 426161
rect 335979 426051 355531 426147
rect 335880 426037 355531 426051
rect 355597 426037 355629 426147
rect 335880 426029 355629 426037
rect 325048 425639 335115 426018
rect 336297 426014 355629 426029
rect 355870 426157 375494 426196
rect 355870 426047 355903 426157
rect 355969 426131 375494 426157
rect 375560 426131 375592 426241
rect 355969 426108 375592 426131
rect 375833 426251 392312 426290
rect 375833 426141 375866 426251
rect 375932 426141 392312 426251
rect 375833 426119 392312 426141
rect 355969 426047 375002 426108
rect 355870 426025 375002 426047
rect 336297 425639 355101 426014
rect 356268 425639 375002 426025
rect 376360 425640 392312 426119
rect 393310 425640 393311 426638
rect 376360 425639 393311 425640
rect 241179 425634 245025 425639
rect 392312 425634 393310 425639
rect 240180 425633 245025 425634
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect 356000 422291 356120 422301
rect 355995 422225 356005 422291
rect 356115 422225 356125 422291
rect 356000 422215 356120 422225
rect 356010 421919 356130 421929
rect 356005 421853 356015 421919
rect 356125 421853 356135 421919
rect 356010 421843 356130 421853
rect -800 421540 480 421652
rect 250982 421100 251980 421105
rect 336048 421100 337048 421106
rect 250981 421099 258214 421100
rect 72633 420888 73631 420893
rect 15289 420887 73632 420888
rect 15289 420470 72633 420887
rect -800 420358 72633 420470
rect 15289 419889 72633 420358
rect 73631 419889 73632 420887
rect 250981 420101 250982 421099
rect 251980 420616 258214 421099
rect 259016 420657 278312 421100
rect 279172 420658 298996 421100
rect 259016 420623 278551 420657
rect 279172 420639 299228 420658
rect 299829 420641 319274 421100
rect 258652 420622 278551 420623
rect 251980 420589 258401 420616
rect 251980 420479 258312 420589
rect 258378 420479 258401 420589
rect 251980 420446 258401 420479
rect 258652 420579 278446 420622
rect 258652 420469 258684 420579
rect 258750 420512 278446 420579
rect 278512 420512 278551 420622
rect 258750 420476 278551 420512
rect 278784 420628 299228 420639
rect 278784 420612 299123 420628
rect 278784 420502 278818 420612
rect 278884 420518 299123 420612
rect 299189 420518 299228 420628
rect 278884 420502 299228 420518
rect 278784 420496 299228 420502
rect 299461 420629 319274 420641
rect 299461 420618 319562 420629
rect 320171 420620 336048 421100
rect 299461 420508 299495 420618
rect 299561 420580 319562 420618
rect 299561 420508 319451 420580
rect 258750 420469 278312 420476
rect 278784 420474 298996 420496
rect 299461 420479 319451 420508
rect 251980 420101 258214 420446
rect 258652 420437 278312 420469
rect 250981 420100 258214 420101
rect 259016 420100 278312 420437
rect 279172 420100 298996 420474
rect 299829 420470 319451 420479
rect 319517 420470 319562 420580
rect 299829 420422 319562 420470
rect 319786 420570 336048 420620
rect 319786 420460 319823 420570
rect 319889 420460 336048 420570
rect 319786 420424 336048 420460
rect 299829 420100 319274 420422
rect 320171 420100 336048 420424
rect 337048 420607 353468 421100
rect 354379 420675 373820 421100
rect 374735 420698 387417 421100
rect 354379 420649 374195 420675
rect 354379 420625 374104 420649
rect 337048 420579 353853 420607
rect 337048 420469 353761 420579
rect 353827 420469 353853 420579
rect 337048 420427 353853 420469
rect 354085 420589 374104 420625
rect 354085 420479 354133 420589
rect 354199 420539 374104 420589
rect 374170 420539 374195 420649
rect 354199 420516 374195 420539
rect 374450 420659 387417 420698
rect 374450 420549 374476 420659
rect 374542 420549 387417 420659
rect 354199 420479 373820 420516
rect 374450 420513 387417 420549
rect 354085 420435 373820 420479
rect 337048 420100 353468 420427
rect 354379 420100 373820 420435
rect 374735 420100 387417 420513
rect 388417 420100 388423 421100
rect 250982 420095 251980 420100
rect 336048 420094 337048 420100
rect 15289 419888 73632 419889
rect 72633 419883 73631 419888
rect 25438 419288 25550 419294
rect -800 419176 25438 419288
rect 25438 419170 25550 419176
rect 324539 417183 324659 417188
rect 324534 417178 324664 417183
rect 324534 417112 324544 417178
rect 324654 417112 324664 417178
rect 324534 417107 324664 417112
rect 336549 417108 336669 417113
rect 324539 417102 324659 417107
rect 336544 417103 336674 417108
rect 336544 417037 336554 417103
rect 336664 417037 336674 417103
rect 336544 417032 336674 417037
rect 336549 417027 336669 417032
rect 324549 416806 324669 416816
rect 324544 416740 324554 416806
rect 324664 416740 324674 416806
rect 324549 416730 324669 416740
rect 336559 416731 336679 416741
rect 336554 416665 336564 416731
rect 336674 416665 336684 416731
rect 336559 416655 336679 416665
rect 345540 416210 345988 416215
rect 319461 415947 319471 415952
rect 252967 415912 252977 415917
rect 242014 415906 242565 415912
rect 252967 415372 252972 415912
rect 252967 415367 252977 415372
rect 253517 415367 253523 415917
rect 258331 415881 258881 415887
rect 255268 415727 255820 415732
rect 255268 415722 255273 415727
rect 255815 415722 255820 415727
rect 242014 415360 242019 415365
rect 242560 415360 242565 415365
rect 242014 415355 242565 415360
rect 278445 415820 278997 415826
rect 258331 415336 258336 415341
rect 258876 415336 258881 415341
rect 258331 415331 258881 415336
rect 272927 415814 273479 415820
rect 272927 415267 272932 415272
rect 273474 415267 273479 415272
rect 299131 415818 299683 415824
rect 278445 415273 278450 415278
rect 278992 415273 278997 415278
rect 278445 415268 278997 415273
rect 293209 415789 293219 415794
rect 272927 415262 273479 415267
rect 293209 415247 293214 415789
rect 293209 415242 293219 415247
rect 293761 415242 293767 415794
rect 313343 415324 313349 415876
rect 313891 415871 313901 415876
rect 313896 415329 313901 415871
rect 319461 415405 319466 415947
rect 319461 415400 319471 415405
rect 320013 415400 320019 415952
rect 328154 415901 328164 415906
rect 328154 415359 328159 415901
rect 328154 415354 328164 415359
rect 328706 415354 328712 415906
rect 339870 415863 339880 415868
rect 313891 415324 313901 415329
rect 339870 415321 339875 415863
rect 339870 415316 339880 415321
rect 340422 415316 340428 415868
rect 299131 415271 299136 415276
rect 299678 415271 299683 415276
rect 299131 415266 299683 415271
rect 255268 415174 255820 415180
rect 345540 414894 345550 416210
rect 345978 414894 345988 416210
rect 393660 415932 394212 415938
rect 346907 415822 347027 415832
rect 346902 415756 346912 415822
rect 347022 415756 347032 415822
rect 353568 415775 354120 415780
rect 353568 415770 353573 415775
rect 354115 415770 354120 415775
rect 346907 415746 347027 415756
rect 346917 415450 347037 415460
rect 346912 415384 346922 415450
rect 347032 415384 347042 415450
rect 346917 415374 347037 415384
rect 373933 415298 373939 415850
rect 374481 415845 374491 415850
rect 374486 415303 374491 415845
rect 388612 415849 388622 415854
rect 374481 415298 374491 415303
rect 375335 415649 375345 415654
rect 353568 415222 354120 415228
rect 375335 415107 375340 415649
rect 375335 415102 375345 415107
rect 375887 415102 375893 415654
rect 388612 415307 388617 415849
rect 388612 415302 388622 415307
rect 389164 415302 389170 415854
rect 393660 415385 393665 415390
rect 394207 415385 394212 415390
rect 393660 415380 394212 415385
rect 345540 414889 345988 414894
rect 560017 411318 560129 411324
rect 560129 411206 584800 411318
rect 560017 411200 560129 411206
rect 583520 410024 584800 410136
rect 549018 409466 550016 409471
rect 549017 409465 567924 409466
rect 549017 408467 549018 409465
rect 550016 409023 567924 409465
rect 550016 408988 568141 409023
rect 568785 409012 579376 409466
rect 550016 408878 568046 408988
rect 568112 408878 568141 408988
rect 550016 408850 568141 408878
rect 568383 408978 579376 409012
rect 568383 408868 568418 408978
rect 568484 408954 579376 408978
rect 568484 408868 584800 408954
rect 550016 408467 567924 408850
rect 568383 408842 584800 408868
rect 568383 408832 579376 408842
rect 568384 408831 568498 408832
rect 549017 408466 567924 408467
rect 568785 408466 579376 408832
rect 549018 408461 550016 408466
rect 583520 407660 584800 407772
rect 549540 407196 549675 407209
rect 549519 407130 549553 407196
rect 549663 407130 549699 407196
rect 549519 407096 549699 407130
rect 549519 406824 549681 406849
rect 549519 406758 549543 406824
rect 549653 406758 549681 406824
rect 549533 406753 549663 406758
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 355989 402256 356109 402266
rect 355984 402190 355994 402256
rect 356104 402190 356114 402256
rect 355989 402180 356109 402190
rect 355999 401884 356119 401894
rect 355994 401818 356004 401884
rect 356114 401818 356124 401884
rect 355999 401808 356119 401818
rect 336574 396455 336694 396460
rect 336569 396450 336699 396455
rect 324537 396393 324657 396398
rect 324532 396388 324662 396393
rect 324532 396322 324542 396388
rect 324652 396322 324662 396388
rect 336569 396384 336579 396450
rect 336689 396384 336699 396450
rect 336569 396379 336699 396384
rect 336574 396374 336694 396379
rect 324532 396317 324662 396322
rect 324537 396312 324657 396317
rect 336584 396078 336704 396088
rect 324547 396016 324667 396026
rect 324542 395950 324552 396016
rect 324662 395950 324672 396016
rect 336579 396012 336589 396078
rect 336699 396012 336709 396078
rect 336584 396002 336704 396012
rect 324547 395940 324667 395950
rect 346935 395144 347055 395154
rect 346930 395078 346940 395144
rect 347050 395078 347060 395144
rect 346935 395068 347055 395078
rect 346945 394772 347065 394782
rect 346940 394706 346950 394772
rect 347060 394706 347070 394772
rect 346945 394696 347065 394706
rect 322884 390800 322890 391352
rect 323432 391347 323442 391352
rect 323437 390805 323442 391347
rect 333081 390820 333087 391372
rect 333629 391367 333639 391372
rect 333634 390825 333639 391367
rect 333629 390820 333639 390825
rect 323432 390800 323442 390805
rect 334868 390762 334874 391314
rect 335416 391309 335426 391314
rect 335421 390767 335426 391309
rect 428496 391302 429048 391308
rect 367479 391193 367489 391198
rect 357685 391157 357695 391162
rect 335416 390762 335426 390767
rect 353560 390944 354112 390950
rect 118329 390495 123445 390500
rect 118328 390494 168402 390495
rect 118328 385378 118329 390494
rect 123445 385378 168402 390494
rect 357685 390615 357690 391157
rect 357685 390610 357695 390615
rect 358237 390610 358243 391162
rect 367479 390651 367484 391193
rect 367479 390646 367489 390651
rect 368031 390646 368037 391198
rect 385258 390622 385264 391174
rect 385806 391169 385816 391174
rect 385811 390627 385816 391169
rect 400426 390642 400432 391194
rect 400974 391189 400984 391194
rect 400979 390647 400984 391189
rect 530380 391147 530390 391152
rect 490264 391105 490274 391110
rect 470022 391055 470032 391060
rect 428496 390755 428501 390760
rect 429043 390755 429048 390760
rect 428496 390750 429048 390755
rect 446390 391049 446400 391054
rect 400974 390642 400984 390647
rect 385806 390622 385816 390627
rect 446390 390507 446395 391049
rect 446390 390502 446400 390507
rect 446942 390502 446948 391054
rect 470022 390513 470027 391055
rect 470022 390508 470032 390513
rect 470574 390508 470580 391060
rect 490264 390563 490269 391105
rect 490264 390558 490274 390563
rect 490816 390558 490822 391110
rect 510718 391075 510728 391080
rect 510718 390533 510723 391075
rect 510718 390528 510728 390533
rect 511270 390528 511276 391080
rect 530380 390605 530385 391147
rect 530380 390600 530390 390605
rect 530932 390600 530938 391152
rect 546392 390674 546398 391246
rect 546960 391241 546970 391246
rect 546965 390679 546970 391241
rect 546960 390674 546970 390679
rect 571222 391205 571232 391210
rect 571222 390643 571227 391205
rect 571222 390638 571232 390643
rect 571794 390638 571800 391210
rect 353560 390397 353565 390402
rect 354107 390397 354112 390402
rect 353560 390392 354112 390397
rect 549557 388152 549692 388169
rect 549536 388086 549570 388152
rect 549680 388086 549716 388152
rect 549536 388052 549716 388086
rect 549536 387780 549698 387805
rect 549536 387714 549560 387780
rect 549670 387714 549698 387780
rect 549550 387709 549680 387714
rect 336049 387271 337047 387276
rect 548986 387271 550037 387302
rect 336048 387270 347327 387271
rect 336048 386272 336049 387270
rect 337047 386748 347327 387270
rect 348153 386777 367375 387271
rect 368146 386777 387149 387271
rect 348153 386753 367553 386777
rect 348153 386748 367462 386753
rect 337047 386724 347537 386748
rect 337047 386614 347446 386724
rect 347512 386614 347537 386724
rect 337047 386586 347537 386614
rect 347784 386714 367462 386748
rect 347784 386604 347818 386714
rect 347884 386643 367462 386714
rect 367528 386643 367553 386753
rect 347884 386615 367553 386643
rect 367800 386767 387149 386777
rect 387979 386767 407371 387271
rect 367800 386743 387365 386767
rect 367800 386633 367834 386743
rect 367900 386633 387274 386743
rect 387340 386633 387365 386743
rect 347884 386604 367375 386615
rect 337047 386272 347327 386586
rect 347784 386568 367375 386604
rect 367800 386605 387365 386633
rect 387612 386765 407371 386767
rect 408304 386820 427584 387271
rect 428599 386820 447787 387271
rect 408304 386796 427900 386820
rect 408304 386765 427809 386796
rect 387612 386741 407624 386765
rect 387612 386733 407533 386741
rect 387612 386623 387646 386733
rect 387712 386631 407533 386733
rect 407599 386631 407624 386741
rect 387712 386623 407624 386631
rect 367800 386597 387149 386605
rect 336048 386271 347327 386272
rect 348153 386271 367375 386568
rect 368146 386271 387149 386597
rect 387612 386603 407624 386623
rect 407871 386731 427809 386765
rect 407871 386621 407905 386731
rect 407971 386686 427809 386731
rect 427875 386686 427900 386796
rect 407971 386658 427900 386686
rect 428147 386800 447787 386820
rect 448703 386800 467834 387271
rect 428147 386786 448059 386800
rect 428147 386676 428181 386786
rect 428247 386776 448059 386786
rect 428247 386676 447968 386776
rect 428147 386666 447968 386676
rect 448034 386666 448059 386776
rect 407971 386621 427584 386658
rect 428147 386640 448059 386666
rect 387612 386587 407371 386603
rect 387979 386271 407371 386587
rect 407871 386585 427584 386621
rect 408304 386271 427584 386585
rect 428599 386638 448059 386640
rect 448306 386795 467834 386800
rect 468687 386795 487823 387271
rect 448306 386771 468061 386795
rect 448306 386766 467970 386771
rect 448306 386656 448340 386766
rect 448406 386661 467970 386766
rect 468036 386661 468061 386771
rect 448406 386656 468061 386661
rect 428599 386271 447787 386638
rect 448306 386633 468061 386656
rect 468308 386779 487823 386795
rect 488884 386802 508078 387271
rect 508976 386816 528135 387271
rect 529141 386816 549017 387271
rect 508976 386802 528418 386816
rect 488884 386779 508309 386802
rect 468308 386761 488179 386779
rect 468308 386651 468342 386761
rect 468408 386755 488179 386761
rect 468408 386651 488088 386755
rect 468308 386645 488088 386651
rect 488154 386645 488179 386755
rect 448306 386620 467834 386633
rect 448703 386271 467834 386620
rect 468308 386617 488179 386645
rect 488426 386778 508309 386779
rect 488426 386745 508218 386778
rect 488426 386635 488460 386745
rect 488526 386668 508218 386745
rect 508284 386668 508309 386778
rect 488526 386640 508309 386668
rect 508556 386792 528418 386802
rect 508556 386768 528327 386792
rect 508556 386658 508590 386768
rect 508656 386682 528327 386768
rect 528393 386682 528418 386792
rect 508656 386658 528418 386682
rect 508556 386654 528418 386658
rect 528665 386782 549017 386816
rect 528665 386672 528699 386782
rect 528765 386672 549017 386782
rect 488526 386635 508078 386640
rect 468308 386616 488049 386617
rect 468308 386615 487823 386616
rect 468687 386271 487823 386615
rect 488426 386599 508078 386635
rect 508556 386622 528135 386654
rect 528665 386636 549017 386672
rect 488884 386271 508078 386599
rect 508976 386271 528135 386622
rect 529141 386271 549017 386636
rect 550017 386271 550037 387271
rect 336049 386266 337047 386271
rect 548986 386232 550037 386271
rect 118328 385377 168402 385378
rect 118329 385372 123445 385377
rect 355969 382192 356089 382202
rect 355964 382126 355974 382192
rect 356084 382126 356094 382192
rect 355969 382116 356089 382126
rect -800 381864 480 381976
rect 355979 381820 356099 381830
rect 355974 381754 355984 381820
rect 356094 381754 356104 381820
rect 355979 381744 356099 381754
rect 324048 381237 332767 381238
rect -800 380682 480 380794
rect 324043 380239 324049 381237
rect 325047 380796 332767 381237
rect 333959 380804 357388 381238
rect 325047 380757 333181 380796
rect 333959 380780 357760 380804
rect 358442 380788 386717 381238
rect 325047 380647 333077 380757
rect 333143 380647 333181 380757
rect 325047 380617 333181 380647
rect 333412 380765 357760 380780
rect 333412 380747 357656 380765
rect 333412 380637 333449 380747
rect 333515 380655 357656 380747
rect 357722 380655 357760 380765
rect 333515 380637 357760 380655
rect 333412 380625 357760 380637
rect 357991 380762 386717 380788
rect 388038 380793 407436 381238
rect 357991 380755 387207 380762
rect 357991 380645 358028 380755
rect 358094 380723 387207 380755
rect 388038 380754 407785 380793
rect 408573 380777 427215 381238
rect 388038 380746 407681 380754
rect 358094 380645 387103 380723
rect 325047 380239 332767 380617
rect 333412 380600 357388 380625
rect 357991 380613 387103 380645
rect 387169 380613 387207 380723
rect 357991 380608 387207 380613
rect 324048 380238 332767 380239
rect 333959 380238 357388 380600
rect 358442 380583 387207 380608
rect 387438 380713 407681 380746
rect 387438 380603 387475 380713
rect 387541 380644 407681 380713
rect 407747 380644 407785 380754
rect 387541 380614 407785 380644
rect 408016 380768 427215 380777
rect 428579 380772 447608 381238
rect 448683 380839 467673 381238
rect 448683 380800 467989 380839
rect 468673 380823 488071 381238
rect 408016 380744 427759 380768
rect 428579 380752 448005 380772
rect 448683 380756 467885 380800
rect 408016 380634 408053 380744
rect 408119 380729 427759 380744
rect 408119 380634 427655 380729
rect 408016 380619 427655 380634
rect 427721 380619 427759 380729
rect 387541 380603 407436 380614
rect 358442 380238 386717 380583
rect 387438 380566 407436 380603
rect 408016 380597 427759 380619
rect 388038 380238 407436 380566
rect 408573 380589 427759 380597
rect 427990 380733 448005 380752
rect 427990 380719 447901 380733
rect 427990 380609 428027 380719
rect 428093 380623 447901 380719
rect 447967 380623 448005 380733
rect 428093 380609 448005 380623
rect 427990 380593 448005 380609
rect 448236 380723 467885 380756
rect 448236 380613 448273 380723
rect 448339 380690 467885 380723
rect 467951 380690 467989 380800
rect 448339 380660 467989 380690
rect 468220 380790 488071 380823
rect 468220 380680 468257 380790
rect 468323 380764 488071 380790
rect 489149 380836 507741 381238
rect 489149 380797 508087 380836
rect 508805 380820 528066 381238
rect 468323 380725 488404 380764
rect 489149 380748 507983 380797
rect 468323 380680 488300 380725
rect 448339 380613 467673 380660
rect 468220 380643 488300 380680
rect 408573 380238 427215 380589
rect 427990 380572 447608 380593
rect 448236 380576 467673 380613
rect 428579 380238 447608 380572
rect 448683 380238 467673 380576
rect 468673 380615 488300 380643
rect 488366 380615 488404 380725
rect 468673 380585 488404 380615
rect 488635 380715 507983 380748
rect 488635 380605 488672 380715
rect 488738 380687 507983 380715
rect 508049 380687 508087 380797
rect 488738 380657 508087 380687
rect 508318 380787 528066 380820
rect 508318 380677 508355 380787
rect 508421 380770 528066 380787
rect 508421 380731 528457 380770
rect 529196 380754 548896 381238
rect 508421 380677 528353 380731
rect 488738 380605 507741 380657
rect 508318 380640 528353 380677
rect 468673 380238 488071 380585
rect 488635 380568 507741 380605
rect 489149 380238 507741 380568
rect 508805 380621 528353 380640
rect 528419 380621 528457 380731
rect 508805 380591 528457 380621
rect 528688 380721 548896 380754
rect 528688 380611 528725 380721
rect 528791 380611 548896 380721
rect 508805 380238 528066 380591
rect 528688 380574 548896 380611
rect 529196 380238 548896 380574
rect 549896 380238 550017 381238
rect -800 379500 480 379612
rect 549358 379494 549488 379499
rect 549358 379428 549368 379494
rect 549478 379428 549488 379494
rect 549358 379423 549488 379428
rect 549368 379122 549498 379127
rect 549368 379056 549378 379122
rect 549488 379056 549498 379122
rect 549368 379051 549498 379056
rect 65787 378990 66785 378995
rect 14217 378989 66786 378990
rect 12758 378524 12868 378529
rect 14217 378524 65787 378989
rect 12757 378523 65787 378524
rect -800 378318 480 378430
rect 12757 378413 12758 378523
rect 12868 378413 65787 378523
rect 12757 378412 65787 378413
rect 12758 378407 12868 378412
rect 14217 377991 65787 378412
rect 66785 377991 66786 378989
rect 14217 377990 66786 377991
rect 65787 377985 66785 377990
rect 12757 377248 12869 377254
rect -800 377136 12757 377248
rect 12757 377130 12869 377136
rect 352320 376280 353848 376285
rect 333085 376214 333637 376220
rect 325760 376095 325770 376100
rect -800 375954 25430 376066
rect 25542 375954 25548 376066
rect 325760 375553 325765 376095
rect 325760 375548 325770 375553
rect 326312 375548 326318 376100
rect 333085 375667 333090 375672
rect 333632 375667 333637 375672
rect 333085 375662 333637 375667
rect 337328 376115 337880 376120
rect 337328 376110 337333 376115
rect 337875 376110 337880 376115
rect 337328 375562 337880 375568
rect 345676 376094 346228 376100
rect 352320 375608 352330 376280
rect 353838 375608 353848 376280
rect 526300 376169 526310 376174
rect 352320 375603 353848 375608
rect 357679 376101 357689 376106
rect 357679 375559 357684 376101
rect 357679 375554 357689 375559
rect 358231 375554 358237 376106
rect 367479 376051 367489 376056
rect 345676 375547 345681 375552
rect 346223 375547 346228 375552
rect 345676 375542 346228 375547
rect 367479 375509 367484 376051
rect 367479 375504 367489 375509
rect 368031 375504 368037 376056
rect 388554 375919 388564 375924
rect 388554 375377 388559 375919
rect 388554 375372 388564 375377
rect 389106 375372 389112 375924
rect 400414 375554 400420 376106
rect 400962 376101 400972 376106
rect 400967 375559 400972 376101
rect 400962 375554 400972 375559
rect 429144 376007 429154 376012
rect 429144 375465 429149 376007
rect 429144 375460 429154 375465
rect 429696 375460 429702 376012
rect 446400 375518 446406 376070
rect 446948 376065 446958 376070
rect 446953 375523 446958 376065
rect 446948 375518 446958 375523
rect 466538 375502 466544 376054
rect 467086 376049 467096 376054
rect 467091 375507 467096 376049
rect 467086 375502 467096 375507
rect 485498 375458 485504 376010
rect 486046 376005 486056 376010
rect 486051 375463 486056 376005
rect 486046 375458 486056 375463
rect 505728 375989 505738 375994
rect 505728 375447 505733 375989
rect 505728 375442 505738 375447
rect 506280 375442 506286 375994
rect 526300 375627 526305 376169
rect 526300 375622 526310 375627
rect 526852 375622 526858 376174
rect 562704 376121 563276 376126
rect 562704 376116 562709 376121
rect 563271 376116 563276 376121
rect 552356 376047 552366 376052
rect 552356 375485 552361 376047
rect 552356 375480 552366 375485
rect 552928 375480 552934 376052
rect 562704 375548 563276 375554
rect 118329 374081 123445 374086
rect 118328 374080 168402 374081
rect 118328 368964 118329 374080
rect 123445 368964 168402 374080
rect 346921 373862 347041 373872
rect 346916 373796 346926 373862
rect 347036 373796 347046 373862
rect 346921 373786 347041 373796
rect 346931 373490 347051 373500
rect 346926 373424 346936 373490
rect 347046 373424 347056 373490
rect 346931 373414 347051 373424
rect 118328 368963 168402 368964
rect 118329 368958 123445 368963
rect 560038 364896 560150 364902
rect 560150 364784 584800 364896
rect 560038 364778 560150 364784
rect 549319 364308 549449 364313
rect 549319 364242 549329 364308
rect 549439 364242 549449 364308
rect 549319 364237 549449 364242
rect 549329 363936 549459 363941
rect 549329 363870 549339 363936
rect 549449 363870 549459 363936
rect 549329 363865 549459 363870
rect 583520 363602 584800 363714
rect 548897 363047 549895 363052
rect 548896 363046 567863 363047
rect 356026 362209 356146 362219
rect 356021 362143 356031 362209
rect 356141 362143 356151 362209
rect 356026 362133 356146 362143
rect 548896 362048 548897 363046
rect 549895 362644 567863 363046
rect 549895 362605 568306 362644
rect 569114 362628 578945 363047
rect 549895 362495 568202 362605
rect 568268 362495 568306 362605
rect 549895 362465 568306 362495
rect 568537 362595 578945 362628
rect 568537 362485 568574 362595
rect 568640 362532 578945 362595
rect 568640 362485 584800 362532
rect 549895 362048 567863 362465
rect 568537 362448 584800 362485
rect 548896 362047 567863 362048
rect 569114 362420 584800 362448
rect 569114 362047 578945 362420
rect 548897 362042 549895 362047
rect 356036 361837 356156 361847
rect 356031 361771 356041 361837
rect 356151 361771 356161 361837
rect 356036 361761 356156 361771
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 118329 359181 123445 359186
rect 118328 359180 168402 359181
rect 118328 354064 118329 359180
rect 123445 354064 168402 359180
rect 583520 358874 584800 358986
rect 118328 354063 168402 354064
rect 118329 354058 123445 354063
rect 346921 353012 347041 353022
rect 346916 352946 346926 353012
rect 347036 352946 347046 353012
rect 346921 352936 347041 352946
rect 346931 352640 347051 352650
rect 346926 352574 346936 352640
rect 347046 352574 347056 352640
rect 346931 352564 347051 352574
rect 356026 342206 356146 342216
rect 356021 342140 356031 342206
rect 356141 342140 356151 342206
rect 356026 342130 356146 342140
rect 356036 341834 356156 341844
rect 356031 341768 356041 341834
rect 356151 341768 356161 341834
rect 356036 341758 356156 341768
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect 14352 335076 59670 335077
rect 14352 334684 58671 335076
rect 13037 334683 58671 334684
rect 13032 334573 13038 334683
rect 13148 334573 58671 334683
rect 13037 334572 58671 334573
rect 14352 334078 58671 334572
rect 59669 334078 59675 335076
rect 14352 334077 59670 334078
rect 13037 334026 13149 334032
rect -800 333914 13037 334026
rect 13037 333908 13149 333914
rect 25372 332844 25484 332850
rect -800 332732 25372 332844
rect 25484 332734 25490 332844
rect 25372 332726 25484 332732
rect 347005 332416 347125 332426
rect 347000 332350 347010 332416
rect 347120 332350 347130 332416
rect 347005 332340 347125 332350
rect 347015 332044 347135 332054
rect 347010 331978 347020 332044
rect 347130 331978 347140 332044
rect 347015 331968 347135 331978
rect 118329 323859 123445 323864
rect 118328 323858 168402 323859
rect 118328 318742 118329 323858
rect 123445 318742 168402 323858
rect 355950 322204 356070 322214
rect 355945 322138 355955 322204
rect 356065 322138 356075 322204
rect 355950 322128 356070 322138
rect 355960 321832 356080 321842
rect 355955 321766 355965 321832
rect 356075 321766 356085 321832
rect 355960 321756 356080 321766
rect 565606 319674 565718 319680
rect 565718 319562 584800 319674
rect 565606 319556 565718 319562
rect 118328 318741 168402 318742
rect 118329 318736 123445 318741
rect 578500 318380 584800 318492
rect 365529 317851 366527 317856
rect 365528 317850 576625 317851
rect 365528 316852 365529 317850
rect 366527 317496 576625 317850
rect 578500 317496 578612 318380
rect 366527 317384 578612 317496
rect 366527 316852 576625 317384
rect 583520 317198 584800 317310
rect 365528 316851 576625 316852
rect 365529 316846 366527 316851
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 346977 310548 347097 310558
rect 346972 310482 346982 310548
rect 347092 310482 347102 310548
rect 346977 310472 347097 310482
rect 346987 310176 347107 310186
rect 346982 310110 346992 310176
rect 347102 310110 347112 310176
rect 118329 310099 123445 310104
rect 346987 310100 347107 310110
rect 118328 310098 168402 310099
rect 118328 304982 118329 310098
rect 123445 304982 168402 310098
rect 348014 307618 348486 307623
rect 348014 305644 348024 307618
rect 348476 305644 348486 307618
rect 490709 307004 490719 307009
rect 390695 306940 391254 306945
rect 390695 306935 390700 306940
rect 391249 306935 391254 306940
rect 370683 306812 371242 306817
rect 370683 306807 370688 306812
rect 371237 306807 371242 306812
rect 357940 306784 358492 306790
rect 390695 306380 391254 306386
rect 400259 306898 400818 306903
rect 400259 306893 400264 306898
rect 400813 306893 400818 306898
rect 445435 306860 445994 306865
rect 445435 306855 445440 306860
rect 445989 306855 445994 306860
rect 400259 306338 400818 306344
rect 430709 306662 431268 306667
rect 430709 306657 430714 306662
rect 431263 306657 431268 306662
rect 370683 306252 371242 306258
rect 357940 306237 357945 306242
rect 358487 306237 358492 306242
rect 357940 306232 358492 306237
rect 445435 306300 445994 306306
rect 470713 306780 470723 306785
rect 470713 306231 470718 306780
rect 470713 306226 470723 306231
rect 471272 306226 471278 306785
rect 490709 306455 490714 307004
rect 490709 306450 490719 306455
rect 491268 306450 491274 307009
rect 510695 306896 510705 306901
rect 510695 306347 510700 306896
rect 510695 306342 510705 306347
rect 511254 306342 511260 306901
rect 569353 306811 569932 306817
rect 530675 306188 530681 306747
rect 531230 306742 531240 306747
rect 531235 306193 531240 306742
rect 531230 306188 531240 306193
rect 552156 306168 552162 306735
rect 552719 306730 552729 306735
rect 552724 306173 552729 306730
rect 569353 306237 569358 306242
rect 569927 306237 569932 306242
rect 569353 306232 569932 306237
rect 552719 306168 552729 306173
rect 430709 306102 431268 306108
rect 348014 305639 348486 305644
rect 118328 304981 168402 304982
rect 118329 304976 123445 304981
rect 355988 302183 356108 302193
rect 355983 302117 355993 302183
rect 356103 302117 356113 302183
rect 355988 302107 356108 302117
rect 355998 301811 356118 301821
rect 355993 301745 356003 301811
rect 356113 301745 356123 301811
rect 355998 301735 356118 301745
rect 355562 296500 356560 296505
rect 549082 296500 550082 296506
rect 355561 296499 370526 296500
rect -800 295420 480 295532
rect 355561 295501 355562 296499
rect 356560 296063 370526 296499
rect 371415 296080 390559 296500
rect 391395 296095 410529 296500
rect 371415 296078 390932 296080
rect 356560 296034 370923 296063
rect 356560 295924 370828 296034
rect 370894 295924 370923 296034
rect 356560 295895 370923 295924
rect 371171 296051 390932 296078
rect 371171 296044 390837 296051
rect 371171 295934 371200 296044
rect 371266 295941 390837 296044
rect 390903 295941 390932 296051
rect 371266 295934 390932 295941
rect 371171 295912 390932 295934
rect 391180 296061 410529 296095
rect 411463 296127 430574 296500
rect 431412 296142 450540 296500
rect 411463 296098 430934 296127
rect 411463 296066 430839 296098
rect 391180 295951 391209 296061
rect 391275 296051 410529 296061
rect 391275 296022 410938 296051
rect 391275 295951 410843 296022
rect 391180 295927 410843 295951
rect 391395 295912 410843 295927
rect 410909 295912 410938 296022
rect 371171 295910 390559 295912
rect 356560 295501 370526 295895
rect 355561 295500 370526 295501
rect 371415 295500 390559 295910
rect 391395 295883 410938 295912
rect 411186 296032 430839 296066
rect 411186 295922 411215 296032
rect 411281 295988 430839 296032
rect 430905 295988 430934 296098
rect 411281 295959 430934 295988
rect 431182 296108 450540 296142
rect 451463 296119 470577 296500
rect 471415 296152 490522 296500
rect 491465 296167 510532 296500
rect 471415 296134 490948 296152
rect 471201 296123 490948 296134
rect 451463 296109 470953 296119
rect 431182 295998 431211 296108
rect 431277 296094 450540 296108
rect 431277 296065 450951 296094
rect 431277 295998 450856 296065
rect 431182 295974 450856 295998
rect 411281 295922 430574 295959
rect 411186 295898 430574 295922
rect 391395 295500 410529 295883
rect 411463 295500 430574 295898
rect 431412 295955 450856 295974
rect 450922 295955 450951 296065
rect 431412 295926 450951 295955
rect 451199 296090 470953 296109
rect 451199 296075 470858 296090
rect 451199 295965 451228 296075
rect 451294 295980 470858 296075
rect 470924 295980 470953 296090
rect 451294 295965 470953 295980
rect 471201 296100 490853 296123
rect 471201 295990 471230 296100
rect 471296 296013 490853 296100
rect 490919 296013 490948 296123
rect 471296 295990 490948 296013
rect 491196 296133 510532 296167
rect 491196 296023 491225 296133
rect 491291 296108 510532 296133
rect 511449 296152 530507 296500
rect 531462 296167 549082 296500
rect 511449 296123 530926 296152
rect 491291 296079 510941 296108
rect 491291 296023 510846 296079
rect 491196 295999 510846 296023
rect 471201 295984 490948 295990
rect 471201 295966 490522 295984
rect 451199 295951 470953 295965
rect 451199 295941 470577 295951
rect 431412 295500 450540 295926
rect 451463 295500 470577 295941
rect 471415 295500 490522 295966
rect 491465 295969 510846 295999
rect 510912 295969 510941 296079
rect 491465 295940 510941 295969
rect 511189 296089 530831 296123
rect 511189 295979 511218 296089
rect 511284 296013 530831 296089
rect 530897 296013 530926 296123
rect 511284 295984 530926 296013
rect 531174 296133 549082 296167
rect 531174 296023 531203 296133
rect 531269 296023 549082 296133
rect 531174 295999 549082 296023
rect 511284 295979 530507 295984
rect 511189 295955 530507 295979
rect 491465 295500 510532 295940
rect 511449 295500 530507 295955
rect 531462 295500 549082 295999
rect 355562 295495 356560 295500
rect 549082 295494 550082 295500
rect -800 294238 480 294350
rect 118329 293773 123445 293778
rect 118328 293772 168402 293773
rect -800 293056 480 293168
rect 49270 292102 50268 292107
rect 14352 292101 50269 292102
rect -800 291874 480 291986
rect 13045 291699 13155 291704
rect 14352 291699 49270 292101
rect 13044 291698 49270 291699
rect 13044 291588 13045 291698
rect 13155 291588 49270 291698
rect 13044 291587 49270 291588
rect 13045 291582 13155 291587
rect 14352 291103 49270 291587
rect 50268 291103 50269 292101
rect 14352 291102 50269 291103
rect 49270 291097 50268 291102
rect 13044 290804 13156 290810
rect -800 290692 13044 290804
rect 13044 290686 13156 290692
rect 25372 289622 25484 289628
rect -800 289510 25372 289622
rect 25372 289504 25484 289510
rect 118328 288656 118329 293772
rect 123445 288656 168402 293772
rect 549537 293441 549667 293446
rect 549537 293375 549547 293441
rect 549657 293375 549667 293441
rect 549537 293370 549667 293375
rect 549547 293069 549677 293074
rect 549547 293003 549557 293069
rect 549667 293003 549677 293069
rect 549547 292998 549677 293003
rect 346935 288890 347055 288900
rect 346930 288824 346940 288890
rect 347050 288824 347060 288890
rect 346935 288814 347055 288824
rect 118328 288655 168402 288656
rect 118329 288650 123445 288655
rect 346945 288518 347065 288528
rect 346940 288452 346950 288518
rect 347060 288452 347070 288518
rect 346945 288442 347065 288452
rect 345700 287588 346172 287593
rect 345700 285614 345710 287588
rect 346162 285614 346172 287588
rect 445447 287026 446006 287032
rect 400175 286908 400734 286914
rect 354030 286266 354036 286818
rect 354578 286813 354588 286818
rect 354583 286271 354588 286813
rect 390695 286696 391254 286702
rect 354578 286266 354588 286271
rect 370683 286607 370693 286612
rect 370683 286058 370688 286607
rect 370683 286053 370693 286058
rect 371242 286053 371248 286612
rect 400175 286354 400180 286359
rect 400729 286354 400734 286359
rect 400175 286349 400734 286354
rect 430709 286814 431268 286820
rect 490709 286883 490719 286888
rect 445447 286472 445452 286477
rect 446001 286472 446006 286477
rect 445447 286467 446006 286472
rect 470713 286753 470723 286758
rect 430709 286260 430714 286265
rect 431263 286260 431268 286265
rect 430709 286255 431268 286260
rect 470713 286204 470718 286753
rect 470713 286199 470723 286204
rect 471272 286199 471278 286758
rect 490709 286334 490714 286883
rect 490709 286329 490719 286334
rect 491268 286329 491274 286888
rect 510695 286819 510705 286824
rect 510695 286270 510700 286819
rect 510695 286265 510705 286270
rect 511254 286265 511260 286824
rect 530681 286807 530691 286812
rect 530681 286258 530686 286807
rect 530681 286253 530691 286258
rect 531240 286253 531246 286812
rect 546309 286421 546315 286988
rect 546872 286983 546882 286988
rect 546877 286426 546882 286983
rect 546872 286421 546882 286426
rect 568313 286887 568892 286893
rect 568313 286313 568318 286318
rect 568887 286313 568892 286318
rect 568313 286308 568892 286313
rect 390695 286142 390700 286147
rect 391249 286142 391254 286147
rect 390695 286137 391254 286142
rect 345700 285609 346172 285614
rect 565650 275140 565656 275252
rect 565768 275140 584800 275252
rect 549072 274464 550093 274475
rect 549072 274463 551155 274464
rect 549072 273465 549083 274463
rect 550081 274045 551155 274463
rect 552079 274060 571543 274464
rect 550081 274016 551544 274045
rect 550081 273906 551449 274016
rect 551515 273906 551544 274016
rect 550081 273877 551544 273906
rect 551792 274026 571543 274060
rect 551792 273916 551821 274026
rect 551887 274005 571543 274026
rect 572548 274070 580774 274464
rect 572548 274020 584800 274070
rect 551887 273976 572007 274005
rect 551887 273916 571912 273976
rect 551792 273892 571912 273916
rect 550081 273465 551155 273877
rect 549072 273464 551155 273465
rect 552079 273866 571912 273892
rect 571978 273866 572007 273976
rect 552079 273837 572007 273866
rect 572255 273986 584800 274020
rect 572255 273876 572284 273986
rect 572350 273958 584800 273986
rect 572350 273876 580774 273958
rect 572255 273852 580774 273876
rect 552079 273464 571543 273837
rect 572548 273464 580774 273852
rect 549072 273450 550093 273464
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 83449 268390 83455 269390
rect 84455 268390 425035 269390
rect 426035 268390 426041 269390
rect 583520 269230 584800 269342
rect 78269 267390 79269 267396
rect 79269 266390 423042 267390
rect 424042 266390 424048 267390
rect 78269 266384 79269 266390
rect 72626 264390 72632 265390
rect 73632 264390 421075 265390
rect 422075 264390 422081 265390
rect 346893 264110 347013 264120
rect 346888 264044 346898 264110
rect 347008 264044 347018 264110
rect 346893 264034 347013 264044
rect 346903 263738 347023 263748
rect 346898 263672 346908 263738
rect 347018 263672 347028 263738
rect 346903 263662 347023 263672
rect 65786 263390 66786 263396
rect 66786 262390 419082 263390
rect 420082 262390 420088 263390
rect 65786 262384 66786 262390
rect 58670 261390 59670 261396
rect 59670 260390 417049 261390
rect 418049 260390 418055 261390
rect 58670 260384 59670 260390
rect 49263 258390 49269 259390
rect 50269 258390 415074 259390
rect 416074 258390 416080 259390
rect 49269 257390 50269 257396
rect 50269 256390 413046 257390
rect 414046 256390 414052 257390
rect 49269 256384 50269 256390
rect 58938 255390 59938 255396
rect 59938 254390 411018 255390
rect 412018 254390 412024 255390
rect 58938 254384 59938 254390
rect 65894 253390 66894 253396
rect -800 252398 480 252510
rect 66894 252390 409097 253390
rect 410097 252390 410103 253390
rect 65894 252384 66894 252390
rect 72906 251390 73906 251396
rect -800 251216 480 251328
rect 73906 250390 407015 251390
rect 408015 250390 408021 251390
rect 72906 250384 73906 250390
rect -800 250034 480 250146
rect 78414 249390 79414 249396
rect -800 248852 480 248964
rect 79414 248390 405094 249390
rect 406094 248390 406100 249390
rect 78414 248384 79414 248390
rect 14889 248052 50269 248053
rect 14889 247782 49270 248052
rect -800 247670 49270 247782
rect 14889 247054 49270 247670
rect 50268 247054 50274 248052
rect 83668 247390 84668 247396
rect 403025 247390 404061 247405
rect 14889 247053 50269 247054
rect 25415 246600 25527 246606
rect -800 246488 25415 246600
rect 25415 246482 25527 246488
rect 84668 247389 404061 247390
rect 84668 246391 403046 247389
rect 404044 246391 404061 247389
rect 84668 246390 404061 246391
rect 83668 246384 84668 246390
rect 403025 246376 404061 246390
rect 346977 242736 347097 242746
rect 346972 242670 346982 242736
rect 347092 242670 347102 242736
rect 346977 242660 347097 242670
rect 346987 242364 347107 242374
rect 346982 242298 346992 242364
rect 347102 242298 347112 242364
rect 346987 242288 347107 242298
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 347005 222860 347125 222870
rect 347000 222794 347010 222860
rect 347120 222794 347130 222860
rect 347005 222784 347125 222794
rect 347015 222488 347135 222498
rect 347010 222422 347020 222488
rect 347130 222422 347140 222488
rect 347015 222412 347135 222422
rect -800 214888 1660 219688
rect 347972 213096 348458 213101
rect -800 204888 1660 209688
rect 347972 208088 347982 213096
rect 348448 208088 348458 213096
rect 347972 208083 348458 208088
rect 346949 201032 347069 201042
rect 346944 200966 346954 201032
rect 347064 200966 347074 201032
rect 346949 200956 347069 200966
rect 346959 200660 347079 200670
rect 346954 200594 346964 200660
rect 347074 200594 347084 200660
rect 346959 200584 347079 200594
rect 570495 191330 570501 196290
rect 575461 196288 580012 196290
rect 575461 196230 583067 196288
rect 575461 191430 584800 196230
rect 575461 191330 583067 191430
rect 578955 191312 583067 191330
rect 570408 181252 570414 186370
rect 575532 186368 580012 186370
rect 575532 186230 583645 186368
rect 575532 181430 584800 186230
rect 575532 181256 583643 181430
rect 575532 181252 580012 181256
rect 346963 179998 347083 180008
rect 346958 179932 346968 179998
rect 347078 179932 347088 179998
rect 346963 179922 347083 179932
rect 346973 179626 347093 179636
rect 346968 179560 346978 179626
rect 347088 179560 347098 179626
rect 346973 179550 347093 179560
rect 990 177688 13066 177860
rect -800 172888 13066 177688
rect 990 172742 13066 172888
rect 18184 172742 18190 177860
rect 345712 177826 346198 177831
rect 345712 172818 345722 177826
rect 346188 172818 346198 177826
rect 345712 172813 346198 172818
rect 808 167688 13374 167862
rect -800 162888 13374 167688
rect 808 162744 13374 162888
rect 18492 162744 18498 167862
rect 345688 167836 346174 167841
rect 345688 162828 345698 167836
rect 346164 162828 346174 167836
rect 345688 162823 346174 162828
rect 346921 158610 347041 158620
rect 346916 158544 346926 158610
rect 347036 158544 347046 158610
rect 346921 158534 347041 158544
rect 346931 158238 347051 158248
rect 346926 158172 346936 158238
rect 347046 158172 347056 158238
rect 346931 158162 347051 158172
rect 582340 146830 584800 151630
rect 334816 136838 334822 137390
rect 335364 137385 335374 137390
rect 335369 136843 335374 137385
rect 358790 137369 358800 137374
rect 346865 137264 346985 137274
rect 346860 137198 346870 137264
rect 346980 137198 346990 137264
rect 346865 137188 346985 137198
rect 346875 136892 346995 136902
rect 335364 136838 335374 136843
rect 346870 136826 346880 136892
rect 346990 136826 347000 136892
rect 358790 136827 358795 137369
rect 346875 136816 346995 136826
rect 358790 136822 358800 136827
rect 359342 136822 359348 137374
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect 58939 120855 59937 120860
rect 14112 120854 59938 120855
rect 14112 120160 58939 120854
rect -800 120048 58939 120160
rect 14112 119856 58939 120048
rect 59937 119856 59938 120854
rect 14112 119855 59938 119856
rect 58939 119850 59937 119855
rect 25403 118978 25515 118984
rect -800 118866 25403 118978
rect 25403 118860 25515 118866
rect 346921 116130 347041 116140
rect 346916 116064 346926 116130
rect 347036 116064 347046 116130
rect 346921 116054 347041 116064
rect 346931 115758 347051 115768
rect 346926 115692 346936 115758
rect 347046 115692 347056 115758
rect 346931 115682 347051 115692
rect 334788 95092 334794 95644
rect 335336 95639 335346 95644
rect 335341 95097 335346 95639
rect 359138 95639 359148 95644
rect 346949 95520 347069 95530
rect 346944 95454 346954 95520
rect 347064 95454 347074 95520
rect 346949 95444 347069 95454
rect 346959 95148 347079 95158
rect 335336 95092 335346 95097
rect 346954 95082 346964 95148
rect 347074 95082 347084 95148
rect 359138 95097 359143 95639
rect 359138 95092 359148 95097
rect 359690 95092 359696 95644
rect 583520 95118 584800 95230
rect 346959 95072 347079 95082
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 14112 79051 66894 79052
rect 12334 78528 12444 78533
rect 14112 78528 65895 79051
rect 12333 78527 65895 78528
rect 12333 78417 12334 78527
rect 12444 78417 65895 78527
rect 12333 78416 65895 78417
rect 12334 78411 12444 78416
rect -800 78008 480 78120
rect 14112 78053 65895 78416
rect 66893 78053 66899 79051
rect 14112 78052 66894 78053
rect 12333 76938 12445 76944
rect -800 76826 12333 76938
rect 12333 76820 12445 76826
rect 25414 75756 25526 75762
rect -800 75644 25414 75756
rect 25414 75638 25526 75644
rect 346935 74838 347055 74848
rect 346930 74772 346940 74838
rect 347050 74772 347060 74838
rect 346935 74762 347055 74772
rect 346945 74466 347065 74476
rect 346940 74400 346950 74466
rect 347060 74400 347070 74466
rect 346945 74390 347065 74400
rect 72894 66137 73915 66152
rect 15445 66136 73915 66137
rect 12619 65629 12729 65634
rect 15445 65629 72907 66136
rect 12618 65628 72907 65629
rect 12618 65518 12619 65628
rect 12729 65518 72907 65628
rect 12618 65517 72907 65518
rect 12619 65512 12729 65517
rect 15445 65138 72907 65517
rect 73905 65138 73915 66136
rect 15445 65137 73915 65138
rect 72894 65128 73915 65137
rect 78386 62396 79436 62431
rect 15445 62395 79436 62396
rect 14459 62017 14569 62022
rect 15445 62017 78415 62395
rect 14458 62016 78415 62017
rect 14458 61906 14459 62016
rect 14569 61906 78415 62016
rect 14458 61905 78415 61906
rect 14459 61900 14569 61905
rect 15445 61397 78415 61905
rect 79413 61397 79436 62395
rect 15445 61396 79436 61397
rect 78386 61367 79436 61396
rect 90274 60006 91548 60011
rect 83660 59107 84676 59115
rect 15445 59106 84676 59107
rect 15445 58593 83669 59106
rect 15445 58483 16146 58593
rect 16256 58483 83669 58593
rect 15445 58108 83669 58483
rect 84667 58108 84676 59106
rect 90274 58752 90284 60006
rect 91538 58752 91548 60006
rect 302574 59503 302584 59508
rect 240070 59386 240622 59392
rect 133044 59376 133596 59382
rect 111722 59366 112274 59372
rect 133044 58829 133049 58834
rect 133591 58829 133596 58834
rect 133044 58824 133596 58829
rect 154602 59332 155154 59338
rect 111722 58819 111727 58824
rect 112269 58819 112274 58824
rect 111722 58814 112274 58819
rect 154602 58785 154607 58790
rect 155149 58785 155154 58790
rect 154602 58780 155154 58785
rect 175808 59332 176360 59338
rect 219084 59310 219636 59316
rect 175808 58785 175813 58790
rect 176355 58785 176360 58790
rect 175808 58780 176360 58785
rect 197190 59288 197742 59294
rect 90274 58747 91548 58752
rect 240070 58839 240075 58844
rect 240617 58839 240622 58844
rect 240070 58834 240622 58839
rect 260572 59379 260582 59384
rect 260572 58837 260577 59379
rect 260572 58832 260582 58837
rect 261124 58832 261130 59384
rect 281384 59135 281394 59140
rect 219084 58763 219089 58768
rect 219631 58763 219636 58768
rect 219084 58758 219636 58763
rect 197190 58741 197195 58746
rect 197737 58741 197742 58746
rect 197190 58736 197742 58741
rect 281384 58593 281389 59135
rect 281384 58588 281394 58593
rect 281936 58588 281942 59140
rect 302574 58961 302579 59503
rect 302574 58956 302584 58961
rect 303126 58956 303132 59508
rect 324116 58956 324122 59508
rect 324664 59503 324674 59508
rect 324669 58961 324674 59503
rect 324664 58956 324674 58961
rect 15445 58107 84676 58108
rect 83660 58099 84676 58107
rect 334718 54530 335270 54536
rect 334718 53983 334723 53988
rect 335265 53983 335270 53988
rect 334718 53978 335270 53983
rect 358800 54525 358810 54530
rect 358800 53983 358805 54525
rect 358800 53978 358810 53983
rect 359352 53978 359358 54530
rect 39900 52866 40872 52872
rect 39900 51899 39905 51904
rect 40867 51899 40872 51904
rect 39900 51894 40872 51899
rect 347005 51258 347125 51268
rect 347000 51192 347010 51258
rect 347120 51192 347130 51258
rect 347005 51182 347125 51192
rect 347015 50886 347135 50896
rect 347010 50820 347020 50886
rect 347130 50820 347140 50886
rect 347015 50810 347135 50820
rect 583520 50460 584800 50572
rect 34106 49302 35106 49308
rect 35106 48906 47892 49302
rect 48726 48966 69174 49302
rect 69998 48982 90482 49302
rect 48726 48946 69374 48966
rect 48726 48922 69284 48946
rect 35106 48886 48080 48906
rect 35106 48776 47990 48886
rect 48056 48776 48080 48886
rect 35106 48752 48080 48776
rect 48332 48896 69284 48922
rect 48332 48786 48362 48896
rect 48428 48836 69284 48896
rect 69350 48836 69374 48946
rect 48428 48812 69374 48836
rect 69626 48956 90482 48982
rect 69626 48846 69656 48956
rect 69722 48892 90482 48956
rect 91386 48936 111558 49302
rect 112450 48980 132872 49302
rect 133768 48996 154450 49302
rect 112450 48960 133122 48980
rect 112450 48952 133032 48960
rect 91386 48916 111800 48936
rect 91386 48908 111710 48916
rect 69722 48872 90740 48892
rect 69722 48846 90650 48872
rect 69626 48828 90650 48846
rect 48428 48786 69174 48812
rect 48332 48768 69174 48786
rect 35106 48302 47892 48752
rect 48726 48302 69174 48768
rect 69998 48762 90650 48828
rect 90716 48762 90740 48872
rect 69998 48738 90740 48762
rect 90992 48882 111710 48908
rect 90992 48772 91022 48882
rect 91088 48806 111710 48882
rect 111776 48806 111800 48916
rect 91088 48782 111800 48806
rect 112052 48926 133032 48952
rect 112052 48816 112082 48926
rect 112148 48850 133032 48926
rect 133098 48850 133122 48960
rect 112148 48826 133122 48850
rect 133374 48970 154450 48996
rect 133374 48860 133404 48970
rect 133470 48950 154450 48970
rect 155320 48966 175654 49302
rect 133470 48930 154680 48950
rect 133470 48860 154590 48930
rect 133374 48842 154590 48860
rect 112148 48816 132872 48826
rect 112052 48798 132872 48816
rect 91088 48772 111558 48782
rect 90992 48754 111558 48772
rect 69998 48302 90482 48738
rect 91386 48302 111558 48754
rect 112450 48302 132872 48798
rect 133768 48820 154590 48842
rect 154656 48820 154680 48930
rect 133768 48796 154680 48820
rect 154932 48940 175654 48966
rect 154932 48830 154962 48940
rect 155028 48922 175654 48940
rect 176512 48980 197072 49302
rect 197864 48996 218938 49302
rect 176512 48960 197268 48980
rect 176512 48938 197178 48960
rect 155028 48902 175886 48922
rect 155028 48830 175796 48902
rect 154932 48812 175796 48830
rect 133768 48302 154450 48796
rect 155320 48792 175796 48812
rect 175862 48792 175886 48902
rect 155320 48768 175886 48792
rect 176138 48912 197178 48938
rect 176138 48802 176168 48912
rect 176234 48850 197178 48912
rect 197244 48850 197268 48960
rect 176234 48826 197268 48850
rect 197520 48970 218938 48996
rect 197520 48860 197550 48970
rect 197616 48892 218938 48970
rect 219830 48908 239926 49302
rect 197616 48872 219162 48892
rect 197616 48860 219072 48872
rect 197520 48842 219072 48860
rect 176234 48802 197072 48826
rect 176138 48784 197072 48802
rect 155320 48302 175654 48768
rect 176512 48302 197072 48784
rect 197864 48762 219072 48842
rect 219138 48762 219162 48872
rect 197864 48738 219162 48762
rect 219414 48882 239926 48908
rect 219414 48772 219444 48882
rect 219510 48862 239926 48882
rect 240788 48922 260446 49302
rect 261264 49024 281258 49302
rect 282082 49040 302450 49302
rect 261264 49004 281462 49024
rect 261264 48938 281372 49004
rect 240788 48902 260650 48922
rect 240788 48878 260560 48902
rect 219510 48842 240148 48862
rect 219510 48772 240058 48842
rect 219414 48754 240058 48772
rect 197864 48302 218938 48738
rect 219830 48732 240058 48754
rect 240124 48732 240148 48842
rect 219830 48708 240148 48732
rect 240400 48852 260560 48878
rect 240400 48742 240430 48852
rect 240496 48792 260560 48852
rect 260626 48792 260650 48902
rect 240496 48768 260650 48792
rect 260902 48912 281372 48938
rect 260902 48802 260932 48912
rect 260998 48894 281372 48912
rect 281438 48894 281462 49004
rect 260998 48870 281462 48894
rect 281714 49014 302450 49040
rect 281714 48904 281744 49014
rect 281810 48904 302450 49014
rect 281714 48886 302450 48904
rect 260998 48802 281258 48870
rect 260902 48784 281258 48802
rect 240496 48742 260446 48768
rect 240400 48724 260446 48742
rect 219830 48302 239926 48708
rect 240788 48302 260446 48724
rect 261264 48302 281258 48784
rect 282082 48818 302450 48886
rect 303290 48854 323962 49302
rect 324824 49301 347574 49302
rect 324824 48870 346575 49301
rect 303290 48834 324200 48854
rect 282082 48798 302652 48818
rect 282082 48688 302562 48798
rect 302628 48688 302652 48798
rect 282082 48664 302652 48688
rect 302904 48808 324110 48834
rect 302904 48698 302934 48808
rect 303000 48724 324110 48808
rect 324176 48724 324200 48834
rect 303000 48700 324200 48724
rect 324452 48844 346575 48870
rect 324452 48734 324482 48844
rect 324548 48734 346575 48844
rect 324452 48716 346575 48734
rect 303000 48698 323962 48700
rect 302904 48680 323962 48698
rect 282082 48302 302450 48664
rect 303290 48302 323962 48680
rect 324824 48303 346575 48716
rect 347573 48303 347579 49301
rect 583520 49278 584800 49390
rect 324824 48302 347574 48303
rect 34106 48296 35106 48302
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 34573 43004 34693 43014
rect 34568 42938 34578 43004
rect 34688 42938 34698 43004
rect 34573 42928 34693 42938
rect 34583 42632 34703 42642
rect 34578 42566 34588 42632
rect 34698 42566 34708 42632
rect 34583 42556 34703 42566
rect 39640 39258 42772 39263
rect -800 38332 480 38444
rect -800 37150 480 37262
rect 39640 36270 39650 39258
rect 42762 36270 42772 39258
rect 69298 38013 69850 38018
rect 69298 38008 69303 38013
rect 69845 38008 69850 38013
rect 48004 37907 48556 37912
rect 48004 37902 48009 37907
rect 48551 37902 48556 37907
rect 197192 37933 197744 37938
rect 197192 37928 197197 37933
rect 197739 37928 197744 37933
rect 154604 37835 155156 37840
rect 154604 37830 154609 37835
rect 155151 37830 155156 37835
rect 111724 37747 112276 37752
rect 111724 37742 111729 37747
rect 112271 37742 112276 37747
rect 69298 37460 69850 37466
rect 90664 37695 91216 37700
rect 90664 37690 90669 37695
rect 91211 37690 91216 37695
rect 48004 37354 48556 37360
rect 111724 37194 112276 37200
rect 133046 37667 133056 37672
rect 90664 37142 91216 37148
rect 133046 37125 133051 37667
rect 133046 37120 133056 37125
rect 133598 37120 133604 37672
rect 154604 37282 155156 37288
rect 175810 37835 176362 37840
rect 175810 37830 175815 37835
rect 176357 37830 176362 37835
rect 197192 37380 197744 37386
rect 219086 37883 219638 37888
rect 219086 37878 219091 37883
rect 219633 37878 219638 37883
rect 219086 37330 219638 37336
rect 175810 37282 176362 37288
rect 240066 37234 240072 37786
rect 240614 37781 240624 37786
rect 240619 37239 240624 37781
rect 240614 37234 240624 37239
rect 260568 37172 260574 37724
rect 261116 37719 261126 37724
rect 261121 37177 261126 37719
rect 281380 37268 281386 37820
rect 281928 37815 281938 37820
rect 281933 37273 281938 37815
rect 302570 37372 302576 37924
rect 303118 37919 303128 37924
rect 303123 37377 303128 37919
rect 303118 37372 303128 37377
rect 324118 37320 324124 37872
rect 324666 37867 324676 37872
rect 324671 37325 324676 37867
rect 324666 37320 324676 37325
rect 281928 37268 281938 37273
rect 261116 37172 261126 37177
rect 39640 36265 42772 36270
rect -800 35968 480 36080
rect -800 34786 480 34898
rect 12618 33716 12730 33722
rect -800 33604 12618 33716
rect 12618 33598 12730 33604
rect -800 32422 25408 32534
rect 25520 32422 25526 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 34573 20906 34693 20916
rect 34568 20840 34578 20906
rect 34688 20840 34698 20906
rect 34573 20830 34693 20840
rect 34583 20534 34703 20544
rect 34578 20468 34588 20534
rect 34698 20468 34708 20534
rect 34583 20458 34703 20468
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 25446 18906 25558 18912
rect 21662 18905 25446 18906
rect 21657 18795 21663 18905
rect 21773 18795 25446 18905
rect 21662 18794 25446 18795
rect 25446 18788 25558 18794
rect 583520 18092 584800 18204
rect 25438 18068 25550 18074
rect 22608 18067 25438 18068
rect 22603 17957 22609 18067
rect 22719 17957 25438 18067
rect 22608 17956 25438 17957
rect 25438 17950 25550 17956
rect 24982 17174 25982 17180
rect 565200 17174 566198 17179
rect -800 16910 480 17022
rect 25982 17173 566199 17174
rect 25982 16175 565200 17173
rect 566198 16175 566199 17173
rect 583520 16910 584800 17022
rect 25982 16174 566199 16175
rect 24982 16168 25982 16174
rect 565200 16169 566198 16174
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect 14458 12294 14570 12300
rect -800 12182 14458 12294
rect 583520 12182 584800 12294
rect 14458 12176 14570 12182
rect 21662 11112 21774 11118
rect -800 11000 21662 11112
rect 583520 11000 584800 11112
rect 21662 10994 21774 11000
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect 338571 8590 338693 8595
rect 344312 8590 344424 8596
rect 338571 8478 338576 8590
rect 338688 8478 344312 8590
rect 338571 8473 338693 8478
rect 344312 8472 344424 8478
rect 350866 8200 350978 8206
rect 356301 8200 356423 8205
rect 350978 8088 356306 8200
rect 356418 8088 356423 8200
rect 350866 8082 350978 8088
rect 356301 8083 356423 8088
rect 342117 7854 342239 7859
rect 345070 7854 345182 7860
rect 342117 7742 342122 7854
rect 342234 7742 345070 7854
rect 342117 7737 342239 7742
rect 345070 7736 345182 7742
rect 16145 7566 16257 7572
rect -800 7454 16145 7566
rect 583520 7454 584800 7566
rect 16145 7448 16257 7454
rect 350238 7296 350350 7302
rect 352755 7296 352877 7301
rect 345663 7256 345785 7261
rect 348884 7256 348996 7262
rect 345663 7144 345668 7256
rect 345780 7144 348884 7256
rect 350350 7184 352760 7296
rect 352872 7184 352877 7296
rect 350238 7178 350350 7184
rect 352755 7179 352877 7184
rect 345663 7139 345785 7144
rect 348884 7138 348996 7144
rect 349579 6633 349701 6639
rect 349579 6516 349584 6521
rect 349696 6516 349701 6521
rect 349579 6511 349701 6516
rect 22608 6384 22720 6390
rect -800 6272 22608 6384
rect 583520 6272 584800 6384
rect 22608 6266 22720 6272
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect 476865 4020 476987 4025
rect 478105 4020 478215 4025
rect 480411 4020 480533 4025
rect -800 3908 480 4020
rect 34107 3948 35105 3953
rect 4138 3582 6352 3948
rect 7356 3642 27596 3948
rect 28538 3947 35106 3948
rect 28538 3658 34107 3947
rect 7356 3622 27830 3642
rect 7356 3598 27740 3622
rect 4138 3562 6638 3582
rect 2637 3494 2747 3499
rect 4138 3494 6548 3562
rect 2636 3493 6548 3494
rect 2636 3383 2637 3493
rect 2747 3452 6548 3493
rect 6614 3452 6638 3562
rect 2747 3428 6638 3452
rect 6890 3572 27740 3598
rect 6890 3462 6920 3572
rect 6986 3512 27740 3572
rect 27806 3512 27830 3622
rect 6986 3488 27830 3512
rect 28082 3632 34107 3658
rect 28082 3522 28112 3632
rect 28178 3522 34107 3632
rect 28082 3504 34107 3522
rect 6986 3462 27596 3488
rect 6890 3444 27596 3462
rect 2747 3383 6352 3428
rect 2636 3382 6352 3383
rect 2637 3377 2747 3382
rect 4138 2948 6352 3382
rect 7356 2948 27596 3444
rect 28538 2949 34107 3504
rect 35105 2949 35106 3947
rect 476865 3908 476870 4020
rect 476982 4019 478216 4020
rect 476982 3909 478105 4019
rect 478215 3909 478216 4019
rect 476982 3908 478216 3909
rect 480411 3908 480416 4020
rect 480528 4014 480533 4020
rect 483957 4024 484079 4029
rect 488006 4024 488116 4029
rect 482770 4014 482880 4019
rect 480528 4013 482881 4014
rect 480528 3908 482770 4013
rect 476865 3903 476987 3908
rect 478105 3903 478215 3908
rect 480411 3903 482770 3908
rect 482880 3903 482881 4013
rect 483957 3912 483962 4024
rect 484074 4023 488116 4024
rect 484074 3913 488006 4023
rect 484074 3912 488116 3913
rect 483957 3907 484079 3912
rect 488006 3907 488116 3912
rect 583520 3908 584800 4020
rect 480412 3902 482881 3903
rect 482770 3897 482880 3902
rect 28538 2948 35106 2949
rect 34107 2943 35105 2948
rect 2636 2838 2748 2844
rect -800 2726 2636 2838
rect 583520 2726 584800 2838
rect 2636 2720 2748 2726
rect 25358 1656 25470 1662
rect -800 1544 25358 1656
rect 583520 1544 584800 1656
rect 25358 1538 25470 1544
<< via3 >>
rect 8383 643688 13471 648776
rect 8391 633670 13463 638742
rect 570818 639592 575920 644694
rect 570873 629638 575909 634674
rect 487607 602558 488607 603558
rect 482433 596090 483433 597090
rect 477776 589077 478776 590077
rect 565585 589472 565697 589584
rect 544392 586294 545390 587292
rect 537804 579323 538406 579328
rect 537804 578721 537809 579323
rect 537809 578721 538406 579323
rect 537804 578716 538406 578721
rect 544736 573153 544846 573219
rect 544726 572781 544836 572847
rect 505085 567274 506083 568272
rect 513276 567273 514276 568273
rect 522152 567444 523150 568442
rect 530514 567443 531514 568443
rect 513762 562597 513872 562663
rect 513752 562225 513862 562291
rect 505449 560504 505559 560570
rect 505439 560132 505549 560198
rect 509408 554242 509938 556160
rect 526608 554236 527208 556182
rect 547182 554212 547758 556178
rect 531032 553043 531142 553109
rect 544746 552904 544856 552970
rect 531022 552671 531132 552737
rect 544736 552532 544846 552598
rect 522511 550426 522621 550492
rect 522501 550054 522611 550120
rect 118329 537740 123445 542856
rect 513742 542155 513852 542221
rect 513732 541783 513842 541849
rect 505559 539916 505669 539982
rect 500438 539631 501050 539636
rect 484633 539557 485235 539562
rect 464242 539447 464844 539452
rect 464242 538845 464839 539447
rect 464839 538845 464844 539447
rect 464242 538840 464844 538845
rect 484633 538955 485230 539557
rect 485230 538955 485235 539557
rect 484633 538950 485235 538955
rect 500438 539034 500443 539631
rect 500443 539034 501045 539631
rect 501045 539034 501050 539631
rect 505549 539544 505659 539610
rect 517874 538396 518574 540212
rect 537834 538328 538410 540294
rect 565238 538344 566160 540236
rect 425730 535325 425794 535389
rect 423449 532885 423513 532949
rect 544751 532678 544861 532744
rect 355561 531597 356561 532597
rect 544741 532306 544851 532372
rect 530987 531798 531097 531864
rect 118329 521230 123445 526346
rect 355991 522045 356101 522111
rect 530977 531426 531087 531492
rect 421586 530323 421650 530387
rect 522560 529649 522670 529715
rect 522550 529277 522660 529343
rect 419511 527883 419575 527947
rect 417545 525321 417609 525385
rect 415545 522881 415609 522945
rect 513739 522184 513849 522250
rect 356001 521673 356111 521739
rect 513729 521812 513839 521878
rect 413516 520319 413580 520383
rect 505084 518692 506084 519692
rect 513277 518804 514275 519802
rect 522151 518803 523151 519803
rect 530515 518804 531513 519802
rect 544391 518792 545391 519792
rect 411487 517879 411551 517943
rect 365528 516349 366528 517349
rect 409483 515317 409547 515381
rect 407542 512877 407606 512941
rect 405502 510315 405566 510379
rect 501674 509564 502674 510564
rect 508549 509565 509547 510563
rect 514542 509484 515542 510484
rect 521017 509485 522015 510483
rect 527090 509404 528090 510404
rect 533845 509405 534843 510403
rect 12230 508776 12340 508886
rect 83456 508248 84454 509246
rect 534334 508886 534444 508952
rect 534344 508514 534454 508580
rect 515038 507867 515148 507933
rect 12229 506802 12341 506914
rect 25370 505620 25482 505732
rect 118329 502694 123445 507810
rect 387914 507753 387978 507817
rect 403541 507753 403605 507817
rect 515028 507495 515138 507561
rect 508942 506459 509052 506525
rect 508932 506087 509042 506153
rect 350839 504704 351065 504930
rect 373642 504702 373712 504707
rect 373642 504642 373647 504702
rect 373647 504642 373707 504702
rect 373707 504642 373712 504702
rect 373642 504637 373712 504642
rect 383216 504757 383280 504762
rect 383216 504697 383275 504757
rect 383275 504697 383280 504757
rect 383216 504692 383280 504697
rect 392784 504716 392848 504721
rect 392784 504656 392843 504716
rect 392843 504656 392848 504716
rect 392784 504651 392848 504656
rect 350185 502752 350411 502978
rect 355956 502136 356066 502202
rect 355966 501764 356076 501830
rect 502178 500260 502288 500326
rect 559955 500050 560067 500162
rect 502168 499888 502278 499954
rect 521392 498333 521502 498399
rect 521382 497961 521492 498027
rect 549986 497325 550984 498323
rect 349515 496736 349741 496962
rect 527466 495935 527576 496001
rect 527456 495563 527566 495629
rect 348839 494692 349065 494918
rect 550466 491990 550576 492056
rect 550456 491618 550566 491684
rect 387905 490687 388015 490753
rect 392808 490701 392918 490767
rect 373616 490608 373726 490674
rect 383268 490606 383378 490672
rect 387915 490315 388025 490381
rect 392818 490329 392928 490395
rect 373626 490236 373736 490302
rect 383278 490234 383388 490300
rect 534344 488486 534454 488552
rect 534354 488114 534464 488180
rect 515001 487666 515111 487732
rect 346574 486302 347574 487302
rect 514991 487294 515101 487360
rect 508954 486408 509064 486474
rect 508944 486036 509054 486102
rect 458514 485307 459126 485312
rect 360438 485147 360990 485152
rect 345009 484496 345235 484722
rect 360438 484610 360443 485147
rect 360443 484610 360985 485147
rect 360985 484610 360990 485147
rect 375484 484747 375489 485284
rect 375489 484747 376031 485284
rect 376031 484747 376036 485284
rect 375484 484742 376036 484747
rect 386090 484671 386095 485208
rect 386095 484671 386637 485208
rect 386637 484671 386642 485208
rect 386090 484666 386642 484671
rect 390324 485211 390876 485216
rect 390324 484674 390329 485211
rect 390329 484674 390871 485211
rect 390871 484674 390876 485211
rect 400218 485181 400770 485186
rect 400218 484644 400223 485181
rect 400223 484644 400765 485181
rect 400765 484644 400770 485181
rect 428636 484679 428641 485216
rect 428641 484679 429183 485216
rect 429183 484679 429188 485216
rect 428636 484674 429188 484679
rect 434800 484627 434805 485224
rect 434805 484627 435407 485224
rect 435407 484627 435412 485224
rect 458514 484710 458519 485307
rect 458519 484710 459121 485307
rect 459121 484710 459126 485307
rect 464285 485157 464897 485162
rect 434800 484622 435412 484627
rect 464285 484560 464290 485157
rect 464290 484560 464892 485157
rect 464892 484560 464897 485157
rect 475004 485127 475616 485132
rect 475004 484530 475009 485127
rect 475009 484530 475611 485127
rect 475611 484530 475616 485127
rect 484623 485195 485225 485200
rect 484623 484593 484628 485195
rect 484628 484593 485225 485195
rect 504622 485165 505234 485170
rect 484623 484588 485225 484593
rect 498498 485111 499100 485116
rect 498498 484509 498503 485111
rect 498503 484509 499100 485111
rect 504622 484568 504627 485165
rect 504627 484568 505229 485165
rect 505229 484568 505234 485165
rect 511839 485215 512441 485220
rect 511839 484613 511844 485215
rect 511844 484613 512441 485215
rect 511839 484608 512441 484613
rect 518208 485215 518838 485220
rect 518208 484585 518213 485215
rect 518213 484585 518838 485215
rect 530384 485173 530996 485178
rect 518208 484580 518838 484585
rect 524295 485159 524897 485164
rect 524295 484557 524892 485159
rect 524892 484557 524897 485159
rect 524295 484552 524897 484557
rect 530384 484576 530389 485173
rect 530389 484576 530991 485173
rect 530991 484576 530996 485173
rect 531886 484591 531891 485216
rect 531891 484591 532521 485216
rect 532521 484591 532526 485216
rect 567854 485171 568484 485176
rect 531886 484586 532526 484591
rect 498498 484504 499100 484509
rect 545779 485127 546409 485132
rect 545779 484497 545784 485127
rect 545784 484497 546409 485127
rect 567854 484541 568479 485171
rect 568479 484541 568484 485171
rect 567854 484536 568484 484541
rect 545779 484492 546409 484497
rect 344281 482178 344507 482404
rect 356018 482192 356128 482258
rect 356028 481820 356138 481886
rect 382735 479110 383733 480108
rect 501675 479115 502673 480113
rect 508548 479114 509548 480114
rect 514543 479115 515541 480113
rect 521016 479114 522016 480114
rect 527091 479115 528089 480113
rect 533844 479116 534844 480116
rect 549985 479109 550985 480109
rect 346982 478252 347092 478318
rect 346992 477880 347102 477946
rect 373156 475017 374154 476015
rect 501707 475012 502705 476010
rect 508580 475011 509580 476011
rect 514575 475012 515573 476010
rect 521048 475011 522048 476011
rect 527123 475012 528121 476010
rect 533876 475009 534876 476009
rect 549890 475016 550890 476016
rect 380562 473159 381104 473164
rect 352776 472981 353318 472986
rect 352776 472439 352781 472981
rect 352781 472439 353318 472981
rect 380562 472617 381099 473159
rect 381099 472617 381104 473159
rect 380562 472612 381104 472617
rect 389486 472541 389491 473078
rect 389491 472541 390033 473078
rect 390033 472541 390038 473078
rect 394692 472615 394697 473152
rect 394697 472615 395239 473152
rect 395239 472615 395244 473152
rect 394692 472610 395244 472615
rect 400586 472567 400591 473104
rect 400591 472567 401133 473104
rect 401133 472567 401138 473104
rect 400586 472562 401138 472567
rect 428290 473109 428842 473114
rect 428290 472572 428295 473109
rect 428295 472572 428837 473109
rect 428837 472572 428842 473109
rect 445478 473047 446090 473052
rect 389486 472536 390038 472541
rect 445478 472450 445483 473047
rect 445483 472450 446085 473047
rect 446085 472450 446090 473047
rect 462130 472457 462135 473054
rect 462135 472457 462737 473054
rect 462737 472457 462742 473054
rect 485292 472501 485297 473098
rect 485297 472501 485899 473098
rect 485899 472501 485904 473098
rect 497347 472566 497352 473189
rect 497352 472566 497980 473189
rect 497980 472566 497985 473189
rect 536948 473163 537550 473168
rect 497347 472561 497985 472566
rect 485292 472496 485904 472501
rect 462130 472452 462742 472457
rect 352776 472434 353318 472439
rect 503855 472370 503860 472993
rect 503860 472370 504488 472993
rect 504488 472370 504493 472993
rect 506690 473001 507292 473006
rect 506690 472399 506695 473001
rect 506695 472399 507292 473001
rect 518230 473087 518832 473092
rect 518230 472485 518235 473087
rect 518235 472485 518832 473087
rect 522944 472495 525127 473097
rect 536948 472561 537545 473163
rect 537545 472561 537550 473163
rect 536948 472556 537550 472561
rect 537962 473141 538592 473146
rect 537962 472511 538587 473141
rect 538587 472511 538592 473141
rect 537962 472506 538592 472511
rect 548148 473207 548778 473212
rect 548148 472577 548153 473207
rect 548153 472577 548778 473207
rect 548148 472572 548778 472577
rect 553168 473131 553798 473136
rect 553168 472501 553793 473131
rect 553793 472501 553798 473131
rect 553168 472496 553798 472501
rect 562798 473059 563438 473064
rect 518230 472480 518832 472485
rect 562798 472434 562803 473059
rect 562803 472434 563433 473059
rect 563433 472434 563438 473059
rect 506690 472394 507292 472399
rect 503855 472365 504493 472370
rect 387914 469723 388024 469789
rect 392806 469723 392916 469789
rect 387924 469351 388034 469417
rect 392816 469351 392926 469417
rect 508976 469023 509086 469089
rect 508986 468651 509096 468717
rect 515023 467765 515133 467831
rect 515033 467393 515143 467459
rect 534386 466945 534496 467011
rect 534376 466573 534486 466639
rect 13363 464658 13473 464768
rect 78270 464203 79268 465201
rect 13362 463580 13474 463692
rect 25407 462398 25519 462510
rect 356026 462172 356136 462238
rect 356036 461800 356146 461866
rect 550370 459665 550480 459731
rect 527531 459536 527641 459602
rect 550360 459293 550470 459359
rect 240180 456761 241180 457761
rect 527521 459164 527631 459230
rect 250981 456761 251981 457761
rect 521414 457098 521524 457164
rect 346996 456998 347106 457064
rect 521424 456726 521534 456792
rect 347006 456626 347116 456692
rect 240701 455849 240811 455915
rect 251423 455827 251533 455893
rect 560008 455628 560120 455740
rect 240711 455477 240821 455543
rect 251433 455455 251543 455521
rect 502200 455171 502310 455237
rect 502210 454799 502320 454865
rect 549891 452861 550889 453859
rect 508964 448972 509074 449038
rect 392796 448771 392906 448837
rect 387875 448703 387985 448769
rect 508974 448600 509084 448666
rect 392806 448399 392916 448465
rect 387885 448331 387995 448397
rect 515060 447564 515170 447630
rect 515070 447192 515180 447258
rect 534376 446545 534486 446611
rect 534366 446173 534476 446239
rect 501706 444561 502706 445561
rect 508581 444562 509579 445560
rect 514574 444641 515574 445641
rect 521049 444642 522047 445640
rect 527122 444721 528122 445721
rect 533877 444722 534875 445720
rect 356000 442179 356110 442245
rect 356010 441807 356120 441873
rect 346968 436390 347078 436456
rect 346978 436018 347088 436084
rect 240621 434332 240731 434398
rect 251406 434046 251516 434112
rect 240631 433960 240741 434026
rect 251416 433674 251526 433740
rect 238861 430259 239402 430264
rect 238861 429718 238866 430259
rect 238866 429718 239402 430259
rect 249230 430379 249772 430384
rect 249230 429837 249235 430379
rect 249235 429837 249772 430379
rect 249230 429832 249772 429837
rect 252975 430363 253527 430368
rect 332864 430371 333416 430376
rect 252975 429826 252980 430363
rect 252980 429826 253522 430363
rect 253522 429826 253527 430363
rect 258343 430362 258883 430367
rect 258343 429822 258878 430362
rect 258878 429822 258883 430362
rect 258343 429817 258883 429822
rect 293219 430355 293761 430360
rect 278455 430343 278997 430348
rect 272935 429757 272940 430294
rect 272940 429757 273482 430294
rect 273482 429757 273487 430294
rect 278455 429801 278992 430343
rect 278992 429801 278997 430343
rect 278455 429796 278997 429801
rect 293219 429813 293756 430355
rect 293756 429813 293761 430355
rect 293219 429808 293761 429813
rect 299167 430255 299709 430260
rect 272935 429752 273487 429757
rect 238861 429713 239402 429718
rect 299167 429713 299704 430255
rect 299704 429713 299709 430255
rect 299167 429708 299709 429713
rect 322090 430215 322632 430220
rect 313343 430191 313895 430196
rect 313343 429654 313348 430191
rect 313348 429654 313890 430191
rect 313890 429654 313895 430191
rect 319481 430157 320023 430162
rect 319481 429615 320018 430157
rect 320018 429615 320023 430157
rect 319481 429610 320023 429615
rect 322090 429673 322627 430215
rect 322627 429673 322632 430215
rect 322090 429668 322632 429673
rect 332864 429834 332869 430371
rect 332869 429834 333411 430371
rect 333411 429834 333416 430371
rect 335399 430253 335941 430258
rect 335399 429711 335936 430253
rect 335936 429711 335941 430253
rect 335399 429706 335941 429711
rect 348094 429382 348522 430698
rect 359996 430439 360548 430444
rect 354352 429727 354357 430264
rect 354357 429727 354899 430264
rect 354899 429727 354904 430264
rect 359996 429902 360001 430439
rect 360001 429902 360543 430439
rect 360543 429902 360548 430439
rect 362166 429901 362171 430438
rect 362171 429901 362713 430438
rect 362713 429901 362718 430438
rect 497205 430398 497843 430403
rect 362166 429896 362718 429901
rect 373955 430191 374497 430196
rect 354352 429722 354904 429727
rect 373955 429649 374492 430191
rect 374492 429649 374497 430191
rect 373955 429644 374497 429649
rect 375347 430195 375899 430200
rect 375347 429658 375352 430195
rect 375352 429658 375894 430195
rect 375894 429658 375899 430195
rect 385928 430287 386470 430292
rect 385928 429745 385933 430287
rect 385933 429745 386470 430287
rect 391200 430371 391742 430376
rect 391200 429829 391205 430371
rect 391205 429829 391742 430371
rect 391200 429824 391742 429829
rect 497205 429775 497210 430398
rect 497210 429775 497838 430398
rect 497838 429775 497843 430398
rect 513062 430335 513674 430340
rect 510278 430285 510890 430290
rect 385928 429740 386470 429745
rect 510278 429688 510283 430285
rect 510283 429688 510885 430285
rect 510885 429688 510890 430285
rect 513062 429738 513067 430335
rect 513067 429738 513669 430335
rect 513669 429738 513674 430335
rect 528964 430329 529594 430334
rect 522306 430301 522908 430306
rect 522306 429699 522311 430301
rect 522311 429699 522908 430301
rect 522306 429694 522908 429699
rect 528964 429699 529589 430329
rect 529589 429699 529594 430329
rect 528964 429694 529594 429699
rect 545778 430403 546408 430408
rect 545778 429773 545783 430403
rect 545783 429773 546408 430403
rect 545778 429768 546408 429773
rect 562796 429699 562801 430324
rect 562801 429699 563431 430324
rect 563431 429699 563436 430324
rect 562796 429694 563436 429699
rect 387904 427660 388014 427726
rect 392828 427679 392938 427745
rect 387914 427288 388024 427354
rect 392838 427307 392948 427373
rect 240181 425634 241179 426632
rect 324048 425639 325048 426639
rect 392312 425640 393310 426638
rect 356005 422225 356115 422291
rect 356015 421853 356125 421919
rect 72633 419889 73631 420887
rect 250982 420101 251980 421099
rect 336048 420100 337048 421100
rect 387417 420100 388417 421100
rect 25438 419176 25550 419288
rect 324544 417112 324654 417178
rect 336554 417037 336664 417103
rect 324554 416740 324664 416806
rect 336564 416665 336674 416731
rect 319471 415947 320013 415952
rect 252977 415912 253517 415917
rect 242014 415901 242565 415906
rect 242014 415365 242019 415901
rect 242019 415365 242560 415901
rect 242560 415365 242565 415901
rect 252977 415372 253512 415912
rect 253512 415372 253517 415912
rect 252977 415367 253517 415372
rect 258331 415876 258881 415881
rect 255268 415185 255273 415722
rect 255273 415185 255815 415722
rect 255815 415185 255820 415722
rect 258331 415341 258336 415876
rect 258336 415341 258876 415876
rect 258876 415341 258881 415876
rect 272927 415809 273479 415814
rect 272927 415272 272932 415809
rect 272932 415272 273474 415809
rect 273474 415272 273479 415809
rect 278445 415815 278997 415820
rect 278445 415278 278450 415815
rect 278450 415278 278992 415815
rect 278992 415278 278997 415815
rect 299131 415813 299683 415818
rect 293219 415789 293761 415794
rect 293219 415247 293756 415789
rect 293756 415247 293761 415789
rect 293219 415242 293761 415247
rect 299131 415276 299136 415813
rect 299136 415276 299678 415813
rect 299678 415276 299683 415813
rect 313349 415871 313891 415876
rect 313349 415329 313354 415871
rect 313354 415329 313891 415871
rect 319471 415405 320008 415947
rect 320008 415405 320013 415947
rect 319471 415400 320013 415405
rect 328164 415901 328706 415906
rect 328164 415359 328701 415901
rect 328701 415359 328706 415901
rect 328164 415354 328706 415359
rect 339880 415863 340422 415868
rect 313349 415324 313891 415329
rect 339880 415321 340417 415863
rect 340417 415321 340422 415863
rect 339880 415316 340422 415321
rect 255268 415180 255820 415185
rect 345550 414894 345978 416210
rect 393660 415927 394212 415932
rect 346912 415756 347022 415822
rect 346922 415384 347032 415450
rect 353568 415233 353573 415770
rect 353573 415233 354115 415770
rect 354115 415233 354120 415770
rect 373939 415845 374481 415850
rect 373939 415303 373944 415845
rect 373944 415303 374481 415845
rect 388622 415849 389164 415854
rect 373939 415298 374481 415303
rect 375345 415649 375887 415654
rect 353568 415228 354120 415233
rect 375345 415107 375882 415649
rect 375882 415107 375887 415649
rect 375345 415102 375887 415107
rect 388622 415307 389159 415849
rect 389159 415307 389164 415849
rect 388622 415302 389164 415307
rect 393660 415390 393665 415927
rect 393665 415390 394207 415927
rect 394207 415390 394212 415927
rect 560017 411206 560129 411318
rect 549018 408467 550016 409465
rect 549553 407130 549663 407196
rect 549543 406758 549653 406824
rect 355994 402190 356104 402256
rect 356004 401818 356114 401884
rect 324542 396322 324652 396388
rect 336579 396384 336689 396450
rect 324552 395950 324662 396016
rect 336589 396012 336699 396078
rect 346940 395078 347050 395144
rect 346950 394706 347060 394772
rect 322890 391347 323432 391352
rect 322890 390805 322895 391347
rect 322895 390805 323432 391347
rect 333087 391367 333629 391372
rect 333087 390825 333092 391367
rect 333092 390825 333629 391367
rect 333087 390820 333629 390825
rect 322890 390800 323432 390805
rect 334874 391309 335416 391314
rect 334874 390767 334879 391309
rect 334879 390767 335416 391309
rect 428496 391297 429048 391302
rect 367489 391193 368031 391198
rect 357695 391157 358237 391162
rect 334874 390762 335416 390767
rect 353560 390939 354112 390944
rect 118329 385378 123445 390494
rect 353560 390402 353565 390939
rect 353565 390402 354107 390939
rect 354107 390402 354112 390939
rect 357695 390615 358232 391157
rect 358232 390615 358237 391157
rect 357695 390610 358237 390615
rect 367489 390651 368026 391193
rect 368026 390651 368031 391193
rect 367489 390646 368031 390651
rect 385264 391169 385806 391174
rect 385264 390627 385269 391169
rect 385269 390627 385806 391169
rect 400432 391189 400974 391194
rect 400432 390647 400437 391189
rect 400437 390647 400974 391189
rect 428496 390760 428501 391297
rect 428501 390760 429043 391297
rect 429043 390760 429048 391297
rect 530390 391147 530932 391152
rect 490274 391105 490816 391110
rect 470032 391055 470574 391060
rect 446400 391049 446942 391054
rect 400432 390642 400974 390647
rect 385264 390622 385806 390627
rect 446400 390507 446937 391049
rect 446937 390507 446942 391049
rect 446400 390502 446942 390507
rect 470032 390513 470569 391055
rect 470569 390513 470574 391055
rect 470032 390508 470574 390513
rect 490274 390563 490811 391105
rect 490811 390563 490816 391105
rect 490274 390558 490816 390563
rect 510728 391075 511270 391080
rect 510728 390533 511265 391075
rect 511265 390533 511270 391075
rect 510728 390528 511270 390533
rect 530390 390605 530927 391147
rect 530927 390605 530932 391147
rect 530390 390600 530932 390605
rect 546398 391241 546960 391246
rect 546398 390679 546403 391241
rect 546403 390679 546960 391241
rect 546398 390674 546960 390679
rect 571232 391205 571794 391210
rect 571232 390643 571789 391205
rect 571789 390643 571794 391205
rect 571232 390638 571794 390643
rect 549570 388086 549680 388152
rect 549560 387714 549670 387780
rect 336049 386272 337047 387270
rect 549017 386271 550017 387271
rect 355974 382126 356084 382192
rect 355984 381754 356094 381820
rect 324049 380239 325047 381237
rect 548896 380238 549896 381238
rect 549368 379428 549478 379494
rect 549378 379056 549488 379122
rect 12758 378413 12868 378523
rect 65787 377991 66785 378989
rect 12757 377136 12869 377248
rect 333085 376209 333637 376214
rect 325770 376095 326312 376100
rect 25430 375954 25542 376066
rect 325770 375553 326307 376095
rect 326307 375553 326312 376095
rect 325770 375548 326312 375553
rect 333085 375672 333090 376209
rect 333090 375672 333632 376209
rect 333632 375672 333637 376209
rect 337328 375573 337333 376110
rect 337333 375573 337875 376110
rect 337875 375573 337880 376110
rect 337328 375568 337880 375573
rect 345676 376089 346228 376094
rect 345676 375552 345681 376089
rect 345681 375552 346223 376089
rect 346223 375552 346228 376089
rect 352330 375608 353838 376280
rect 526310 376169 526852 376174
rect 357689 376101 358231 376106
rect 357689 375559 358226 376101
rect 358226 375559 358231 376101
rect 357689 375554 358231 375559
rect 367489 376051 368031 376056
rect 367489 375509 368026 376051
rect 368026 375509 368031 376051
rect 367489 375504 368031 375509
rect 388564 375919 389106 375924
rect 388564 375377 389101 375919
rect 389101 375377 389106 375919
rect 388564 375372 389106 375377
rect 400420 376101 400962 376106
rect 400420 375559 400425 376101
rect 400425 375559 400962 376101
rect 400420 375554 400962 375559
rect 429154 376007 429696 376012
rect 429154 375465 429691 376007
rect 429691 375465 429696 376007
rect 429154 375460 429696 375465
rect 446406 376065 446948 376070
rect 446406 375523 446411 376065
rect 446411 375523 446948 376065
rect 446406 375518 446948 375523
rect 466544 376049 467086 376054
rect 466544 375507 466549 376049
rect 466549 375507 467086 376049
rect 466544 375502 467086 375507
rect 485504 376005 486046 376010
rect 485504 375463 485509 376005
rect 485509 375463 486046 376005
rect 485504 375458 486046 375463
rect 505738 375989 506280 375994
rect 505738 375447 506275 375989
rect 506275 375447 506280 375989
rect 505738 375442 506280 375447
rect 526310 375627 526847 376169
rect 526847 375627 526852 376169
rect 526310 375622 526852 375627
rect 552366 376047 552928 376052
rect 552366 375485 552923 376047
rect 552923 375485 552928 376047
rect 552366 375480 552928 375485
rect 562704 375559 562709 376116
rect 562709 375559 563271 376116
rect 563271 375559 563276 376116
rect 562704 375554 563276 375559
rect 118329 368964 123445 374080
rect 346926 373796 347036 373862
rect 346936 373424 347046 373490
rect 560038 364784 560150 364896
rect 549329 364242 549439 364308
rect 549339 363870 549449 363936
rect 356031 362143 356141 362209
rect 548897 362048 549895 363046
rect 356041 361771 356151 361837
rect 118329 354064 123445 359180
rect 346926 352946 347036 353012
rect 346936 352574 347046 352640
rect 356031 342140 356141 342206
rect 356041 341768 356151 341834
rect 13038 334573 13148 334683
rect 58671 334078 59669 335076
rect 13037 333914 13149 334026
rect 25372 332732 25484 332844
rect 347010 332350 347120 332416
rect 347020 331978 347130 332044
rect 118329 318742 123445 323858
rect 355955 322138 356065 322204
rect 355965 321766 356075 321832
rect 565606 319562 565718 319674
rect 365529 316852 366527 317850
rect 346982 310482 347092 310548
rect 346992 310110 347102 310176
rect 118329 304982 123445 310098
rect 348024 305644 348476 307618
rect 490719 307004 491268 307009
rect 357940 306779 358492 306784
rect 357940 306242 357945 306779
rect 357945 306242 358487 306779
rect 358487 306242 358492 306779
rect 370683 306263 370688 306807
rect 370688 306263 371237 306807
rect 371237 306263 371242 306807
rect 390695 306391 390700 306935
rect 390700 306391 391249 306935
rect 391249 306391 391254 306935
rect 390695 306386 391254 306391
rect 400259 306349 400264 306893
rect 400264 306349 400813 306893
rect 400813 306349 400818 306893
rect 400259 306344 400818 306349
rect 370683 306258 371242 306263
rect 430709 306113 430714 306657
rect 430714 306113 431263 306657
rect 431263 306113 431268 306657
rect 445435 306311 445440 306855
rect 445440 306311 445989 306855
rect 445989 306311 445994 306855
rect 445435 306306 445994 306311
rect 470723 306780 471272 306785
rect 470723 306231 471267 306780
rect 471267 306231 471272 306780
rect 470723 306226 471272 306231
rect 490719 306455 491263 307004
rect 491263 306455 491268 307004
rect 490719 306450 491268 306455
rect 510705 306896 511254 306901
rect 510705 306347 511249 306896
rect 511249 306347 511254 306896
rect 510705 306342 511254 306347
rect 569353 306806 569932 306811
rect 530681 306742 531230 306747
rect 530681 306193 530686 306742
rect 530686 306193 531230 306742
rect 530681 306188 531230 306193
rect 552162 306730 552719 306735
rect 552162 306173 552167 306730
rect 552167 306173 552719 306730
rect 569353 306242 569358 306806
rect 569358 306242 569927 306806
rect 569927 306242 569932 306806
rect 552162 306168 552719 306173
rect 430709 306108 431268 306113
rect 355993 302117 356103 302183
rect 356003 301745 356113 301811
rect 355562 295501 356560 296499
rect 549082 295500 550082 296500
rect 13045 291588 13155 291698
rect 49270 291103 50268 292101
rect 13044 290692 13156 290804
rect 25372 289510 25484 289622
rect 118329 288656 123445 293772
rect 549547 293375 549657 293441
rect 549557 293003 549667 293069
rect 346940 288824 347050 288890
rect 346950 288452 347060 288518
rect 345710 285614 346162 287588
rect 445447 287021 446006 287026
rect 400175 286903 400734 286908
rect 354036 286813 354578 286818
rect 354036 286271 354041 286813
rect 354041 286271 354578 286813
rect 390695 286691 391254 286696
rect 354036 286266 354578 286271
rect 370693 286607 371242 286612
rect 370693 286058 371237 286607
rect 371237 286058 371242 286607
rect 370693 286053 371242 286058
rect 390695 286147 390700 286691
rect 390700 286147 391249 286691
rect 391249 286147 391254 286691
rect 400175 286359 400180 286903
rect 400180 286359 400729 286903
rect 400729 286359 400734 286903
rect 430709 286809 431268 286814
rect 430709 286265 430714 286809
rect 430714 286265 431263 286809
rect 431263 286265 431268 286809
rect 445447 286477 445452 287021
rect 445452 286477 446001 287021
rect 446001 286477 446006 287021
rect 490719 286883 491268 286888
rect 470723 286753 471272 286758
rect 470723 286204 471267 286753
rect 471267 286204 471272 286753
rect 470723 286199 471272 286204
rect 490719 286334 491263 286883
rect 491263 286334 491268 286883
rect 490719 286329 491268 286334
rect 510705 286819 511254 286824
rect 510705 286270 511249 286819
rect 511249 286270 511254 286819
rect 510705 286265 511254 286270
rect 530691 286807 531240 286812
rect 530691 286258 531235 286807
rect 531235 286258 531240 286807
rect 530691 286253 531240 286258
rect 546315 286983 546872 286988
rect 546315 286426 546320 286983
rect 546320 286426 546872 286983
rect 546315 286421 546872 286426
rect 568313 286882 568892 286887
rect 568313 286318 568318 286882
rect 568318 286318 568887 286882
rect 568887 286318 568892 286882
rect 565656 275140 565768 275252
rect 549083 273465 550081 274463
rect 83455 268390 84455 269390
rect 425035 268390 426035 269390
rect 78269 266390 79269 267390
rect 423042 266390 424042 267390
rect 72632 264390 73632 265390
rect 421075 264390 422075 265390
rect 346898 264044 347008 264110
rect 346908 263672 347018 263738
rect 65786 262390 66786 263390
rect 419082 262390 420082 263390
rect 58670 260390 59670 261390
rect 417049 260390 418049 261390
rect 49269 258390 50269 259390
rect 415074 258390 416074 259390
rect 49269 256390 50269 257390
rect 413046 256390 414046 257390
rect 58938 254390 59938 255390
rect 411018 254390 412018 255390
rect 65894 252390 66894 253390
rect 409097 252390 410097 253390
rect 72906 250390 73906 251390
rect 407015 250390 408015 251390
rect 78414 248390 79414 249390
rect 405094 248390 406094 249390
rect 49270 247054 50268 248052
rect 25415 246488 25527 246600
rect 83668 246390 84668 247390
rect 403046 246391 404044 247389
rect 346982 242670 347092 242736
rect 346992 242298 347102 242364
rect 347010 222794 347120 222860
rect 347020 222422 347130 222488
rect 347982 208088 348448 213096
rect 346954 200966 347064 201032
rect 346964 200594 347074 200660
rect 570501 191330 575461 196290
rect 570414 181252 575532 186370
rect 346968 179932 347078 179998
rect 346978 179560 347088 179626
rect 13066 172742 18184 177860
rect 345722 172818 346188 177826
rect 13374 162744 18492 167862
rect 345698 162828 346164 167836
rect 346926 158544 347036 158610
rect 346936 158172 347046 158238
rect 334822 137385 335364 137390
rect 334822 136843 334827 137385
rect 334827 136843 335364 137385
rect 358800 137369 359342 137374
rect 346870 137198 346980 137264
rect 334822 136838 335364 136843
rect 346880 136826 346990 136892
rect 358800 136827 359337 137369
rect 359337 136827 359342 137369
rect 358800 136822 359342 136827
rect 58939 119856 59937 120854
rect 25403 118866 25515 118978
rect 346926 116064 347036 116130
rect 346936 115692 347046 115758
rect 334794 95639 335336 95644
rect 334794 95097 334799 95639
rect 334799 95097 335336 95639
rect 359148 95639 359690 95644
rect 346954 95454 347064 95520
rect 334794 95092 335336 95097
rect 346964 95082 347074 95148
rect 359148 95097 359685 95639
rect 359685 95097 359690 95639
rect 359148 95092 359690 95097
rect 12334 78417 12444 78527
rect 65895 78053 66893 79051
rect 12333 76826 12445 76938
rect 25414 75644 25526 75756
rect 346940 74772 347050 74838
rect 346950 74400 347060 74466
rect 12619 65518 12729 65628
rect 72907 65138 73905 66136
rect 14459 61906 14569 62016
rect 78415 61397 79413 62395
rect 16146 58483 16256 58593
rect 83669 58108 84667 59106
rect 90284 58752 91538 60006
rect 302584 59503 303126 59508
rect 111722 59361 112274 59366
rect 111722 58824 111727 59361
rect 111727 58824 112269 59361
rect 112269 58824 112274 59361
rect 133044 59371 133596 59376
rect 133044 58834 133049 59371
rect 133049 58834 133591 59371
rect 133591 58834 133596 59371
rect 240070 59381 240622 59386
rect 154602 59327 155154 59332
rect 154602 58790 154607 59327
rect 154607 58790 155149 59327
rect 155149 58790 155154 59327
rect 175808 59327 176360 59332
rect 175808 58790 175813 59327
rect 175813 58790 176355 59327
rect 176355 58790 176360 59327
rect 219084 59305 219636 59310
rect 197190 59283 197742 59288
rect 197190 58746 197195 59283
rect 197195 58746 197737 59283
rect 197737 58746 197742 59283
rect 219084 58768 219089 59305
rect 219089 58768 219631 59305
rect 219631 58768 219636 59305
rect 240070 58844 240075 59381
rect 240075 58844 240617 59381
rect 240617 58844 240622 59381
rect 260582 59379 261124 59384
rect 260582 58837 261119 59379
rect 261119 58837 261124 59379
rect 260582 58832 261124 58837
rect 281394 59135 281936 59140
rect 281394 58593 281931 59135
rect 281931 58593 281936 59135
rect 281394 58588 281936 58593
rect 302584 58961 303121 59503
rect 303121 58961 303126 59503
rect 302584 58956 303126 58961
rect 324122 59503 324664 59508
rect 324122 58961 324127 59503
rect 324127 58961 324664 59503
rect 324122 58956 324664 58961
rect 334718 54525 335270 54530
rect 334718 53988 334723 54525
rect 334723 53988 335265 54525
rect 335265 53988 335270 54525
rect 358810 54525 359352 54530
rect 358810 53983 359347 54525
rect 359347 53983 359352 54525
rect 358810 53978 359352 53983
rect 39900 52861 40872 52866
rect 39900 51904 39905 52861
rect 39905 51904 40867 52861
rect 40867 51904 40872 52861
rect 347010 51192 347120 51258
rect 347020 50820 347130 50886
rect 34106 48302 35106 49302
rect 346575 48303 347573 49301
rect 34578 42938 34688 43004
rect 34588 42566 34698 42632
rect 39650 36270 42762 39258
rect 48004 37365 48009 37902
rect 48009 37365 48551 37902
rect 48551 37365 48556 37902
rect 69298 37471 69303 38008
rect 69303 37471 69845 38008
rect 69845 37471 69850 38008
rect 69298 37466 69850 37471
rect 48004 37360 48556 37365
rect 90664 37153 90669 37690
rect 90669 37153 91211 37690
rect 91211 37153 91216 37690
rect 111724 37205 111729 37742
rect 111729 37205 112271 37742
rect 112271 37205 112276 37742
rect 111724 37200 112276 37205
rect 133056 37667 133598 37672
rect 90664 37148 91216 37153
rect 133056 37125 133593 37667
rect 133593 37125 133598 37667
rect 133056 37120 133598 37125
rect 154604 37293 154609 37830
rect 154609 37293 155151 37830
rect 155151 37293 155156 37830
rect 154604 37288 155156 37293
rect 175810 37293 175815 37830
rect 175815 37293 176357 37830
rect 176357 37293 176362 37830
rect 197192 37391 197197 37928
rect 197197 37391 197739 37928
rect 197739 37391 197744 37928
rect 197192 37386 197744 37391
rect 219086 37341 219091 37878
rect 219091 37341 219633 37878
rect 219633 37341 219638 37878
rect 219086 37336 219638 37341
rect 175810 37288 176362 37293
rect 240072 37781 240614 37786
rect 240072 37239 240077 37781
rect 240077 37239 240614 37781
rect 240072 37234 240614 37239
rect 260574 37719 261116 37724
rect 260574 37177 260579 37719
rect 260579 37177 261116 37719
rect 281386 37815 281928 37820
rect 281386 37273 281391 37815
rect 281391 37273 281928 37815
rect 302576 37919 303118 37924
rect 302576 37377 302581 37919
rect 302581 37377 303118 37919
rect 302576 37372 303118 37377
rect 324124 37867 324666 37872
rect 324124 37325 324129 37867
rect 324129 37325 324666 37867
rect 324124 37320 324666 37325
rect 281386 37268 281928 37273
rect 260574 37172 261116 37177
rect 12618 33604 12730 33716
rect 25408 32422 25520 32534
rect 34578 20840 34688 20906
rect 34588 20468 34698 20534
rect 21663 18795 21773 18905
rect 25446 18794 25558 18906
rect 22609 17957 22719 18067
rect 25438 17956 25550 18068
rect 24982 16174 25982 17174
rect 565200 16175 566198 17173
rect 14458 12182 14570 12294
rect 21662 11000 21774 11112
rect 344312 8478 344424 8590
rect 350866 8088 350978 8200
rect 345070 7742 345182 7854
rect 16145 7454 16257 7566
rect 348884 7144 348996 7256
rect 350238 7184 350350 7296
rect 349579 6628 349701 6633
rect 349579 6521 349584 6628
rect 349584 6521 349696 6628
rect 349696 6521 349701 6628
rect 22608 6272 22720 6384
rect 2637 3383 2747 3493
rect 34107 2949 35105 3947
rect 478105 3909 478215 4019
rect 482770 3903 482880 4013
rect 488006 3913 488116 4023
rect 2636 2726 2748 2838
rect 25358 1544 25470 1656
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 131021 648752 136109 649974
rect 131021 643712 131219 648752
rect 131021 638718 136109 643712
rect 131021 633694 131043 638718
rect 136067 633694 136109 638718
rect 118328 614123 123446 614371
rect 118328 580341 123446 609005
rect 131021 584235 136109 633694
rect 559614 644687 560614 645250
rect 559614 639595 559620 644687
rect 559614 634721 560614 639595
rect 560609 629629 560614 634721
rect 437075 605496 442175 629601
rect 449668 609029 449681 612029
rect 454751 609029 454786 612029
rect 378807 584076 379427 584275
rect 437075 584137 442163 605496
rect 396631 584080 397251 584136
rect 118328 577835 118354 580341
rect 123274 577835 123446 580341
rect 118328 542856 123446 577835
rect 118328 537740 118329 542856
rect 123445 537740 123446 542856
rect 118328 526346 123446 537740
rect 118328 521230 118329 526346
rect 123445 521230 123446 526346
rect 12229 508886 12341 508887
rect 12229 508776 12230 508886
rect 12340 508776 12341 508886
rect 12229 506915 12341 508776
rect 12228 506914 12342 506915
rect 12228 506802 12229 506914
rect 12341 506802 12342 506914
rect 12228 506801 12342 506802
rect 24982 505732 25982 520014
rect 24982 505620 25370 505732
rect 25482 505620 25982 505732
rect 13362 464768 13474 464769
rect 13362 464658 13363 464768
rect 13473 464658 13474 464768
rect 13362 463693 13474 464658
rect 13361 463692 13475 463693
rect 13361 463580 13362 463692
rect 13474 463580 13475 463692
rect 13361 463579 13475 463580
rect 24982 462510 25982 505620
rect 83455 509246 84455 509247
rect 83455 508248 83456 509246
rect 84454 508248 84455 509246
rect 24982 462398 25407 462510
rect 25519 462398 25982 462510
rect 24982 419288 25982 462398
rect 78269 465201 79269 465202
rect 78269 464203 78270 465201
rect 79268 464203 79269 465201
rect 24982 419176 25438 419288
rect 25550 419176 25982 419288
rect 12757 378523 12869 378524
rect 12757 378413 12758 378523
rect 12868 378413 12869 378523
rect 12757 377249 12869 378413
rect 12756 377248 12870 377249
rect 12756 377136 12757 377248
rect 12869 377136 12870 377248
rect 12756 377135 12870 377136
rect 24982 376066 25982 419176
rect 72632 420887 73632 420888
rect 72632 419889 72633 420887
rect 73631 419889 73632 420887
rect 24982 375954 25430 376066
rect 25542 375954 25982 376066
rect 13037 334683 13149 334684
rect 13037 334573 13038 334683
rect 13148 334573 13149 334683
rect 13037 334027 13149 334573
rect 13036 334026 13150 334027
rect 13036 333914 13037 334026
rect 13149 333914 13150 334026
rect 13036 333913 13150 333914
rect 24982 332844 25982 375954
rect 65786 378989 66786 378990
rect 65786 377991 65787 378989
rect 66785 377991 66786 378989
rect 24982 332732 25372 332844
rect 25484 332732 25982 332844
rect 13044 291698 13156 291699
rect 13044 291588 13045 291698
rect 13155 291588 13156 291698
rect 13044 290805 13156 291588
rect 13043 290804 13157 290805
rect 13043 290692 13044 290804
rect 13156 290692 13157 290804
rect 13043 290691 13157 290692
rect 24982 289622 25982 332732
rect 58670 335076 59670 335345
rect 58670 334078 58671 335076
rect 59669 334078 59670 335076
rect 24982 289510 25372 289622
rect 25484 289510 25982 289622
rect 24982 246600 25982 289510
rect 49269 292101 50269 292102
rect 49269 291103 49270 292101
rect 50268 291103 50269 292101
rect 49269 259391 50269 291103
rect 58670 261391 59670 334078
rect 65786 263391 66786 377991
rect 72632 265391 73632 419889
rect 78269 267391 79269 464203
rect 83455 269391 84455 508248
rect 118328 507810 123446 521230
rect 118328 502694 118329 507810
rect 123445 502694 123446 507810
rect 118328 467391 123446 502694
rect 131021 542664 136109 581875
rect 131021 537576 148716 542664
rect 131021 526232 136109 537576
rect 377567 534554 378187 578103
rect 378807 534486 379427 582061
rect 396631 534614 397251 582065
rect 397871 580068 398491 580202
rect 437075 578606 442163 581960
rect 449668 580116 454786 609029
rect 487606 603558 488608 603559
rect 487606 602558 487607 603558
rect 488607 602558 488608 603558
rect 487606 602557 488608 602558
rect 482432 597090 483434 597091
rect 482432 596090 482433 597090
rect 483433 596090 483434 597090
rect 482432 596089 483434 596090
rect 477775 590077 478777 590078
rect 477775 589077 477776 590077
rect 478776 589077 478777 590077
rect 477775 589076 478777 589077
rect 397871 534943 398491 578053
rect 437075 556351 442175 578606
rect 425729 535389 425795 535390
rect 425729 535325 425730 535389
rect 425794 535325 425795 535389
rect 425729 535324 425795 535325
rect 425732 533985 425792 535324
rect 423448 532949 423514 532950
rect 423448 532885 423449 532949
rect 423513 532885 423514 532949
rect 423448 532884 423514 532885
rect 355560 532597 356562 532598
rect 355560 531597 355561 532597
rect 356561 531597 356562 532597
rect 355560 531596 356562 531597
rect 131021 521144 148590 526232
rect 355561 522496 356561 531596
rect 423451 531548 423511 532884
rect 421585 530387 421651 530388
rect 421585 530323 421586 530387
rect 421650 530323 421651 530387
rect 421585 530322 421651 530323
rect 421588 528704 421648 530322
rect 419510 527947 419576 527948
rect 419510 527883 419511 527947
rect 419575 527883 419576 527947
rect 419510 527882 419576 527883
rect 419513 526413 419573 527882
rect 417544 525385 417610 525386
rect 417544 525321 417545 525385
rect 417609 525321 417610 525385
rect 417544 525320 417610 525321
rect 417547 523744 417607 525320
rect 415544 522945 415610 522946
rect 415544 522881 415545 522945
rect 415609 522881 415610 522945
rect 415544 522880 415610 522881
rect 355960 522111 356134 522496
rect 355960 522045 355991 522111
rect 356101 522045 356134 522111
rect 355960 522016 356134 522045
rect 355969 521739 356143 521771
rect 355969 521673 356001 521739
rect 356111 521725 356143 521739
rect 356111 521673 356144 521725
rect 355969 521420 356144 521673
rect 131021 507796 136109 521144
rect 131021 502708 148488 507796
rect 350838 504930 351066 504931
rect 350838 504704 350839 504930
rect 351065 504704 351066 504930
rect 350838 504703 351066 504704
rect 350184 502978 350412 502979
rect 350184 502752 350185 502978
rect 350411 502752 350412 502978
rect 350184 502751 350412 502752
rect 118328 416703 123446 465128
rect 131021 463295 136109 502708
rect 349514 496962 349742 496963
rect 349514 496736 349515 496962
rect 349741 496736 349742 496962
rect 349514 496735 349742 496736
rect 348838 494918 349066 494919
rect 348838 494692 348839 494918
rect 349065 494692 349066 494918
rect 348838 494691 349066 494692
rect 346573 487302 347575 487303
rect 346573 486302 346574 487302
rect 347574 486302 347575 487302
rect 346573 486301 347575 486302
rect 345008 484722 345236 484723
rect 345008 484496 345009 484722
rect 345235 484496 345236 484722
rect 345008 484495 345236 484496
rect 344280 482404 344508 482405
rect 344280 482178 344281 482404
rect 344507 482178 344508 482404
rect 344280 482177 344508 482178
rect 136035 461032 136109 463295
rect 131021 431115 136109 461032
rect 240179 457761 241181 457762
rect 240179 456761 240180 457761
rect 241180 456761 241181 457761
rect 240179 456760 241181 456761
rect 250980 457761 251982 457762
rect 250980 456761 250981 457761
rect 251981 456761 251982 457761
rect 250980 456760 251982 456761
rect 240180 456221 241180 456760
rect 240669 455915 240843 456221
rect 250981 456066 251981 456760
rect 240669 455849 240701 455915
rect 240811 455849 240843 455915
rect 240669 455817 240843 455849
rect 251391 455893 251565 456066
rect 251391 455827 251423 455893
rect 251533 455827 251565 455893
rect 251391 455795 251565 455827
rect 240678 455543 240852 455572
rect 240678 455477 240711 455543
rect 240821 455477 240852 455543
rect 240678 455053 240852 455477
rect 251400 455521 251574 455550
rect 251400 455455 251433 455521
rect 251543 455455 251574 455521
rect 251400 455081 251574 455455
rect 240180 434580 241180 455053
rect 240589 434398 240763 434580
rect 240589 434332 240621 434398
rect 240731 434332 240763 434398
rect 240589 434300 240763 434332
rect 250981 434199 251981 455081
rect 251374 434112 251548 434199
rect 240598 434026 240772 434055
rect 240598 433960 240631 434026
rect 240741 433960 240772 434026
rect 251374 434046 251406 434112
rect 251516 434046 251548 434112
rect 251374 434014 251548 434046
rect 240598 433653 240772 433960
rect 251383 433740 251557 433769
rect 251383 433674 251416 433740
rect 251526 433674 251557 433740
rect 136102 428852 136109 431115
rect 239401 430264 239403 430265
rect 239402 429713 239403 430264
rect 239401 429712 239403 429713
rect 118328 390494 123446 414440
rect 118328 385378 118329 390494
rect 123445 385378 123446 390494
rect 118328 374080 123446 385378
rect 118328 368964 118329 374080
rect 123445 368964 123446 374080
rect 118328 359180 123446 368964
rect 118328 354064 118329 359180
rect 123445 354064 123446 359180
rect 118328 323858 123446 354064
rect 118328 318742 118329 323858
rect 123445 318742 123446 323858
rect 118328 310098 123446 318742
rect 118328 304982 118329 310098
rect 123445 304982 123446 310098
rect 118328 293772 123446 304982
rect 118328 288656 118329 293772
rect 123445 288656 123446 293772
rect 83454 269390 84456 269391
rect 83454 268390 83455 269390
rect 84455 268390 84456 269390
rect 83454 268389 84456 268390
rect 78268 267390 79270 267391
rect 78268 266390 78269 267390
rect 79269 266390 79270 267390
rect 78268 266389 79270 266390
rect 72631 265390 73633 265391
rect 72631 264390 72632 265390
rect 73632 264390 73633 265390
rect 72631 264389 73633 264390
rect 65785 263390 66787 263391
rect 65785 262390 65786 263390
rect 66786 262390 66787 263390
rect 65785 262389 66787 262390
rect 58669 261390 59671 261391
rect 58669 260390 58670 261390
rect 59670 260390 59671 261390
rect 58669 260389 59671 260390
rect 49268 259390 50270 259391
rect 49268 258390 49269 259390
rect 50269 258390 50270 259390
rect 49268 258389 50270 258390
rect 49268 257390 50270 257391
rect 49268 256390 49269 257390
rect 50269 256390 50270 257390
rect 49268 256389 50270 256390
rect 49269 248052 50269 256389
rect 58937 255390 59939 255391
rect 58937 254390 58938 255390
rect 59938 254390 59939 255390
rect 58937 254389 59939 254390
rect 49269 247054 49270 248052
rect 50268 247054 50269 248052
rect 49269 247053 50269 247054
rect 24982 246488 25415 246600
rect 25527 246488 25982 246600
rect 24982 177806 25982 246488
rect 24982 167760 25982 172855
rect 24982 162809 25000 167760
rect 24982 118978 25982 162809
rect 58938 120854 59938 254389
rect 65893 253390 66895 253391
rect 65893 252390 65894 253390
rect 66894 252390 66895 253390
rect 65893 252389 66895 252390
rect 58938 119856 58939 120854
rect 59937 119856 59938 120854
rect 58938 119855 59938 119856
rect 24982 118866 25403 118978
rect 25515 118866 25982 118978
rect 12333 78527 12445 78528
rect 12333 78417 12334 78527
rect 12444 78417 12445 78527
rect 12333 76939 12445 78417
rect 12332 76938 12446 76939
rect 12332 76826 12333 76938
rect 12445 76826 12446 76938
rect 12332 76825 12446 76826
rect 24982 75756 25982 118866
rect 65894 79051 66894 252389
rect 72905 251390 73907 251391
rect 72905 250390 72906 251390
rect 73906 250390 73907 251390
rect 72905 250389 73907 250390
rect 65894 78053 65895 79051
rect 66893 78053 66894 79051
rect 65894 78052 66894 78053
rect 24982 75644 25414 75756
rect 25526 75644 25982 75756
rect 12618 65628 12730 65629
rect 12618 65518 12619 65628
rect 12729 65518 12730 65628
rect 12618 33717 12730 65518
rect 14458 62016 14570 62017
rect 14458 61906 14459 62016
rect 14569 61906 14570 62016
rect 12617 33716 12731 33717
rect 12617 33604 12618 33716
rect 12730 33604 12731 33716
rect 12617 33603 12731 33604
rect 14458 12295 14570 61906
rect 16145 58593 16257 58594
rect 16145 58483 16146 58593
rect 16256 58483 16257 58593
rect 14457 12294 14571 12295
rect 14457 12182 14458 12294
rect 14570 12182 14571 12294
rect 14457 12181 14571 12182
rect 16145 7567 16257 58483
rect 24982 32534 25982 75644
rect 72906 66152 73906 250389
rect 78413 249390 79415 249391
rect 78413 248390 78414 249390
rect 79414 248390 79415 249390
rect 78413 248389 79415 248390
rect 72894 66136 73915 66152
rect 72894 65138 72907 66136
rect 73905 65138 73915 66136
rect 72894 65128 73915 65138
rect 72906 65038 73906 65128
rect 78414 62431 79414 248389
rect 83667 247390 84669 247391
rect 83667 246390 83668 247390
rect 84668 246390 84669 247390
rect 83667 246389 84669 246390
rect 78386 62395 79436 62431
rect 78386 61397 78415 62395
rect 79413 61397 79436 62395
rect 78386 61367 79436 61397
rect 78414 61319 79414 61367
rect 83668 59115 84668 246389
rect 118328 177836 123446 288656
rect 131021 390412 136109 428852
rect 240180 426632 241180 433653
rect 251383 433419 251557 433674
rect 249229 429832 249230 429843
rect 249772 429832 249773 429843
rect 249229 429831 249773 429832
rect 240180 425634 240181 426632
rect 241179 425634 241180 426632
rect 240180 425633 241180 425634
rect 250981 421099 251981 433419
rect 252974 429826 252975 429827
rect 253527 429826 253528 429827
rect 252974 429825 253528 429826
rect 258342 430367 258344 430368
rect 258342 429817 258343 430367
rect 293218 430360 293220 430361
rect 278454 430348 278456 430349
rect 258342 429816 258344 429817
rect 272934 430294 273488 430295
rect 272934 430293 272935 430294
rect 273487 430293 273488 430294
rect 278454 429796 278455 430348
rect 293218 429808 293219 430360
rect 293218 429807 293220 429808
rect 299166 430260 299168 430261
rect 278454 429795 278456 429796
rect 299166 429708 299167 430260
rect 322089 430220 322091 430221
rect 299166 429707 299168 429708
rect 313342 429654 313343 429655
rect 313895 429654 313896 429655
rect 313342 429653 313896 429654
rect 319480 430162 319482 430163
rect 319480 429610 319481 430162
rect 322089 429668 322090 430220
rect 332863 429834 332864 429835
rect 333416 429834 333417 429835
rect 332863 429833 333417 429834
rect 335398 430258 335400 430259
rect 335398 429706 335399 430258
rect 335398 429705 335400 429706
rect 322089 429667 322091 429668
rect 319480 429609 319482 429610
rect 324047 426639 325049 426640
rect 324047 425639 324048 426639
rect 325048 425639 325049 426639
rect 324047 425638 325049 425639
rect 250981 420101 250982 421099
rect 251980 420101 251981 421099
rect 250981 420100 251981 420101
rect 324048 417422 325048 425638
rect 336047 421100 337049 421101
rect 336047 420100 336048 421100
rect 337048 420100 337049 421100
rect 336047 420099 337049 420100
rect 324512 417178 324686 417422
rect 336048 417263 337048 420099
rect 324512 417112 324544 417178
rect 324654 417112 324686 417178
rect 324512 417080 324686 417112
rect 336522 417103 336696 417263
rect 336522 417037 336554 417103
rect 336664 417037 336696 417103
rect 336522 417005 336696 417037
rect 324521 416806 324695 416835
rect 324521 416740 324554 416806
rect 324664 416740 324695 416806
rect 324521 416333 324695 416740
rect 336531 416731 336705 416760
rect 336531 416665 336564 416731
rect 336674 416665 336705 416731
rect 336531 416377 336705 416665
rect 319470 415952 319472 415953
rect 252976 415917 252978 415918
rect 252976 415367 252977 415917
rect 252976 415366 252978 415367
rect 255267 415722 255821 415723
rect 255267 415721 255268 415722
rect 255820 415721 255821 415722
rect 242013 415365 242014 415366
rect 242565 415365 242566 415366
rect 242013 415364 242566 415365
rect 313890 415876 313892 415877
rect 258330 415341 258331 415342
rect 258881 415341 258882 415342
rect 258330 415340 258882 415341
rect 278444 415278 278445 415279
rect 278997 415278 278998 415279
rect 278444 415277 278998 415278
rect 293218 415794 293220 415795
rect 272926 415272 272927 415273
rect 273479 415272 273480 415273
rect 272926 415271 273480 415272
rect 293218 415242 293219 415794
rect 313891 415324 313892 415876
rect 319470 415400 319471 415952
rect 319470 415399 319472 415400
rect 313890 415323 313892 415324
rect 299130 415276 299131 415277
rect 299683 415276 299684 415277
rect 299130 415275 299684 415276
rect 293218 415241 293220 415242
rect 324048 396630 325048 416333
rect 328163 415906 328165 415907
rect 328163 415354 328164 415906
rect 328163 415353 328165 415354
rect 324510 396388 324684 396630
rect 336048 396599 337048 416377
rect 339879 415868 339881 415869
rect 339879 415316 339880 415868
rect 339879 415315 339881 415316
rect 324510 396322 324542 396388
rect 324652 396322 324684 396388
rect 336547 396450 336721 396599
rect 336547 396384 336579 396450
rect 336689 396384 336721 396450
rect 336547 396352 336721 396384
rect 324510 396290 324684 396322
rect 336556 396078 336730 396107
rect 324519 396016 324693 396045
rect 324519 395950 324552 396016
rect 324662 395950 324693 396016
rect 324519 395566 324693 395950
rect 336556 396012 336589 396078
rect 336699 396012 336730 396078
rect 336556 395728 336730 396012
rect 323431 391352 323433 391353
rect 323432 390800 323433 391352
rect 323431 390799 323433 390800
rect 131021 385324 168402 390412
rect 131021 374300 136109 385324
rect 324048 381237 325048 395566
rect 333628 391372 333630 391373
rect 333629 390820 333630 391372
rect 333628 390819 333630 390820
rect 335415 391314 335417 391315
rect 335416 390762 335417 391314
rect 335415 390761 335417 390762
rect 336048 387270 337048 395728
rect 336048 386272 336049 387270
rect 337047 386272 337048 387270
rect 336048 386271 337048 386272
rect 324048 380239 324049 381237
rect 325047 380239 325048 381237
rect 324048 380238 325048 380239
rect 325769 376100 325771 376101
rect 325769 375548 325770 376100
rect 333084 375672 333085 375673
rect 333637 375672 333638 375673
rect 333084 375671 333638 375672
rect 337327 376110 337881 376111
rect 337327 376109 337328 376110
rect 337880 376109 337881 376110
rect 325769 375547 325771 375548
rect 131021 369212 168402 374300
rect 131021 359400 136109 369212
rect 131021 354312 168402 359400
rect 131021 323844 136109 354312
rect 131021 318756 168402 323844
rect 131021 310084 136109 318756
rect 131021 304996 168402 310084
rect 131021 293990 136109 304996
rect 131021 288902 168402 293990
rect 131021 213150 136109 288902
rect 123398 172766 123446 177836
rect 118328 167838 123446 172766
rect 123264 162768 123446 167838
rect 118328 160061 123446 162768
rect 332563 177836 337681 177860
rect 332563 172766 332587 177836
rect 337657 172766 337681 177836
rect 332563 137390 337681 172766
rect 332563 136838 334822 137390
rect 335364 136838 337681 137390
rect 332563 95644 337681 136838
rect 332563 95092 334794 95644
rect 335336 95092 337681 95644
rect 332563 61843 337681 95092
rect 90283 60006 91539 60007
rect 83660 59106 84676 59115
rect 83660 58108 83669 59106
rect 84667 58108 84676 59106
rect 90283 58752 90284 60006
rect 91538 58752 91539 60006
rect 302583 59508 302585 59509
rect 133043 58834 133044 58835
rect 133596 58834 133597 58835
rect 133043 58833 133597 58834
rect 111721 58824 111722 58825
rect 112274 58824 112275 58825
rect 111721 58823 112275 58824
rect 154601 58790 154602 58791
rect 155154 58790 155155 58791
rect 154601 58789 155155 58790
rect 175807 58790 175808 58791
rect 176360 58790 176361 58791
rect 175807 58789 176361 58790
rect 90283 58751 91539 58752
rect 240069 58844 240070 58845
rect 240622 58844 240623 58845
rect 240069 58843 240623 58844
rect 260581 59384 260583 59385
rect 260581 58832 260582 59384
rect 260581 58831 260583 58832
rect 281393 59140 281395 59141
rect 219083 58768 219084 58769
rect 219636 58768 219637 58769
rect 219083 58767 219637 58768
rect 197189 58746 197190 58747
rect 197742 58746 197743 58747
rect 197189 58745 197743 58746
rect 281393 58588 281394 59140
rect 302583 58956 302584 59508
rect 302583 58955 302585 58956
rect 324663 59508 324665 59509
rect 324664 58956 324665 59508
rect 324663 58955 324665 58956
rect 281393 58587 281395 58588
rect 83660 58099 84676 58108
rect 332563 54530 337681 56725
rect 332563 53988 334718 54530
rect 335270 53988 337681 54530
rect 332563 52541 337681 53988
rect 39899 51904 39900 51905
rect 40872 51904 40873 51905
rect 39899 51903 40873 51904
rect 34105 49302 35107 49303
rect 34105 48302 34106 49302
rect 35106 48302 35107 49302
rect 34105 48301 35107 48302
rect 34106 43300 35106 48301
rect 34547 43004 34721 43300
rect 34547 42938 34578 43004
rect 34688 42938 34721 43004
rect 34547 42909 34721 42938
rect 34556 42632 34730 42664
rect 34556 42566 34588 42632
rect 34698 42618 34730 42632
rect 34698 42566 34731 42618
rect 34556 42468 34731 42566
rect 24982 32422 25408 32534
rect 25520 32422 25982 32534
rect 24982 18906 25982 32422
rect 34106 21194 35106 42468
rect 39649 39258 42763 39259
rect 39649 36270 39650 39258
rect 42762 36270 42763 39258
rect 69297 38008 69851 38009
rect 69297 38007 69298 38008
rect 69850 38007 69851 38008
rect 48003 37902 48557 37903
rect 48003 37901 48004 37902
rect 48556 37901 48557 37902
rect 197191 37928 197745 37929
rect 197191 37927 197192 37928
rect 197744 37927 197745 37928
rect 154603 37830 155157 37831
rect 154603 37829 154604 37830
rect 155156 37829 155157 37830
rect 111723 37742 112277 37743
rect 111723 37741 111724 37742
rect 112276 37741 112277 37742
rect 90663 37690 91217 37691
rect 90663 37689 90664 37690
rect 91216 37689 91217 37690
rect 133055 37672 133057 37673
rect 133055 37120 133056 37672
rect 175809 37830 176363 37831
rect 175809 37829 175810 37830
rect 176362 37829 176363 37830
rect 303117 37924 303119 37925
rect 219085 37878 219639 37879
rect 219085 37877 219086 37878
rect 219638 37877 219639 37878
rect 281927 37820 281929 37821
rect 240613 37786 240615 37787
rect 240614 37234 240615 37786
rect 240613 37233 240615 37234
rect 261115 37724 261117 37725
rect 261116 37172 261117 37724
rect 281928 37268 281929 37820
rect 303118 37372 303119 37924
rect 303117 37371 303119 37372
rect 324665 37872 324667 37873
rect 324666 37320 324667 37872
rect 324665 37319 324667 37320
rect 281927 37267 281929 37268
rect 261115 37171 261117 37172
rect 133055 37119 133057 37120
rect 39649 36269 42763 36270
rect 34547 20906 34721 21194
rect 34547 20840 34578 20906
rect 34688 20840 34721 20906
rect 34547 20811 34721 20840
rect 34556 20534 34730 20566
rect 34556 20468 34588 20534
rect 34698 20520 34730 20534
rect 34698 20468 34731 20520
rect 34556 20368 34731 20468
rect 21662 18905 21774 18906
rect 21662 18795 21663 18905
rect 21773 18795 21774 18905
rect 21662 11113 21774 18795
rect 24982 18794 25446 18906
rect 25558 18794 25982 18906
rect 24982 18068 25982 18794
rect 22608 18067 22720 18068
rect 22608 17957 22609 18067
rect 22719 17957 22720 18067
rect 21661 11112 21775 11113
rect 21661 11000 21662 11112
rect 21774 11000 21775 11112
rect 21661 10999 21775 11000
rect 16144 7566 16258 7567
rect 16144 7454 16145 7566
rect 16257 7454 16258 7566
rect 16144 7453 16258 7454
rect 22608 6385 22720 17957
rect 24982 17956 25438 18068
rect 25550 17956 25982 18068
rect 24982 17175 25982 17956
rect 24981 17174 25983 17175
rect 24981 16174 24982 17174
rect 25982 16174 25983 17174
rect 24981 16173 25983 16174
rect 22607 6384 22721 6385
rect 22607 6272 22608 6384
rect 22720 6272 22721 6384
rect 22607 6271 22721 6272
rect 2636 3493 2748 3494
rect 2636 3383 2637 3493
rect 2747 3383 2748 3493
rect 2636 2839 2748 3383
rect 2635 2838 2749 2839
rect 2635 2726 2636 2838
rect 2748 2726 2749 2838
rect 2635 2725 2749 2726
rect 25358 1657 25470 16173
rect 34106 3947 35106 20368
rect 344281 12006 344507 482177
rect 345009 12006 345235 484495
rect 346574 478576 347574 486301
rect 346951 478318 347125 478576
rect 346951 478252 346982 478318
rect 347092 478252 347125 478318
rect 346951 478223 347125 478252
rect 346960 477946 347134 477978
rect 346960 477880 346992 477946
rect 347102 477932 347134 477946
rect 347102 477880 347135 477932
rect 346960 477688 347135 477880
rect 346574 457342 347574 477688
rect 346965 457064 347139 457342
rect 346965 456998 346996 457064
rect 347106 456998 347139 457064
rect 346965 456969 347139 456998
rect 346974 456692 347148 456724
rect 346974 456626 347006 456692
rect 347116 456678 347148 456692
rect 347116 456626 347149 456678
rect 346974 456454 347149 456626
rect 346574 436728 347574 456454
rect 346937 436456 347111 436728
rect 346937 436390 346968 436456
rect 347078 436390 347111 436456
rect 346937 436361 347111 436390
rect 346946 436084 347120 436116
rect 346946 436018 346978 436084
rect 347088 436070 347120 436084
rect 347088 436018 347121 436070
rect 346946 435840 347121 436018
rect 345549 416210 345979 416211
rect 345549 414894 345550 416210
rect 345978 414894 345979 416210
rect 346574 416116 347574 435840
rect 348093 430698 348523 430699
rect 348093 429382 348094 430698
rect 348522 429382 348523 430698
rect 348093 429381 348523 429382
rect 346881 415822 347055 416116
rect 346881 415756 346912 415822
rect 347022 415756 347055 415822
rect 346881 415727 347055 415756
rect 346890 415450 347064 415482
rect 346890 415384 346922 415450
rect 347032 415436 347064 415450
rect 347032 415384 347065 415436
rect 346890 415228 347065 415384
rect 345549 414893 345979 414894
rect 346574 395422 347574 415228
rect 346909 395144 347083 395422
rect 346909 395078 346940 395144
rect 347050 395078 347083 395144
rect 346909 395049 347083 395078
rect 346918 394772 347092 394804
rect 346918 394706 346950 394772
rect 347060 394758 347092 394772
rect 347060 394706 347093 394758
rect 346918 394534 347093 394706
rect 345675 375552 345676 375553
rect 346228 375552 346229 375553
rect 345675 375551 346229 375552
rect 346574 374160 347574 394534
rect 346895 373862 347069 374160
rect 346895 373796 346926 373862
rect 347036 373796 347069 373862
rect 346895 373767 347069 373796
rect 346904 373490 347078 373522
rect 346904 373424 346936 373490
rect 347046 373476 347078 373490
rect 347046 373424 347079 373476
rect 346904 373272 347079 373424
rect 346574 353278 347574 373272
rect 346895 353012 347069 353278
rect 346895 352946 346926 353012
rect 347036 352946 347069 353012
rect 346895 352917 347069 352946
rect 346904 352640 347078 352672
rect 346904 352574 346936 352640
rect 347046 352626 347078 352640
rect 347046 352574 347079 352626
rect 346904 352390 347079 352574
rect 346574 332692 347574 352390
rect 346979 332416 347153 332692
rect 346979 332350 347010 332416
rect 347120 332350 347153 332416
rect 346979 332321 347153 332350
rect 346988 332044 347162 332076
rect 346988 331978 347020 332044
rect 347130 332030 347162 332044
rect 347130 331978 347163 332030
rect 346988 331804 347163 331978
rect 346574 310824 347574 331804
rect 346951 310548 347125 310824
rect 346951 310482 346982 310548
rect 347092 310482 347125 310548
rect 346951 310453 347125 310482
rect 346960 310176 347134 310208
rect 346960 310110 346992 310176
rect 347102 310162 347134 310176
rect 347102 310110 347135 310162
rect 346960 309936 347135 310110
rect 346574 289160 347574 309936
rect 348023 307618 348477 307619
rect 348023 305644 348024 307618
rect 348476 305644 348477 307618
rect 348023 305643 348477 305644
rect 346909 288890 347083 289160
rect 346909 288824 346940 288890
rect 347050 288824 347083 288890
rect 346909 288795 347083 288824
rect 346918 288518 347092 288550
rect 346918 288452 346950 288518
rect 347060 288504 347092 288518
rect 347060 288452 347093 288504
rect 346918 288272 347093 288452
rect 345709 287588 346163 287589
rect 345709 285614 345710 287588
rect 346162 285614 346163 287588
rect 345709 285613 346163 285614
rect 346574 264386 347574 288272
rect 346867 264110 347041 264386
rect 346867 264044 346898 264110
rect 347008 264044 347041 264110
rect 346867 264015 347041 264044
rect 346876 263738 347050 263770
rect 346876 263672 346908 263738
rect 347018 263724 347050 263738
rect 347018 263672 347051 263724
rect 346876 263498 347051 263672
rect 346574 243026 347574 263498
rect 346951 242736 347125 243026
rect 346951 242670 346982 242736
rect 347092 242670 347125 242736
rect 346951 242641 347125 242670
rect 346960 242364 347134 242396
rect 346960 242298 346992 242364
rect 347102 242350 347134 242364
rect 347102 242298 347135 242350
rect 346960 242138 347135 242298
rect 346574 223146 347574 242138
rect 346979 222860 347153 223146
rect 346979 222794 347010 222860
rect 347120 222794 347153 222860
rect 346979 222765 347153 222794
rect 346988 222488 347162 222520
rect 346988 222422 347020 222488
rect 347130 222474 347162 222488
rect 347130 222422 347163 222474
rect 346988 222258 347163 222422
rect 346574 201336 347574 222258
rect 347981 213096 348449 213097
rect 347981 208088 347982 213096
rect 348448 208088 348449 213096
rect 347981 208087 348449 208088
rect 346923 201032 347097 201336
rect 346923 200966 346954 201032
rect 347064 200966 347097 201032
rect 346923 200937 347097 200966
rect 346932 200660 347106 200692
rect 346932 200594 346964 200660
rect 347074 200646 347106 200660
rect 347074 200594 347107 200646
rect 346932 200448 347107 200594
rect 346574 180300 347574 200448
rect 346937 179998 347111 180300
rect 346937 179932 346968 179998
rect 347078 179932 347111 179998
rect 346937 179903 347111 179932
rect 346946 179626 347120 179658
rect 346946 179560 346978 179626
rect 347088 179612 347120 179626
rect 347088 179560 347121 179612
rect 346946 179412 347121 179560
rect 345721 177826 346189 177827
rect 345721 172818 345722 177826
rect 346188 172818 346189 177826
rect 345721 172817 346189 172818
rect 345697 167836 346165 167837
rect 345697 162828 345698 167836
rect 346164 162828 346165 167836
rect 345697 162827 346165 162828
rect 346574 158876 347574 179412
rect 346895 158610 347069 158876
rect 346895 158544 346926 158610
rect 347036 158544 347069 158610
rect 346895 158515 347069 158544
rect 346904 158238 347078 158270
rect 346904 158172 346936 158238
rect 347046 158224 347078 158238
rect 347046 158172 347079 158224
rect 346904 157988 347079 158172
rect 346574 137564 347574 157988
rect 346839 137264 347013 137564
rect 346839 137198 346870 137264
rect 346980 137198 347013 137264
rect 346839 137169 347013 137198
rect 346848 136892 347022 136924
rect 346848 136826 346880 136892
rect 346990 136878 347022 136892
rect 346990 136826 347023 136878
rect 346848 136676 347023 136826
rect 346574 116416 347574 136676
rect 346895 116130 347069 116416
rect 346895 116064 346926 116130
rect 347036 116064 347069 116130
rect 346895 116035 347069 116064
rect 346904 115758 347078 115790
rect 346904 115692 346936 115758
rect 347046 115744 347078 115758
rect 347046 115692 347079 115744
rect 346904 115528 347079 115692
rect 346574 95818 347574 115528
rect 346923 95520 347097 95818
rect 346923 95454 346954 95520
rect 347064 95454 347097 95520
rect 346923 95425 347097 95454
rect 346932 95148 347106 95180
rect 346932 95082 346964 95148
rect 347074 95134 347106 95148
rect 347074 95082 347107 95134
rect 346932 94930 347107 95082
rect 346574 75112 347574 94930
rect 346909 74838 347083 75112
rect 346909 74772 346940 74838
rect 347050 74772 347083 74838
rect 346909 74743 347083 74772
rect 346918 74466 347092 74498
rect 346918 74400 346950 74466
rect 347060 74452 347092 74466
rect 347060 74400 347093 74452
rect 346918 74224 347093 74400
rect 346574 51540 347574 74224
rect 346979 51258 347153 51540
rect 346979 51192 347010 51258
rect 347120 51192 347153 51258
rect 346979 51163 347153 51192
rect 346988 50886 347162 50918
rect 346988 50820 347020 50886
rect 347130 50872 347162 50886
rect 347130 50820 347163 50872
rect 346988 50652 347163 50820
rect 346574 49301 347574 50652
rect 346574 48303 346575 49301
rect 347573 48303 347574 49301
rect 346574 48302 347574 48303
rect 348839 12006 349065 494691
rect 349515 12006 349741 496735
rect 350185 12006 350411 502751
rect 350839 12006 351065 504703
rect 355561 502549 356561 521420
rect 415547 521278 415607 522880
rect 413515 520383 413581 520384
rect 413515 520319 413516 520383
rect 413580 520319 413581 520383
rect 413515 520318 413581 520319
rect 413518 518914 413578 520318
rect 411486 517943 411552 517944
rect 411486 517879 411487 517943
rect 411551 517879 411552 517943
rect 411486 517878 411552 517879
rect 365527 517349 366529 517350
rect 365527 516349 365528 517349
rect 366528 516349 366529 517349
rect 365527 516348 366529 516349
rect 355925 502202 356099 502549
rect 355925 502136 355956 502202
rect 356066 502136 356099 502202
rect 355925 502107 356099 502136
rect 355934 501830 356108 501862
rect 355934 501764 355966 501830
rect 356076 501816 356108 501830
rect 356076 501764 356109 501816
rect 355934 501569 356109 501764
rect 355561 482593 356561 501569
rect 360437 484610 360438 484611
rect 360990 484610 360991 484611
rect 360437 484609 360991 484610
rect 355987 482258 356161 482593
rect 355987 482192 356018 482258
rect 356128 482192 356161 482258
rect 355987 482163 356161 482192
rect 355996 481886 356170 481918
rect 355996 481820 356028 481886
rect 356138 481872 356170 481886
rect 356138 481820 356171 481872
rect 355996 481593 356171 481820
rect 353317 472986 353319 472987
rect 353318 472434 353319 472986
rect 353317 472433 353319 472434
rect 355561 462516 356561 481593
rect 355995 462238 356169 462516
rect 355995 462172 356026 462238
rect 356136 462172 356169 462238
rect 355995 462143 356169 462172
rect 356004 461866 356178 461898
rect 356004 461800 356036 461866
rect 356146 461852 356178 461866
rect 356146 461800 356179 461852
rect 356004 461614 356179 461800
rect 355561 442547 356561 461614
rect 355969 442245 356143 442547
rect 355969 442179 356000 442245
rect 356110 442179 356143 442245
rect 355969 442150 356143 442179
rect 355978 441873 356152 441905
rect 355978 441807 356010 441873
rect 356120 441859 356152 441873
rect 356120 441807 356153 441859
rect 355978 441628 356153 441807
rect 354351 430264 354905 430265
rect 354351 430263 354352 430264
rect 354904 430263 354905 430264
rect 355561 422597 356561 441628
rect 359995 429902 359996 429903
rect 360548 429902 360549 429903
rect 359995 429901 360549 429902
rect 362165 430438 362719 430439
rect 362165 430437 362166 430438
rect 362718 430437 362719 430438
rect 355969 422291 356148 422597
rect 355969 422225 356005 422291
rect 356115 422225 356148 422291
rect 355969 422196 356148 422225
rect 355969 422187 356144 422196
rect 355983 421919 356157 421951
rect 355983 421853 356015 421919
rect 356125 421905 356157 421919
rect 356125 421853 356158 421905
rect 355983 421667 356158 421853
rect 353567 415770 354121 415771
rect 353567 415769 353568 415770
rect 354120 415769 354121 415770
rect 355561 402555 356561 421667
rect 355958 402256 356137 402555
rect 355958 402190 355994 402256
rect 356104 402190 356137 402256
rect 355958 402161 356137 402190
rect 355958 402139 356133 402161
rect 355972 401884 356146 401916
rect 355972 401818 356004 401884
rect 356114 401870 356146 401884
rect 356114 401818 356147 401870
rect 355972 401602 356147 401818
rect 353559 390402 353560 390403
rect 354112 390402 354113 390403
rect 353559 390401 354113 390402
rect 355561 382488 356561 401602
rect 357694 391162 357696 391163
rect 357694 390610 357695 391162
rect 357694 390609 357696 390610
rect 355938 382192 356117 382488
rect 355938 382126 355974 382192
rect 356084 382126 356117 382192
rect 355938 382098 356117 382126
rect 355952 381820 356126 381852
rect 355952 381754 355984 381820
rect 356094 381806 356126 381820
rect 356094 381754 356127 381806
rect 355952 381590 356127 381754
rect 352329 376280 353839 376281
rect 352329 375608 352330 376280
rect 353838 375608 353839 376280
rect 352329 375607 353839 375608
rect 355561 362485 356561 381590
rect 357688 376106 357690 376107
rect 357688 375554 357689 376106
rect 357688 375553 357690 375554
rect 355995 362209 356174 362485
rect 355995 362143 356031 362209
rect 356141 362143 356174 362209
rect 355995 362122 356174 362143
rect 356009 361837 356183 361869
rect 356009 361771 356041 361837
rect 356151 361823 356183 361837
rect 356151 361771 356184 361823
rect 356009 361624 356184 361771
rect 355561 342536 356561 361624
rect 355995 342206 356174 342536
rect 355995 342140 356031 342206
rect 356141 342140 356174 342206
rect 355995 342122 356174 342140
rect 356009 341834 356183 341866
rect 356009 341768 356041 341834
rect 356151 341820 356183 341834
rect 356151 341768 356184 341820
rect 356009 341633 356184 341768
rect 355561 322489 356561 341633
rect 355919 322204 356098 322489
rect 355919 322138 355955 322204
rect 356065 322138 356098 322204
rect 355919 322119 356098 322138
rect 355933 321832 356107 321864
rect 355933 321766 355965 321832
rect 356075 321818 356107 321832
rect 356075 321766 356108 321818
rect 355933 321626 356108 321766
rect 355561 302545 356561 321626
rect 365528 317850 366528 516348
rect 411489 516312 411549 517878
rect 409482 515381 409548 515382
rect 409482 515317 409483 515381
rect 409547 515317 409548 515381
rect 409482 515316 409548 515317
rect 409485 513846 409545 515316
rect 407541 512941 407607 512942
rect 407541 512877 407542 512941
rect 407606 512877 407607 512941
rect 407541 512876 407607 512877
rect 407544 511313 407604 512876
rect 405501 510379 405567 510380
rect 405501 510315 405502 510379
rect 405566 510315 405567 510379
rect 405501 510314 405567 510315
rect 405504 508779 405564 510314
rect 373152 504829 374155 504968
rect 373155 504707 374155 504829
rect 373155 504637 373642 504707
rect 373712 504637 374155 504707
rect 373155 490885 374155 504637
rect 373583 490674 373758 490885
rect 373583 490622 373616 490674
rect 373584 490608 373616 490622
rect 373726 490608 373758 490674
rect 373584 490576 373758 490608
rect 373593 490302 373767 490331
rect 373593 490236 373626 490302
rect 373736 490236 373767 490302
rect 373593 489858 373767 490236
rect 373155 476015 374155 489858
rect 375483 485284 376037 485285
rect 375483 485283 375484 485284
rect 376036 485283 376037 485284
rect 373155 475017 373156 476015
rect 374154 475017 374155 476015
rect 373155 475016 374155 475017
rect 377567 467291 378187 508101
rect 377567 465237 378187 465285
rect 378807 463289 379427 508379
rect 387913 507817 387979 507818
rect 387913 507753 387914 507817
rect 387978 507753 387979 507817
rect 387913 507752 387979 507753
rect 382734 504762 383734 505017
rect 387916 504968 387976 507752
rect 382734 504692 383216 504762
rect 383280 504692 383734 504762
rect 382734 490881 383734 504692
rect 387425 490889 388425 504968
rect 392312 504721 393312 504968
rect 392312 504651 392784 504721
rect 392848 504651 393312 504721
rect 392312 504631 393312 504651
rect 392311 504474 393312 504631
rect 392311 490902 393311 504474
rect 383235 490672 383410 490881
rect 383235 490620 383268 490672
rect 383236 490606 383268 490620
rect 383378 490606 383410 490672
rect 387873 490753 388047 490889
rect 387873 490687 387905 490753
rect 388015 490687 388047 490753
rect 387873 490655 388047 490687
rect 392776 490767 392950 490902
rect 392776 490701 392808 490767
rect 392918 490701 392950 490767
rect 392776 490669 392950 490701
rect 383236 490574 383410 490606
rect 387882 490381 388056 490410
rect 383245 490300 383419 490329
rect 383245 490234 383278 490300
rect 383388 490234 383419 490300
rect 383245 489881 383419 490234
rect 387882 490315 387915 490381
rect 388025 490315 388056 490381
rect 387882 490003 388056 490315
rect 392785 490395 392959 490424
rect 392785 490329 392818 490395
rect 392928 490329 392959 490395
rect 392785 490010 392959 490329
rect 382734 480108 383734 489881
rect 387425 485346 388425 490003
rect 386089 485208 386643 485209
rect 386089 485207 386090 485208
rect 386642 485207 386643 485208
rect 387423 484741 388425 485346
rect 382734 479110 382735 480108
rect 383733 479110 383734 480108
rect 382734 479109 383734 479110
rect 380561 473164 380563 473165
rect 380561 472612 380562 473164
rect 380561 472611 380563 472612
rect 387423 469942 388423 484741
rect 390323 484674 390324 484675
rect 390876 484674 390877 484675
rect 390323 484673 390877 484674
rect 389485 473078 390039 473079
rect 389485 473077 389486 473078
rect 390038 473077 390039 473078
rect 392311 469962 393311 490010
rect 394691 473152 395245 473153
rect 394691 473151 394692 473152
rect 395244 473151 395245 473152
rect 387882 469789 388056 469942
rect 387882 469723 387914 469789
rect 388024 469723 388056 469789
rect 387882 469691 388056 469723
rect 392774 469789 392948 469962
rect 392774 469723 392806 469789
rect 392916 469723 392948 469789
rect 392774 469691 392948 469723
rect 387891 469417 388065 469446
rect 387891 469351 387924 469417
rect 388034 469351 388065 469417
rect 387891 468965 388065 469351
rect 392783 469417 392957 469446
rect 392783 469351 392816 469417
rect 392926 469351 392957 469417
rect 387423 448891 388423 468965
rect 392783 468944 392957 469351
rect 392311 449136 393311 468944
rect 396631 463277 397251 507704
rect 397871 467290 398491 507962
rect 403540 507817 403606 507818
rect 403540 507753 403541 507817
rect 403605 507753 403606 507817
rect 403540 507752 403606 507753
rect 403543 506068 403603 507752
rect 400217 484644 400218 484645
rect 400770 484644 400771 484645
rect 400217 484643 400771 484644
rect 400585 473104 401139 473105
rect 400585 473103 400586 473104
rect 401138 473103 401139 473104
rect 387843 448769 388017 448891
rect 387843 448703 387875 448769
rect 387985 448703 388017 448769
rect 392747 448837 392944 449136
rect 392747 448771 392796 448837
rect 392906 448771 392944 448837
rect 392747 448733 392944 448771
rect 387843 448671 388017 448703
rect 392773 448465 392947 448494
rect 387852 448397 388026 448426
rect 387852 448331 387885 448397
rect 387995 448331 388026 448397
rect 387852 448061 388026 448331
rect 392773 448399 392806 448465
rect 392916 448399 392947 448465
rect 386469 430292 386471 430293
rect 373954 430196 373956 430197
rect 373954 429644 373955 430196
rect 386470 429740 386471 430292
rect 386469 429739 386471 429740
rect 375346 429658 375347 429659
rect 375899 429658 375900 429659
rect 375346 429657 375900 429658
rect 373954 429643 373956 429644
rect 387423 427905 388423 448061
rect 392773 447981 392947 448399
rect 391741 430376 391743 430377
rect 391742 429824 391743 430376
rect 391741 429823 391743 429824
rect 392311 427912 393311 447981
rect 387872 427726 388046 427905
rect 387872 427660 387904 427726
rect 388014 427660 388046 427726
rect 387872 427628 388046 427660
rect 392779 427745 392976 427912
rect 392779 427679 392828 427745
rect 392938 427679 392976 427745
rect 392779 427641 392976 427679
rect 387881 427354 388055 427383
rect 387881 427288 387914 427354
rect 388024 427288 388055 427354
rect 387881 426943 388055 427288
rect 392805 427373 392979 427402
rect 392805 427307 392838 427373
rect 392948 427307 392979 427373
rect 387423 421101 388423 426943
rect 392805 426938 392979 427307
rect 392311 426638 393311 426938
rect 392311 425640 392312 426638
rect 393310 425640 393311 426638
rect 392311 425639 393311 425640
rect 387416 421100 388423 421101
rect 387416 420100 387417 421100
rect 388417 420100 388418 421100
rect 387416 420099 388418 420100
rect 388621 415854 388623 415855
rect 374480 415850 374482 415851
rect 374481 415298 374482 415850
rect 374480 415297 374482 415298
rect 375344 415654 375346 415655
rect 375344 415102 375345 415654
rect 388621 415302 388622 415854
rect 393659 415390 393660 415391
rect 394212 415390 394213 415391
rect 393659 415389 394213 415390
rect 388621 415301 388623 415302
rect 375344 415101 375346 415102
rect 367488 391198 367490 391199
rect 367488 390646 367489 391198
rect 400973 391194 400975 391195
rect 367488 390645 367490 390646
rect 385805 391174 385807 391175
rect 385806 390622 385807 391174
rect 400974 390642 400975 391194
rect 400973 390641 400975 390642
rect 385805 390621 385807 390622
rect 400961 376106 400963 376107
rect 367488 376056 367490 376057
rect 367488 375504 367489 376056
rect 367488 375503 367490 375504
rect 388563 375924 388565 375925
rect 388563 375372 388564 375924
rect 400962 375554 400963 376106
rect 400961 375553 400963 375554
rect 388563 375371 388565 375372
rect 365528 316852 365529 317850
rect 366527 316852 366528 317850
rect 365528 316851 366528 316852
rect 390694 306935 391255 306936
rect 390694 306934 390695 306935
rect 391254 306934 391255 306935
rect 370682 306807 371243 306808
rect 370682 306806 370683 306807
rect 371242 306806 371243 306807
rect 400258 306893 400819 306894
rect 400258 306892 400259 306893
rect 400818 306892 400819 306893
rect 357939 306242 357940 306243
rect 358492 306242 358493 306243
rect 357939 306241 358493 306242
rect 355957 302183 356136 302545
rect 355957 302117 355993 302183
rect 356103 302117 356136 302183
rect 355957 302102 356136 302117
rect 355971 301811 356145 301843
rect 355971 301745 356003 301811
rect 356113 301797 356145 301811
rect 356113 301745 356146 301797
rect 355971 301598 356146 301745
rect 355561 296499 356561 301598
rect 355561 295501 355562 296499
rect 356560 295501 356561 296499
rect 355561 295500 356561 295501
rect 354577 286818 354579 286819
rect 354578 286266 354579 286818
rect 354577 286265 354579 286266
rect 370692 286612 370694 286613
rect 370692 286053 370693 286612
rect 400174 286359 400175 286360
rect 400734 286359 400735 286360
rect 400174 286358 400735 286359
rect 390694 286147 390695 286148
rect 391254 286147 391255 286148
rect 390694 286146 391255 286147
rect 370692 286052 370694 286053
rect 403045 247405 404045 506068
rect 405045 249391 406045 508779
rect 407045 251391 408045 511313
rect 409045 253391 410045 513846
rect 411045 255391 412045 516312
rect 413045 257391 414045 518914
rect 415045 259391 416045 521278
rect 417045 261391 418045 523744
rect 419045 263391 420045 526413
rect 421045 265391 422045 528704
rect 423045 267391 424045 531548
rect 425045 269391 426045 533985
rect 437075 530351 442175 554088
rect 449668 540461 454786 577998
rect 464241 539452 464243 539453
rect 464241 538840 464242 539452
rect 464241 538839 464243 538840
rect 442149 529681 442175 530351
rect 437075 513406 442175 529681
rect 449668 531568 454786 538198
rect 449668 530898 449712 531568
rect 437075 512736 437103 513406
rect 437075 486137 442175 512736
rect 449668 512175 454786 530898
rect 449668 511505 449671 512175
rect 454772 511505 454786 512175
rect 434799 485224 435413 485225
rect 434799 485223 434800 485224
rect 435412 485223 435413 485224
rect 428635 485216 429189 485217
rect 428635 485215 428636 485216
rect 429188 485215 429189 485216
rect 428289 472572 428290 472573
rect 428842 472572 428843 472573
rect 428289 472571 428843 472572
rect 437075 463376 442175 483874
rect 449668 474001 454786 511505
rect 458513 484710 458514 484711
rect 459126 484710 459127 484711
rect 458513 484709 459127 484710
rect 464284 484560 464285 484561
rect 464897 484560 464898 484561
rect 464284 484559 464898 484560
rect 475003 484530 475004 484531
rect 475616 484530 475617 484531
rect 475003 484529 475617 484530
rect 445477 472450 445478 472451
rect 446090 472450 446091 472451
rect 445477 472449 446091 472450
rect 462129 473054 462743 473055
rect 462129 473053 462130 473054
rect 462742 473053 462743 473054
rect 449668 467421 454786 471738
rect 449668 465158 449674 467421
rect 437075 431177 442175 461113
rect 437075 392083 442175 428914
rect 449668 416727 454786 465158
rect 428495 390760 428496 390761
rect 429048 390760 429049 390761
rect 428495 390759 429049 390760
rect 446399 391054 446401 391055
rect 446399 390502 446400 391054
rect 446399 390501 446401 390502
rect 429153 376012 429155 376013
rect 429153 375460 429154 376012
rect 429153 375459 429155 375460
rect 437075 307769 442175 389820
rect 449668 377007 454786 414464
rect 470031 391060 470033 391061
rect 470031 390508 470032 391060
rect 470031 390507 470033 390508
rect 446947 376070 446949 376071
rect 446948 375518 446949 376070
rect 446947 375517 446949 375518
rect 467085 376054 467087 376055
rect 467086 375502 467087 376054
rect 467085 375501 467087 375502
rect 430708 306657 431269 306658
rect 430708 306656 430709 306657
rect 431268 306656 431269 306657
rect 445434 306855 445995 306856
rect 445434 306854 445435 306855
rect 445994 306854 445995 306855
rect 430708 286265 430709 286266
rect 431268 286265 431269 286266
rect 430708 286264 431269 286265
rect 425034 269390 426045 269391
rect 425034 268390 425035 269390
rect 426035 268390 426045 269390
rect 425034 268389 426045 268390
rect 425045 268228 426045 268389
rect 423041 267390 424045 267391
rect 423041 266390 423042 267390
rect 424042 266390 424045 267390
rect 423041 266389 424045 266390
rect 423045 266279 424045 266389
rect 421045 265390 422076 265391
rect 421045 264390 421075 265390
rect 422075 264390 422076 265390
rect 421045 264389 422076 264390
rect 421045 264274 422045 264389
rect 419045 263390 420083 263391
rect 419045 262390 419082 263390
rect 420082 262390 420083 263390
rect 419045 262389 420083 262390
rect 419045 262214 420045 262389
rect 417045 261390 418050 261391
rect 417045 260390 417049 261390
rect 418049 260390 418050 261390
rect 417045 260389 418050 260390
rect 417045 260265 418045 260389
rect 415045 259390 416075 259391
rect 415045 258390 415074 259390
rect 416074 258390 416075 259390
rect 415045 258389 416075 258390
rect 415045 258205 416045 258389
rect 413045 257390 414047 257391
rect 413045 256390 413046 257390
rect 414046 256390 414047 257390
rect 413045 256389 414047 256390
rect 413045 256256 414045 256389
rect 411017 255390 412045 255391
rect 411017 254390 411018 255390
rect 412018 254390 412045 255390
rect 411017 254389 412045 254390
rect 411045 254252 412045 254389
rect 409045 253390 410098 253391
rect 409045 252390 409097 253390
rect 410097 252390 410098 253390
rect 409045 252389 410098 252390
rect 409045 252247 410045 252389
rect 407014 251390 408045 251391
rect 407014 250390 407015 251390
rect 408015 250390 408045 251390
rect 407014 250389 408045 250390
rect 407045 250197 408045 250389
rect 405045 249390 406095 249391
rect 405045 248390 405094 249390
rect 406094 248390 406095 249390
rect 405045 248389 406095 248390
rect 405045 248355 406045 248389
rect 403025 247389 404061 247405
rect 403025 246391 403046 247389
rect 404044 246391 404061 247389
rect 403025 246376 404061 246391
rect 356446 213126 361534 213150
rect 356446 208086 356470 213126
rect 361510 208086 361534 213126
rect 437075 213126 442175 305506
rect 449668 287781 454786 374744
rect 470722 306785 470724 306786
rect 470722 306226 470723 306785
rect 470722 306225 470724 306226
rect 445446 286477 445447 286478
rect 446006 286477 446007 286478
rect 445446 286476 446007 286477
rect 470722 286758 470724 286759
rect 470722 286199 470723 286758
rect 470722 286198 470724 286199
rect 437075 208170 437112 213126
rect 442152 208170 442175 213126
rect 356446 137374 361534 208086
rect 449668 196266 454786 285518
rect 454435 191354 454786 196266
rect 449668 186346 454786 191354
rect 454514 181276 454786 186346
rect 449668 177836 454786 181276
rect 449668 172766 449876 177836
rect 449668 167838 454786 172766
rect 449668 162995 449738 167838
rect 356446 136822 358800 137374
rect 359342 136822 361534 137374
rect 356446 95644 361534 136822
rect 356446 95092 359148 95644
rect 359690 95092 361534 95644
rect 356446 54530 361534 95092
rect 356446 53978 358810 54530
rect 359352 53978 361534 54530
rect 477776 54057 478776 589076
rect 482433 54057 483433 596089
rect 484632 539562 484634 539563
rect 484632 538950 484633 539562
rect 484632 538949 484634 538950
rect 485224 485200 485226 485201
rect 485225 484588 485226 485200
rect 485224 484587 485226 484588
rect 485291 473098 485905 473099
rect 485291 473097 485292 473098
rect 485904 473097 485905 473098
rect 486045 376010 486047 376011
rect 486046 375458 486047 376010
rect 486045 375457 486047 375458
rect 487607 54057 488607 602557
rect 544391 587292 545391 587293
rect 544391 586294 544392 587292
rect 545390 586294 545391 587292
rect 538405 579328 538407 579329
rect 538406 578716 538407 579328
rect 538405 578715 538407 578716
rect 544391 573515 545391 586294
rect 544690 573219 544888 573515
rect 544690 573153 544736 573219
rect 544846 573153 544888 573219
rect 544690 573113 544888 573153
rect 544684 572847 544874 572889
rect 544684 572781 544726 572847
rect 544836 572781 544874 572847
rect 544684 572442 544874 572781
rect 530513 568443 531515 568444
rect 522151 568442 523151 568443
rect 513275 568273 514277 568274
rect 505084 568272 506084 568273
rect 505084 567274 505085 568272
rect 506083 567274 506084 568272
rect 505084 560842 506084 567274
rect 513275 567273 513276 568273
rect 514276 567273 514277 568273
rect 513275 567272 514277 567273
rect 522151 567444 522152 568442
rect 523150 567444 523151 568442
rect 513276 563131 514276 567272
rect 513724 562663 513914 563131
rect 513724 562597 513762 562663
rect 513872 562597 513914 562663
rect 513724 562555 513914 562597
rect 513710 562291 513906 562328
rect 513710 562225 513752 562291
rect 513862 562225 513906 562291
rect 513710 561895 513906 562225
rect 505408 560570 505598 560842
rect 505408 560504 505449 560570
rect 505559 560504 505598 560570
rect 505408 560469 505598 560504
rect 505397 560198 505587 560240
rect 505397 560132 505439 560198
rect 505549 560132 505587 560198
rect 505397 559638 505587 560132
rect 505084 540151 506084 559638
rect 509407 556160 509939 556161
rect 509407 554242 509408 556160
rect 509938 554242 509939 556160
rect 509407 554241 509939 554242
rect 513276 542492 514276 561895
rect 522151 550736 523151 567444
rect 530513 567443 530514 568443
rect 531514 567443 531515 568443
rect 530513 567442 531515 567443
rect 526607 556182 527209 556183
rect 526607 554236 526608 556182
rect 527208 554236 527209 556182
rect 526607 554235 527209 554236
rect 530514 553436 531514 567442
rect 530994 553109 531184 553436
rect 530994 553043 531032 553109
rect 531142 553043 531184 553109
rect 544391 553095 545391 572442
rect 547181 556178 547759 556179
rect 547181 554212 547182 556178
rect 547758 554212 547759 556178
rect 547181 554211 547759 554212
rect 559614 556132 560614 629629
rect 559614 554240 559640 556132
rect 560562 554240 560614 556132
rect 530994 553001 531184 553043
rect 544705 552970 544895 553095
rect 544705 552904 544746 552970
rect 544856 552904 544895 552970
rect 544705 552869 544895 552904
rect 530982 552737 531180 552777
rect 530982 552671 531022 552737
rect 531132 552671 531180 552737
rect 530982 552449 531180 552671
rect 544694 552598 544884 552640
rect 544694 552532 544736 552598
rect 544846 552532 544884 552598
rect 522463 550492 522664 550736
rect 522463 550426 522511 550492
rect 522621 550426 522664 550492
rect 522463 550386 522664 550426
rect 522459 550120 522649 550162
rect 522459 550054 522501 550120
rect 522611 550054 522649 550120
rect 522459 549532 522649 550054
rect 513704 542221 513894 542492
rect 513704 542155 513742 542221
rect 513852 542155 513894 542221
rect 513704 542113 513894 542155
rect 513693 541849 513883 541884
rect 513693 541783 513732 541849
rect 513842 541783 513883 541849
rect 513693 541542 513883 541783
rect 505518 539982 505708 540151
rect 505518 539916 505559 539982
rect 505669 539916 505708 539982
rect 505518 539881 505708 539916
rect 505507 539610 505697 539652
rect 505507 539544 505549 539610
rect 505659 539544 505697 539610
rect 505507 539168 505697 539544
rect 500437 539034 500438 539035
rect 501050 539034 501051 539035
rect 500437 539033 501051 539034
rect 505084 519693 506084 539168
rect 513276 522651 514276 541542
rect 517873 540212 518575 540213
rect 517873 538396 517874 540212
rect 518574 538396 518575 540212
rect 517873 538395 518575 538396
rect 522151 529967 523151 549532
rect 530514 532158 531514 552449
rect 544694 552193 544884 552532
rect 537833 540294 538411 540295
rect 537833 538328 537834 540294
rect 538410 538328 538411 540294
rect 537833 538327 538411 538328
rect 544391 532856 545391 552193
rect 544710 532744 544900 532856
rect 544710 532678 544751 532744
rect 544861 532678 544900 532744
rect 544710 532643 544900 532678
rect 544699 532372 544889 532414
rect 544699 532306 544741 532372
rect 544851 532306 544889 532372
rect 530949 531864 531139 532158
rect 544699 532011 544889 532306
rect 530949 531798 530987 531864
rect 531097 531798 531139 531864
rect 530949 531756 531139 531798
rect 530938 531492 531128 531527
rect 530938 531426 530977 531492
rect 531087 531426 531128 531492
rect 530938 531309 531128 531426
rect 522519 529715 522709 529967
rect 522519 529649 522560 529715
rect 522670 529649 522709 529715
rect 522519 529614 522709 529649
rect 522508 529343 522698 529385
rect 522508 529277 522550 529343
rect 522660 529277 522698 529343
rect 522508 528963 522698 529277
rect 513701 522250 513891 522651
rect 513701 522184 513739 522250
rect 513849 522184 513891 522250
rect 513701 522142 513891 522184
rect 513690 521878 513880 521913
rect 513690 521812 513729 521878
rect 513839 521812 513880 521878
rect 513690 521600 513880 521812
rect 513276 519802 514276 521600
rect 522151 519804 523151 528963
rect 505083 519692 506085 519693
rect 505083 518692 505084 519692
rect 506084 518692 506085 519692
rect 513276 518804 513277 519802
rect 514275 518804 514276 519802
rect 513276 518803 514276 518804
rect 522150 519803 523152 519804
rect 522150 518803 522151 519803
rect 523151 518803 523152 519803
rect 530514 519802 531514 531309
rect 530514 518804 530515 519802
rect 531513 518804 531514 519802
rect 544391 519793 545391 532011
rect 530514 518803 531514 518804
rect 544390 519792 545392 519793
rect 522150 518802 523152 518803
rect 544390 518792 544391 519792
rect 545391 518792 545392 519792
rect 544390 518791 545392 518792
rect 505083 518691 506085 518692
rect 501673 510564 502675 510565
rect 501673 509564 501674 510564
rect 502674 509564 502675 510564
rect 501673 509563 502675 509564
rect 508548 510563 509548 510564
rect 508548 509565 508549 510563
rect 509547 509565 509548 510563
rect 501674 500723 502674 509563
rect 508548 506656 509548 509565
rect 514541 510484 515543 510485
rect 514541 509484 514542 510484
rect 515542 509484 515543 510484
rect 514541 509483 515543 509484
rect 521016 510483 522016 510484
rect 521016 509485 521017 510483
rect 522015 509485 522016 510483
rect 514542 508375 515542 509483
rect 514997 507933 515190 508375
rect 514997 507867 515038 507933
rect 515148 507867 515190 507933
rect 514997 507839 515190 507867
rect 514988 507561 515178 507600
rect 514988 507495 515028 507561
rect 515138 507495 515178 507561
rect 514988 507222 515178 507495
rect 508904 506525 509082 506656
rect 508904 506459 508942 506525
rect 509052 506459 509082 506525
rect 508904 506417 509082 506459
rect 508902 506153 509080 506190
rect 508902 506087 508932 506153
rect 509042 506087 509080 506153
rect 508902 505754 509080 506087
rect 502143 500326 502324 500723
rect 502143 500260 502178 500326
rect 502288 500260 502324 500326
rect 502143 500230 502324 500260
rect 502126 499954 502307 499986
rect 502126 499888 502168 499954
rect 502278 499888 502307 499954
rect 502126 499618 502307 499888
rect 499099 485116 499101 485117
rect 499100 484504 499101 485116
rect 499099 484503 499101 484504
rect 501674 480113 502674 499618
rect 508548 486751 509548 505754
rect 514542 488076 515542 507222
rect 521016 498750 522016 509485
rect 527089 510404 528091 510405
rect 527089 509404 527090 510404
rect 528090 509404 528091 510404
rect 527089 509403 528091 509404
rect 533844 510403 534844 510404
rect 533844 509405 533845 510403
rect 534843 509405 534844 510403
rect 521355 498399 521536 498750
rect 521355 498333 521392 498399
rect 521502 498333 521536 498399
rect 521355 498294 521536 498333
rect 521348 498027 521529 498071
rect 521348 497961 521382 498027
rect 521492 497961 521529 498027
rect 521348 497493 521529 497961
rect 514965 487732 515151 488076
rect 514965 487666 515001 487732
rect 515111 487666 515151 487732
rect 514965 487633 515151 487666
rect 514955 487360 515144 487395
rect 514955 487294 514991 487360
rect 515101 487294 515144 487360
rect 514955 486997 515144 487294
rect 508919 486474 509091 486751
rect 508919 486408 508954 486474
rect 509064 486408 509091 486474
rect 508919 486363 509091 486408
rect 508911 486102 509083 486135
rect 508911 486036 508944 486102
rect 509054 486036 509083 486102
rect 508911 485689 509083 486036
rect 504621 484568 504622 484569
rect 505234 484568 505235 484569
rect 504621 484567 505235 484568
rect 508548 480115 509548 485689
rect 512440 485220 512442 485221
rect 512441 484608 512442 485220
rect 512440 484607 512442 484608
rect 501674 479115 501675 480113
rect 502673 479115 502674 480113
rect 501674 479114 502674 479115
rect 508547 480114 509549 480115
rect 508547 479114 508548 480114
rect 509548 479114 509549 480114
rect 514542 480113 515542 486997
rect 518837 485220 518839 485221
rect 518838 484580 518839 485220
rect 518837 484579 518839 484580
rect 521016 480115 522016 497493
rect 527090 496411 528090 509403
rect 533844 509082 534844 509405
rect 534303 508952 534478 509082
rect 534303 508886 534334 508952
rect 534444 508886 534478 508952
rect 534303 508848 534478 508886
rect 534307 508580 534482 508609
rect 534307 508514 534344 508580
rect 534454 508514 534482 508580
rect 534307 508193 534482 508514
rect 527429 496001 527610 496411
rect 527429 495935 527466 496001
rect 527576 495935 527610 496001
rect 527429 495891 527610 495935
rect 527422 495629 527603 495668
rect 527422 495563 527456 495629
rect 527566 495563 527603 495629
rect 527422 495154 527603 495563
rect 524294 485164 524296 485165
rect 524294 484552 524295 485164
rect 524294 484551 524296 484552
rect 514542 479115 514543 480113
rect 515541 479115 515542 480113
rect 514542 479114 515542 479115
rect 521015 480114 522017 480115
rect 521015 479114 521016 480114
rect 522016 479114 522017 480114
rect 527090 480113 528090 495154
rect 533844 488880 534844 508193
rect 559614 500162 560614 554240
rect 559614 500050 559955 500162
rect 560067 500050 560614 500162
rect 549985 498323 550985 498324
rect 549985 497325 549986 498323
rect 550984 497325 550985 498323
rect 549985 492479 550985 497325
rect 550417 492056 550622 492479
rect 550417 491990 550466 492056
rect 550576 491990 550622 492056
rect 550417 491953 550622 491990
rect 550408 491684 550613 491715
rect 550408 491618 550456 491684
rect 550566 491618 550613 491684
rect 550408 491319 550613 491618
rect 534289 488552 534495 488880
rect 534289 488486 534344 488552
rect 534454 488486 534495 488552
rect 534289 488461 534495 488486
rect 534317 488180 534492 488209
rect 534317 488114 534354 488180
rect 534464 488114 534492 488180
rect 534317 487739 534492 488114
rect 531885 485216 532527 485217
rect 531885 485215 531886 485216
rect 532526 485215 532527 485216
rect 530383 484576 530384 484577
rect 530996 484576 530997 484577
rect 530383 484575 530997 484576
rect 533844 480117 534844 487739
rect 546408 485132 546410 485133
rect 546409 484492 546410 485132
rect 546408 484491 546410 484492
rect 527090 479115 527091 480113
rect 528089 479115 528090 480113
rect 533843 480116 534845 480117
rect 533843 479116 533844 480116
rect 534844 479116 534845 480116
rect 549985 480110 550985 491319
rect 559614 485896 560614 500050
rect 559614 484004 559636 485896
rect 560558 484004 560614 485896
rect 533843 479115 534845 479116
rect 549984 480109 550986 480110
rect 527090 479114 528090 479115
rect 508547 479113 509549 479114
rect 521015 479113 522017 479114
rect 549984 479109 549985 480109
rect 550985 479109 550986 480109
rect 549984 479108 550986 479109
rect 549889 476016 550891 476017
rect 508579 476011 509581 476012
rect 521047 476011 522049 476012
rect 501706 476010 502706 476011
rect 501706 475012 501707 476010
rect 502705 475012 502706 476010
rect 497346 473189 497986 473190
rect 497346 473188 497347 473189
rect 497985 473188 497986 473189
rect 501706 455507 502706 475012
rect 508579 475011 508580 476011
rect 509580 475011 509581 476011
rect 508579 475010 509581 475011
rect 514574 476010 515574 476011
rect 514574 475012 514575 476010
rect 515573 475012 515574 476010
rect 507291 473006 507293 473007
rect 503854 472993 504494 472994
rect 503854 472992 503855 472993
rect 504493 472992 504494 472993
rect 507292 472394 507293 473006
rect 507291 472393 507293 472394
rect 508580 469436 509580 475010
rect 508943 469089 509115 469436
rect 508943 469023 508976 469089
rect 509086 469023 509115 469089
rect 508943 468990 509115 469023
rect 508951 468717 509123 468762
rect 508951 468651 508986 468717
rect 509096 468651 509123 468717
rect 508951 468374 509123 468651
rect 502158 455237 502339 455507
rect 502158 455171 502200 455237
rect 502310 455171 502339 455237
rect 502158 455139 502339 455171
rect 502175 454865 502356 454895
rect 502175 454799 502210 454865
rect 502320 454799 502356 454865
rect 502175 454402 502356 454799
rect 501706 445562 502706 454402
rect 508580 449371 509580 468374
rect 514574 468128 515574 475012
rect 521047 475011 521048 476011
rect 522048 475011 522049 476011
rect 521047 475010 522049 475011
rect 527122 476010 528122 476011
rect 527122 475012 527123 476010
rect 528121 475012 528122 476010
rect 518831 473092 518833 473093
rect 518832 472480 518833 473092
rect 518831 472479 518833 472480
rect 514987 467831 515176 468128
rect 514987 467765 515023 467831
rect 515133 467765 515176 467831
rect 514987 467730 515176 467765
rect 514997 467459 515183 467492
rect 514997 467393 515033 467459
rect 515143 467393 515183 467459
rect 514997 467049 515183 467393
rect 508934 449038 509112 449371
rect 508934 448972 508964 449038
rect 509074 448972 509112 449038
rect 508934 448935 509112 448972
rect 508936 448666 509114 448708
rect 508936 448600 508974 448666
rect 509084 448600 509114 448666
rect 508936 448469 509114 448600
rect 501705 445561 502707 445562
rect 501705 444561 501706 445561
rect 502706 444561 502707 445561
rect 508580 445560 509580 448469
rect 514574 447903 515574 467049
rect 521048 457632 522048 475010
rect 522943 473097 525128 473098
rect 522943 472495 522944 473097
rect 525127 472495 525128 473097
rect 522943 472494 525128 472495
rect 527122 459880 528122 475012
rect 533875 476009 534877 476010
rect 533875 475009 533876 476009
rect 534876 475009 534877 476009
rect 549889 475016 549890 476016
rect 550890 475016 550891 476016
rect 549889 475015 550891 475016
rect 533875 475008 534877 475009
rect 533876 467386 534876 475008
rect 548777 473212 548779 473213
rect 536947 473168 536949 473169
rect 536947 472556 536948 473168
rect 536947 472555 536949 472556
rect 537961 473146 537963 473147
rect 537961 472506 537962 473146
rect 548778 472572 548779 473212
rect 548777 472571 548779 472572
rect 537961 472505 537963 472506
rect 534349 467011 534524 467386
rect 534349 466945 534386 467011
rect 534496 466945 534524 467011
rect 534349 466916 534524 466945
rect 534321 466639 534527 466664
rect 534321 466573 534376 466639
rect 534486 466573 534527 466639
rect 534321 466245 534527 466573
rect 527497 459602 527672 459880
rect 527497 459536 527531 459602
rect 527641 459536 527672 459602
rect 527497 459498 527672 459536
rect 527493 459230 527668 459259
rect 527493 459164 527521 459230
rect 527631 459164 527668 459230
rect 527493 458758 527668 459164
rect 521380 457164 521561 457632
rect 521380 457098 521414 457164
rect 521524 457098 521561 457164
rect 521380 457054 521561 457098
rect 521387 456792 521568 456831
rect 521387 456726 521424 456792
rect 521534 456726 521568 456792
rect 521387 456375 521568 456726
rect 515020 447630 515210 447903
rect 515020 447564 515060 447630
rect 515170 447564 515210 447630
rect 515020 447525 515210 447564
rect 515029 447258 515222 447286
rect 515029 447192 515070 447258
rect 515180 447192 515222 447258
rect 515029 446750 515222 447192
rect 514574 445642 515574 446750
rect 508580 444562 508581 445560
rect 509579 444562 509580 445560
rect 514573 445641 515575 445642
rect 514573 444641 514574 445641
rect 515574 444641 515575 445641
rect 521048 445640 522048 456375
rect 527122 445722 528122 458758
rect 533876 446932 534876 466245
rect 549890 460018 550890 475015
rect 553167 473136 553169 473137
rect 553167 472496 553168 473136
rect 553167 472495 553169 472496
rect 549890 460016 550187 460018
rect 550329 460016 550890 460018
rect 550329 459731 550535 460016
rect 550329 459665 550370 459731
rect 550480 459665 550535 459731
rect 550329 459640 550535 459665
rect 550332 459359 550507 459388
rect 550332 459293 550360 459359
rect 550470 459293 550507 459359
rect 550332 458808 550507 459293
rect 549890 453859 550890 458808
rect 549890 452861 549891 453859
rect 550889 452861 550890 453859
rect 549890 452860 550890 452861
rect 559614 455740 560614 484004
rect 565199 589584 566199 604185
rect 565199 589472 565585 589584
rect 565697 589472 566199 589584
rect 565199 540236 566199 589472
rect 565199 538344 565238 540236
rect 566160 538344 566199 540236
rect 565199 473748 566199 538344
rect 567853 485176 567855 485177
rect 567853 484536 567854 485176
rect 567853 484535 567855 484536
rect 562797 472434 562798 472435
rect 563438 472434 563439 472435
rect 562797 472433 563439 472434
rect 559614 455628 560008 455740
rect 560120 455628 560614 455740
rect 534339 446611 534514 446932
rect 534339 446545 534376 446611
rect 534486 446545 534514 446611
rect 534339 446516 534514 446545
rect 534335 446239 534510 446277
rect 534335 446173 534366 446239
rect 534476 446173 534510 446239
rect 534335 446043 534510 446173
rect 521048 444642 521049 445640
rect 522047 444642 522048 445640
rect 527121 445721 528123 445722
rect 527121 444721 527122 445721
rect 528122 444721 528123 445721
rect 533876 445720 534876 446043
rect 533876 444722 533877 445720
rect 534875 444722 534876 445720
rect 533876 444721 534876 444722
rect 527121 444720 528123 444721
rect 521048 444641 522048 444642
rect 514573 444640 515575 444641
rect 508580 444561 509580 444562
rect 501705 444560 502707 444561
rect 559614 431014 560614 455628
rect 546407 430408 546409 430409
rect 497204 429775 497205 429776
rect 497843 429775 497844 429776
rect 497204 429774 497844 429775
rect 528963 430334 528965 430335
rect 513061 429738 513062 429739
rect 513674 429738 513675 429739
rect 513061 429737 513675 429738
rect 522907 430306 522909 430307
rect 522908 429694 522909 430306
rect 522907 429693 522909 429694
rect 528963 429694 528964 430334
rect 546408 429768 546409 430408
rect 546407 429767 546409 429768
rect 528963 429693 528965 429694
rect 510277 429688 510278 429689
rect 510890 429688 510891 429689
rect 510277 429687 510891 429688
rect 559614 429122 559662 431014
rect 560584 429122 560614 431014
rect 565199 471856 565224 473748
rect 566146 471856 566199 473748
rect 562795 430324 563437 430325
rect 562795 430323 562796 430324
rect 563436 430323 563437 430324
rect 559614 411318 560614 429122
rect 559614 411206 560017 411318
rect 560129 411206 560614 411318
rect 549017 409465 550017 409466
rect 549017 408467 549018 409465
rect 550016 408467 550017 409465
rect 549017 407568 550017 408467
rect 549518 407196 549702 407568
rect 549518 407130 549553 407196
rect 549663 407130 549702 407196
rect 549518 407096 549702 407130
rect 549532 406824 549662 406831
rect 549532 406758 549543 406824
rect 549653 406758 549662 406824
rect 549532 406605 549662 406758
rect 546959 391246 546961 391247
rect 530389 391152 530391 391153
rect 490273 391110 490275 391111
rect 490273 390558 490274 391110
rect 490273 390557 490275 390558
rect 510727 391080 510729 391081
rect 510727 390528 510728 391080
rect 530389 390600 530390 391152
rect 546960 390674 546961 391246
rect 546959 390673 546961 390674
rect 530389 390599 530391 390600
rect 510727 390527 510729 390528
rect 549017 388403 550017 406605
rect 559614 391876 560614 411206
rect 559614 389984 559660 391876
rect 560582 389984 560614 391876
rect 549535 388152 549719 388403
rect 549535 388086 549570 388152
rect 549680 388086 549719 388152
rect 549535 388052 549719 388086
rect 549549 387780 549679 387787
rect 549549 387714 549560 387780
rect 549670 387714 549679 387780
rect 549549 387589 549679 387714
rect 549017 387302 550017 387589
rect 548986 387271 550037 387302
rect 548986 386271 549017 387271
rect 550017 386271 550037 387271
rect 548986 386232 550037 386271
rect 548895 381238 549897 381239
rect 548895 380238 548896 381238
rect 549896 380238 549897 381238
rect 548895 380237 549897 380238
rect 548896 379726 549896 380237
rect 549338 379494 549517 379726
rect 549338 379428 549368 379494
rect 549478 379428 549517 379494
rect 549338 379407 549517 379428
rect 549334 379122 549528 379156
rect 549334 379056 549378 379122
rect 549488 379056 549528 379122
rect 549334 378588 549528 379056
rect 526309 376174 526311 376175
rect 505737 375994 505739 375995
rect 505737 375442 505738 375994
rect 526309 375622 526310 376174
rect 526309 375621 526311 375622
rect 505737 375441 505739 375442
rect 548896 364616 549896 378588
rect 552365 376052 552367 376053
rect 552365 375480 552366 376052
rect 552365 375479 552367 375480
rect 559614 364896 560614 389984
rect 565199 416560 566199 471856
rect 565199 414668 565236 416560
rect 566158 414668 566199 416560
rect 565199 376796 566199 414668
rect 571231 391210 571233 391211
rect 571231 390638 571232 391210
rect 571231 390637 571233 390638
rect 562703 376116 563277 376117
rect 562703 376115 562704 376116
rect 563276 376115 563277 376116
rect 559614 364784 560038 364896
rect 560150 364784 560614 364896
rect 549298 364308 549480 364616
rect 549298 364242 549329 364308
rect 549439 364242 549480 364308
rect 549298 364208 549480 364242
rect 549310 363936 549498 363972
rect 549310 363870 549339 363936
rect 549449 363870 549498 363936
rect 549310 363442 549498 363870
rect 548896 363046 549896 363442
rect 548896 362048 548897 363046
rect 549895 362048 549896 363046
rect 548896 362047 549896 362048
rect 559614 307562 560614 364784
rect 490718 307009 490720 307010
rect 490718 306450 490719 307009
rect 490718 306449 490720 306450
rect 510704 306901 510706 306902
rect 510704 306342 510705 306901
rect 510704 306341 510706 306342
rect 531229 306747 531231 306748
rect 531230 306188 531231 306747
rect 531229 306187 531231 306188
rect 552718 306735 552720 306736
rect 552719 306168 552720 306735
rect 552718 306167 552720 306168
rect 559614 305670 559644 307562
rect 560566 305670 560614 307562
rect 549081 296500 550083 296501
rect 549081 295500 549082 296500
rect 550082 295500 550083 296500
rect 549081 295499 550083 295500
rect 549082 293761 550082 295499
rect 549514 293441 549688 293761
rect 549514 293375 549547 293441
rect 549657 293375 549688 293441
rect 549514 293351 549688 293375
rect 549527 293069 549701 293096
rect 549527 293003 549557 293069
rect 549667 293003 549701 293069
rect 549527 292839 549701 293003
rect 546871 286988 546873 286989
rect 490718 286888 490720 286889
rect 490718 286329 490719 286888
rect 490718 286328 490720 286329
rect 510704 286824 510706 286825
rect 510704 286265 510705 286824
rect 510704 286264 510706 286265
rect 530690 286812 530692 286813
rect 530690 286253 530691 286812
rect 546872 286421 546873 286988
rect 546871 286420 546873 286421
rect 530690 286252 530692 286253
rect 549082 274475 550082 292839
rect 559614 283514 560614 305670
rect 565199 374904 565224 376796
rect 566146 374904 566199 376796
rect 565199 319674 566199 374904
rect 565199 319562 565606 319674
rect 565718 319562 566199 319674
rect 565199 287548 566199 319562
rect 569352 306242 569353 306243
rect 569932 306242 569933 306243
rect 569352 306241 569933 306242
rect 565199 285656 565232 287548
rect 566154 285656 566199 287548
rect 568312 286318 568313 286319
rect 568892 286318 568893 286319
rect 568312 286317 568893 286318
rect 565199 275252 566199 285656
rect 565199 275140 565656 275252
rect 565768 275140 566199 275252
rect 549072 274463 550093 274475
rect 549072 273465 549083 274463
rect 550081 273465 550093 274463
rect 549072 273450 550093 273465
rect 549082 273312 550082 273450
rect 565199 196299 566199 275140
rect 566194 191348 566199 196299
rect 565199 186266 566199 191348
rect 575460 196290 575462 196291
rect 575461 191330 575462 196290
rect 575460 191329 575462 191330
rect 565199 181315 565206 186266
rect 356446 40402 361534 53978
rect 344312 8591 344424 12006
rect 344311 8590 344425 8591
rect 344311 8478 344312 8590
rect 344424 8478 344425 8590
rect 344311 8477 344425 8478
rect 345070 7855 345182 12006
rect 345069 7854 345183 7855
rect 345069 7742 345070 7854
rect 345182 7742 345183 7854
rect 345069 7741 345183 7742
rect 348884 7257 348996 12006
rect 348883 7256 348997 7257
rect 348883 7144 348884 7256
rect 348996 7144 348997 7256
rect 348883 7143 348997 7144
rect 349584 6634 349696 12006
rect 350238 7297 350350 12006
rect 350866 8201 350978 12006
rect 350865 8200 350979 8201
rect 350865 8088 350866 8200
rect 350978 8088 350979 8200
rect 350865 8087 350979 8088
rect 350237 7296 350351 7297
rect 350237 7184 350238 7296
rect 350350 7184 350351 7296
rect 350237 7183 350351 7184
rect 349578 6633 349702 6634
rect 349578 6521 349579 6633
rect 349701 6521 349702 6633
rect 349578 6520 349702 6521
rect 34106 2949 34107 3947
rect 35105 2949 35106 3947
rect 478104 4019 478216 54057
rect 478104 3909 478105 4019
rect 478215 3909 478216 4019
rect 478104 3908 478216 3909
rect 482769 4013 482881 54057
rect 482769 3903 482770 4013
rect 482880 3903 482881 4013
rect 488005 4023 488117 54057
rect 565199 17173 566199 181315
rect 565199 16175 565200 17173
rect 566198 16175 566199 17173
rect 565199 16174 566199 16175
rect 488005 3913 488006 4023
rect 488116 3913 488117 4023
rect 488005 3912 488117 3913
rect 482769 3902 482881 3903
rect 34106 2948 35106 2949
rect 25357 1656 25471 1657
rect 25357 1544 25358 1656
rect 25470 1544 25471 1656
rect 25357 1543 25471 1544
<< via4 >>
rect 8382 648776 13472 648777
rect 8382 643688 8383 648776
rect 8383 643688 13471 648776
rect 13471 643688 13472 648776
rect 8382 643687 13472 643688
rect 131219 643712 136259 648752
rect 8390 638742 13464 638743
rect 8390 633670 8391 638742
rect 8391 633670 13463 638742
rect 13463 633670 13464 638742
rect 8390 633669 13464 633670
rect 131043 633694 136067 638718
rect 118328 609005 123446 614123
rect 437023 629601 442234 648802
rect 570817 644694 575921 644695
rect 559620 639595 560618 644687
rect 570817 639592 570818 644694
rect 570818 639592 575920 644694
rect 575920 639592 575921 644694
rect 570817 639591 575921 639592
rect 559611 629629 560609 634721
rect 570872 634674 575910 634675
rect 570872 629638 570873 634674
rect 570873 629638 575909 634674
rect 575909 629638 575910 634674
rect 570872 629637 575910 629638
rect 449681 609029 454751 614099
rect 130984 581875 136121 584235
rect 378792 582061 379469 584076
rect 396584 582065 397261 584080
rect 118354 577835 123274 580341
rect 377445 578103 378296 580049
rect 437037 581960 442172 584137
rect 397858 578053 398535 580068
rect 449647 577998 454787 580116
rect 437056 554088 442208 556351
rect 118302 465128 123454 467391
rect 130883 461032 136035 463295
rect 130950 428852 136102 431115
rect 238860 430264 239401 430265
rect 238860 429713 238861 430264
rect 238861 429713 239401 430264
rect 238860 429712 239401 429713
rect 118304 414440 123456 416703
rect 13065 177860 18185 177861
rect 13065 172742 13066 177860
rect 13066 172742 18184 177860
rect 18184 172742 18185 177860
rect 24981 172855 25988 177806
rect 13065 172741 18185 172742
rect 13373 167862 18493 167863
rect 13373 162744 13374 167862
rect 13374 162744 18492 167862
rect 18492 162744 18493 167862
rect 13373 162743 18493 162744
rect 25000 162809 26007 167760
rect 249229 430384 249773 430385
rect 249229 429843 249230 430384
rect 249230 429843 249772 430384
rect 249772 429843 249773 430384
rect 332863 430376 333417 430377
rect 252974 430368 253528 430369
rect 252974 429827 252975 430368
rect 252975 429827 253527 430368
rect 253527 429827 253528 430368
rect 258344 430367 258884 430368
rect 258344 429817 258883 430367
rect 258883 429817 258884 430367
rect 293220 430360 293762 430361
rect 278456 430348 278998 430349
rect 258344 429816 258884 429817
rect 272934 429752 272935 430293
rect 272935 429752 273487 430293
rect 273487 429752 273488 430293
rect 278456 429796 278997 430348
rect 278997 429796 278998 430348
rect 293220 429808 293761 430360
rect 293761 429808 293762 430360
rect 293220 429807 293762 429808
rect 299168 430260 299710 430261
rect 278456 429795 278998 429796
rect 272934 429751 273488 429752
rect 299168 429708 299709 430260
rect 299709 429708 299710 430260
rect 322091 430220 322633 430221
rect 299168 429707 299710 429708
rect 313342 430196 313896 430197
rect 313342 429655 313343 430196
rect 313343 429655 313895 430196
rect 313895 429655 313896 430196
rect 319482 430162 320024 430163
rect 319482 429610 320023 430162
rect 320023 429610 320024 430162
rect 322091 429668 322632 430220
rect 322632 429668 322633 430220
rect 332863 429835 332864 430376
rect 332864 429835 333416 430376
rect 333416 429835 333417 430376
rect 335400 430258 335942 430259
rect 335400 429706 335941 430258
rect 335941 429706 335942 430258
rect 335400 429705 335942 429706
rect 322091 429667 322633 429668
rect 319482 429609 320024 429610
rect 319472 415952 320014 415953
rect 252978 415917 253518 415918
rect 242013 415906 242566 415907
rect 242013 415366 242014 415906
rect 242014 415366 242565 415906
rect 242565 415366 242566 415906
rect 252978 415367 253517 415917
rect 253517 415367 253518 415917
rect 258330 415881 258882 415882
rect 252978 415366 253518 415367
rect 255267 415180 255268 415721
rect 255268 415180 255820 415721
rect 255820 415180 255821 415721
rect 258330 415342 258331 415881
rect 258331 415342 258881 415881
rect 258881 415342 258882 415881
rect 313348 415876 313890 415877
rect 278444 415820 278998 415821
rect 272926 415814 273480 415815
rect 272926 415273 272927 415814
rect 272927 415273 273479 415814
rect 273479 415273 273480 415814
rect 278444 415279 278445 415820
rect 278445 415279 278997 415820
rect 278997 415279 278998 415820
rect 299130 415818 299684 415819
rect 293220 415794 293762 415795
rect 293220 415242 293761 415794
rect 293761 415242 293762 415794
rect 299130 415277 299131 415818
rect 299131 415277 299683 415818
rect 299683 415277 299684 415818
rect 313348 415324 313349 415876
rect 313349 415324 313890 415876
rect 319472 415400 320013 415952
rect 320013 415400 320014 415952
rect 319472 415399 320014 415400
rect 313348 415323 313890 415324
rect 293220 415241 293762 415242
rect 255267 415179 255821 415180
rect 328165 415906 328707 415907
rect 328165 415354 328706 415906
rect 328706 415354 328707 415906
rect 328165 415353 328707 415354
rect 339881 415868 340423 415869
rect 339881 415316 340422 415868
rect 340422 415316 340423 415868
rect 339881 415315 340423 415316
rect 322889 391352 323431 391353
rect 322889 390800 322890 391352
rect 322890 390800 323431 391352
rect 322889 390799 323431 390800
rect 333086 391372 333628 391373
rect 333086 390820 333087 391372
rect 333087 390820 333628 391372
rect 333086 390819 333628 390820
rect 334873 391314 335415 391315
rect 334873 390762 334874 391314
rect 334874 390762 335415 391314
rect 334873 390761 335415 390762
rect 333084 376214 333638 376215
rect 325771 376100 326313 376101
rect 325771 375548 326312 376100
rect 326312 375548 326313 376100
rect 333084 375673 333085 376214
rect 333085 375673 333637 376214
rect 333637 375673 333638 376214
rect 337327 375568 337328 376109
rect 337328 375568 337880 376109
rect 337880 375568 337881 376109
rect 337327 375567 337881 375568
rect 325771 375547 326313 375548
rect 131021 208062 136109 213150
rect 118328 172766 123398 177836
rect 118194 162768 123264 167838
rect 332587 172766 337657 177836
rect 90284 58752 91538 60006
rect 302585 59508 303127 59509
rect 240069 59386 240623 59387
rect 133043 59376 133597 59377
rect 111721 59366 112275 59367
rect 111721 58825 111722 59366
rect 111722 58825 112274 59366
rect 112274 58825 112275 59366
rect 133043 58835 133044 59376
rect 133044 58835 133596 59376
rect 133596 58835 133597 59376
rect 154601 59332 155155 59333
rect 154601 58791 154602 59332
rect 154602 58791 155154 59332
rect 155154 58791 155155 59332
rect 175807 59332 176361 59333
rect 175807 58791 175808 59332
rect 175808 58791 176360 59332
rect 176360 58791 176361 59332
rect 219083 59310 219637 59311
rect 197189 59288 197743 59289
rect 197189 58747 197190 59288
rect 197190 58747 197742 59288
rect 197742 58747 197743 59288
rect 219083 58769 219084 59310
rect 219084 58769 219636 59310
rect 219636 58769 219637 59310
rect 240069 58845 240070 59386
rect 240070 58845 240622 59386
rect 240622 58845 240623 59386
rect 260583 59384 261125 59385
rect 260583 58832 261124 59384
rect 261124 58832 261125 59384
rect 260583 58831 261125 58832
rect 281395 59140 281937 59141
rect 281395 58588 281936 59140
rect 281936 58588 281937 59140
rect 302585 58956 303126 59508
rect 303126 58956 303127 59508
rect 302585 58955 303127 58956
rect 324121 59508 324663 59509
rect 324121 58956 324122 59508
rect 324122 58956 324663 59508
rect 324121 58955 324663 58956
rect 281395 58587 281937 58588
rect 332563 56725 337681 61843
rect 39899 52866 40873 52867
rect 39899 51905 39900 52866
rect 39900 51905 40872 52866
rect 40872 51905 40873 52866
rect 39650 36270 42762 39258
rect 48003 37360 48004 37901
rect 48004 37360 48556 37901
rect 48556 37360 48557 37901
rect 69297 37466 69298 38007
rect 69298 37466 69850 38007
rect 69850 37466 69851 38007
rect 69297 37465 69851 37466
rect 48003 37359 48557 37360
rect 90663 37148 90664 37689
rect 90664 37148 91216 37689
rect 91216 37148 91217 37689
rect 111723 37200 111724 37741
rect 111724 37200 112276 37741
rect 112276 37200 112277 37741
rect 111723 37199 112277 37200
rect 133057 37672 133599 37673
rect 90663 37147 91217 37148
rect 133057 37120 133598 37672
rect 133598 37120 133599 37672
rect 154603 37288 154604 37829
rect 154604 37288 155156 37829
rect 155156 37288 155157 37829
rect 154603 37287 155157 37288
rect 175809 37288 175810 37829
rect 175810 37288 176362 37829
rect 176362 37288 176363 37829
rect 197191 37386 197192 37927
rect 197192 37386 197744 37927
rect 197744 37386 197745 37927
rect 302575 37924 303117 37925
rect 197191 37385 197745 37386
rect 219085 37336 219086 37877
rect 219086 37336 219638 37877
rect 219638 37336 219639 37877
rect 281385 37820 281927 37821
rect 219085 37335 219639 37336
rect 240071 37786 240613 37787
rect 175809 37287 176363 37288
rect 240071 37234 240072 37786
rect 240072 37234 240613 37786
rect 240071 37233 240613 37234
rect 260573 37724 261115 37725
rect 260573 37172 260574 37724
rect 260574 37172 261115 37724
rect 281385 37268 281386 37820
rect 281386 37268 281927 37820
rect 302575 37372 302576 37924
rect 302576 37372 303117 37924
rect 302575 37371 303117 37372
rect 324123 37872 324665 37873
rect 324123 37320 324124 37872
rect 324124 37320 324665 37872
rect 324123 37319 324665 37320
rect 281385 37267 281927 37268
rect 260573 37171 261115 37172
rect 133057 37119 133599 37120
rect 345550 414894 345978 416210
rect 348094 429382 348522 430698
rect 345675 376094 346229 376095
rect 345675 375553 345676 376094
rect 345676 375553 346228 376094
rect 346228 375553 346229 376094
rect 348024 305644 348476 307618
rect 345710 285614 346162 287588
rect 347982 208088 348448 213096
rect 345722 172818 346188 177826
rect 345698 162828 346164 167836
rect 360437 485152 360991 485153
rect 360437 484611 360438 485152
rect 360438 484611 360990 485152
rect 360990 484611 360991 485152
rect 352775 472986 353317 472987
rect 352775 472434 352776 472986
rect 352776 472434 353317 472986
rect 352775 472433 353317 472434
rect 354351 429722 354352 430263
rect 354352 429722 354904 430263
rect 354904 429722 354905 430263
rect 354351 429721 354905 429722
rect 359995 430444 360549 430445
rect 359995 429903 359996 430444
rect 359996 429903 360548 430444
rect 360548 429903 360549 430444
rect 362165 429896 362166 430437
rect 362166 429896 362718 430437
rect 362718 429896 362719 430437
rect 362165 429895 362719 429896
rect 353567 415228 353568 415769
rect 353568 415228 354120 415769
rect 354120 415228 354121 415769
rect 353567 415227 354121 415228
rect 353559 390944 354113 390945
rect 353559 390403 353560 390944
rect 353560 390403 354112 390944
rect 354112 390403 354113 390944
rect 357696 391162 358238 391163
rect 357696 390610 358237 391162
rect 358237 390610 358238 391162
rect 357696 390609 358238 390610
rect 352330 375608 353838 376280
rect 357690 376106 358232 376107
rect 357690 375554 358231 376106
rect 358231 375554 358232 376106
rect 357690 375553 358232 375554
rect 375483 484742 375484 485283
rect 375484 484742 376036 485283
rect 376036 484742 376037 485283
rect 375483 484741 376037 484742
rect 377512 465285 378229 467291
rect 386089 484666 386090 485207
rect 386090 484666 386642 485207
rect 386642 484666 386643 485207
rect 386089 484665 386643 484666
rect 390323 485216 390877 485217
rect 380563 473164 381105 473165
rect 380563 472612 381104 473164
rect 381104 472612 381105 473164
rect 380563 472611 381105 472612
rect 390323 484675 390324 485216
rect 390324 484675 390876 485216
rect 390876 484675 390877 485216
rect 389485 472536 389486 473077
rect 389486 472536 390038 473077
rect 390038 472536 390039 473077
rect 389485 472535 390039 472536
rect 394691 472610 394692 473151
rect 394692 472610 395244 473151
rect 395244 472610 395245 473151
rect 394691 472609 395245 472610
rect 378782 461283 379499 463289
rect 400217 485186 400771 485187
rect 400217 484645 400218 485186
rect 400218 484645 400770 485186
rect 400770 484645 400771 485186
rect 400585 472562 400586 473103
rect 400586 472562 401138 473103
rect 401138 472562 401139 473103
rect 400585 472561 401139 472562
rect 397854 465284 398571 467290
rect 396581 461271 397298 463277
rect 385927 430292 386469 430293
rect 375346 430200 375900 430201
rect 373956 430196 374498 430197
rect 373956 429644 374497 430196
rect 374497 429644 374498 430196
rect 375346 429659 375347 430200
rect 375347 429659 375899 430200
rect 375899 429659 375900 430200
rect 385927 429740 385928 430292
rect 385928 429740 386469 430292
rect 385927 429739 386469 429740
rect 373956 429643 374498 429644
rect 391199 430376 391741 430377
rect 391199 429824 391200 430376
rect 391200 429824 391741 430376
rect 391199 429823 391741 429824
rect 393659 415932 394213 415933
rect 388623 415854 389165 415855
rect 373938 415850 374480 415851
rect 373938 415298 373939 415850
rect 373939 415298 374480 415850
rect 373938 415297 374480 415298
rect 375346 415654 375888 415655
rect 375346 415102 375887 415654
rect 375887 415102 375888 415654
rect 388623 415302 389164 415854
rect 389164 415302 389165 415854
rect 393659 415391 393660 415932
rect 393660 415391 394212 415932
rect 394212 415391 394213 415932
rect 388623 415301 389165 415302
rect 375346 415101 375888 415102
rect 367490 391198 368032 391199
rect 367490 390646 368031 391198
rect 368031 390646 368032 391198
rect 400431 391194 400973 391195
rect 367490 390645 368032 390646
rect 385263 391174 385805 391175
rect 385263 390622 385264 391174
rect 385264 390622 385805 391174
rect 400431 390642 400432 391194
rect 400432 390642 400973 391194
rect 400431 390641 400973 390642
rect 385263 390621 385805 390622
rect 400419 376106 400961 376107
rect 367490 376056 368032 376057
rect 367490 375504 368031 376056
rect 368031 375504 368032 376056
rect 367490 375503 368032 375504
rect 388565 375924 389107 375925
rect 388565 375372 389106 375924
rect 389106 375372 389107 375924
rect 400419 375554 400420 376106
rect 400420 375554 400961 376106
rect 400419 375553 400961 375554
rect 388565 375371 389107 375372
rect 357939 306784 358493 306785
rect 357939 306243 357940 306784
rect 357940 306243 358492 306784
rect 358492 306243 358493 306784
rect 370682 306258 370683 306806
rect 370683 306258 371242 306806
rect 371242 306258 371243 306806
rect 390694 306386 390695 306934
rect 390695 306386 391254 306934
rect 391254 306386 391255 306934
rect 390694 306385 391255 306386
rect 400258 306344 400259 306892
rect 400259 306344 400818 306892
rect 400818 306344 400819 306892
rect 400258 306343 400819 306344
rect 370682 306257 371243 306258
rect 400174 286908 400735 286909
rect 354035 286818 354577 286819
rect 354035 286266 354036 286818
rect 354036 286266 354577 286818
rect 390694 286696 391255 286697
rect 354035 286265 354577 286266
rect 370694 286612 371243 286613
rect 370694 286053 371242 286612
rect 371242 286053 371243 286612
rect 390694 286148 390695 286696
rect 390695 286148 391254 286696
rect 391254 286148 391255 286696
rect 400174 286360 400175 286908
rect 400175 286360 400734 286908
rect 400734 286360 400735 286908
rect 370694 286052 371243 286053
rect 449636 538198 454788 540461
rect 464243 539452 464845 539453
rect 464243 538840 464844 539452
rect 464844 538840 464845 539452
rect 464243 538839 464845 538840
rect 437048 529681 442149 530351
rect 449712 530898 454813 531568
rect 437103 512736 442204 513406
rect 449671 511505 454772 512175
rect 428635 484674 428636 485215
rect 428636 484674 429188 485215
rect 429188 484674 429189 485215
rect 428635 484673 429189 484674
rect 434799 484622 434800 485223
rect 434800 484622 435412 485223
rect 435412 484622 435413 485223
rect 434799 484621 435413 484622
rect 437052 483874 442204 486137
rect 428289 473114 428843 473115
rect 428289 472573 428290 473114
rect 428290 472573 428842 473114
rect 428842 472573 428843 473114
rect 458513 485312 459127 485313
rect 458513 484711 458514 485312
rect 458514 484711 459126 485312
rect 459126 484711 459127 485312
rect 464284 485162 464898 485163
rect 464284 484561 464285 485162
rect 464285 484561 464897 485162
rect 464897 484561 464898 485162
rect 475003 485132 475617 485133
rect 475003 484531 475004 485132
rect 475004 484531 475616 485132
rect 475616 484531 475617 485132
rect 445477 473052 446091 473053
rect 445477 472451 445478 473052
rect 445478 472451 446090 473052
rect 446090 472451 446091 473052
rect 449642 471738 454794 474001
rect 462129 472452 462130 473053
rect 462130 472452 462742 473053
rect 462742 472452 462743 473053
rect 462129 472451 462743 472452
rect 449674 465158 454826 467421
rect 437058 461113 442210 463376
rect 437048 428914 442200 431177
rect 449634 414464 454786 416727
rect 428495 391302 429049 391303
rect 428495 390761 428496 391302
rect 428496 390761 429048 391302
rect 429048 390761 429049 391302
rect 437044 389820 442196 392083
rect 446401 391054 446943 391055
rect 446401 390502 446942 391054
rect 446942 390502 446943 391054
rect 446401 390501 446943 390502
rect 429155 376012 429697 376013
rect 429155 375460 429696 376012
rect 429696 375460 429697 376012
rect 429155 375459 429697 375460
rect 470033 391060 470575 391061
rect 470033 390508 470574 391060
rect 470574 390508 470575 391060
rect 470033 390507 470575 390508
rect 446405 376070 446947 376071
rect 446405 375518 446406 376070
rect 446406 375518 446947 376070
rect 446405 375517 446947 375518
rect 449644 374744 454796 377007
rect 466543 376054 467085 376055
rect 466543 375502 466544 376054
rect 466544 375502 467085 376054
rect 466543 375501 467085 375502
rect 430708 306108 430709 306656
rect 430709 306108 431268 306656
rect 431268 306108 431269 306656
rect 430708 306107 431269 306108
rect 437034 305506 442186 307769
rect 445434 306306 445435 306854
rect 445435 306306 445994 306854
rect 445994 306306 445995 306854
rect 445434 306305 445995 306306
rect 430708 286814 431269 286815
rect 430708 286266 430709 286814
rect 430709 286266 431268 286814
rect 431268 286266 431269 286814
rect 356470 208086 361510 213126
rect 470724 306785 471273 306786
rect 470724 306226 471272 306785
rect 471272 306226 471273 306785
rect 470724 306225 471273 306226
rect 445446 287026 446007 287027
rect 445446 286478 445447 287026
rect 445447 286478 446006 287026
rect 446006 286478 446007 287026
rect 449650 285518 454802 287781
rect 470724 286758 471273 286759
rect 470724 286199 471272 286758
rect 471272 286199 471273 286758
rect 470724 286198 471273 286199
rect 437112 208086 442152 213126
rect 449523 191354 454435 196266
rect 449444 181276 454514 186346
rect 449876 172766 454946 177836
rect 449738 162768 454808 167838
rect 484634 539562 485236 539563
rect 484634 538950 485235 539562
rect 485235 538950 485236 539562
rect 484634 538949 485236 538950
rect 484622 485200 485224 485201
rect 484622 484588 484623 485200
rect 484623 484588 485224 485200
rect 484622 484587 485224 484588
rect 485291 472496 485292 473097
rect 485292 472496 485904 473097
rect 485904 472496 485905 473097
rect 485291 472495 485905 472496
rect 485503 376010 486045 376011
rect 485503 375458 485504 376010
rect 485504 375458 486045 376010
rect 485503 375457 486045 375458
rect 537803 579328 538405 579329
rect 537803 578716 537804 579328
rect 537804 578716 538405 579328
rect 537803 578715 538405 578716
rect 509408 554242 509938 556160
rect 526608 554236 527208 556182
rect 547182 554212 547758 556178
rect 559640 554240 560562 556132
rect 500437 539636 501051 539637
rect 500437 539035 500438 539636
rect 500438 539035 501050 539636
rect 501050 539035 501051 539636
rect 517874 538396 518574 540212
rect 537834 538328 538410 540294
rect 498497 485116 499099 485117
rect 498497 484504 498498 485116
rect 498498 484504 499099 485116
rect 498497 484503 499099 484504
rect 504621 485170 505235 485171
rect 504621 484569 504622 485170
rect 504622 484569 505234 485170
rect 505234 484569 505235 485170
rect 511838 485220 512440 485221
rect 511838 484608 511839 485220
rect 511839 484608 512440 485220
rect 511838 484607 512440 484608
rect 518207 485220 518837 485221
rect 518207 484580 518208 485220
rect 518208 484580 518837 485220
rect 518207 484579 518837 484580
rect 524296 485164 524898 485165
rect 524296 484552 524897 485164
rect 524897 484552 524898 485164
rect 524296 484551 524898 484552
rect 530383 485178 530997 485179
rect 530383 484577 530384 485178
rect 530384 484577 530996 485178
rect 530996 484577 530997 485178
rect 531885 484586 531886 485215
rect 531886 484586 532526 485215
rect 532526 484586 532527 485215
rect 531885 484585 532527 484586
rect 545778 485132 546408 485133
rect 545778 484492 545779 485132
rect 545779 484492 546408 485132
rect 545778 484491 546408 484492
rect 559636 484004 560558 485896
rect 497346 472561 497347 473188
rect 497347 472561 497985 473188
rect 497985 472561 497986 473188
rect 497346 472560 497986 472561
rect 506689 473006 507291 473007
rect 503854 472365 503855 472992
rect 503855 472365 504493 472992
rect 504493 472365 504494 472992
rect 506689 472394 506690 473006
rect 506690 472394 507291 473006
rect 506689 472393 507291 472394
rect 503854 472364 504494 472365
rect 518229 473092 518831 473093
rect 518229 472480 518230 473092
rect 518230 472480 518831 473092
rect 518229 472479 518831 472480
rect 522944 472495 525127 473097
rect 548147 473212 548777 473213
rect 536949 473168 537551 473169
rect 536949 472556 537550 473168
rect 537550 472556 537551 473168
rect 536949 472555 537551 472556
rect 537963 473146 538593 473147
rect 537963 472506 538592 473146
rect 538592 472506 538593 473146
rect 548147 472572 548148 473212
rect 548148 472572 548777 473212
rect 548147 472571 548777 472572
rect 537963 472505 538593 472506
rect 553169 473136 553799 473137
rect 553169 472496 553798 473136
rect 553798 472496 553799 473136
rect 553169 472495 553799 472496
rect 565238 538344 566160 540236
rect 567855 485176 568485 485177
rect 567855 484536 568484 485176
rect 568484 484536 568485 485176
rect 567855 484535 568485 484536
rect 562797 473064 563439 473065
rect 562797 472435 562798 473064
rect 562798 472435 563438 473064
rect 563438 472435 563439 473064
rect 545777 430408 546407 430409
rect 497204 430403 497844 430404
rect 497204 429776 497205 430403
rect 497205 429776 497843 430403
rect 497843 429776 497844 430403
rect 513061 430340 513675 430341
rect 510277 430290 510891 430291
rect 510277 429689 510278 430290
rect 510278 429689 510890 430290
rect 510890 429689 510891 430290
rect 513061 429739 513062 430340
rect 513062 429739 513674 430340
rect 513674 429739 513675 430340
rect 528965 430334 529595 430335
rect 522305 430306 522907 430307
rect 522305 429694 522306 430306
rect 522306 429694 522907 430306
rect 522305 429693 522907 429694
rect 528965 429694 529594 430334
rect 529594 429694 529595 430334
rect 545777 429768 545778 430408
rect 545778 429768 546407 430408
rect 545777 429767 546407 429768
rect 528965 429693 529595 429694
rect 559662 429122 560584 431014
rect 565224 471856 566146 473748
rect 562795 429694 562796 430323
rect 562796 429694 563436 430323
rect 563436 429694 563437 430323
rect 562795 429693 563437 429694
rect 546397 391246 546959 391247
rect 530391 391152 530933 391153
rect 490275 391110 490817 391111
rect 490275 390558 490816 391110
rect 490816 390558 490817 391110
rect 490275 390557 490817 390558
rect 510729 391080 511271 391081
rect 510729 390528 511270 391080
rect 511270 390528 511271 391080
rect 530391 390600 530932 391152
rect 530932 390600 530933 391152
rect 546397 390674 546398 391246
rect 546398 390674 546959 391246
rect 546397 390673 546959 390674
rect 530391 390599 530933 390600
rect 510729 390527 511271 390528
rect 559660 389984 560582 391876
rect 526311 376174 526853 376175
rect 505739 375994 506281 375995
rect 505739 375442 506280 375994
rect 506280 375442 506281 375994
rect 526311 375622 526852 376174
rect 526852 375622 526853 376174
rect 526311 375621 526853 375622
rect 505739 375441 506281 375442
rect 552367 376052 552929 376053
rect 552367 375480 552928 376052
rect 552928 375480 552929 376052
rect 552367 375479 552929 375480
rect 565236 414668 566158 416560
rect 571233 391210 571795 391211
rect 571233 390638 571794 391210
rect 571794 390638 571795 391210
rect 571233 390637 571795 390638
rect 562703 375554 562704 376115
rect 562704 375554 563276 376115
rect 563276 375554 563277 376115
rect 562703 375553 563277 375554
rect 490720 307009 491269 307010
rect 490720 306450 491268 307009
rect 491268 306450 491269 307009
rect 490720 306449 491269 306450
rect 510706 306901 511255 306902
rect 510706 306342 511254 306901
rect 511254 306342 511255 306901
rect 510706 306341 511255 306342
rect 530680 306747 531229 306748
rect 530680 306188 530681 306747
rect 530681 306188 531229 306747
rect 530680 306187 531229 306188
rect 552161 306735 552718 306736
rect 552161 306168 552162 306735
rect 552162 306168 552718 306735
rect 552161 306167 552718 306168
rect 559644 305670 560566 307562
rect 546314 286988 546871 286989
rect 490720 286888 491269 286889
rect 490720 286329 491268 286888
rect 491268 286329 491269 286888
rect 490720 286328 491269 286329
rect 510706 286824 511255 286825
rect 510706 286265 511254 286824
rect 511254 286265 511255 286824
rect 510706 286264 511255 286265
rect 530692 286812 531241 286813
rect 530692 286253 531240 286812
rect 531240 286253 531241 286812
rect 546314 286421 546315 286988
rect 546315 286421 546871 286988
rect 546314 286420 546871 286421
rect 530692 286252 531241 286253
rect 565224 374904 566146 376796
rect 569352 306811 569933 306812
rect 569352 306243 569353 306811
rect 569353 306243 569932 306811
rect 569932 306243 569933 306811
rect 565232 285656 566154 287548
rect 568312 286887 568893 286888
rect 568312 286319 568313 286887
rect 568313 286319 568892 286887
rect 568892 286319 568893 286887
rect 565187 191348 566194 196299
rect 570500 196290 575460 196291
rect 570500 191330 570501 196290
rect 570501 191330 575460 196290
rect 570500 191329 575460 191330
rect 570413 186370 575533 186371
rect 565206 181315 566213 186266
rect 356446 35314 361534 40402
rect 570413 181252 570414 186370
rect 570414 181252 575532 186370
rect 575532 181252 575533 186370
rect 570413 181251 575533 181252
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 436999 648802 442258 648826
rect 8358 648777 13496 648801
rect 8358 643687 8382 648777
rect 13472 648776 13496 648777
rect 436999 648776 437023 648802
rect 13472 648752 437023 648776
rect 13472 643712 131219 648752
rect 136259 643712 437023 648752
rect 13472 643688 437023 643712
rect 13472 643687 13496 643688
rect 8358 643663 13496 643687
rect 8366 638743 13488 638767
rect 8366 633669 8390 638743
rect 13464 638742 13488 638743
rect 436999 638742 437023 643688
rect 13464 638718 437023 638742
rect 13464 633694 131043 638718
rect 136067 633694 437023 638718
rect 13464 633670 437023 633694
rect 13464 633669 13488 633670
rect 8366 633645 13488 633669
rect 436999 629601 437023 633670
rect 442234 644694 442258 648802
rect 559596 644694 560642 644711
rect 570793 644695 575945 644719
rect 570793 644694 570817 644695
rect 442234 644687 570817 644694
rect 442234 639595 559620 644687
rect 560618 639595 570817 644687
rect 442234 639592 570817 639595
rect 442234 634674 442258 639592
rect 559596 639571 560642 639592
rect 570793 639591 570817 639592
rect 575921 639591 575945 644695
rect 570793 639567 575945 639591
rect 559587 634721 560633 634745
rect 559587 634674 559611 634721
rect 442234 629638 559611 634674
rect 442234 629601 442258 629638
rect 559587 629629 559611 629638
rect 560609 634674 560633 634721
rect 570848 634675 575934 634699
rect 570848 634674 570872 634675
rect 560609 629638 570872 634674
rect 560609 629629 560633 629638
rect 559587 629605 560633 629629
rect 570848 629637 570872 629638
rect 575910 629637 575934 634675
rect 570848 629613 575934 629637
rect 436999 629577 442258 629601
rect 118304 614123 123470 614147
rect 118304 609005 118328 614123
rect 123446 614099 454775 614123
rect 123446 609029 449681 614099
rect 454751 609029 454775 614099
rect 123446 609005 454775 609029
rect 118304 608981 123470 609005
rect 130960 584235 136145 584259
rect 130960 581875 130984 584235
rect 136121 584062 136145 584235
rect 437013 584137 442196 584161
rect 378768 584076 379493 584100
rect 378768 584062 378792 584076
rect 136121 582062 181559 584062
rect 338673 582062 378792 584062
rect 136121 581875 136145 582062
rect 378768 582061 378792 582062
rect 379469 584062 379493 584076
rect 396560 584080 397285 584104
rect 396560 584062 396584 584080
rect 379469 582065 396584 584062
rect 397261 584062 397285 584080
rect 437013 584062 437037 584137
rect 397261 582065 437037 584062
rect 379469 582062 437037 582065
rect 379469 582061 379493 582062
rect 378768 582037 379493 582061
rect 396560 582041 397285 582062
rect 437013 581960 437037 582062
rect 442172 581960 442196 584137
rect 437013 581936 442196 581960
rect 130960 581851 136145 581875
rect 118330 580341 123298 580365
rect 118330 577835 118354 580341
rect 123274 580062 123298 580341
rect 449623 580116 454811 580140
rect 377421 580062 378320 580073
rect 397834 580068 398559 580092
rect 397834 580062 397858 580068
rect 123274 578062 179747 580062
rect 338673 580049 397858 580062
rect 338673 578103 377445 580049
rect 378296 578103 397858 580049
rect 338673 578062 397858 578103
rect 123274 577835 123298 578062
rect 397834 578053 397858 578062
rect 398535 580062 398559 580068
rect 449623 580062 449647 580116
rect 398535 578062 449647 580062
rect 398535 578053 398559 578062
rect 397834 578029 398559 578053
rect 449623 577998 449647 578062
rect 454787 580062 454811 580116
rect 454787 579329 539492 580062
rect 454787 578715 537803 579329
rect 538405 578715 539492 579329
rect 454787 578062 539492 578715
rect 454787 577998 454811 578062
rect 449623 577974 454811 577998
rect 118330 577811 123298 577835
rect 437032 556351 442232 556375
rect 437032 556202 437056 556351
rect 409002 554202 437056 556202
rect 437032 554088 437056 554202
rect 442208 556202 442232 556351
rect 526584 556202 527232 556206
rect 442208 556182 571610 556202
rect 442208 556160 526608 556182
rect 442208 554242 509408 556160
rect 509938 554242 526608 556160
rect 442208 554236 526608 554242
rect 527208 556178 571610 556182
rect 527208 554236 547182 556178
rect 442208 554212 547182 554236
rect 547758 556132 571610 556178
rect 547758 554240 559640 556132
rect 560562 554240 571610 556132
rect 547758 554212 571610 554240
rect 442208 554202 571610 554212
rect 442208 554088 442232 554202
rect 547158 554188 547782 554202
rect 437032 554064 442232 554088
rect 449612 540461 454812 540485
rect 449612 540310 449636 540461
rect 408468 538310 449636 540310
rect 449612 538198 449636 538310
rect 454788 540310 454812 540461
rect 537810 540310 538434 540318
rect 454788 540294 571610 540310
rect 454788 540212 537834 540294
rect 454788 539637 517874 540212
rect 454788 539563 500437 539637
rect 454788 539453 484634 539563
rect 454788 538839 464243 539453
rect 464845 538949 484634 539453
rect 485236 539035 500437 539563
rect 501051 539035 517874 539637
rect 485236 538949 517874 539035
rect 464845 538839 517874 538949
rect 454788 538396 517874 538839
rect 518574 538396 537834 540212
rect 454788 538328 537834 538396
rect 538410 540236 571610 540294
rect 538410 538344 565238 540236
rect 566160 538344 571610 540236
rect 538410 538328 571610 538344
rect 454788 538310 571610 538328
rect 454788 538198 454812 538310
rect 537810 538304 538434 538310
rect 449612 538174 454812 538198
rect 449688 531568 454837 531592
rect 449688 531548 449712 531568
rect 401948 530928 449712 531548
rect 449688 530898 449712 530928
rect 454813 530898 454837 531568
rect 449688 530874 454837 530898
rect 437024 530351 442173 530375
rect 437024 530308 437048 530351
rect 401922 529688 437048 530308
rect 437024 529681 437048 529688
rect 442149 529681 442173 530351
rect 437024 529657 442173 529681
rect 437079 513406 442228 513430
rect 437079 513368 437103 513406
rect 402069 512748 437103 513368
rect 437079 512736 437103 512748
rect 442204 512736 442228 513406
rect 437079 512712 442228 512736
rect 449647 512175 454796 512199
rect 449647 512128 449671 512175
rect 401970 511508 449671 512128
rect 449647 511505 449671 511508
rect 454772 511505 454796 512175
rect 449647 511481 454796 511505
rect 437028 486137 442228 486161
rect 437028 485956 437052 486137
rect 352292 485283 437052 485956
rect 352292 485153 375483 485283
rect 352292 484611 360437 485153
rect 360991 484741 375483 485153
rect 376037 485223 437052 485283
rect 376037 485217 434799 485223
rect 376037 485207 390323 485217
rect 376037 484741 386089 485207
rect 360991 484665 386089 484741
rect 386643 484675 390323 485207
rect 390877 485215 434799 485217
rect 390877 485187 428635 485215
rect 390877 484675 400217 485187
rect 386643 484665 400217 484675
rect 360991 484645 400217 484665
rect 400771 484673 428635 485187
rect 429189 484673 434799 485215
rect 400771 484645 434799 484673
rect 360991 484621 434799 484645
rect 435413 484621 437052 485223
rect 360991 484611 437052 484621
rect 352292 483956 437052 484611
rect 437028 483874 437052 483956
rect 442204 485956 442228 486137
rect 442204 485896 569028 485956
rect 442204 485313 559636 485896
rect 442204 484711 458513 485313
rect 459127 485221 559636 485313
rect 459127 485201 511838 485221
rect 459127 485163 484622 485201
rect 459127 484711 464284 485163
rect 442204 484561 464284 484711
rect 464898 485133 484622 485163
rect 464898 484561 475003 485133
rect 442204 484531 475003 484561
rect 475617 484587 484622 485133
rect 485224 485171 511838 485201
rect 485224 485117 504621 485171
rect 485224 484587 498497 485117
rect 475617 484531 498497 484587
rect 442204 484503 498497 484531
rect 499099 484569 504621 485117
rect 505235 484607 511838 485171
rect 512440 484607 518207 485221
rect 505235 484579 518207 484607
rect 518837 485215 559636 485221
rect 518837 485179 531885 485215
rect 518837 485165 530383 485179
rect 518837 484579 524296 485165
rect 505235 484569 524296 484579
rect 499099 484551 524296 484569
rect 524898 484577 530383 485165
rect 530997 484585 531885 485179
rect 532527 485133 559636 485215
rect 532527 484585 545778 485133
rect 530997 484577 545778 484585
rect 524898 484551 545778 484577
rect 499099 484503 545778 484551
rect 442204 484491 545778 484503
rect 546408 484491 559636 485133
rect 442204 484004 559636 484491
rect 560558 485177 569028 485896
rect 560558 484535 567855 485177
rect 568485 484535 569028 485177
rect 560558 484004 569028 484535
rect 442204 483956 569028 484004
rect 442204 483874 442228 483956
rect 437028 483850 442228 483874
rect 449618 474001 454818 474025
rect 449618 473822 449642 474001
rect 352440 473165 449642 473822
rect 352440 472987 380563 473165
rect 352440 472433 352775 472987
rect 353317 472611 380563 472987
rect 381105 473151 449642 473165
rect 381105 473077 394691 473151
rect 381105 472611 389485 473077
rect 353317 472535 389485 472611
rect 390039 472609 394691 473077
rect 395245 473115 449642 473151
rect 395245 473103 428289 473115
rect 395245 472609 400585 473103
rect 390039 472561 400585 472609
rect 401139 472573 428289 473103
rect 428843 473053 449642 473115
rect 428843 472573 445477 473053
rect 401139 472561 445477 472573
rect 390039 472535 445477 472561
rect 353317 472451 445477 472535
rect 446091 472451 449642 473053
rect 353317 472433 449642 472451
rect 352440 471822 449642 472433
rect 449618 471738 449642 471822
rect 454794 473822 454818 474001
rect 454794 473748 569028 473822
rect 454794 473213 565224 473748
rect 454794 473188 548147 473213
rect 454794 473097 497346 473188
rect 454794 473053 485291 473097
rect 454794 472451 462129 473053
rect 462743 472495 485291 473053
rect 485905 472560 497346 473097
rect 497986 473169 548147 473188
rect 497986 473097 536949 473169
rect 497986 473093 522944 473097
rect 497986 473007 518229 473093
rect 497986 472992 506689 473007
rect 497986 472560 503854 472992
rect 485905 472495 503854 472560
rect 462743 472451 503854 472495
rect 454794 472364 503854 472451
rect 504494 472393 506689 472992
rect 507291 472479 518229 473007
rect 518831 472495 522944 473093
rect 525127 472555 536949 473097
rect 537551 473147 548147 473169
rect 537551 472555 537963 473147
rect 525127 472505 537963 472555
rect 538593 472571 548147 473147
rect 548777 473137 565224 473213
rect 548777 472571 553169 473137
rect 538593 472505 553169 472571
rect 525127 472495 553169 472505
rect 553799 473065 565224 473137
rect 553799 472495 562797 473065
rect 518831 472479 562797 472495
rect 507291 472435 562797 472479
rect 563439 472435 565224 473065
rect 507291 472393 565224 472435
rect 504494 472364 565224 472393
rect 454794 471856 565224 472364
rect 566146 471856 569028 473748
rect 454794 471822 569028 471856
rect 454794 471738 454818 471822
rect 449618 471714 454818 471738
rect 449650 467421 454850 467445
rect 118278 467391 123478 467415
rect 118278 467280 118302 467391
rect 118170 465280 118302 467280
rect 118278 465128 118302 465280
rect 123454 467280 123478 467391
rect 377488 467291 378253 467315
rect 377488 467280 377512 467291
rect 123454 465280 180364 467280
rect 338673 465285 377512 467280
rect 378229 467280 378253 467291
rect 397830 467290 398595 467314
rect 397830 467280 397854 467290
rect 378229 465285 397854 467280
rect 338673 465284 397854 465285
rect 398571 467280 398595 467290
rect 449650 467280 449674 467421
rect 398571 465284 449674 467280
rect 338673 465280 449674 465284
rect 123454 465128 123478 465280
rect 377488 465261 378253 465280
rect 397830 465260 398595 465280
rect 449650 465158 449674 465280
rect 454826 465158 454850 467421
rect 449650 465134 454850 465158
rect 118278 465104 123478 465128
rect 437034 463376 442234 463400
rect 130859 463295 136059 463319
rect 130859 463280 130883 463295
rect 130434 461280 130883 463280
rect 130859 461032 130883 461280
rect 136035 463280 136059 463295
rect 378758 463289 379523 463313
rect 378758 463280 378782 463289
rect 136035 461280 180216 463280
rect 338673 461283 378782 463280
rect 379499 463280 379523 463289
rect 396557 463280 397322 463301
rect 437034 463280 437058 463376
rect 379499 463277 437058 463280
rect 379499 461283 396581 463277
rect 338673 461280 396581 461283
rect 136035 461032 136059 461280
rect 378758 461259 379523 461280
rect 396557 461271 396581 461280
rect 397298 461280 437058 463277
rect 397298 461271 397322 461280
rect 396557 461247 397322 461271
rect 437034 461113 437058 461280
rect 442210 463280 442234 463376
rect 442210 461280 442485 463280
rect 442210 461113 442234 461280
rect 437034 461089 442234 461113
rect 130859 461008 136059 461032
rect 437024 431177 442224 431201
rect 130926 431115 136126 431139
rect 130926 428852 130950 431115
rect 136102 431050 136126 431115
rect 437024 431050 437048 431177
rect 136102 430698 437048 431050
rect 136102 430385 348094 430698
rect 136102 430265 249229 430385
rect 136102 429712 238860 430265
rect 239401 429843 249229 430265
rect 249773 430377 348094 430385
rect 249773 430369 332863 430377
rect 249773 429843 252974 430369
rect 239401 429827 252974 429843
rect 253528 430368 332863 430369
rect 253528 429827 258344 430368
rect 239401 429816 258344 429827
rect 258884 430361 332863 430368
rect 258884 430349 293220 430361
rect 258884 430293 278456 430349
rect 258884 429816 272934 430293
rect 239401 429751 272934 429816
rect 273488 429795 278456 430293
rect 278998 429807 293220 430349
rect 293762 430261 332863 430361
rect 293762 429807 299168 430261
rect 278998 429795 299168 429807
rect 273488 429751 299168 429795
rect 239401 429712 299168 429751
rect 136102 429707 299168 429712
rect 299710 430221 332863 430261
rect 299710 430197 322091 430221
rect 299710 429707 313342 430197
rect 136102 429655 313342 429707
rect 313896 430163 322091 430197
rect 313896 429655 319482 430163
rect 136102 429609 319482 429655
rect 320024 429667 322091 430163
rect 322633 429835 332863 430221
rect 333417 430259 348094 430377
rect 333417 429835 335400 430259
rect 322633 429705 335400 429835
rect 335942 429705 348094 430259
rect 322633 429667 348094 429705
rect 320024 429609 348094 429667
rect 136102 429382 348094 429609
rect 348522 430445 437048 430698
rect 348522 430263 359995 430445
rect 348522 429721 354351 430263
rect 354905 429903 359995 430263
rect 360549 430437 437048 430445
rect 360549 429903 362165 430437
rect 354905 429895 362165 429903
rect 362719 430377 437048 430437
rect 362719 430293 391199 430377
rect 362719 430201 385927 430293
rect 362719 430197 375346 430201
rect 362719 429895 373956 430197
rect 354905 429721 373956 429895
rect 348522 429643 373956 429721
rect 374498 429659 375346 430197
rect 375900 429739 385927 430201
rect 386469 429823 391199 430293
rect 391741 429823 437048 430377
rect 386469 429739 437048 429823
rect 375900 429659 437048 429739
rect 374498 429643 437048 429659
rect 348522 429382 437048 429643
rect 136102 429050 437048 429382
rect 136102 428852 136126 429050
rect 437024 428914 437048 429050
rect 442200 431050 442224 431177
rect 442200 431014 568562 431050
rect 442200 430409 559662 431014
rect 442200 430404 545777 430409
rect 442200 429776 497204 430404
rect 497844 430341 545777 430404
rect 497844 430291 513061 430341
rect 497844 429776 510277 430291
rect 442200 429689 510277 429776
rect 510891 429739 513061 430291
rect 513675 430335 545777 430341
rect 513675 430307 528965 430335
rect 513675 429739 522305 430307
rect 510891 429693 522305 429739
rect 522907 429693 528965 430307
rect 529595 429767 545777 430335
rect 546407 429767 559662 430409
rect 529595 429693 559662 429767
rect 510891 429689 559662 429693
rect 442200 429122 559662 429689
rect 560584 430323 568562 431014
rect 560584 429693 562795 430323
rect 563437 429693 568562 430323
rect 560584 429122 568562 429693
rect 442200 429050 568562 429122
rect 442200 428914 442224 429050
rect 437024 428890 442224 428914
rect 130926 428828 136126 428852
rect 449610 416727 454810 416751
rect 118280 416703 123480 416727
rect 118280 414440 118304 416703
rect 123456 416606 123480 416703
rect 449610 416606 449634 416727
rect 123456 416210 449634 416606
rect 123456 415953 345550 416210
rect 123456 415918 319472 415953
rect 123456 415907 252978 415918
rect 123456 415366 242013 415907
rect 242566 415366 252978 415907
rect 253518 415882 319472 415918
rect 253518 415721 258330 415882
rect 253518 415366 255267 415721
rect 123456 415179 255267 415366
rect 255821 415342 258330 415721
rect 258882 415877 319472 415882
rect 258882 415821 313348 415877
rect 258882 415815 278444 415821
rect 258882 415342 272926 415815
rect 255821 415273 272926 415342
rect 273480 415279 278444 415815
rect 278998 415819 313348 415821
rect 278998 415795 299130 415819
rect 278998 415279 293220 415795
rect 273480 415273 293220 415279
rect 255821 415241 293220 415273
rect 293762 415277 299130 415795
rect 299684 415323 313348 415819
rect 313890 415399 319472 415877
rect 320014 415907 345550 415953
rect 320014 415399 328165 415907
rect 313890 415353 328165 415399
rect 328707 415869 345550 415907
rect 328707 415353 339881 415869
rect 313890 415323 339881 415353
rect 299684 415315 339881 415323
rect 340423 415315 345550 415869
rect 299684 415277 345550 415315
rect 293762 415241 345550 415277
rect 255821 415179 345550 415241
rect 123456 414894 345550 415179
rect 345978 415933 449634 416210
rect 345978 415855 393659 415933
rect 345978 415851 388623 415855
rect 345978 415769 373938 415851
rect 345978 415227 353567 415769
rect 354121 415297 373938 415769
rect 374480 415655 388623 415851
rect 374480 415297 375346 415655
rect 354121 415227 375346 415297
rect 345978 415101 375346 415227
rect 375888 415301 388623 415655
rect 389165 415391 393659 415855
rect 394213 415391 449634 415933
rect 389165 415301 449634 415391
rect 375888 415101 449634 415301
rect 345978 414894 449634 415101
rect 123456 414606 449634 414894
rect 123456 414440 123480 414606
rect 449610 414464 449634 414606
rect 454786 416606 454810 416727
rect 454786 416560 568562 416606
rect 454786 414668 565236 416560
rect 566158 414668 568562 416560
rect 454786 414606 568562 414668
rect 454786 414464 454810 414606
rect 449610 414440 454810 414464
rect 118280 414416 123480 414440
rect 437020 392083 442220 392107
rect 437020 391948 437044 392083
rect 318284 391373 437044 391948
rect 318284 391353 333086 391373
rect 318284 390799 322889 391353
rect 323431 390819 333086 391353
rect 333628 391315 437044 391373
rect 333628 390819 334873 391315
rect 323431 390799 334873 390819
rect 318284 390761 334873 390799
rect 335415 391303 437044 391315
rect 335415 391199 428495 391303
rect 335415 391163 367490 391199
rect 335415 390945 357696 391163
rect 335415 390761 353559 390945
rect 318284 390403 353559 390761
rect 354113 390609 357696 390945
rect 358238 390645 367490 391163
rect 368032 391195 428495 391199
rect 368032 391175 400431 391195
rect 368032 390645 385263 391175
rect 358238 390621 385263 390645
rect 385805 390641 400431 391175
rect 400973 390761 428495 391195
rect 429049 390761 437044 391303
rect 400973 390641 437044 390761
rect 385805 390621 437044 390641
rect 358238 390609 437044 390621
rect 354113 390403 437044 390609
rect 318284 389948 437044 390403
rect 437020 389820 437044 389948
rect 442196 391948 442220 392083
rect 442196 391876 571940 391948
rect 442196 391247 559660 391876
rect 442196 391153 546397 391247
rect 442196 391111 530391 391153
rect 442196 391061 490275 391111
rect 442196 391055 470033 391061
rect 442196 390501 446401 391055
rect 446943 390507 470033 391055
rect 470575 390557 490275 391061
rect 490817 391081 530391 391111
rect 490817 390557 510729 391081
rect 470575 390527 510729 390557
rect 511271 390599 530391 391081
rect 530933 390673 546397 391153
rect 546959 390673 559660 391247
rect 530933 390599 559660 390673
rect 511271 390527 559660 390599
rect 470575 390507 559660 390527
rect 446943 390501 559660 390507
rect 442196 389984 559660 390501
rect 560582 391211 571940 391876
rect 560582 390637 571233 391211
rect 571795 390637 571940 391211
rect 560582 389984 571940 390637
rect 442196 389948 571940 389984
rect 442196 389820 442220 389948
rect 437020 389796 442220 389820
rect 449620 377007 454820 377031
rect 449620 376832 449644 377007
rect 318676 376280 449644 376832
rect 318676 376215 352330 376280
rect 318676 376101 333084 376215
rect 318676 375547 325771 376101
rect 326313 375673 333084 376101
rect 333638 376109 352330 376215
rect 333638 375673 337327 376109
rect 326313 375567 337327 375673
rect 337881 376095 352330 376109
rect 337881 375567 345675 376095
rect 326313 375553 345675 375567
rect 346229 375608 352330 376095
rect 353838 376107 449644 376280
rect 353838 375608 357690 376107
rect 346229 375553 357690 375608
rect 358232 376057 400419 376107
rect 358232 375553 367490 376057
rect 326313 375547 367490 375553
rect 318676 375503 367490 375547
rect 368032 375925 400419 376057
rect 368032 375503 388565 375925
rect 318676 375371 388565 375503
rect 389107 375553 400419 375925
rect 400961 376071 449644 376107
rect 400961 376013 446405 376071
rect 400961 375553 429155 376013
rect 389107 375459 429155 375553
rect 429697 375517 446405 376013
rect 446947 375517 449644 376071
rect 429697 375459 449644 375517
rect 389107 375371 449644 375459
rect 318676 374832 449644 375371
rect 449620 374744 449644 374832
rect 454796 376832 454820 377007
rect 454796 376796 572106 376832
rect 454796 376175 565224 376796
rect 454796 376055 526311 376175
rect 454796 375501 466543 376055
rect 467085 376011 526311 376055
rect 467085 375501 485503 376011
rect 454796 375457 485503 375501
rect 486045 375995 526311 376011
rect 486045 375457 505739 375995
rect 454796 375441 505739 375457
rect 506281 375621 526311 375995
rect 526853 376115 565224 376175
rect 526853 376053 562703 376115
rect 526853 375621 552367 376053
rect 506281 375479 552367 375621
rect 552929 375553 562703 376053
rect 563277 375553 565224 376115
rect 552929 375479 565224 375553
rect 506281 375441 565224 375479
rect 454796 374904 565224 375441
rect 566146 374904 572106 376796
rect 454796 374832 572106 374904
rect 454796 374744 454820 374832
rect 449620 374720 454820 374744
rect 437010 307769 442210 307793
rect 348000 307624 348500 307642
rect 437010 307624 437034 307769
rect 344000 307618 437034 307624
rect 344000 305644 348024 307618
rect 348476 306934 437034 307618
rect 348476 306806 390694 306934
rect 348476 306785 370682 306806
rect 348476 306243 357939 306785
rect 358493 306257 370682 306785
rect 371243 306385 390694 306806
rect 391255 306892 437034 306934
rect 391255 306385 400258 306892
rect 371243 306343 400258 306385
rect 400819 306656 437034 306892
rect 400819 306343 430708 306656
rect 371243 306257 430708 306343
rect 358493 306243 430708 306257
rect 348476 306107 430708 306243
rect 431269 306107 437034 306656
rect 348476 305644 437034 306107
rect 344000 305624 437034 305644
rect 348000 305620 348500 305624
rect 437010 305506 437034 305624
rect 442186 307624 442210 307769
rect 442186 307562 570998 307624
rect 442186 307010 559644 307562
rect 442186 306854 490720 307010
rect 442186 306305 445434 306854
rect 445995 306786 490720 306854
rect 445995 306305 470724 306786
rect 442186 306225 470724 306305
rect 471273 306449 490720 306786
rect 491269 306902 559644 307010
rect 491269 306449 510706 306902
rect 471273 306341 510706 306449
rect 511255 306748 559644 306902
rect 511255 306341 530680 306748
rect 471273 306225 530680 306341
rect 442186 306187 530680 306225
rect 531229 306736 559644 306748
rect 531229 306187 552161 306736
rect 442186 306167 552161 306187
rect 552718 306167 559644 306736
rect 442186 305670 559644 306167
rect 560566 306812 570998 307562
rect 560566 306243 569352 306812
rect 569933 306243 570998 306812
rect 560566 305670 570998 306243
rect 442186 305624 570998 305670
rect 442186 305506 442210 305624
rect 437010 305482 442210 305506
rect 449626 287781 454826 287805
rect 345686 287600 346186 287612
rect 449626 287600 449650 287781
rect 343250 287588 449650 287600
rect 343250 285614 345710 287588
rect 346162 287027 449650 287588
rect 346162 286909 445446 287027
rect 346162 286819 400174 286909
rect 346162 286265 354035 286819
rect 354577 286697 400174 286819
rect 354577 286613 390694 286697
rect 354577 286265 370694 286613
rect 346162 286052 370694 286265
rect 371243 286148 390694 286613
rect 391255 286360 400174 286697
rect 400735 286815 445446 286909
rect 400735 286360 430708 286815
rect 391255 286266 430708 286360
rect 431269 286478 445446 286815
rect 446007 286478 449650 287027
rect 431269 286266 449650 286478
rect 391255 286148 449650 286266
rect 371243 286052 449650 286148
rect 346162 285614 449650 286052
rect 343250 285600 449650 285614
rect 345686 285590 346186 285600
rect 449626 285518 449650 285600
rect 454802 287600 454826 287781
rect 454802 287548 570476 287600
rect 454802 286989 565232 287548
rect 454802 286889 546314 286989
rect 454802 286759 490720 286889
rect 454802 286198 470724 286759
rect 471273 286328 490720 286759
rect 491269 286825 546314 286889
rect 491269 286328 510706 286825
rect 471273 286264 510706 286328
rect 511255 286813 546314 286825
rect 511255 286264 530692 286813
rect 471273 286252 530692 286264
rect 531241 286420 546314 286813
rect 546871 286420 565232 286989
rect 531241 286252 565232 286420
rect 471273 286198 565232 286252
rect 454802 285656 565232 286198
rect 566154 286888 570476 287548
rect 566154 286319 568312 286888
rect 568893 286319 570476 286888
rect 566154 285656 570476 286319
rect 454802 285600 570476 285656
rect 454802 285518 454826 285600
rect 449626 285494 454826 285518
rect 130997 213150 136133 213174
rect 130997 208062 131021 213150
rect 136109 213126 442176 213150
rect 136109 213096 356470 213126
rect 136109 208088 347982 213096
rect 348448 208088 356470 213096
rect 136109 208086 356470 208088
rect 361510 208086 437112 213126
rect 442152 208086 442176 213126
rect 136109 208062 442176 208086
rect 130997 208038 136133 208062
rect 565163 196299 566218 196323
rect 565163 196290 565187 196299
rect 449499 196266 565187 196290
rect 449499 191354 449523 196266
rect 454435 191354 565187 196266
rect 449499 191348 565187 191354
rect 566194 196290 566218 196299
rect 570476 196291 575484 196315
rect 570476 196290 570500 196291
rect 566194 191348 570500 196290
rect 449499 191330 570500 191348
rect 565163 191324 566218 191330
rect 570476 191329 570500 191330
rect 575460 191329 575484 196291
rect 570476 191305 575484 191329
rect 570389 186371 575557 186395
rect 570389 186370 570413 186371
rect 449420 186346 570413 186370
rect 449420 181276 449444 186346
rect 454514 186266 570413 186346
rect 454514 181315 565206 186266
rect 566213 181315 570413 186266
rect 454514 181276 570413 181315
rect 449420 181252 570413 181276
rect 570389 181251 570413 181252
rect 575533 181251 575557 186371
rect 570389 181227 575557 181251
rect 13041 177861 18209 177885
rect 13041 172741 13065 177861
rect 18185 177860 18209 177861
rect 18185 177836 454970 177860
rect 18185 177806 118328 177836
rect 18185 172855 24981 177806
rect 25988 172855 118328 177806
rect 18185 172766 118328 172855
rect 123398 172766 332587 177836
rect 337657 177826 449876 177836
rect 337657 172818 345722 177826
rect 346188 172818 449876 177826
rect 337657 172766 449876 172818
rect 454946 172766 454970 177836
rect 18185 172742 454970 172766
rect 18185 172741 18209 172742
rect 13041 172717 18209 172741
rect 13349 167863 18517 167887
rect 13349 162743 13373 167863
rect 18493 167862 18517 167863
rect 18493 167838 454832 167862
rect 18493 167760 118194 167838
rect 18493 162809 25000 167760
rect 26007 162809 118194 167760
rect 18493 162768 118194 162809
rect 123264 167836 449738 167838
rect 123264 162828 345698 167836
rect 346164 162828 449738 167836
rect 123264 162768 449738 162828
rect 454808 162768 454832 167838
rect 18493 162744 454832 162768
rect 18493 162743 18517 162744
rect 13349 162719 18517 162743
rect 332539 61843 337705 61867
rect 38445 60006 332563 61843
rect 38445 58752 90284 60006
rect 91538 59509 332563 60006
rect 91538 59387 302585 59509
rect 91538 59377 240069 59387
rect 91538 59367 133043 59377
rect 91538 58825 111721 59367
rect 112275 58835 133043 59367
rect 133597 59333 240069 59377
rect 133597 58835 154601 59333
rect 112275 58825 154601 58835
rect 91538 58791 154601 58825
rect 155155 58791 175807 59333
rect 176361 59311 240069 59333
rect 176361 59289 219083 59311
rect 176361 58791 197189 59289
rect 91538 58752 197189 58791
rect 38445 58747 197189 58752
rect 197743 58769 219083 59289
rect 219637 58845 240069 59311
rect 240623 59385 302585 59387
rect 240623 58845 260583 59385
rect 219637 58831 260583 58845
rect 261125 59141 302585 59385
rect 261125 58831 281395 59141
rect 219637 58769 281395 58831
rect 197743 58747 281395 58769
rect 38445 58587 281395 58747
rect 281937 58955 302585 59141
rect 303127 58955 324121 59509
rect 324663 58955 332563 59509
rect 281937 58587 332563 58955
rect 38445 56725 332563 58587
rect 337681 56725 337705 61843
rect 39905 52891 40867 56725
rect 332539 56701 337705 56725
rect 39875 52867 40897 52891
rect 39875 51905 39899 52867
rect 40873 51905 40897 52867
rect 39875 51881 40897 51905
rect 356422 40402 361558 40426
rect 38042 39258 356446 40402
rect 38042 36270 39650 39258
rect 42762 38007 356446 39258
rect 42762 37901 69297 38007
rect 42762 37359 48003 37901
rect 48557 37465 69297 37901
rect 69851 37927 356446 38007
rect 69851 37829 197191 37927
rect 69851 37741 154603 37829
rect 69851 37689 111723 37741
rect 69851 37465 90663 37689
rect 48557 37359 90663 37465
rect 42762 37147 90663 37359
rect 91217 37199 111723 37689
rect 112277 37673 154603 37741
rect 112277 37199 133057 37673
rect 91217 37147 133057 37199
rect 42762 37119 133057 37147
rect 133599 37287 154603 37673
rect 155157 37287 175809 37829
rect 176363 37385 197191 37829
rect 197745 37925 356446 37927
rect 197745 37877 302575 37925
rect 197745 37385 219085 37877
rect 176363 37335 219085 37385
rect 219639 37821 302575 37877
rect 219639 37787 281385 37821
rect 219639 37335 240071 37787
rect 176363 37287 240071 37335
rect 133599 37233 240071 37287
rect 240613 37725 281385 37787
rect 240613 37233 260573 37725
rect 133599 37171 260573 37233
rect 261115 37267 281385 37725
rect 281927 37371 302575 37821
rect 303117 37873 356446 37925
rect 303117 37371 324123 37873
rect 281927 37319 324123 37371
rect 324665 37319 356446 37873
rect 281927 37267 356446 37319
rect 261115 37171 356446 37267
rect 133599 37119 356446 37171
rect 42762 36270 356446 37119
rect 38042 35314 356446 36270
rect 361534 35314 361558 40402
rect 356422 35290 361558 35314
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use analog_top  analog_top_0
timestamp 1655456512
transform 1 0 173490 0 1 497666
box 4703 -40917 166970 91353
use digital_filter  digital_filter_0
timestamp 1655456512
transform 1 0 373631 0 1 507651
box 0 0 28796 27744
use sky130_fd_pr__cap_mim_m3_1_PXTAZD  sky130_fd_pr__cap_mim_m3_1_PXTAZD_0
timestamp 1655456512
transform 1 0 155484 0 1 524150
box -12624 -25192 12470 25192
use sky130_fd_pr__cap_mim_m3_1_PXTAZD  sky130_fd_pr__cap_mim_m3_1_PXTAZD_1
timestamp 1655456512
transform 1 0 155188 0 1 374916
box -12624 -25192 12470 25192
use sky130_fd_pr__cap_mim_m3_1_PXTAZD  sky130_fd_pr__cap_mim_m3_1_PXTAZD_2
timestamp 1655456512
transform 1 0 155188 0 1 308808
box -12624 -25192 12470 25192
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655456512
transform 0 -1 251696 1 0 455368
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_1
timestamp 1655456512
transform 0 -1 251679 1 0 433587
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_2
timestamp 1655456512
transform -1 0 278971 0 1 420349
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_3
timestamp 1655456512
transform -1 0 258837 0 1 420316
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_4
timestamp 1655456512
transform -1 0 319976 0 1 420307
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_5
timestamp 1655456512
transform -1 0 299648 0 1 420355
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_6
timestamp 1655456512
transform 0 -1 336827 1 0 416578
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_7
timestamp 1655456512
transform 1 0 353674 0 1 420316
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_8
timestamp 1655456512
transform 1 0 374017 0 1 420386
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_9
timestamp 1655456512
transform 0 -1 388177 1 0 427201
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_10
timestamp 1655456512
transform 0 -1 388148 1 0 448244
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_11
timestamp 1655456512
transform 0 -1 388187 1 0 469264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_12
timestamp 1655456512
transform 0 -1 388178 1 0 490228
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_13
timestamp 1655456512
transform 0 -1 336852 1 0 395925
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_14
timestamp 1655456512
transform -1 0 347971 0 1 386451
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_15
timestamp 1655456512
transform -1 0 367987 0 1 386480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_16
timestamp 1655456512
transform -1 0 387799 0 1 386470
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_17
timestamp 1655456512
transform -1 0 408058 0 1 386468
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_18
timestamp 1655456512
transform -1 0 428334 0 1 386523
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_19
timestamp 1655456512
transform -1 0 448493 0 1 386503
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_20
timestamp 1655456512
transform -1 0 468495 0 1 386498
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_21
timestamp 1655456512
transform -1 0 488613 0 1 386482
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_22
timestamp 1655456512
transform -1 0 508743 0 1 386505
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_23
timestamp 1655456512
transform -1 0 528852 0 1 386519
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_24
timestamp 1655456512
transform 0 -1 549833 -1 0 388239
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_25
timestamp 1655456512
transform 0 -1 549816 -1 0 407283
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_26
timestamp 1655456512
transform -1 0 568571 0 1 408715
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_27
timestamp 1655456512
transform 0 -1 240974 1 0 455390
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_28
timestamp 1655456512
transform 0 -1 240894 1 0 433873
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_29
timestamp 1655456512
transform -1 0 253483 0 1 425814
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_30
timestamp 1655456512
transform -1 0 273429 0 1 425879
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_31
timestamp 1655456512
transform -1 0 293710 0 1 425913
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_32
timestamp 1655456512
transform -1 0 313859 0 1 425903
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_33
timestamp 1655456512
transform 1 0 355444 0 1 425884
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_34
timestamp 1655456512
transform 1 0 335454 0 1 425888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_35
timestamp 1655456512
transform 1 0 375407 0 1 425978
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_36
timestamp 1655456512
transform 0 -1 393101 1 0 427220
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_37
timestamp 1655456512
transform 0 -1 393069 1 0 448312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_38
timestamp 1655456512
transform 0 -1 393079 1 0 469264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_39
timestamp 1655456512
transform 0 -1 393081 1 0 490242
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_40
timestamp 1655456512
transform 0 -1 324817 1 0 416653
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_41
timestamp 1655456512
transform 0 -1 324815 1 0 395863
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_42
timestamp 1655456512
transform -1 0 333602 0 1 380484
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_43
timestamp 1655456512
transform -1 0 358181 0 1 380492
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_44
timestamp 1655456512
transform -1 0 387628 0 1 380450
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_45
timestamp 1655456512
transform -1 0 408206 0 1 380481
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_46
timestamp 1655456512
transform -1 0 428180 0 1 380456
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_47
timestamp 1655456512
transform -1 0 448426 0 1 380460
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_48
timestamp 1655456512
transform -1 0 468410 0 1 380527
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_49
timestamp 1655456512
transform -1 0 488825 0 1 380452
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_50
timestamp 1655456512
transform -1 0 508508 0 1 380524
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_51
timestamp 1655456512
transform -1 0 528878 0 1 380458
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_52
timestamp 1655456512
transform 0 -1 549641 1 0 378969
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_53
timestamp 1655456512
transform 0 -1 549602 1 0 363783
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_54
timestamp 1655456512
transform -1 0 568727 0 1 362332
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_55
timestamp 1655456512
transform 0 -1 383541 1 0 490147
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_56
timestamp 1655456512
transform 0 -1 373889 1 0 490149
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_57
timestamp 1655456512
transform -1 0 379576 0 -1 475772
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_58
timestamp 1655456512
transform -1 0 400066 0 -1 475805
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_59
timestamp 1655456512
transform -1 0 420308 0 -1 475745
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_60
timestamp 1655456512
transform -1 0 460846 0 -1 475786
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_61
timestamp 1655456512
transform -1 0 440546 0 -1 475774
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_62
timestamp 1655456512
transform -1 0 481028 0 -1 475764
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_63
timestamp 1655456512
transform -1 0 501016 0 -1 475782
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_64
timestamp 1655456512
transform 0 1 521261 -1 0 457251
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_65
timestamp 1655456512
transform 0 -1 502473 1 0 454712
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_66
timestamp 1655456512
transform 0 1 508811 -1 0 449125
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_67
timestamp 1655456512
transform 0 1 508823 -1 0 469176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_68
timestamp 1655456512
transform 0 -1 515296 1 0 467306
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_69
timestamp 1655456512
transform -1 0 523466 0 1 475219
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_70
timestamp 1655456512
transform 0 -1 515333 1 0 447105
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_71
timestamp 1655456512
transform 0 1 527368 1 0 459077
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_72
timestamp 1655456512
transform 0 -1 534639 -1 0 446698
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_73
timestamp 1655456512
transform 0 -1 534649 -1 0 467098
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_74
timestamp 1655456512
transform -1 0 546380 0 1 475255
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_75
timestamp 1655456512
transform 0 1 550207 1 0 459206
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_76
timestamp 1655456512
transform -1 0 564689 0 -1 453558
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_77
timestamp 1655456512
transform -1 0 523434 0 -1 479906
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_78
timestamp 1655456512
transform -1 0 500984 0 1 479343
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_79
timestamp 1655456512
transform 0 -1 534617 1 0 488027
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_80
timestamp 1655456512
transform 0 -1 515264 -1 0 487819
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_81
timestamp 1655456512
transform 0 1 508791 1 0 485949
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_82
timestamp 1655456512
transform 0 -1 534607 1 0 508427
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_83
timestamp 1655456512
transform 0 -1 515301 -1 0 508020
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_84
timestamp 1655456512
transform 0 1 521229 1 0 497874
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_85
timestamp 1655456512
transform 0 1 508779 1 0 506000
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_86
timestamp 1655456512
transform 0 -1 502441 -1 0 500413
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_87
timestamp 1655456512
transform -1 0 546327 0 1 479347
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_88
timestamp 1655456512
transform 0 -1 527729 -1 0 496088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_89
timestamp 1655456512
transform 0 -1 550729 -1 0 492143
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_90
timestamp 1655456512
transform -1 0 564755 0 1 497597
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_91
timestamp 1655456512
transform 1 0 424172 0 -1 519341
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_92
timestamp 1655456512
transform 1 0 444185 0 -1 519400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_93
timestamp 1655456512
transform 1 0 464368 0 -1 519483
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_94
timestamp 1655456512
transform 1 0 484700 0 -1 519444
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_95
timestamp 1655456512
transform 1 0 504174 0 -1 519451
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_96
timestamp 1655456512
transform 0 1 505396 1 0 539457
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_97
timestamp 1655456512
transform 0 1 505286 1 0 560045
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_98
timestamp 1655456512
transform 0 -1 514025 -1 0 562750
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_99
timestamp 1655456512
transform 0 1 522348 1 0 549967
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_100
timestamp 1655456512
transform 0 -1 514005 -1 0 542308
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_101
timestamp 1655456512
transform 0 -1 514002 -1 0 522337
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_102
timestamp 1655456512
transform 0 1 522397 1 0 529190
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_103
timestamp 1655456512
transform 1 0 525233 0 -1 568134
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_104
timestamp 1655456512
transform 0 -1 531295 -1 0 553196
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_105
timestamp 1655456512
transform 0 -1 531250 -1 0 531951
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_106
timestamp 1655456512
transform 1 0 537603 0 -1 519596
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_107
timestamp 1655456512
transform 0 1 544588 1 0 532219
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_108
timestamp 1655456512
transform 0 1 544583 1 0 552445
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_109
timestamp 1655456512
transform 0 1 544573 1 0 572694
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_110
timestamp 1655456512
transform 1 0 550784 0 -1 587014
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_111
timestamp 1655456512
transform 1 0 571795 0 -1 587045
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_112
timestamp 1655456512
transform -1 0 481028 0 -1 479857
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_113
timestamp 1655456512
transform -1 0 440546 0 -1 479867
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_114
timestamp 1655456512
transform -1 0 460846 0 -1 479879
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_115
timestamp 1655456512
transform -1 0 420308 0 -1 479838
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_116
timestamp 1655456512
transform -1 0 400066 0 -1 479898
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_117
timestamp 1655456512
transform -1 0 384611 0 -1 479873
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_118
timestamp 1655456512
transform 0 1 355865 -1 0 482345
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_119
timestamp 1655456512
transform 0 1 355803 -1 0 502289
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_120
timestamp 1655456512
transform 0 1 355838 -1 0 522198
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_121
timestamp 1655456512
transform 0 1 355873 -1 0 462325
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_122
timestamp 1655456512
transform 0 1 355847 -1 0 442332
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_123
timestamp 1655456512
transform 0 1 355852 -1 0 422378
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_124
timestamp 1655456512
transform 0 1 355841 -1 0 402343
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_125
timestamp 1655456512
transform 0 1 355821 -1 0 382279
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_126
timestamp 1655456512
transform 0 1 355878 -1 0 362296
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_127
timestamp 1655456512
transform 0 1 355878 -1 0 342293
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_128
timestamp 1655456512
transform 0 1 355802 -1 0 322291
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_129
timestamp 1655456512
transform 0 1 355840 -1 0 302270
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_130
timestamp 1655456512
transform 1 0 370741 0 1 295771
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_131
timestamp 1655456512
transform 1 0 390750 0 1 295788
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_132
timestamp 1655456512
transform 1 0 410756 0 1 295759
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_133
timestamp 1655456512
transform 1 0 430752 0 1 295835
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_134
timestamp 1655456512
transform 1 0 450769 0 1 295802
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_135
timestamp 1655456512
transform 1 0 470771 0 1 295827
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_136
timestamp 1655456512
transform 1 0 490766 0 1 295860
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_137
timestamp 1655456512
transform 1 0 510759 0 1 295816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_138
timestamp 1655456512
transform 1 0 530744 0 1 295860
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_139
timestamp 1655456512
transform 1 0 551362 0 1 273753
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_140
timestamp 1655456512
transform 1 0 571825 0 1 273713
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_141
timestamp 1655456512
transform 0 1 549394 -1 0 293528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_142
timestamp 1655456512
transform 0 1 346829 -1 0 478405
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_143
timestamp 1655456512
transform 0 1 346843 -1 0 457151
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_144
timestamp 1655456512
transform 0 1 346815 -1 0 436543
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_145
timestamp 1655456512
transform 0 1 346759 -1 0 415909
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_146
timestamp 1655456512
transform 0 1 346787 -1 0 395231
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_147
timestamp 1655456512
transform 0 1 346773 -1 0 373949
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_148
timestamp 1655456512
transform 0 1 346773 -1 0 353099
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_149
timestamp 1655456512
transform 0 1 346857 -1 0 332503
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_150
timestamp 1655456512
transform 0 1 346829 -1 0 310635
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_151
timestamp 1655456512
transform 0 1 346787 -1 0 288977
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_152
timestamp 1655456512
transform 0 1 346745 -1 0 264197
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_153
timestamp 1655456512
transform 0 1 346829 -1 0 242823
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_154
timestamp 1655456512
transform 0 1 346857 -1 0 222947
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_155
timestamp 1655456512
transform 0 1 346801 -1 0 201119
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_156
timestamp 1655456512
transform 0 1 346815 -1 0 180085
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_157
timestamp 1655456512
transform 0 1 346773 -1 0 158697
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_158
timestamp 1655456512
transform 0 1 346717 -1 0 137351
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_159
timestamp 1655456512
transform 0 1 346773 -1 0 116217
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_160
timestamp 1655456512
transform 0 1 346801 -1 0 95607
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_161
timestamp 1655456512
transform 0 1 346787 -1 0 74925
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_162
timestamp 1655456512
transform 0 1 346857 -1 0 51345
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_163
timestamp 1655456512
transform -1 0 324635 0 -1 48997
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_164
timestamp 1655456512
transform -1 0 303087 0 -1 48961
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_165
timestamp 1655456512
transform -1 0 281897 0 -1 49167
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_166
timestamp 1655456512
transform -1 0 261085 0 -1 49065
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_167
timestamp 1655456512
transform -1 0 240583 0 -1 49005
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_168
timestamp 1655456512
transform -1 0 219597 0 -1 49035
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_169
timestamp 1655456512
transform -1 0 197703 0 -1 49123
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_170
timestamp 1655456512
transform -1 0 176321 0 -1 49065
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_171
timestamp 1655456512
transform -1 0 155115 0 -1 49093
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_172
timestamp 1655456512
transform -1 0 133557 0 -1 49123
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_173
timestamp 1655456512
transform -1 0 112235 0 -1 49079
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_174
timestamp 1655456512
transform -1 0 91175 0 -1 49035
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_175
timestamp 1655456512
transform -1 0 69809 0 -1 49109
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_176
timestamp 1655456512
transform -1 0 48515 0 -1 49049
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_177
timestamp 1655456512
transform 0 1 34425 -1 0 43091
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_178
timestamp 1655456512
transform 0 1 34425 -1 0 20993
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_179
timestamp 1655456512
transform -1 0 28265 0 -1 3785
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_180
timestamp 1655456512
transform -1 0 7073 0 -1 3725
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655456512
transform 0 -1 251696 1 0 455276
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1655456512
transform 0 -1 251679 1 0 433495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1655456512
transform -1 0 279063 0 1 420349
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1655456512
transform -1 0 258929 0 1 420316
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1655456512
transform -1 0 320068 0 1 420307
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1655456512
transform -1 0 299740 0 1 420355
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1655456512
transform 0 -1 336827 1 0 416486
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1655456512
transform 1 0 353582 0 1 420316
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1655456512
transform 1 0 373925 0 1 420386
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1655456512
transform 0 -1 388177 1 0 427109
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1655456512
transform 0 -1 388148 1 0 448152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1655456512
transform 0 -1 388187 1 0 469172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1655456512
transform 0 -1 388178 1 0 490136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1655456512
transform 0 -1 336852 1 0 395833
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1655456512
transform -1 0 348063 0 1 386451
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1655456512
transform -1 0 368079 0 1 386480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1655456512
transform -1 0 387891 0 1 386470
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1655456512
transform -1 0 408150 0 1 386468
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1655456512
transform -1 0 428426 0 1 386523
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1655456512
transform -1 0 448585 0 1 386503
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1655456512
transform -1 0 468587 0 1 386498
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1655456512
transform -1 0 488705 0 1 386482
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1655456512
transform -1 0 508835 0 1 386505
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1655456512
transform -1 0 528944 0 1 386519
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1655456512
transform 0 -1 549833 -1 0 388331
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1655456512
transform 0 -1 549816 -1 0 407375
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1655456512
transform -1 0 568663 0 1 408715
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1655456512
transform 0 -1 240974 1 0 455298
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1655456512
transform 0 -1 240894 1 0 433781
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1655456512
transform -1 0 253575 0 1 425814
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1655456512
transform -1 0 273521 0 1 425879
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1655456512
transform -1 0 293802 0 1 425913
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1655456512
transform -1 0 313951 0 1 425903
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1655456512
transform 1 0 355352 0 1 425884
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1655456512
transform 1 0 335362 0 1 425888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1655456512
transform 1 0 375315 0 1 425978
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1655456512
transform 0 -1 393101 1 0 427128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1655456512
transform 0 -1 393069 1 0 448220
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1655456512
transform 0 -1 393079 1 0 469172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1655456512
transform 0 -1 393081 1 0 490150
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1655456512
transform 0 -1 324817 1 0 416561
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1655456512
transform 0 -1 324815 1 0 395771
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1655456512
transform -1 0 333694 0 1 380484
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1655456512
transform -1 0 358273 0 1 380492
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1655456512
transform -1 0 387720 0 1 380450
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1655456512
transform -1 0 408298 0 1 380481
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1655456512
transform -1 0 428272 0 1 380456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1655456512
transform -1 0 448518 0 1 380460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1655456512
transform -1 0 468502 0 1 380527
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1655456512
transform -1 0 488917 0 1 380452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1655456512
transform -1 0 508600 0 1 380524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1655456512
transform -1 0 528970 0 1 380458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1655456512
transform 0 -1 549641 1 0 378877
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1655456512
transform 0 -1 549602 1 0 363691
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1655456512
transform -1 0 568819 0 1 362332
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1655456512
transform 0 -1 383541 1 0 490055
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1655456512
transform 0 -1 373889 1 0 490057
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1655456512
transform -1 0 379668 0 -1 475772
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1655456512
transform -1 0 400158 0 -1 475805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1655456512
transform -1 0 420400 0 -1 475745
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1655456512
transform -1 0 460938 0 -1 475786
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1655456512
transform -1 0 440638 0 -1 475774
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1655456512
transform -1 0 481120 0 -1 475764
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1655456512
transform -1 0 501108 0 -1 475782
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1655456512
transform 0 1 521261 -1 0 457343
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1655456512
transform 0 -1 502473 1 0 454620
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1655456512
transform 0 1 508811 -1 0 449217
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1655456512
transform 0 1 508823 -1 0 469268
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1655456512
transform 0 -1 515296 1 0 467214
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1655456512
transform -1 0 523558 0 1 475219
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1655456512
transform 0 -1 515333 1 0 447013
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1655456512
transform 0 1 527368 1 0 458985
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1655456512
transform 0 -1 534639 -1 0 446790
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1655456512
transform 0 -1 534649 -1 0 467190
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1655456512
transform -1 0 546472 0 1 475255
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1655456512
transform 0 1 550207 1 0 459114
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1655456512
transform -1 0 564781 0 -1 453558
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1655456512
transform -1 0 523526 0 -1 479906
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1655456512
transform -1 0 501076 0 1 479343
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1655456512
transform 0 -1 534617 1 0 487935
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1655456512
transform 0 -1 515264 -1 0 487911
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1655456512
transform 0 1 508791 1 0 485857
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1655456512
transform 0 -1 534607 1 0 508335
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1655456512
transform 0 -1 515301 -1 0 508112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1655456512
transform 0 1 521229 1 0 497782
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1655456512
transform 0 1 508779 1 0 505908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1655456512
transform 0 -1 502441 -1 0 500505
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1655456512
transform -1 0 546419 0 1 479347
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1655456512
transform 0 -1 527729 -1 0 496180
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1655456512
transform 0 -1 550729 -1 0 492235
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1655456512
transform -1 0 564847 0 1 497597
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1655456512
transform 1 0 424080 0 -1 519341
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1655456512
transform 1 0 444093 0 -1 519400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1655456512
transform 1 0 464276 0 -1 519483
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1655456512
transform 1 0 484608 0 -1 519444
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1655456512
transform 1 0 504082 0 -1 519451
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1655456512
transform 0 1 505396 1 0 539365
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1655456512
transform 0 1 505286 1 0 559953
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1655456512
transform 0 -1 514025 -1 0 562842
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1655456512
transform 0 1 522348 1 0 549875
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1655456512
transform 0 -1 514005 -1 0 542400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1655456512
transform 0 -1 514002 -1 0 522429
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1655456512
transform 0 1 522397 1 0 529098
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1655456512
transform 1 0 525141 0 -1 568134
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1655456512
transform 0 -1 531295 -1 0 553288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1655456512
transform 0 -1 531250 -1 0 532043
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1655456512
transform 1 0 537511 0 -1 519596
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1655456512
transform 0 1 544588 1 0 532127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1655456512
transform 0 1 544583 1 0 552353
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1655456512
transform 0 1 544573 1 0 572602
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1655456512
transform 1 0 550692 0 -1 587014
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1655456512
transform 1 0 571703 0 -1 587045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1655456512
transform -1 0 481120 0 -1 479857
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1655456512
transform -1 0 440638 0 -1 479867
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1655456512
transform -1 0 460938 0 -1 479879
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1655456512
transform -1 0 420400 0 -1 479838
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1655456512
transform -1 0 400158 0 -1 479898
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1655456512
transform -1 0 384703 0 -1 479873
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1655456512
transform 0 1 355865 -1 0 482437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1655456512
transform 0 1 355803 -1 0 502381
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1655456512
transform 0 1 355838 -1 0 522290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1655456512
transform 0 1 355873 -1 0 462417
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1655456512
transform 0 1 355847 -1 0 442424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1655456512
transform 0 1 355852 -1 0 422470
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1655456512
transform 0 1 355841 -1 0 402435
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1655456512
transform 0 1 355821 -1 0 382371
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1655456512
transform 0 1 355878 -1 0 362388
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1655456512
transform 0 1 355878 -1 0 342385
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1655456512
transform 0 1 355802 -1 0 322383
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1655456512
transform 0 1 355840 -1 0 302362
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1655456512
transform 1 0 370649 0 1 295771
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1655456512
transform 1 0 390658 0 1 295788
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1655456512
transform 1 0 410664 0 1 295759
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1655456512
transform 1 0 430660 0 1 295835
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1655456512
transform 1 0 450677 0 1 295802
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1655456512
transform 1 0 470679 0 1 295827
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1655456512
transform 1 0 490674 0 1 295860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1655456512
transform 1 0 510667 0 1 295816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1655456512
transform 1 0 530652 0 1 295860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1655456512
transform 1 0 551270 0 1 273753
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1655456512
transform 1 0 571733 0 1 273713
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1655456512
transform 0 1 549394 -1 0 293620
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1655456512
transform 0 1 346829 -1 0 478497
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1655456512
transform 0 1 346843 -1 0 457243
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1655456512
transform 0 1 346815 -1 0 436635
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1655456512
transform 0 1 346759 -1 0 416001
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1655456512
transform 0 1 346787 -1 0 395323
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1655456512
transform 0 1 346773 -1 0 374041
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1655456512
transform 0 1 346773 -1 0 353191
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1655456512
transform 0 1 346857 -1 0 332595
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1655456512
transform 0 1 346829 -1 0 310727
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1655456512
transform 0 1 346787 -1 0 289069
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1655456512
transform 0 1 346745 -1 0 264289
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1655456512
transform 0 1 346829 -1 0 242915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1655456512
transform 0 1 346857 -1 0 223039
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1655456512
transform 0 1 346801 -1 0 201211
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1655456512
transform 0 1 346815 -1 0 180177
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1655456512
transform 0 1 346773 -1 0 158789
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1655456512
transform 0 1 346717 -1 0 137443
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1655456512
transform 0 1 346773 -1 0 116309
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1655456512
transform 0 1 346801 -1 0 95699
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1655456512
transform 0 1 346787 -1 0 75017
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1655456512
transform 0 1 346857 -1 0 51437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1655456512
transform -1 0 324727 0 -1 48997
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1655456512
transform -1 0 303179 0 -1 48961
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1655456512
transform -1 0 281989 0 -1 49167
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1655456512
transform -1 0 261177 0 -1 49065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1655456512
transform -1 0 240675 0 -1 49005
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1655456512
transform -1 0 219689 0 -1 49035
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1655456512
transform -1 0 197795 0 -1 49123
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1655456512
transform -1 0 176413 0 -1 49065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1655456512
transform -1 0 155207 0 -1 49093
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1655456512
transform -1 0 133649 0 -1 49123
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1655456512
transform -1 0 112327 0 -1 49079
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1655456512
transform -1 0 91267 0 -1 49035
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1655456512
transform -1 0 69901 0 -1 49109
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1655456512
transform -1 0 48607 0 -1 49049
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1655456512
transform 0 1 34425 -1 0 43183
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1655456512
transform 0 1 34425 -1 0 21085
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1655456512
transform -1 0 28357 0 -1 3785
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1655456512
transform -1 0 7165 0 -1 3725
box -38 -48 130 592
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
<< end >>
