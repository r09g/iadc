magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< pwell >>
rect -116 3990 7122 4864
rect 13289 3990 22069 5305
rect -116 1 22069 3990
<< locali >>
rect 6609 19960 6865 20216
rect -61 8576 5805 8582
rect -61 8332 5555 8576
rect 5799 8332 5805 8576
rect -61 8326 5805 8332
rect 23491 8569 23747 8575
rect -61 379 195 8326
rect 23491 8325 23497 8569
rect 23741 8325 23747 8569
rect 7193 6918 7449 7996
rect 11584 6968 11840 7996
rect 16315 6980 16571 7996
rect 21581 6945 21837 8022
rect -60 18 195 379
rect 23491 280 23747 8325
rect 21894 24 23747 280
<< viali >>
rect 8715 8761 8971 9017
rect 19650 8749 19906 9005
rect 5555 8332 5799 8576
rect 23497 8325 23741 8569
<< metal1 >>
rect 6805 13640 6815 14159
rect 6910 13640 6920 14159
rect 6338 11097 6348 11637
rect 6458 11097 6468 11637
rect 21875 11225 21885 11732
rect 21996 11539 22006 11732
rect 21997 11429 22006 11539
rect 21996 11225 22006 11429
rect 5728 9289 5738 9829
rect 5848 9289 5858 9829
rect 22389 9295 22399 9835
rect 22509 9295 22519 9835
rect 8703 9017 8983 9023
rect 8703 8761 8715 9017
rect 8971 8761 8983 9017
rect 8703 8755 8983 8761
rect 19638 9005 19918 9011
rect 8715 8582 8971 8755
rect 19638 8749 19650 9005
rect 19906 8749 19918 9005
rect 19638 8743 19918 8749
rect 5543 8576 8971 8582
rect 5543 8332 5555 8576
rect 5799 8332 8971 8576
rect 5543 8326 8971 8332
rect 19650 8575 19906 8743
rect 19650 8569 23753 8575
rect 19650 8325 23497 8569
rect 23741 8325 23753 8569
rect 19650 8319 23753 8325
rect 2937 4263 2993 5118
rect 4720 4263 4776 5118
rect 647 3692 657 3802
rect 767 3692 777 3802
rect 21251 1092 22312 1220
<< via1 >>
rect 6815 13640 6910 14159
rect 6348 11097 6458 11637
rect 21885 11539 21996 11732
rect 21885 11429 21997 11539
rect 21885 11225 21996 11429
rect 5738 9289 5848 9829
rect 22399 9295 22509 9835
rect 657 3692 767 3802
<< metal2 >>
rect 6815 14159 6910 14169
rect 613 13772 6815 13978
rect 613 3802 819 13772
rect 6910 13772 6912 13978
rect 6815 13630 6910 13640
rect 21885 11732 21996 11742
rect 6331 11637 6537 11649
rect 6331 11443 6348 11637
rect 6342 11105 6348 11443
rect 6334 11097 6348 11105
rect 6458 11534 6537 11637
rect 23475 11592 23656 11602
rect 6458 11097 6540 11534
rect 21881 11429 21885 11539
rect 21997 11429 23475 11539
rect 23475 11363 23656 11373
rect 21885 11215 21996 11225
rect 6334 10899 6540 11097
rect 5666 9829 5872 9846
rect 5666 9738 5738 9829
rect 5664 9289 5738 9738
rect 5848 9640 5872 9829
rect 5848 9289 5870 9640
rect 5664 4245 5870 9289
rect 5664 4000 5870 4039
rect 613 3692 657 3802
rect 767 3692 819 3802
rect 613 3682 819 3692
rect 6342 3859 6540 10899
rect 22387 9835 22593 9877
rect 22387 9295 22399 9835
rect 22509 9295 22593 9835
rect 8757 4244 8881 4254
rect 8757 4029 8881 4039
rect 6342 3849 6541 3859
rect 6342 3675 6343 3849
rect 6343 3665 6541 3675
rect 11452 3848 11558 3855
rect 11452 3845 11561 3848
rect 11558 3839 11561 3845
rect 11558 3730 11561 3739
rect 11452 3632 11558 3642
rect 17433 3017 17535 3018
rect 17432 3008 17542 3017
rect 17432 3007 17433 3008
rect 17535 3007 17542 3008
rect 17432 2887 17433 2897
rect 17535 2887 17542 2897
rect 22387 3004 22593 9295
rect 17433 2793 17535 2803
rect 22387 2788 22593 2798
<< via2 >>
rect 23475 11373 23656 11592
rect 5664 4039 5870 4245
rect 8757 4039 8881 4244
rect 6343 3675 6541 3849
rect 11452 3839 11558 3845
rect 11452 3739 11561 3839
rect 11452 3642 11558 3739
rect 17433 3007 17535 3008
rect 17432 2897 17542 3007
rect 17433 2803 17535 2897
rect 22387 2798 22593 3004
<< metal3 >>
rect 23462 11592 23668 11618
rect 23462 11373 23475 11592
rect 23656 11373 23668 11592
rect 5654 4245 5880 4250
rect 8747 4245 8891 4249
rect 5654 4039 5664 4245
rect 5870 4244 8891 4245
rect 5870 4039 8757 4244
rect 8881 4039 8891 4244
rect 5654 4034 5880 4039
rect 8747 4034 8891 4039
rect 6333 3849 6551 3854
rect 6333 3675 6343 3849
rect 6541 3845 6551 3849
rect 11442 3845 11568 3850
rect 6541 3675 11452 3845
rect 11558 3839 11579 3845
rect 11561 3739 11579 3839
rect 23462 3833 23668 11373
rect 6333 3670 11452 3675
rect 6342 3642 11452 3670
rect 11558 3642 11579 3739
rect 6342 3640 11579 3642
rect 6434 3639 11579 3640
rect 11442 3637 11568 3639
rect 13209 3627 23668 3833
rect 13209 2681 13415 3627
rect 17423 3012 17545 3013
rect 17422 3008 17552 3012
rect 17422 3007 17433 3008
rect 17535 3007 17552 3008
rect 17422 2897 17432 3007
rect 17542 3006 17552 3007
rect 22377 3006 22603 3009
rect 17542 3004 22603 3006
rect 17542 2897 22387 3004
rect 17422 2892 17433 2897
rect 17423 2803 17433 2892
rect 17535 2803 22387 2897
rect 17423 2800 22387 2803
rect 17423 2798 17545 2800
rect 22377 2798 22387 2800
rect 22593 2798 22603 3004
rect 22377 2793 22603 2798
rect -170 2475 13415 2681
<< metal4 >>
rect 7353 20556 21191 20620
rect 7272 20156 7581 20220
rect 7272 19756 7872 19820
rect 7272 19356 8182 19420
use ota_v2_without_cmfb  ota_v2_without_cmfb_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/ota_v2
timestamp 1655484843
transform -1 0 21026 0 1 335
box -1054 -334 21142 6713
use sc_cmfb  sc_cmfb_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/sc_cmfb
timestamp 1655484843
transform 1 0 11071 0 1 10659
box -5376 -2919 11546 9969
<< labels >>
flabel metal1 2965 4960 2965 4960 1 FreeSans 800 0 0 0 in
port 2 n
flabel metal1 4751 4964 4751 4964 1 FreeSans 800 0 0 0 ip
port 1 n
flabel metal4 7524 20588 7524 20588 1 FreeSans 800 0 0 0 p2_b
port 6 n
flabel metal4 7520 20183 7520 20183 1 FreeSans 800 0 0 0 p2
port 5 n
flabel metal4 7522 19788 7522 19788 1 FreeSans 800 0 0 0 p1_b
port 4 n
flabel metal4 7522 19380 7522 19380 1 FreeSans 800 0 0 0 p1
port 3 n
flabel metal2 5790 8141 5790 8141 1 FreeSans 800 0 0 0 op
port 7 n
flabel metal2 6403 8150 6403 8150 1 FreeSans 800 0 0 0 on
port 8 n
flabel metal1 22248 1153 22248 1153 1 FreeSans 800 0 0 0 i_bias
port 9 n
flabel metal3 -153 2588 -153 2588 1 FreeSans 800 0 0 0 cm
port 10 n
flabel locali 6730 20089 6730 20089 1 FreeSans 800 0 0 0 VDD
port 11 n power bidirectional
flabel locali 11 93 11 93 1 FreeSans 800 0 0 0 VSS
port 12 n power bidirectional
<< end >>
