* analog_top

.include "../sky130_fd_sc_hd.spice"

.subckt analog_top ip in rst_n i_bias_1 i_bias_2 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1 debug op
+ a_probe_0 a_probe_1 a_probe_2 a_probe_3 clk d_probe_0 d_probe_1 d_probe_2 d_probe_3 d_clk_grp_1_ctrl_0
+ d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VDD VSS
*.ipin ip
*.ipin in
*.ipin rst_n
*.ipin i_bias_1
*.ipin i_bias_2
*.ipin a_mod_grp_ctrl_0
*.ipin a_mod_grp_ctrl_1
*.ipin debug
*.opin op
*.opin a_probe_0
*.opin a_probe_1
*.opin a_probe_2
*.opin a_probe_3
*.ipin clk
*.opin d_probe_0
*.opin d_probe_1
*.opin d_probe_2
*.opin d_probe_3
*.ipin d_clk_grp_1_ctrl_0
*.ipin d_clk_grp_1_ctrl_1
*.ipin d_clk_grp_2_ctrl_0
*.ipin d_clk_grp_2_ctrl_1
x1 ip in A A_b Ad Ad_b B B_b Bd Bd_b p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b rst_n rst_n_b i_bias_1
+ i_bias_2 op bias_a bias_b bias_c bias_d cm1 cmc op2 op1 on1 on2 VDD VSS modulator_w_test
x2 a_mod_grp_ctrl_1 a_mod_grp_ctrl_0 debug cm1 bias_b cmc net1 a_probe_2 VDD VSS a_mux4_en
x3 a_mod_grp_ctrl_1 a_mod_grp_ctrl_0 debug bias_a bias_c bias_d net2 a_probe_3 VDD VSS a_mux4_en
x4 a_mod_grp_ctrl_0 debug op1 on1 a_probe_0 VDD VSS a_mux2_en
x5 a_mod_grp_ctrl_0 debug op2 on2 a_probe_1 VDD VSS a_mux2_en
x8 a_probe_0 VDD VSS esd_cell
x9 a_probe_1 VDD VSS esd_cell
x10 a_probe_2 VDD VSS esd_cell
x11 a_probe_3 VDD VSS esd_cell
x12 i_bias_1 VDD VSS esd_cell
x13 i_bias_2 VDD VSS esd_cell
x14 ip VDD VSS esd_cell
x15 in VDD VSS esd_cell
x6 A A_b Ad Ad_b Bd_b Bd B_b B p2 p2_b p2d clk p2d_b p1d_b p1d p1_b p1 VDD VSS clock_v2
x16 p1 A p1_b A_b d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 VSS VSS VDD VDD net3 sky130_fd_sc_hd__mux4_1
x17 p2 B p2_b B_b d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 VSS VSS VDD VDD net4 sky130_fd_sc_hd__mux4_1
x18 p1d Ad p1d_b Ad_b d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VSS VDD VDD net5
+ sky130_fd_sc_hd__mux4_1
x19 p2d Bd p2d_b Bd_b d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VSS VDD VDD net6
+ sky130_fd_sc_hd__mux4_1
x20 net3 VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkinv_4
x21 net7 VSS VSS VDD VDD d_probe_0 sky130_fd_sc_hd__clkinv_16
x22 net4 VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkinv_4
x23 net8 VSS VSS VDD VDD d_probe_1 sky130_fd_sc_hd__clkinv_16
x24 net5 VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkinv_4
x25 net9 VSS VSS VDD VDD d_probe_2 sky130_fd_sc_hd__clkinv_16
x26 net6 VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkinv_4
x27 net10 VSS VSS VDD VDD d_probe_3 sky130_fd_sc_hd__clkinv_16
x7 rst_n VSS VSS VDD VDD rst_n_b sky130_fd_sc_hd__clkinv_4
xDC1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
xDC2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
xDC3 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
xDC4 VSS VSS VDD VDD sky130_fd_sc_hd__decap_12
.ends

* expanding   symbol:  modulator_w_test.sym # of pins=33
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/modulator_w_test.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/modulator_w_test.sch
.subckt modulator_w_test  ip in A A_b Ad Ad_b B B_b Bd Bd_b p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b
+ rst_n rst_n_b i_bias_1 i_bias_2 op bias_a bias_b bias_c bias_d cm1 cmc op2 op1 on1 on2  VDD  VSS
*.ipin ip
*.ipin in
*.ipin A
*.ipin A_b
*.ipin Ad
*.ipin Ad_b
*.ipin B
*.ipin B_b
*.ipin Bd
*.ipin Bd_b
*.ipin p1
*.ipin p1_b
*.ipin p1d
*.ipin p1d_b
*.ipin p2
*.ipin p2_b
*.ipin p2d
*.ipin p2d_b
*.ipin rst_n
*.ipin rst_n_b
*.ipin i_bias_1
*.ipin i_bias_2
*.opin op
*.opin bias_a
*.opin bias_b
*.opin bias_c
*.opin bias_d
*.opin cm1
*.opin cmc
*.opin op1
*.opin on1
*.opin op2
*.opin on2
x4 c1r in1 p2 p2_b VDD VSS transmission_gate
x5 net1 ip1 p2 p2_b VDD VSS transmission_gate
x2 c1r cm1 p1 p1_b VDD VSS transmission_gate
x3 net1 cm1 p1 p1_b VDD VSS transmission_gate
x10 ip c1l p1d p1d_b VDD VSS transmission_gate
x11 dac_n net2 p2d p2d_b VDD VSS transmission_gate
x12 VDD VSS op dac_p on VDD VSS 1b_dac
x13 dac_p c1l p2d p2d_b VDD VSS transmission_gate
x14 in net2 p1d p1d_b VDD VSS transmission_gate
x19 on1 op1 rst_n_b rst_n VDD VSS transmission_gate
x20 cm1 in1 rst_n_b rst_n VDD VSS transmission_gate
x21 cm1 ip1 rst_n_b rst_n VDD VSS transmission_gate
x22 op1 c3l p1d p1d_b VDD VSS transmission_gate
x23 on1 net3 p1d p1d_b VDD VSS transmission_gate
x24 net3 c3l p2d p2d_b VDD VSS transmission_gate
x25 c3r cm2 p1 p1_b VDD VSS transmission_gate
x26 net4 cm2 p1 p1_b VDD VSS transmission_gate
x27 ip c4l p1d p1d_b VDD VSS transmission_gate
x28 dac_p c4l p2d p2d_b VDD VSS transmission_gate
x29 c3r in2 p2 p2_b VDD VSS transmission_gate
x30 net4 ip2 p2 p2_b VDD VSS transmission_gate
x32 cm2 in2 rst_n_b rst_n VDD VSS transmission_gate
x33 cm2 ip2 rst_n_b rst_n VDD VSS transmission_gate
x34 on2 op2 rst_n_b rst_n VDD VSS transmission_gate
x36 VSS VDD op dac_n on VDD VSS 1b_dac
x37 in net5 p1d p1d_b VDD VSS transmission_gate
x38 dac_n net5 p2d p2d_b VDD VSS transmission_gate
XC11 c1l c1r sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=2 m=2
XC1 net2 net1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=2 m=2
XC2 op1 in1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=10 m=10
XC3 on1 ip1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=10 m=10
XC4 c3r c4l sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=1 m=1
XC5 c3r c3l sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=2 m=2
XC6 net4 net3 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=2 m=2
XC7 net4 net5 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=1 m=1
XC8 op2 in2 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=14 m=14
XC9 on2 ip2 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=14 m=14
XC10 op2 VSS sky130_fd_pr__cap_mim_m3_1 W=11.6 L=11.6 MF=1 m=1
XC12 on2 VSS sky130_fd_pr__cap_mim_m3_1 W=11.6 L=11.6 MF=1 m=1
x6 in1 in1_c A A_b VDD VSS transmission_gate
x8 ip1 in1_c B B_b VDD VSS transmission_gate
x15 op1_c op1 Ad Ad_b VDD VSS transmission_gate
x16 on1_c on1 Ad Ad_b VDD VSS transmission_gate
x17 op1_c on1 Bd Bd_b VDD VSS transmission_gate
x18 on1_c op1 Bd Bd_b VDD VSS transmission_gate
x7 ip1 ip1_c A A_b VDD VSS transmission_gate
x9 in1 ip1_c B B_b VDD VSS transmission_gate
XC13 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=24 m=24
XC14 __UNCONNECTED_PIN__2 __UNCONNECTED_PIN__3 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=38 m=38
x35 op2 on2 op p1_b on VDD VSS comparator
XM2 VSS on VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM3 VDD on VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
x1 i_bias_1 ip1_c in1_c p1 p1_b p2 p2_b op1_c on1_c cm1 bias_a bias_b bias_c bias_d cmc VDD VSS
+ ota_w_test
x31 i_bias_2 ip2 in2 p1 p1_b p2 p2_b op2 on2 cm2 VDD VSS ota
.ends


* expanding   symbol:  a_mux4_en.sym # of pins=8
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux4_en.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux4_en.sch
.subckt a_mux4_en  s0 s1 en in0 in1 in2 in3 out  VDD  VSS
*.ipin en
*.ipin s1
*.ipin s0
*.ipin in0
*.ipin in1
*.ipin in2
*.ipin in3
*.opin out
x1 net4 out net5 en3_b VDD VSS switch_5t
x2 net3 out net6 en2_b VDD VSS switch_5t
x3 net2 out net7 en1_b VDD VSS switch_5t
x4 net1 out net8 en0_b VDD VSS switch_5t
x5 en3_b VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x6 en2_b VSS VSS VDD VDD net6 sky130_fd_sc_hd__inv_1
x7 en1_b VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
x8 en0_b VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_1
x13 s0 VSS VSS VDD VDD s0_b sky130_fd_sc_hd__inv_1
x14 s1 VSS VSS VDD VDD s1_b sky130_fd_sc_hd__inv_1
x9 s1_b s0_b VSS VSS VDD VDD en0_b sky130_fd_sc_hd__nand2_1
x10 s1 s0_b VSS VSS VDD VDD en1_b sky130_fd_sc_hd__nand2_1
x11 s0 s1_b VSS VSS VDD VDD en2_b sky130_fd_sc_hd__nand2_1
x12 s0 s1 VSS VSS VDD VDD en3_b sky130_fd_sc_hd__nand2_1
x15 in0 net1 en en_b VDD VSS transmission_gate
x16 in1 net2 en en_b VDD VSS transmission_gate
x17 in2 net3 en en_b VDD VSS transmission_gate
x18 in3 net4 en en_b VDD VSS transmission_gate
x19 en VSS VSS VDD VDD en_b sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  a_mux2_en.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux2_en.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux2_en.sch
.subckt a_mux2_en  s0 en in0 in1 out  VDD  VSS
*.ipin en
*.ipin s0
*.ipin in0
*.ipin in1
*.opin out
x3 net2 out s0 s0_b VDD VSS switch_5t
x4 net1 out s0_b s0 VDD VSS switch_5t
x15 in0 net1 en en_b VDD VSS transmission_gate
x16 in1 net2 en en_b VDD VSS transmission_gate
x19 en VSS VSS VDD VDD en_b sky130_fd_sc_hd__inv_1
x1 s0 VSS VSS VDD VDD s0_b sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  esd_cell.sym # of pins=1
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/esd_cell.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/esd_cell.sch
.subckt esd_cell  esd  VDD  VSS
*.iopin esd
XM1 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM2 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
.ends


* expanding   symbol:  clock_v2.sym # of pins=17
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/clock_v2.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/clock_v2.sch
.subckt clock_v2  A A_b Ad Ad_b Bd_b Bd B_b B p2 p2_b p2d clk p2d_b p1d_b p1d p1_b p1  VDD  VSS
*.ipin clk
*.opin p2d_b
*.opin p2d
*.opin p2_b
*.opin p2
*.opin p1d_b
*.opin p1d
*.opin p1_b
*.opin p1
*.opin Ad_b
*.opin Ad
*.opin A_b
*.opin A
*.opin Bd_b
*.opin Bd
*.opin B_b
*.opin B
xDC1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
xDC2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
xDC3 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
xDC4 VSS VSS VDD VDD sky130_fd_sc_hd__decap_12
x2 latch_out clk VSS VSS VDD VDD net1 sky130_fd_sc_hd__nand2_1
x3 net3 net6 VSS VSS VDD VDD net4 sky130_fd_sc_hd__nand2_1
x4 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__clkinv_4
x6 net2 VSS VSS VDD VDD net34 sky130_fd_sc_hd__clkinv_1
x9 net4 VSS VSS VDD VDD net5 sky130_fd_sc_hd__clkinv_4
x11 net5 VSS VSS VDD VDD net35 sky130_fd_sc_hd__clkinv_1
x1 clk VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkinv_1
x20 net36 VSS VSS VDD VDD latch_in sky130_fd_sc_hd__clkdlybuf4s50_1
x21 net37 VSS VSS VDD VDD net6 sky130_fd_sc_hd__clkdlybuf4s50_1
x22 net34 VSS VSS VDD VDD net38 sky130_fd_sc_hd__clkdlybuf4s50_1
x25 net35 VSS VSS VDD VDD net39 sky130_fd_sc_hd__clkdlybuf4s50_1
x7 net40 VSS VSS VDD VDD net36 sky130_fd_sc_hd__clkdlybuf4s50_1
x12 net41 VSS VSS VDD VDD net37 sky130_fd_sc_hd__clkdlybuf4s50_1
x14 net38 VSS VSS VDD VDD net42 sky130_fd_sc_hd__clkdlybuf4s50_1
x15 net39 VSS VSS VDD VDD net43 sky130_fd_sc_hd__clkdlybuf4s50_1
x16 net44 VSS VSS VDD VDD net40 sky130_fd_sc_hd__clkdlybuf4s50_1
x17 net45 VSS VSS VDD VDD net41 sky130_fd_sc_hd__clkdlybuf4s50_1
x18 net42 VSS VSS VDD VDD net46 sky130_fd_sc_hd__clkdlybuf4s50_1
x19 net43 VSS VSS VDD VDD net47 sky130_fd_sc_hd__clkdlybuf4s50_1
x23 net48 VSS VSS VDD VDD net44 sky130_fd_sc_hd__clkdlybuf4s50_1
x24 net49 VSS VSS VDD VDD net45 sky130_fd_sc_hd__clkdlybuf4s50_1
x26 net46 VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkdlybuf4s50_1
x27 net47 VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkdlybuf4s50_1
x28 net50 VSS VSS VDD VDD net48 sky130_fd_sc_hd__clkdlybuf4s50_1
x29 net51 VSS VSS VDD VDD net49 sky130_fd_sc_hd__clkdlybuf4s50_1
x32 net52 VSS VSS VDD VDD net50 sky130_fd_sc_hd__clkdlybuf4s50_1
x33 net53 VSS VSS VDD VDD net51 sky130_fd_sc_hd__clkdlybuf4s50_1
x36 net54 VSS VSS VDD VDD net52 sky130_fd_sc_hd__clkdlybuf4s50_1
x37 net55 VSS VSS VDD VDD net53 sky130_fd_sc_hd__clkdlybuf4s50_1
x40 net56 VSS VSS VDD VDD net54 sky130_fd_sc_hd__clkdlybuf4s50_1
x41 net57 VSS VSS VDD VDD net55 sky130_fd_sc_hd__clkdlybuf4s50_1
x44 net58 VSS VSS VDD VDD net56 sky130_fd_sc_hd__clkdlybuf4s50_1
x45 net59 VSS VSS VDD VDD net57 sky130_fd_sc_hd__clkdlybuf4s50_1
x48 net60 VSS VSS VDD VDD net58 sky130_fd_sc_hd__clkdlybuf4s50_1
x49 net61 VSS VSS VDD VDD net59 sky130_fd_sc_hd__clkdlybuf4s50_1
x52 net62 VSS VSS VDD VDD net60 sky130_fd_sc_hd__clkdlybuf4s50_1
x53 net63 VSS VSS VDD VDD net61 sky130_fd_sc_hd__clkdlybuf4s50_1
x56 net64 VSS VSS VDD VDD net62 sky130_fd_sc_hd__clkdlybuf4s50_1
x57 net65 VSS VSS VDD VDD net63 sky130_fd_sc_hd__clkdlybuf4s50_1
x60 net66 VSS VSS VDD VDD net64 sky130_fd_sc_hd__clkdlybuf4s50_1
x61 net67 VSS VSS VDD VDD net65 sky130_fd_sc_hd__clkdlybuf4s50_1
x64 net68 VSS VSS VDD VDD net66 sky130_fd_sc_hd__clkdlybuf4s50_1
x65 net69 VSS VSS VDD VDD net67 sky130_fd_sc_hd__clkdlybuf4s50_1
x68 net70 VSS VSS VDD VDD net68 sky130_fd_sc_hd__clkdlybuf4s50_1
x69 net71 VSS VSS VDD VDD net69 sky130_fd_sc_hd__clkdlybuf4s50_1
x72 net72 VSS VSS VDD VDD net70 sky130_fd_sc_hd__clkdlybuf4s50_1
x73 net73 VSS VSS VDD VDD net71 sky130_fd_sc_hd__clkdlybuf4s50_1
x76 net74 VSS VSS VDD VDD net72 sky130_fd_sc_hd__clkdlybuf4s50_1
x77 net75 VSS VSS VDD VDD net73 sky130_fd_sc_hd__clkdlybuf4s50_1
x80 net76 VSS VSS VDD VDD net74 sky130_fd_sc_hd__clkdlybuf4s50_1
x81 net77 VSS VSS VDD VDD net75 sky130_fd_sc_hd__clkdlybuf4s50_1
x84 net78 VSS VSS VDD VDD net79 sky130_fd_sc_hd__clkdlybuf4s50_1
x85 net80 VSS VSS VDD VDD net81 sky130_fd_sc_hd__clkdlybuf4s50_1
x86 net82 VSS VSS VDD VDD net78 sky130_fd_sc_hd__clkdlybuf4s50_1
x87 net83 VSS VSS VDD VDD net80 sky130_fd_sc_hd__clkdlybuf4s50_1
x88 net29 VSS VSS VDD VDD net82 sky130_fd_sc_hd__clkdlybuf4s50_1
x89 net28 VSS VSS VDD VDD net83 sky130_fd_sc_hd__clkdlybuf4s50_1
x30 clk_div net17 VSS VSS VDD VDD net9 sky130_fd_sc_hd__nand2_1
x31 net16 net12 VSS VSS VDD VDD net13 sky130_fd_sc_hd__nand2_1
x34 net9 VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkinv_4
x35 net10 VSS VSS VDD VDD net84 sky130_fd_sc_hd__clkinv_1
x38 net13 VSS VSS VDD VDD net14 sky130_fd_sc_hd__clkinv_4
x39 net14 VSS VSS VDD VDD net85 sky130_fd_sc_hd__clkinv_1
x42 clk_div VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkinv_1
x43 net86 VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkdlybuf4s50_1
x46 net87 VSS VSS VDD VDD net16 sky130_fd_sc_hd__clkdlybuf4s50_1
x47 net84 VSS VSS VDD VDD net88 sky130_fd_sc_hd__clkdlybuf4s50_1
x50 net85 VSS VSS VDD VDD net89 sky130_fd_sc_hd__clkdlybuf4s50_1
x51 net90 VSS VSS VDD VDD net86 sky130_fd_sc_hd__clkdlybuf4s50_1
x54 net91 VSS VSS VDD VDD net87 sky130_fd_sc_hd__clkdlybuf4s50_1
x55 net88 VSS VSS VDD VDD net92 sky130_fd_sc_hd__clkdlybuf4s50_1
x58 net89 VSS VSS VDD VDD net93 sky130_fd_sc_hd__clkdlybuf4s50_1
x59 net94 VSS VSS VDD VDD net90 sky130_fd_sc_hd__clkdlybuf4s50_1
x62 net95 VSS VSS VDD VDD net91 sky130_fd_sc_hd__clkdlybuf4s50_1
x63 net92 VSS VSS VDD VDD net96 sky130_fd_sc_hd__clkdlybuf4s50_1
x66 net93 VSS VSS VDD VDD net97 sky130_fd_sc_hd__clkdlybuf4s50_1
x67 net98 VSS VSS VDD VDD net94 sky130_fd_sc_hd__clkdlybuf4s50_1
x70 net99 VSS VSS VDD VDD net95 sky130_fd_sc_hd__clkdlybuf4s50_1
x71 net96 VSS VSS VDD VDD net18 sky130_fd_sc_hd__clkdlybuf4s50_1
x74 net97 VSS VSS VDD VDD net20 sky130_fd_sc_hd__clkdlybuf4s50_1
x75 net100 VSS VSS VDD VDD net98 sky130_fd_sc_hd__clkdlybuf4s50_1
x136 net101 VSS VSS VDD VDD net99 sky130_fd_sc_hd__clkdlybuf4s50_1
x137 net102 VSS VSS VDD VDD net100 sky130_fd_sc_hd__clkdlybuf4s50_1
x138 net103 VSS VSS VDD VDD net101 sky130_fd_sc_hd__clkdlybuf4s50_1
x139 net104 VSS VSS VDD VDD net102 sky130_fd_sc_hd__clkdlybuf4s50_1
x140 net105 VSS VSS VDD VDD net103 sky130_fd_sc_hd__clkdlybuf4s50_1
x141 net106 VSS VSS VDD VDD net104 sky130_fd_sc_hd__clkdlybuf4s50_1
x142 net107 VSS VSS VDD VDD net105 sky130_fd_sc_hd__clkdlybuf4s50_1
x143 net108 VSS VSS VDD VDD net106 sky130_fd_sc_hd__clkdlybuf4s50_1
x144 net109 VSS VSS VDD VDD net107 sky130_fd_sc_hd__clkdlybuf4s50_1
x145 net110 VSS VSS VDD VDD net108 sky130_fd_sc_hd__clkdlybuf4s50_1
x146 net111 VSS VSS VDD VDD net109 sky130_fd_sc_hd__clkdlybuf4s50_1
x147 net112 VSS VSS VDD VDD net110 sky130_fd_sc_hd__clkdlybuf4s50_1
x148 net113 VSS VSS VDD VDD net111 sky130_fd_sc_hd__clkdlybuf4s50_1
x149 net114 VSS VSS VDD VDD net112 sky130_fd_sc_hd__clkdlybuf4s50_1
x150 net115 VSS VSS VDD VDD net113 sky130_fd_sc_hd__clkdlybuf4s50_1
x151 net116 VSS VSS VDD VDD net114 sky130_fd_sc_hd__clkdlybuf4s50_1
x152 net117 VSS VSS VDD VDD net115 sky130_fd_sc_hd__clkdlybuf4s50_1
x153 net118 VSS VSS VDD VDD net116 sky130_fd_sc_hd__clkdlybuf4s50_1
x154 net119 VSS VSS VDD VDD net117 sky130_fd_sc_hd__clkdlybuf4s50_1
x155 net120 VSS VSS VDD VDD net118 sky130_fd_sc_hd__clkdlybuf4s50_1
x156 net121 VSS VSS VDD VDD net119 sky130_fd_sc_hd__clkdlybuf4s50_1
x157 net122 VSS VSS VDD VDD net120 sky130_fd_sc_hd__clkdlybuf4s50_1
x158 net123 VSS VSS VDD VDD net121 sky130_fd_sc_hd__clkdlybuf4s50_1
x195 net9 net18 VSS VSS VDD VDD net23 sky130_fd_sc_hd__nand2_4
x196 net10 VSS VSS VDD VDD net22 sky130_fd_sc_hd__clkinv_4
x197 net14 VSS VSS VDD VDD net21 sky130_fd_sc_hd__clkinv_4
x198 net13 net20 VSS VSS VDD VDD net19 sky130_fd_sc_hd__nand2_4
x223 clk net24 VSS VSS VDD VDD clk_div net24 sky130_fd_sc_hd__dfxbp_1
x224 p2 clk_div VSS VSS VDD VDD net25 net124 sky130_fd_sc_hd__dfxbp_1
x225 Ad_b Bd_b net25 VSS VSS VDD VDD net26 sky130_fd_sc_hd__mux2_1
x226 net26 latch_in VSS VSS VDD VDD net27 sky130_fd_sc_hd__nand2_1
x227 net27 VSS VSS VDD VDD latch_out sky130_fd_sc_hd__clkinv_1
x232 net22 VSS VSS VDD VDD A_b sky130_fd_sc_hd__clkbuf_16
x233 net10 VSS VSS VDD VDD A sky130_fd_sc_hd__clkbuf_16
x234 net11 VSS VSS VDD VDD Ad_b sky130_fd_sc_hd__clkbuf_16
x235 net23 VSS VSS VDD VDD Ad sky130_fd_sc_hd__clkbuf_16
x236 net19 VSS VSS VDD VDD Bd sky130_fd_sc_hd__clkbuf_16
x237 net15 VSS VSS VDD VDD Bd_b sky130_fd_sc_hd__clkbuf_16
x238 net14 VSS VSS VDD VDD B sky130_fd_sc_hd__clkbuf_16
x239 net21 VSS VSS VDD VDD B_b sky130_fd_sc_hd__clkbuf_16
x228 net23 VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkinv_4
x229 net19 VSS VSS VDD VDD net15 sky130_fd_sc_hd__clkinv_4
x5 net1 net7 VSS VSS VDD VDD net33 sky130_fd_sc_hd__nand2_4
x10 net2 VSS VSS VDD VDD net32 sky130_fd_sc_hd__clkinv_4
x116 net5 VSS VSS VDD VDD net31 sky130_fd_sc_hd__clkinv_4
x117 net4 net8 VSS VSS VDD VDD net30 sky130_fd_sc_hd__nand2_4
x230 net32 VSS VSS VDD VDD p2_b sky130_fd_sc_hd__clkbuf_16
x231 net2 VSS VSS VDD VDD p2 sky130_fd_sc_hd__clkbuf_16
x240 net28 VSS VSS VDD VDD p2d_b sky130_fd_sc_hd__clkbuf_16
x241 net33 VSS VSS VDD VDD p2d sky130_fd_sc_hd__clkbuf_16
x242 net30 VSS VSS VDD VDD p1d sky130_fd_sc_hd__clkbuf_16
x243 net29 VSS VSS VDD VDD p1d_b sky130_fd_sc_hd__clkbuf_16
x244 net5 VSS VSS VDD VDD p1 sky130_fd_sc_hd__clkbuf_16
x245 net31 VSS VSS VDD VDD p1_b sky130_fd_sc_hd__clkbuf_16
x246 net33 VSS VSS VDD VDD net28 sky130_fd_sc_hd__clkinv_4
x247 net30 VSS VSS VDD VDD net29 sky130_fd_sc_hd__clkinv_4
x8 net125 VSS VSS VDD VDD net123 sky130_fd_sc_hd__clkdlybuf4s50_1
x13 net126 VSS VSS VDD VDD net122 sky130_fd_sc_hd__clkdlybuf4s50_1
x78 net127 VSS VSS VDD VDD net125 sky130_fd_sc_hd__clkdlybuf4s50_1
x79 net128 VSS VSS VDD VDD net126 sky130_fd_sc_hd__clkdlybuf4s50_1
x82 net129 VSS VSS VDD VDD net130 sky130_fd_sc_hd__clkdlybuf4s50_1
x83 net131 VSS VSS VDD VDD net132 sky130_fd_sc_hd__clkdlybuf4s50_1
x90 net133 VSS VSS VDD VDD net129 sky130_fd_sc_hd__clkdlybuf4s50_1
x91 net134 VSS VSS VDD VDD net131 sky130_fd_sc_hd__clkdlybuf4s50_1
x92 net11 VSS VSS VDD VDD net133 sky130_fd_sc_hd__clkdlybuf4s50_1
x93 net15 VSS VSS VDD VDD net134 sky130_fd_sc_hd__clkdlybuf4s50_1
x94 net135 VSS VSS VDD VDD net128 sky130_fd_sc_hd__clkdlybuf4s50_1
x95 net136 VSS VSS VDD VDD net127 sky130_fd_sc_hd__clkdlybuf4s50_1
x96 net137 VSS VSS VDD VDD net135 sky130_fd_sc_hd__clkdlybuf4s50_1
x97 net138 VSS VSS VDD VDD net136 sky130_fd_sc_hd__clkdlybuf4s50_1
x98 net139 VSS VSS VDD VDD net137 sky130_fd_sc_hd__clkdlybuf4s50_1
x99 net140 VSS VSS VDD VDD net138 sky130_fd_sc_hd__clkdlybuf4s50_1
x100 net141 VSS VSS VDD VDD net140 sky130_fd_sc_hd__clkdlybuf4s50_1
x101 net142 VSS VSS VDD VDD net139 sky130_fd_sc_hd__clkdlybuf4s50_1
x102 net130 VSS VSS VDD VDD net141 sky130_fd_sc_hd__clkdlybuf4s50_1
x103 net132 VSS VSS VDD VDD net142 sky130_fd_sc_hd__clkdlybuf4s50_1
x104 net143 VSS VSS VDD VDD net77 sky130_fd_sc_hd__clkdlybuf4s50_1
x105 net144 VSS VSS VDD VDD net76 sky130_fd_sc_hd__clkdlybuf4s50_1
x106 net145 VSS VSS VDD VDD net143 sky130_fd_sc_hd__clkdlybuf4s50_1
x107 net146 VSS VSS VDD VDD net144 sky130_fd_sc_hd__clkdlybuf4s50_1
x108 net147 VSS VSS VDD VDD net145 sky130_fd_sc_hd__clkdlybuf4s50_1
x109 net148 VSS VSS VDD VDD net146 sky130_fd_sc_hd__clkdlybuf4s50_1
x110 net149 VSS VSS VDD VDD net148 sky130_fd_sc_hd__clkdlybuf4s50_1
x111 net150 VSS VSS VDD VDD net147 sky130_fd_sc_hd__clkdlybuf4s50_1
x112 net79 VSS VSS VDD VDD net149 sky130_fd_sc_hd__clkdlybuf4s50_1
x113 net81 VSS VSS VDD VDD net150 sky130_fd_sc_hd__clkdlybuf4s50_1
.ends


* expanding   symbol:  transmission_gate.sym # of pins=4
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/transmission_gate.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/transmission_gate.sch
.subckt transmission_gate  in out en en_b  VDD  VSS     N=1 W_N=5.3 L_N=0.15 W_P=13.7 L_P=0.15
*.iopin in
*.iopin out
*.ipin en
*.ipin en_b
XM1 out en in VSS sky130_fd_pr__nfet_01v8 L='L_N' W='W_N' nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='N' m='N' 
XM2 out en_b in VDD sky130_fd_pr__pfet_01v8 L='L_P' W='W_P' nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='N' m='N' 
.ends


* expanding   symbol:  1b_dac.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/1b_dac.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/1b_dac.sch
.subckt 1b_dac  v_hi v_lo v out v_b  VDD  VSS
*.ipin v_hi
*.ipin v_lo
*.ipin v
*.ipin v_b
*.opin out
x1 v_hi out v v_b VDD VSS transmission_gate
x2 v_lo out v_b v VDD VSS transmission_gate
.ends


* expanding   symbol:  comparator.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator.sch
.subckt comparator  ip in outp clk outn  VDD  VSS
*.ipin clk
*.ipin ip
*.ipin in
*.opin outp
*.opin outn
x2 s_b VSS VSS VDD VDD s_b_buf sky130_fd_sc_hd__buf_2
x3 r_b VSS VSS VDD VDD r_b_buf sky130_fd_sc_hd__buf_2
x4 s_b_buf r_b_buf outp outn VDD VSS rs_b_latch
x1 ip in s_b clk r_b VDD VSS comparator_core_large
.ends


* expanding   symbol:  ota_w_test.sym # of pins=15
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota_w_test.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota_w_test.sch
.subckt ota_w_test  i_bias ip in phi1 phi1_b phi2 phi2_b op on cm bias_a bias_b bias_c bias_d cmc
+  VDD  VSS
*.ipin ip
*.ipin in
*.ipin phi1
*.ipin phi1_b
*.ipin phi2
*.ipin phi2_b
*.opin op
*.opin on
*.ipin i_bias
*.opin cm
*.opin bias_a
*.opin bias_b
*.opin bias_c
*.opin bias_d
*.opin cmc
x1 bias_a bias_b bias_c bias_d cm i_bias VDD VSS folded_cascode_3_bias
x3 phi1 phi1_b op on cm bias_a cmc phi2 phi2_b VDD VSS sc_cmfb
x2 cmc ip in bias_a bias_b bias_c bias_d op on VDD VSS folded_cascode_3_core
XM43 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM45 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=23 m=23 
.ends


* expanding   symbol:  ota.sym # of pins=10
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota.sch
.subckt ota  i_bias ip in phi1 phi1_b phi2 phi2_b op on cm  VDD  VSS
*.ipin ip
*.ipin in
*.ipin phi1
*.ipin phi1_b
*.ipin phi2
*.ipin phi2_b
*.opin op
*.opin on
*.ipin i_bias
*.opin cm
x1 bias_a bias_b bias_c bias_d cm i_bias VDD VSS folded_cascode_3_bias
x3 phi1 phi1_b op on cm bias_a cmc phi2 phi2_b VDD VSS sc_cmfb
x2 cmc ip in bias_a bias_b bias_c bias_d op on VDD VSS folded_cascode_3_core
XM43 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM45 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=23 m=23 
.ends


* expanding   symbol:  switch_5t.sym # of pins=4
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/switch_5t.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/switch_5t.sch
.subckt switch_5t  in out en en_b  VDD  VSS
*.iopin in
*.iopin out
*.ipin en
*.ipin en_b
x1 in net1 en en_b VDD VSS transmission_gate
x2 net1 out en en_b VDD VSS transmission_gate
XM1 net1 en_b VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  rs_b_latch.sym # of pins=4
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/rs_b_latch.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/rs_b_latch.sch
.subckt rs_b_latch  s_b r_b q q_b  VDD  VSS
*.ipin s_b
*.ipin r_b
*.opin q
*.opin q_b
x1 s_b q_b VSS VSS VDD VDD q sky130_fd_sc_hd__nand2_4
x2 r_b q VSS VSS VDD VDD q_b sky130_fd_sc_hd__nand2_4
.ends


* expanding   symbol:  comparator_core_large.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator_core_large.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator_core_large.sch
.subckt comparator_core_large  ip in s_b clk r_b  VDD  VSS
*.ipin clk
*.ipin ip
*.ipin in
*.opin s_b
*.opin r_b
XM1 tail_d clk VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=32 m=32 
XM2 p ip tail_d VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=160 m=160 
XM3 q in tail_d VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=160 m=160 
XM4 s_b r_b p VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=80 m=80 
XM5 r_b s_b q VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=80 m=80 
XM6 s_b r_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=40 m=40 
XM7 r_b s_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=40 m=40 
XM8 s_b clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM9 r_b clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM10 p clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM11 q clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM12 tail_d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM13 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=24 m=24 
XM17 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM14 q VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM15 p VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM16 r_b VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM18 s_b VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  folded_cascode_3_bias.sym # of pins=6
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_bias.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_bias.sch
.subckt folded_cascode_3_bias  bias_a bias_b bias_c bias_d bias_e i_bias  VDD  VSS
*.opin bias_a
*.opin bias_b
*.opin bias_c
*.opin bias_d
*.opin bias_e
*.ipin i_bias
XM22 bias_b bias_c m21d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM26 m2d bias_c m25d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM32 bias_e bias_c m31d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM21 m21d bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM25 m25d bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM31 m31d bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM1 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=56 m=56 
XM2 m2d m2d bias_d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=50 m=50 
XM3 bias_d m2d bias_a VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM4 bias_a bias_d m5d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM5 m5d bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM6 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM7 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM33 bias_e bias_e net1 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM49 net1 bias_e net2 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM50 net2 bias_e net3 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM63 net3 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM68 bias_e bias_e net4 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM69 net4 bias_e net5 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM70 net5 bias_e net6 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM71 net6 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM72 bias_e bias_e net7 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM73 net7 bias_e net8 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM74 net8 bias_e net9 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM75 net9 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM76 bias_e bias_e net10 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM77 net10 bias_e net11 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM78 net11 bias_e net12 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM79 net12 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM64 bias_e bias_e net13 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM65 net13 bias_e net14 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM66 net14 bias_e net15 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM67 net15 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM57 bias_b VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM58 m2d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM59 bias_e VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM60 m31d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM42 m5d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM44 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM34 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM35 m2d m2d m2d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM36 bias_a bias_a bias_a VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4 
XM37 bias_e bias_e bias_e VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM54 m25d m25d m25d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM29 m5d m5d m5d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM8 i_bias i_bias i_bias VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM10 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM27 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM46 m21d m21d m21d VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM47 m25d m25d m25d VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM48 m31d m31d m31d VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM51 m21d m21d m21d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  sc_cmfb.sym # of pins=9
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/sc_cmfb.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/sc_cmfb.sch
.subckt sc_cmfb  phi1 phi1_b op on cm bias_a cmc phi2 phi2_b  VDD  VSS
*.ipin on
*.ipin cm
*.ipin bias_a
*.ipin op
*.opin cmc
*.ipin phi2_b
*.ipin phi2
*.ipin phi1_b
*.ipin phi1
XC3 op cmc sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=4 m=4
XC4 on cmc sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=4 m=4
x1 net1 op phi2 phi2_b VDD VSS transmission_gate
x2 net2 cmc phi2 phi2_b VDD VSS transmission_gate
x3 net3 on phi2 phi2_b VDD VSS transmission_gate
x4 cm net1 phi1 phi1_b VDD VSS transmission_gate
x5 bias_a net2 phi1 phi1_b VDD VSS transmission_gate
x6 cm net3 phi1 phi1_b VDD VSS transmission_gate
XC1 net1 net2 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
XC2 net3 net2 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
x7 cm net4 phi2 phi2_b VDD VSS transmission_gate
x8 bias_a net5 phi2 phi2_b VDD VSS transmission_gate
x9 cm net6 phi2 phi2_b VDD VSS transmission_gate
x10 net4 op phi1 phi1_b VDD VSS transmission_gate
x11 net5 cmc phi1 phi1_b VDD VSS transmission_gate
x12 net6 on phi1 phi1_b VDD VSS transmission_gate
XC5 net4 net5 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
XC6 net6 net5 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
XCdummy __UNCONNECTED_PIN__4 __UNCONNECTED_PIN__5 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=20 m=20
.ends


* expanding   symbol:  folded_cascode_3_core.sym # of pins=9
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_core.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_core.sch
.subckt folded_cascode_3_core  cmc ip in bias_a bias_b bias_c bias_d op on  VDD  VSS
*.ipin cmc
*.ipin ip
*.ipin in
*.ipin bias_a
*.ipin bias_b
*.ipin bias_c
*.ipin bias_d
*.opin op
*.opin on
XM1 foldp ip tail VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM2 foldn in tail VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM6 tail cmc VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=96 m=96 
XM5 tail bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=96 m=96 
XM11 foldp bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24 
XM12 foldn bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24 
XM1A on bias_c foldp VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM8 op bias_c foldn VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM3A on bias_d m3d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM7 op bias_d m4d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM3 m3d bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM4 m4d bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM82 foldn foldn foldn VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM83 foldp foldp foldp VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM55 foldn VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM56 op VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM61 foldp VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM62 on VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM40 m4d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM41 m3d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM38 op op op VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM39 on on on VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM30 tail VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM23 foldp foldp foldp VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM24 foldn foldn foldn VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM80 op VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM81 on VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM28 tail tail tail VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
.ends

