magic
tech sky130A
magscale 1 2
timestamp 1655456512
<< nwell >>
rect 1090 2797 1136 2843
rect 1406 2797 1452 2843
rect 1722 2797 1768 2843
rect 2038 2797 2084 2843
rect 2354 2797 2400 2843
rect 2670 2797 2716 2843
rect 2986 2797 3032 2843
rect 3302 2797 3348 2843
rect 142 1712 188 1815
rect 3302 1758 3348 1799
rect 3141 1502 3193 1545
<< pwell >>
rect 3141 1441 3193 1452
rect 3302 1190 3348 1235
rect 142 116 188 206
rect 458 116 504 206
rect 774 116 820 206
rect 1090 116 1136 206
rect 1406 116 1452 206
rect 1722 116 1768 206
rect 2038 116 2084 206
rect 2354 116 2400 206
rect 2670 116 2716 206
rect 2986 116 3032 206
rect 3302 159 3348 205
<< mvndiff >>
rect 142 194 188 206
rect 458 194 504 206
rect 774 194 820 206
rect 1090 194 1136 206
rect 1406 194 1452 206
rect 1722 194 1768 206
rect 2038 194 2084 206
rect 2354 194 2400 206
rect 2670 194 2716 206
rect 2986 194 3032 206
<< mvpdiff >>
rect 1090 2797 1136 2799
rect 1406 2797 1452 2799
rect 1722 2797 1768 2799
rect 2038 2797 2084 2799
rect 2354 2797 2400 2799
rect 2670 2797 2716 2799
rect 2986 2797 3032 2799
rect 3302 2797 3348 2799
<< locali >>
rect 1096 2797 1130 2803
rect 1412 2797 1446 2803
rect 1728 2797 1762 2803
rect 2044 2797 2078 2803
rect 2360 2797 2394 2803
rect 2676 2797 2710 2803
rect 2992 2797 3026 2803
rect 3308 2797 3342 2803
rect 148 190 182 206
rect 464 190 498 206
rect 780 190 814 206
rect 1096 190 1130 206
rect 1412 190 1446 206
rect 1728 190 1762 206
rect 2044 190 2078 206
rect 2360 190 2394 206
rect 2676 190 2710 206
rect 2992 190 3026 206
<< viali >>
rect 110 2984 3380 3018
rect 14 1676 48 2922
rect 3442 1676 3476 2922
rect 14 80 48 1308
rect 3442 80 3476 1308
rect 110 -16 3380 18
<< metal1 >>
rect 8 3018 3482 3024
rect 8 2984 110 3018
rect 3380 2984 3482 3018
rect 8 2922 3482 2984
rect 8 1676 14 2922
rect 48 2840 3442 2922
rect 48 1758 60 2840
rect 142 2790 188 2840
rect 458 2796 504 2840
rect 774 2797 820 2840
rect 1090 2797 1136 2840
rect 1406 2797 1452 2840
rect 1722 2797 1768 2840
rect 2038 2797 2084 2840
rect 2354 2797 2400 2840
rect 2670 2797 2716 2840
rect 2986 2797 3032 2840
rect 3302 2797 3348 2840
rect 142 1758 188 1815
rect 287 1811 297 2787
rect 349 1811 359 2787
rect 603 1811 613 2787
rect 665 1811 675 2787
rect 919 1811 929 2787
rect 981 1811 991 2787
rect 1235 1811 1245 2787
rect 1297 1811 1307 2787
rect 1551 1811 1561 2787
rect 1613 1811 1623 2787
rect 1867 1811 1877 2787
rect 1929 1811 1939 2787
rect 2183 1811 2193 2787
rect 2245 1811 2255 2787
rect 2499 1811 2509 2787
rect 2561 1811 2571 2787
rect 2815 1811 2825 2787
rect 2877 1811 2887 2787
rect 3131 1811 3141 2787
rect 3193 1811 3203 2787
rect 3302 1758 3348 1799
rect 3430 1758 3442 2840
rect 48 1712 3442 1758
rect 48 1676 54 1712
rect 8 1664 54 1676
rect 3436 1676 3442 1712
rect 3476 1676 3482 2922
rect 3436 1664 3482 1676
rect -64 1545 3554 1556
rect -64 1441 297 1545
rect 349 1441 613 1545
rect 665 1441 929 1545
rect 981 1441 1245 1545
rect 1297 1441 1561 1545
rect 1613 1441 1877 1545
rect 1929 1441 2193 1545
rect 2245 1441 2509 1545
rect 2561 1441 2825 1545
rect 2877 1441 3141 1545
rect 3193 1441 3554 1545
rect -64 1428 3554 1441
rect 8 1308 54 1320
rect 8 80 14 1308
rect 48 1272 54 1308
rect 3436 1308 3482 1320
rect 3436 1272 3442 1308
rect 48 1226 3442 1272
rect 48 162 54 1226
rect 3302 1190 3348 1226
rect 287 206 297 1182
rect 349 206 359 1182
rect 603 206 613 1182
rect 665 206 675 1182
rect 919 206 929 1182
rect 981 206 991 1182
rect 1235 206 1245 1182
rect 1297 206 1307 1182
rect 1551 206 1561 1182
rect 1613 206 1623 1182
rect 1867 206 1877 1182
rect 1929 206 1939 1182
rect 2183 206 2193 1182
rect 2245 206 2255 1182
rect 2499 206 2509 1182
rect 2561 206 2571 1182
rect 2815 206 2825 1182
rect 2877 206 2887 1182
rect 3131 206 3141 1182
rect 3193 206 3203 1182
rect 142 162 188 206
rect 458 162 504 206
rect 774 162 820 206
rect 1090 162 1136 206
rect 1406 162 1452 206
rect 1722 162 1768 206
rect 2038 162 2084 206
rect 2354 162 2400 206
rect 2670 162 2716 206
rect 2986 162 3032 206
rect 3302 162 3348 205
rect 3436 162 3442 1226
rect 48 80 3442 162
rect 3476 80 3482 1308
rect 8 18 3482 80
rect 8 -16 110 18
rect 3380 -16 3482 18
rect 8 -22 3482 -16
<< via1 >>
rect 297 1811 349 2787
rect 613 1811 665 2787
rect 929 1811 981 2787
rect 1245 1811 1297 2787
rect 1561 1811 1613 2787
rect 1877 1811 1929 2787
rect 2193 1811 2245 2787
rect 2509 1811 2561 2787
rect 2825 1811 2877 2787
rect 3141 1811 3193 2787
rect 297 1441 349 1545
rect 613 1441 665 1545
rect 929 1441 981 1545
rect 1245 1441 1297 1545
rect 1561 1441 1613 1545
rect 1877 1441 1929 1545
rect 2193 1441 2245 1545
rect 2509 1441 2561 1545
rect 2825 1441 2877 1545
rect 3141 1441 3193 1545
rect 297 206 349 1182
rect 613 206 665 1182
rect 929 206 981 1182
rect 1245 206 1297 1182
rect 1561 206 1613 1182
rect 1877 206 1929 1182
rect 2193 206 2245 1182
rect 2509 206 2561 1182
rect 2825 206 2877 1182
rect 3141 206 3193 1182
<< metal2 >>
rect 297 2787 349 2797
rect 297 1545 349 1811
rect 297 1182 349 1441
rect 297 196 349 206
rect 613 2787 665 2797
rect 613 1545 665 1811
rect 613 1182 665 1441
rect 613 196 665 206
rect 929 2787 981 2797
rect 929 1545 981 1811
rect 929 1182 981 1441
rect 929 196 981 206
rect 1245 2787 1297 2797
rect 1245 1545 1297 1811
rect 1245 1182 1297 1441
rect 1245 196 1297 206
rect 1561 2787 1613 2797
rect 1561 1545 1613 1811
rect 1561 1182 1613 1441
rect 1561 196 1613 206
rect 1877 2787 1929 2797
rect 1877 1545 1929 1811
rect 1877 1182 1929 1441
rect 1877 196 1929 206
rect 2193 2787 2245 2797
rect 2193 1545 2245 1811
rect 2193 1182 2245 1441
rect 2193 196 2245 206
rect 2509 2787 2561 2797
rect 2509 1545 2561 1811
rect 2509 1182 2561 1441
rect 2509 196 2561 206
rect 2825 2787 2877 2797
rect 2825 1545 2877 1811
rect 2825 1182 2877 1441
rect 2825 196 2877 206
rect 3141 2787 3193 2797
rect 3141 1545 3193 1811
rect 3141 1182 3193 1441
rect 3141 196 3193 206
use sky130_fd_pr__nfet_g5v0d10v5_BRTJC6  sky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0
timestamp 1655456512
transform 1 0 1745 0 1 694
box -1779 -758 1779 758
use sky130_fd_pr__pfet_g5v0d10v5_CADZ46  sky130_fd_pr__pfet_g5v0d10v5_CADZ46_0
timestamp 1655456512
transform 1 0 1745 0 1 2299
box -1809 -797 1809 797
<< labels >>
flabel metal1 -53 1488 -53 1488 1 FreeSans 400 0 0 0 esd
port 1 n
flabel metal1 31 2928 31 2928 1 FreeSans 400 0 0 0 VDD
port 2 n power bidirectional
flabel metal1 31 72 31 72 1 FreeSans 400 0 0 0 VSS
port 3 n power bidirectional
<< end >>
