magic
tech sky130A
magscale 1 2
timestamp 1654898484
<< locali >>
rect 1171 993 1205 1027
rect 81 883 97 933
rect 81 72 97 122
rect 1171 -13 1205 19
<< metal1 >>
rect -53 993 995 1027
rect -53 19 -19 993
rect 193 832 227 993
rect 385 832 419 993
rect 577 832 611 993
rect 769 832 803 993
rect 961 832 995 993
rect 97 430 131 608
rect 289 430 323 608
rect 481 430 515 608
rect 673 430 707 608
rect 865 430 899 608
rect 1057 430 1091 608
rect 97 396 1091 430
rect 97 253 131 396
rect 289 253 323 396
rect 481 253 515 396
rect 673 253 707 396
rect 865 253 899 396
rect 1057 253 1091 396
rect 193 19 227 180
rect 385 19 419 180
rect 577 19 611 180
rect 769 19 803 180
rect 961 19 995 180
rect -53 -15 995 19
use nmos_tgate  nmos_tgate_0
timestamp 1654898484
transform 1 0 593 0 1 213
box -646 -262 648 200
use pmos_tgate  pmos_tgate_0
timestamp 1654898484
transform -1 0 595 0 -1 707
box -646 -356 648 294
<< labels >>
flabel locali 1188 2 1188 2 1 FreeSans 400 0 0 0 VSS
port 6 n ground bidirectional
flabel locali 1188 1010 1188 1010 1 FreeSans 400 0 0 0 VDD
port 5 n power bidirectional
flabel metal1 -34 410 -34 410 1 FreeSans 400 0 0 0 in
port 1 n
flabel metal1 1074 412 1074 412 1 FreeSans 400 0 0 0 out
port 2 n
flabel locali 88 98 88 98 1 FreeSans 400 0 0 0 en
port 3 n
flabel locali 88 910 88 910 1 FreeSans 400 0 0 0 en_b
port 4 n
<< end >>
