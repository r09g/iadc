magic
tech sky130A
magscale 1 2
timestamp 1654898484
<< locali >>
rect -4462 9301 10769 9557
rect -4462 8125 -4206 9301
rect 10513 8595 10769 9301
rect -2356 8339 8835 8595
rect -4462 7869 -3864 8125
rect -4462 6324 -4206 7869
rect -2356 7546 -2100 8339
rect -2679 7290 -2100 7546
rect -4462 6068 -3875 6324
rect -4462 4529 -4206 6068
rect -2356 5768 -2100 7290
rect -2672 5512 -2100 5768
rect -4462 4273 -3867 4529
rect -4462 2728 -4206 4273
rect -2356 3970 -2100 5512
rect -2682 3714 -2100 3970
rect -4462 2472 -3859 2728
rect -4462 893 -4206 2472
rect -2356 2169 -2100 3714
rect -2682 1913 -2100 2169
rect -4462 637 -3867 893
rect -4462 -880 -4206 637
rect -2356 360 -2100 1913
rect -2669 104 -2100 360
rect -4462 -1136 -3856 -880
rect -4462 -1791 -4206 -1136
rect -2356 -1420 -2100 104
rect -2674 -1669 -2100 -1420
rect 8579 7562 8835 8339
rect 10510 8307 10769 8595
rect 10510 8118 10766 8307
rect 10264 7862 10766 8118
rect 8579 7306 9067 7562
rect 8579 5758 8835 7306
rect 10510 6335 10766 7862
rect 10251 6079 10766 6335
rect 8579 5502 9064 5758
rect 8579 3970 8835 5502
rect 10510 4521 10766 6079
rect 10257 4265 10766 4521
rect 8579 3714 9067 3970
rect 8579 2166 8835 3714
rect 10510 2720 10766 4265
rect 10251 2464 10766 2720
rect 8579 1910 9054 2166
rect 8579 355 8835 1910
rect 10510 921 10766 2464
rect 10259 665 10766 921
rect 8579 99 9072 355
rect 8579 -1430 8835 99
rect 10510 -864 10766 665
rect 10262 -1120 10766 -864
rect 8579 -1669 9061 -1430
rect -2674 -1676 9061 -1669
rect -2356 -1686 9061 -1676
rect -4462 -1925 -4203 -1791
rect -2356 -1925 8835 -1686
rect -4459 -2663 -4203 -1925
rect 10510 -2663 10766 -1120
rect -4459 -2919 10766 -2663
<< viali >>
rect -3768 8142 -3734 8176
rect -2809 8142 -2775 8176
rect -3768 7330 -3734 7364
rect -2807 7331 -2773 7365
rect -3768 6343 -3734 6377
rect -2808 6342 -2774 6376
rect -3767 5530 -3733 5564
rect -2810 5530 -2776 5564
rect -3770 4542 -3736 4576
rect -2806 4542 -2772 4576
rect -3767 3730 -3733 3764
rect -2808 3731 -2774 3765
rect -3767 2743 -3733 2777
rect -2809 2743 -2775 2777
rect -3770 1930 -3736 1964
rect -2807 1930 -2773 1964
rect -3770 942 -3736 976
rect -2809 943 -2775 977
rect -3771 130 -3737 164
rect -2809 130 -2775 164
rect -3769 -859 -3735 -825
rect -2809 -856 -2775 -822
rect -3768 -1667 -3734 -1633
rect -2811 -1667 -2777 -1633
rect 9153 8144 9187 8178
rect 10121 8142 10155 8176
rect 9162 7331 9196 7365
rect 10125 7333 10159 7367
rect 9158 6346 9192 6380
rect 10123 6342 10157 6376
rect 9158 5533 9192 5567
rect 10123 5535 10157 5569
rect 9164 4542 9198 4576
rect 10125 4542 10159 4576
rect 9160 3729 9194 3763
rect 10129 3733 10163 3767
rect 9160 2746 9194 2780
rect 10121 2746 10155 2780
rect 9158 1931 9192 1965
rect 10125 1927 10159 1961
rect 9160 946 9194 980
rect 10125 940 10159 974
rect 9160 126 9194 160
rect 10119 131 10153 165
rect 9162 -858 9196 -824
rect 10123 -854 10157 -820
rect 9166 -1670 9200 -1636
rect 10125 -1672 10159 -1638
<< metal1 >>
rect -3795 8124 -3785 8188
rect -3721 8124 -3711 8188
rect -2835 8124 -2825 8188
rect -2761 8124 -2751 8188
rect 9135 8128 9145 8192
rect 9209 8128 9219 8192
rect 10099 8131 10109 8195
rect 10173 8131 10183 8195
rect -5376 7701 -4004 7773
rect -5376 7637 -3748 7701
rect -2635 7697 -335 7701
rect -5376 7566 -4004 7637
rect -2852 7631 -2842 7695
rect -2778 7631 -2768 7695
rect -2635 7637 2411 7697
rect -485 7633 2411 7637
rect 6851 7633 6861 7697
rect 6925 7633 9170 7697
rect -5376 -1267 -5169 7566
rect -3789 7318 -3779 7382
rect -3715 7318 -3705 7382
rect -2834 7314 -2824 7378
rect -2760 7314 -2750 7378
rect 1708 6396 1757 6398
rect -3794 6328 -3784 6392
rect -3720 6328 -3710 6392
rect -2832 6331 -2822 6395
rect -2758 6331 -2748 6395
rect 531 6334 1757 6396
rect 1821 6334 1827 6398
rect 531 6332 1807 6334
rect -4764 5899 -3996 5953
rect -4764 5835 -3748 5899
rect -4764 5746 -3996 5835
rect -2858 5831 -2848 5895
rect -2784 5831 -2774 5895
rect -2637 5893 -431 5894
rect -2637 5830 -477 5893
rect -487 5829 -477 5830
rect -413 5829 -403 5893
rect -4764 577 -4557 5746
rect -3791 5517 -3781 5581
rect -3717 5517 -3707 5581
rect -2833 5517 -2823 5581
rect -2759 5517 -2749 5581
rect 531 4777 595 6332
rect 531 4707 595 4713
rect -3795 4527 -3785 4591
rect -3721 4527 -3711 4591
rect -2834 4527 -2824 4591
rect -2760 4527 -2750 4591
rect 2347 4563 2411 7633
rect 10290 7561 11546 7768
rect 9134 7312 9144 7376
rect 9208 7312 9218 7376
rect 10101 7315 10111 7379
rect 10175 7315 10185 7379
rect 9138 6332 9148 6396
rect 9212 6332 9222 6396
rect 10098 6330 10108 6394
rect 10172 6330 10182 6394
rect 6728 5895 6822 5896
rect 6694 5831 6704 5895
rect 6768 5893 6822 5895
rect 6768 5831 9181 5893
rect 6728 5829 9181 5831
rect 10294 5758 10980 5965
rect 9137 5516 9147 5580
rect 9211 5516 9221 5580
rect 10096 5515 10106 5579
rect 10170 5515 10180 5579
rect 2347 4499 3106 4563
rect 3170 4499 3180 4563
rect 9137 4530 9147 4594
rect 9211 4530 9221 4594
rect 10098 4529 10108 4593
rect 10172 4529 10182 4593
rect -4279 4100 -4072 4168
rect 3249 4148 3259 4212
rect 3323 4148 3333 4212
rect 10773 4159 10980 5758
rect -4279 4036 -3746 4100
rect -4279 2301 -4072 4036
rect -2854 4031 -2844 4095
rect -2780 4031 -2770 4095
rect -2627 4094 -374 4098
rect -2627 4034 -434 4094
rect -444 4030 -434 4034
rect -370 4030 -360 4094
rect 3259 4085 3323 4148
rect -3793 3714 -3783 3778
rect -3719 3714 -3709 3778
rect -2831 3717 -2821 3781
rect -2757 3717 -2747 3781
rect -3796 2725 -3786 2789
rect -3722 2725 -3712 2789
rect -2829 2727 -2819 2791
rect -2755 2727 -2745 2791
rect -4279 2237 -3737 2301
rect -4279 2193 -4072 2237
rect -2857 2231 -2847 2295
rect -2783 2231 -2773 2295
rect -2634 2291 -387 2298
rect -2634 2234 -434 2291
rect -444 2227 -434 2234
rect -370 2227 -360 2291
rect 3259 2223 3322 4085
rect 6749 4031 6759 4095
rect 6823 4031 9191 4095
rect 10287 3952 10980 4159
rect 9136 3714 9146 3778
rect 9210 3714 9220 3778
rect 10099 3719 10109 3783
rect 10173 3719 10183 3783
rect 9137 2727 9147 2791
rect 9211 2727 9221 2791
rect 10097 2727 10107 2791
rect 10171 2727 10181 2791
rect 10773 2355 10980 3952
rect 6754 2233 6764 2297
rect 6828 2233 9179 2297
rect 3249 2159 3259 2223
rect 3323 2159 3333 2223
rect 10290 2148 10980 2355
rect -3794 1917 -3784 1981
rect -3720 1917 -3710 1981
rect -2828 1919 -2818 1983
rect -2754 1919 -2744 1983
rect 9134 1913 9144 1977
rect 9208 1913 9218 1977
rect 10099 1915 10109 1979
rect 10173 1915 10183 1979
rect 6473 1822 6537 1828
rect 5418 1704 5482 1710
rect -364 1576 2330 1640
rect 2394 1576 2404 1640
rect -3794 928 -3784 992
rect -3720 928 -3710 992
rect -2831 928 -2821 992
rect -2757 928 -2747 992
rect -4764 497 -4115 577
rect -4764 433 -3751 497
rect -2850 433 -2840 497
rect -2776 433 -2766 497
rect -364 494 -300 1576
rect 157 1341 221 1347
rect 221 1277 1802 1341
rect 157 1271 221 1277
rect 1738 1041 1802 1277
rect 5418 1206 5482 1640
rect 5418 1136 5482 1142
rect 4720 897 4805 908
rect 6473 897 6537 1758
rect 9136 926 9146 990
rect 9210 926 9220 990
rect 10101 927 10111 991
rect 10175 927 10185 991
rect 4720 833 4731 897
rect 4795 833 6537 897
rect 4720 822 4805 833
rect 10773 602 10980 2148
rect -4764 370 -4115 433
rect -2631 430 -299 494
rect 6722 493 9180 497
rect 6690 429 6700 493
rect 6764 433 9180 493
rect 6764 429 6774 433
rect 10283 395 10980 602
rect -3794 114 -3784 178
rect -3720 114 -3710 178
rect -2831 118 -2821 182
rect -2757 118 -2747 182
rect 9136 115 9146 179
rect 9210 115 9220 179
rect 10098 116 10108 180
rect 10172 116 10182 180
rect -3794 -872 -3784 -808
rect -3720 -872 -3710 -808
rect -2833 -871 -2823 -807
rect -2759 -871 -2749 -807
rect 9138 -873 9148 -809
rect 9212 -873 9222 -809
rect 10098 -873 10108 -809
rect 10172 -873 10182 -809
rect 11339 -1197 11546 7561
rect -5376 -1301 -4113 -1267
rect -5376 -1365 -3759 -1301
rect -512 -1302 -502 -1301
rect -5376 -1474 -4113 -1365
rect -2849 -1368 -2839 -1304
rect -2775 -1368 -2765 -1304
rect -2638 -1365 -502 -1302
rect -438 -1365 -428 -1301
rect 6807 -1363 6817 -1299
rect 6881 -1300 6891 -1299
rect 6881 -1363 9185 -1300
rect 6866 -1364 9185 -1363
rect -2638 -1366 -440 -1365
rect 10286 -1404 11546 -1197
rect -3791 -1686 -3781 -1622
rect -3717 -1686 -3707 -1622
rect -2834 -1684 -2824 -1620
rect -2760 -1684 -2750 -1620
rect 9135 -1683 9145 -1619
rect 9209 -1683 9219 -1619
rect 10100 -1684 10110 -1620
rect 10174 -1684 10184 -1620
<< via1 >>
rect -3785 8176 -3721 8188
rect -3785 8142 -3768 8176
rect -3768 8142 -3734 8176
rect -3734 8142 -3721 8176
rect -3785 8124 -3721 8142
rect -2825 8176 -2761 8188
rect -2825 8142 -2809 8176
rect -2809 8142 -2775 8176
rect -2775 8142 -2761 8176
rect -2825 8124 -2761 8142
rect 9145 8178 9209 8192
rect 9145 8144 9153 8178
rect 9153 8144 9187 8178
rect 9187 8144 9209 8178
rect 9145 8128 9209 8144
rect 10109 8176 10173 8195
rect 10109 8142 10121 8176
rect 10121 8142 10155 8176
rect 10155 8142 10173 8176
rect 10109 8131 10173 8142
rect -2842 7631 -2778 7695
rect 6861 7633 6925 7697
rect -3779 7364 -3715 7382
rect -3779 7330 -3768 7364
rect -3768 7330 -3734 7364
rect -3734 7330 -3715 7364
rect -3779 7318 -3715 7330
rect -2824 7365 -2760 7378
rect -2824 7331 -2807 7365
rect -2807 7331 -2773 7365
rect -2773 7331 -2760 7365
rect -2824 7314 -2760 7331
rect -3784 6377 -3720 6392
rect -3784 6343 -3768 6377
rect -3768 6343 -3734 6377
rect -3734 6343 -3720 6377
rect -3784 6328 -3720 6343
rect -2822 6376 -2758 6395
rect -2822 6342 -2808 6376
rect -2808 6342 -2774 6376
rect -2774 6342 -2758 6376
rect -2822 6331 -2758 6342
rect 1757 6334 1821 6398
rect -2848 5831 -2784 5895
rect -477 5829 -413 5893
rect -3781 5564 -3717 5581
rect -3781 5530 -3767 5564
rect -3767 5530 -3733 5564
rect -3733 5530 -3717 5564
rect -3781 5517 -3717 5530
rect -2823 5564 -2759 5581
rect -2823 5530 -2810 5564
rect -2810 5530 -2776 5564
rect -2776 5530 -2759 5564
rect -2823 5517 -2759 5530
rect 531 4713 595 4777
rect -3785 4576 -3721 4591
rect -3785 4542 -3770 4576
rect -3770 4542 -3736 4576
rect -3736 4542 -3721 4576
rect -3785 4527 -3721 4542
rect -2824 4576 -2760 4591
rect -2824 4542 -2806 4576
rect -2806 4542 -2772 4576
rect -2772 4542 -2760 4576
rect -2824 4527 -2760 4542
rect 9144 7365 9208 7376
rect 9144 7331 9162 7365
rect 9162 7331 9196 7365
rect 9196 7331 9208 7365
rect 9144 7312 9208 7331
rect 10111 7367 10175 7379
rect 10111 7333 10125 7367
rect 10125 7333 10159 7367
rect 10159 7333 10175 7367
rect 10111 7315 10175 7333
rect 9148 6380 9212 6396
rect 9148 6346 9158 6380
rect 9158 6346 9192 6380
rect 9192 6346 9212 6380
rect 9148 6332 9212 6346
rect 10108 6376 10172 6394
rect 10108 6342 10123 6376
rect 10123 6342 10157 6376
rect 10157 6342 10172 6376
rect 10108 6330 10172 6342
rect 6704 5831 6768 5895
rect 9147 5567 9211 5580
rect 9147 5533 9158 5567
rect 9158 5533 9192 5567
rect 9192 5533 9211 5567
rect 9147 5516 9211 5533
rect 10106 5569 10170 5579
rect 10106 5535 10123 5569
rect 10123 5535 10157 5569
rect 10157 5535 10170 5569
rect 10106 5515 10170 5535
rect 3106 4499 3170 4563
rect 9147 4576 9211 4594
rect 9147 4542 9164 4576
rect 9164 4542 9198 4576
rect 9198 4542 9211 4576
rect 9147 4530 9211 4542
rect 10108 4576 10172 4593
rect 10108 4542 10125 4576
rect 10125 4542 10159 4576
rect 10159 4542 10172 4576
rect 10108 4529 10172 4542
rect 3259 4148 3323 4212
rect -2844 4031 -2780 4095
rect -434 4030 -370 4094
rect -3783 3764 -3719 3778
rect -3783 3730 -3767 3764
rect -3767 3730 -3733 3764
rect -3733 3730 -3719 3764
rect -3783 3714 -3719 3730
rect -2821 3765 -2757 3781
rect -2821 3731 -2808 3765
rect -2808 3731 -2774 3765
rect -2774 3731 -2757 3765
rect -2821 3717 -2757 3731
rect -3786 2777 -3722 2789
rect -3786 2743 -3767 2777
rect -3767 2743 -3733 2777
rect -3733 2743 -3722 2777
rect -3786 2725 -3722 2743
rect -2819 2777 -2755 2791
rect -2819 2743 -2809 2777
rect -2809 2743 -2775 2777
rect -2775 2743 -2755 2777
rect -2819 2727 -2755 2743
rect -2847 2231 -2783 2295
rect -434 2227 -370 2291
rect 6759 4031 6823 4095
rect 9146 3763 9210 3778
rect 9146 3729 9160 3763
rect 9160 3729 9194 3763
rect 9194 3729 9210 3763
rect 9146 3714 9210 3729
rect 10109 3767 10173 3783
rect 10109 3733 10129 3767
rect 10129 3733 10163 3767
rect 10163 3733 10173 3767
rect 10109 3719 10173 3733
rect 9147 2780 9211 2791
rect 9147 2746 9160 2780
rect 9160 2746 9194 2780
rect 9194 2746 9211 2780
rect 9147 2727 9211 2746
rect 10107 2780 10171 2791
rect 10107 2746 10121 2780
rect 10121 2746 10155 2780
rect 10155 2746 10171 2780
rect 10107 2727 10171 2746
rect 6764 2233 6828 2297
rect 3259 2159 3323 2223
rect -3784 1964 -3720 1981
rect -3784 1930 -3770 1964
rect -3770 1930 -3736 1964
rect -3736 1930 -3720 1964
rect -3784 1917 -3720 1930
rect -2818 1964 -2754 1983
rect -2818 1930 -2807 1964
rect -2807 1930 -2773 1964
rect -2773 1930 -2754 1964
rect -2818 1919 -2754 1930
rect 9144 1965 9208 1977
rect 9144 1931 9158 1965
rect 9158 1931 9192 1965
rect 9192 1931 9208 1965
rect 9144 1913 9208 1931
rect 10109 1961 10173 1979
rect 10109 1927 10125 1961
rect 10125 1927 10159 1961
rect 10159 1927 10173 1961
rect 10109 1915 10173 1927
rect 6473 1758 6537 1822
rect 5418 1640 5482 1704
rect 2330 1576 2394 1640
rect -3784 976 -3720 992
rect -3784 942 -3770 976
rect -3770 942 -3736 976
rect -3736 942 -3720 976
rect -3784 928 -3720 942
rect -2821 977 -2757 992
rect -2821 943 -2809 977
rect -2809 943 -2775 977
rect -2775 943 -2757 977
rect -2821 928 -2757 943
rect -2840 433 -2776 497
rect 157 1277 221 1341
rect 5418 1142 5482 1206
rect 9146 980 9210 990
rect 9146 946 9160 980
rect 9160 946 9194 980
rect 9194 946 9210 980
rect 9146 926 9210 946
rect 10111 974 10175 991
rect 10111 940 10125 974
rect 10125 940 10159 974
rect 10159 940 10175 974
rect 10111 927 10175 940
rect 4731 833 4795 897
rect 6700 429 6764 493
rect -3784 164 -3720 178
rect -3784 130 -3771 164
rect -3771 130 -3737 164
rect -3737 130 -3720 164
rect -3784 114 -3720 130
rect -2821 164 -2757 182
rect -2821 130 -2809 164
rect -2809 130 -2775 164
rect -2775 130 -2757 164
rect -2821 118 -2757 130
rect 9146 160 9210 179
rect 9146 126 9160 160
rect 9160 126 9194 160
rect 9194 126 9210 160
rect 9146 115 9210 126
rect 10108 165 10172 180
rect 10108 131 10119 165
rect 10119 131 10153 165
rect 10153 131 10172 165
rect 10108 116 10172 131
rect -3784 -825 -3720 -808
rect -3784 -859 -3769 -825
rect -3769 -859 -3735 -825
rect -3735 -859 -3720 -825
rect -3784 -872 -3720 -859
rect -2823 -822 -2759 -807
rect -2823 -856 -2809 -822
rect -2809 -856 -2775 -822
rect -2775 -856 -2759 -822
rect -2823 -871 -2759 -856
rect 9148 -824 9212 -809
rect 9148 -858 9162 -824
rect 9162 -858 9196 -824
rect 9196 -858 9212 -824
rect 9148 -873 9212 -858
rect 10108 -820 10172 -809
rect 10108 -854 10123 -820
rect 10123 -854 10157 -820
rect 10157 -854 10172 -820
rect 10108 -873 10172 -854
rect -2839 -1368 -2775 -1304
rect -502 -1365 -438 -1301
rect 6817 -1363 6881 -1299
rect -3781 -1633 -3717 -1622
rect -3781 -1667 -3768 -1633
rect -3768 -1667 -3734 -1633
rect -3734 -1667 -3717 -1633
rect -3781 -1686 -3717 -1667
rect -2824 -1633 -2760 -1620
rect -2824 -1667 -2811 -1633
rect -2811 -1667 -2777 -1633
rect -2777 -1667 -2760 -1633
rect -2824 -1684 -2760 -1667
rect 9145 -1636 9209 -1619
rect 9145 -1670 9166 -1636
rect 9166 -1670 9200 -1636
rect 9200 -1670 9209 -1636
rect 9145 -1683 9209 -1670
rect 10110 -1638 10174 -1620
rect 10110 -1672 10125 -1638
rect 10125 -1672 10159 -1638
rect 10159 -1672 10174 -1638
rect 10110 -1684 10174 -1672
<< metal2 >>
rect 10121 8205 10185 8206
rect -3785 8188 -3721 8198
rect -2825 8188 -2761 8198
rect -3787 8186 -3785 8187
rect -3794 8134 -3785 8186
rect -3787 8131 -3785 8134
rect -3721 8186 -3713 8187
rect -3721 8134 -2825 8186
rect -3721 8131 -3713 8134
rect -3785 8114 -3721 8124
rect 9145 8192 9209 8202
rect -2761 8134 -2758 8186
rect -2825 8114 -2761 8124
rect 10109 8196 10185 8205
rect 10109 8195 10121 8196
rect 9209 8134 10109 8186
rect 9145 8118 9209 8128
rect 10185 8134 10201 8186
rect 10173 8131 10185 8132
rect 10109 8122 10185 8131
rect 10109 8121 10173 8122
rect -2842 7855 2060 7919
rect -2842 7695 -2778 7855
rect -2842 7621 -2778 7631
rect -3779 7382 -3715 7392
rect -3794 7326 -3779 7378
rect -3484 7378 -3428 7387
rect -2824 7378 -2760 7388
rect -3715 7377 -2824 7378
rect -3715 7326 -3484 7377
rect -3779 7308 -3715 7318
rect -3428 7326 -2824 7377
rect -3484 7311 -3428 7321
rect -2824 7304 -2760 7314
rect 1996 6756 2060 7855
rect 6861 7697 6925 7707
rect 6861 7623 6925 7633
rect 9796 7387 9860 7397
rect 9144 7379 9208 7386
rect 9144 7376 9796 7379
rect 9208 7327 9796 7376
rect 10111 7379 10175 7389
rect 9860 7327 10111 7379
rect 9796 7313 9860 7323
rect 10175 7327 10201 7379
rect 9144 7302 9208 7312
rect 10111 7305 10175 7315
rect 1996 6682 2060 6692
rect -3784 6392 -3720 6402
rect -2822 6395 -2758 6405
rect -3794 6334 -3784 6386
rect -3720 6334 -2822 6386
rect -3784 6318 -3720 6328
rect 1745 6398 1834 6412
rect -2758 6334 -2756 6386
rect 1745 6334 1757 6398
rect 1821 6334 1834 6398
rect 9148 6396 9212 6406
rect -2822 6321 -2758 6331
rect 1745 6322 1834 6334
rect 4715 6297 4724 6361
rect 4788 6297 6497 6361
rect 9133 6334 9148 6386
rect 10108 6402 10172 6404
rect 10108 6394 10184 6402
rect 10172 6392 10184 6394
rect 9212 6334 10108 6386
rect 9148 6322 9212 6332
rect 10184 6334 10201 6386
rect 10108 6328 10120 6330
rect 10108 6320 10184 6328
rect 10120 6318 10184 6320
rect -2848 5895 -2784 5905
rect -2848 5726 -2784 5831
rect -477 5893 -413 5903
rect -477 5819 -413 5829
rect 3410 5781 3474 5791
rect -2848 5662 -133 5726
rect -3781 5581 -3717 5591
rect -3794 5526 -3781 5578
rect -3482 5578 -3426 5588
rect -2823 5581 -2759 5591
rect -3717 5526 -3482 5578
rect -3781 5507 -3717 5517
rect -3426 5526 -2823 5578
rect -3482 5512 -3426 5522
rect -2759 5526 -2747 5578
rect -2823 5507 -2759 5517
rect -197 5170 -133 5662
rect 1162 5616 1226 5622
rect 1162 5612 1346 5616
rect 1226 5552 1346 5612
rect 1162 5537 1226 5548
rect -197 5096 -133 5106
rect 520 4777 606 4789
rect 520 4713 531 4777
rect 595 4713 606 4777
rect 520 4700 606 4713
rect -3785 4591 -3721 4601
rect -3794 4534 -3785 4586
rect -2824 4591 -2760 4601
rect -3721 4534 -2824 4586
rect -3785 4517 -3721 4527
rect -2760 4534 -2756 4586
rect -2824 4517 -2760 4527
rect 1282 4219 1346 5552
rect 1630 5613 1694 5623
rect -434 4155 1429 4219
rect 1493 4155 1502 4219
rect -2844 4095 -2780 4105
rect -2844 3923 -2780 4031
rect -434 4094 -370 4155
rect -434 4020 -370 4030
rect -2844 3859 -369 3923
rect -3783 3778 -3719 3788
rect -3487 3779 -3431 3789
rect -3794 3726 -3783 3778
rect -3719 3726 -3487 3778
rect -3783 3704 -3719 3714
rect -2821 3781 -2757 3791
rect -3431 3726 -2821 3778
rect -3487 3713 -3431 3723
rect -2757 3726 -2752 3778
rect -2821 3707 -2757 3717
rect -433 3327 -369 3859
rect 333 3483 397 3493
rect 333 3409 397 3419
rect 765 3483 829 3493
rect 1408 3483 1472 3493
rect 829 3419 1408 3483
rect 765 3409 829 3419
rect 1408 3409 1472 3419
rect 333 3327 397 3337
rect -433 3307 333 3327
rect -434 3263 333 3307
rect 397 3263 402 3327
rect -3786 2789 -3722 2799
rect -3794 2734 -3786 2786
rect -3192 2787 -3136 2797
rect -3722 2734 -3192 2786
rect -3786 2715 -3722 2725
rect -2819 2791 -2755 2801
rect -3136 2734 -2819 2786
rect -3192 2721 -3136 2731
rect -2755 2734 -2743 2786
rect -2819 2717 -2755 2727
rect -434 2536 -370 3263
rect 333 3253 397 3263
rect 764 3153 828 3163
rect 1630 3153 1694 5549
rect 3410 5169 3474 5717
rect 3410 5095 3474 5105
rect 4658 5106 4722 5116
rect 5418 5106 5482 5116
rect 4722 5042 5418 5106
rect 4658 5032 4722 5042
rect 5418 5032 5482 5042
rect 4084 4928 4148 4938
rect 5706 4928 5770 4938
rect 4148 4864 5706 4928
rect 4084 4854 4148 4864
rect 5706 4854 5770 4864
rect 6433 4764 6497 6297
rect 6704 5895 6768 5905
rect 6704 5821 6768 5831
rect 9147 5580 9211 5590
rect 9130 5527 9147 5579
rect 9792 5582 9856 5592
rect 9211 5527 9792 5579
rect 9147 5506 9211 5516
rect 10106 5579 10170 5589
rect 9856 5527 10106 5579
rect 9792 5508 9856 5518
rect 10170 5527 10201 5579
rect 10106 5505 10170 5515
rect 6424 4700 6433 4764
rect 6497 4700 6506 4764
rect 9147 4594 9211 4604
rect 10120 4603 10184 4607
rect 3106 4563 3170 4573
rect 9144 4534 9147 4586
rect 10108 4597 10184 4603
rect 10108 4593 10120 4597
rect 9211 4534 10108 4586
rect 9147 4520 9211 4530
rect 10184 4534 10201 4586
rect 10172 4529 10184 4533
rect 10108 4523 10184 4529
rect 10108 4519 10172 4523
rect 3106 4489 3170 4499
rect 3259 4212 3323 4222
rect 3259 4138 3323 4148
rect 6759 4095 6823 4105
rect 5952 4031 6759 4095
rect 4876 3980 4940 3990
rect 5206 3980 5270 3990
rect 4940 3916 5206 3980
rect 4876 3906 4940 3916
rect 5206 3906 5270 3916
rect 828 3089 1694 3153
rect 764 3079 828 3089
rect 1630 3088 1694 3089
rect 3257 3862 3321 3872
rect -2847 2472 -370 2536
rect 2052 2507 2116 2791
rect 3257 2623 3321 3798
rect 4510 3462 4574 3472
rect 5952 3462 6016 4031
rect 6759 4021 6823 4031
rect 9146 3779 9210 3788
rect 9793 3783 9857 3793
rect 9146 3778 9793 3779
rect 9210 3727 9793 3778
rect 9146 3704 9210 3714
rect 10109 3783 10173 3793
rect 9857 3727 10109 3779
rect 9793 3709 9857 3719
rect 10173 3727 10201 3779
rect 10109 3709 10173 3719
rect 4574 3398 6016 3462
rect 4510 3388 4574 3398
rect 4508 3151 4572 3161
rect 4572 3087 6011 3151
rect 4508 3077 4572 3087
rect 3257 2549 3321 2559
rect -2847 2295 -2783 2472
rect 2052 2443 2671 2507
rect -2847 2221 -2783 2231
rect -434 2291 -370 2301
rect -3784 1981 -3720 1991
rect -3794 1926 -3784 1978
rect -2891 1983 -2754 1993
rect -2891 1979 -2818 1983
rect -2891 1978 -2884 1979
rect -3720 1926 -2884 1978
rect -3784 1907 -3720 1917
rect -2891 1923 -2884 1926
rect -2828 1923 -2818 1979
rect -2891 1919 -2818 1923
rect -2754 1926 -2725 1978
rect -2891 1909 -2754 1919
rect -434 1674 -370 2227
rect 1830 1674 1894 1684
rect -434 1610 1830 1674
rect 157 1513 221 1522
rect 157 1341 221 1449
rect 542 1513 606 1610
rect 1830 1600 1894 1610
rect 2330 1640 2394 1650
rect 2330 1566 2394 1576
rect 542 1457 544 1513
rect 600 1457 606 1513
rect 542 1418 606 1457
rect 2607 1528 2671 2443
rect 5947 2297 6011 3087
rect 9147 2791 9211 2801
rect 9144 2734 9147 2786
rect 9504 2792 9568 2802
rect 9211 2734 9504 2786
rect 9147 2717 9211 2727
rect 10107 2791 10171 2801
rect 9568 2734 10107 2786
rect 9504 2718 9568 2728
rect 10171 2734 10201 2786
rect 10107 2717 10171 2727
rect 6764 2297 6828 2307
rect 5947 2233 6764 2297
rect 3259 2223 3323 2233
rect 6764 2223 6828 2233
rect 3259 2149 3323 2159
rect 9193 1987 9257 1992
rect 9144 1982 9257 1987
rect 9144 1979 9193 1982
rect 9133 1977 9193 1979
rect 10109 1979 10173 1989
rect 9133 1927 9144 1977
rect 9257 1927 10109 1979
rect 9208 1913 9257 1918
rect 9144 1908 9257 1913
rect 10173 1927 10201 1979
rect 9144 1903 9208 1908
rect 10109 1905 10173 1915
rect 6461 1822 6549 1839
rect 4659 1811 4723 1820
rect 4659 1704 4723 1747
rect 6461 1758 6473 1822
rect 6537 1758 6549 1822
rect 6461 1742 6549 1758
rect 4659 1640 5418 1704
rect 5482 1640 5488 1704
rect 2607 1455 2671 1464
rect 3894 1522 3958 1532
rect 5736 1522 5800 1532
rect 3958 1458 5736 1522
rect 3894 1448 3958 1458
rect 5736 1448 5800 1458
rect 930 1341 994 1351
rect 3943 1341 4007 1351
rect 151 1277 157 1341
rect 221 1277 227 1341
rect 994 1277 3943 1341
rect 930 1267 994 1277
rect 3943 1267 4007 1277
rect 5403 1206 5499 1224
rect 5403 1142 5418 1206
rect 5482 1142 5499 1206
rect 5403 1127 5499 1142
rect -3784 992 -3720 1002
rect -3794 934 -3784 986
rect -3193 988 -3137 998
rect -3720 934 -3193 986
rect -3784 918 -3720 928
rect -2821 992 -2757 1002
rect -3137 934 -2821 986
rect -3193 922 -3137 932
rect 9146 990 9210 1000
rect -2757 934 -2755 986
rect 9144 934 9146 986
rect -2821 918 -2757 928
rect 9503 993 9567 1003
rect 9210 934 9503 986
rect 9146 916 9210 926
rect 10111 991 10175 1001
rect 9567 934 10111 986
rect 9503 919 9567 929
rect 10175 934 10201 986
rect 10111 917 10175 927
rect 4720 897 4805 908
rect 4720 833 4731 897
rect 4795 833 4805 897
rect 4720 822 4805 833
rect -2840 497 -2776 507
rect -2840 348 -2776 433
rect 6700 493 6764 503
rect 6700 419 6764 429
rect 1423 349 1487 359
rect -2840 285 1423 348
rect -2840 284 1487 285
rect 1423 275 1487 284
rect -2876 190 -2751 193
rect -3784 178 -3720 188
rect -2879 182 -2751 190
rect -2879 180 -2821 182
rect -3794 126 -3784 178
rect -3720 126 -2879 178
rect -2823 124 -2821 180
rect -2879 118 -2821 124
rect -2757 118 -2751 182
rect -2879 114 -2751 118
rect -3784 104 -3720 114
rect -2876 106 -2751 114
rect 9146 185 9210 189
rect 9146 179 9262 185
rect 10108 180 10172 190
rect 9210 175 10108 179
rect 9262 127 10108 175
rect 9146 111 9198 115
rect 9146 105 9262 111
rect 10172 127 10201 179
rect 10108 106 10172 116
rect 9198 101 9262 105
rect 160 -218 224 -208
rect -3784 -808 -3720 -798
rect -3794 -866 -3784 -814
rect -3200 -801 -3136 -791
rect -3720 -865 -3200 -814
rect -2823 -807 -2759 -797
rect -3136 -865 -2823 -814
rect -3720 -866 -2823 -865
rect -3784 -882 -3720 -872
rect -3200 -875 -3136 -866
rect -2759 -866 -2753 -814
rect -2823 -881 -2759 -871
rect -364 -1074 -300 -1064
rect -2839 -1138 -364 -1074
rect -2839 -1304 -2775 -1138
rect -364 -1148 -300 -1138
rect -2839 -1378 -2775 -1368
rect -502 -1301 -438 -1291
rect 160 -1301 224 -282
rect 9148 -809 9212 -799
rect 9145 -866 9148 -814
rect 9503 -811 9567 -801
rect 9212 -866 9503 -814
rect 9148 -883 9212 -873
rect 10108 -809 10172 -799
rect 9567 -866 10108 -814
rect 9503 -885 9567 -875
rect 10172 -866 10201 -814
rect 10108 -883 10172 -873
rect -438 -1365 224 -1301
rect 6817 -1299 6881 -1289
rect -502 -1375 -438 -1365
rect 6817 -1373 6881 -1363
rect -3781 -1622 -3717 -1612
rect -2885 -1620 -2760 -1610
rect -3794 -1674 -3781 -1622
rect -3717 -1674 -2885 -1622
rect -3781 -1696 -3717 -1686
rect 9145 -1612 9209 -1609
rect 9145 -1619 9261 -1612
rect 9209 -1621 9261 -1619
rect 10110 -1620 10174 -1610
rect 9209 -1622 10110 -1621
rect -2760 -1674 -2759 -1622
rect -2885 -1694 -2760 -1684
rect 9261 -1673 10110 -1622
rect 9145 -1686 9197 -1683
rect 9145 -1693 9261 -1686
rect 9197 -1696 9261 -1693
rect 10174 -1673 10201 -1621
rect 10110 -1694 10174 -1684
<< via2 >>
rect -3778 8131 -3722 8187
rect 10121 8195 10185 8196
rect 10121 8132 10173 8195
rect 10173 8132 10185 8195
rect -3484 7321 -3428 7377
rect 6861 7633 6925 7697
rect 9796 7323 9860 7387
rect 1996 6692 2060 6756
rect -3780 6330 -3724 6386
rect 1757 6334 1821 6398
rect 4724 6297 4788 6361
rect 10120 6330 10172 6392
rect 10172 6330 10184 6392
rect 10120 6328 10184 6330
rect -477 5829 -413 5893
rect -3482 5522 -3426 5578
rect 3410 5717 3474 5781
rect 1162 5548 1226 5612
rect -197 5106 -133 5170
rect 531 4713 595 4777
rect -3780 4531 -3724 4587
rect 1630 5549 1694 5613
rect 1429 4155 1493 4219
rect -3487 3723 -3431 3779
rect 333 3419 397 3483
rect 765 3419 829 3483
rect 1408 3419 1472 3483
rect 333 3263 397 3327
rect -3192 2731 -3136 2787
rect 3410 5105 3474 5169
rect 4658 5042 4722 5106
rect 5418 5042 5482 5106
rect 4084 4864 4148 4928
rect 5706 4864 5770 4928
rect 6704 5831 6768 5895
rect 9792 5518 9856 5582
rect 6433 4700 6497 4764
rect 3106 4499 3170 4563
rect 10120 4593 10184 4597
rect 10120 4533 10172 4593
rect 10172 4533 10184 4593
rect 3259 4148 3323 4212
rect 4876 3916 4940 3980
rect 5206 3916 5270 3980
rect 764 3089 828 3153
rect 3257 3798 3321 3862
rect 9793 3719 9857 3783
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3257 2559 3321 2623
rect -2884 1923 -2828 1979
rect 1830 1610 1894 1674
rect 157 1449 221 1513
rect 2330 1576 2394 1640
rect 544 1457 600 1513
rect 9504 2728 9568 2792
rect 3259 2159 3323 2223
rect 9193 1977 9257 1982
rect 9193 1918 9208 1977
rect 9208 1918 9257 1977
rect 4659 1747 4723 1811
rect 6473 1758 6537 1822
rect 2607 1464 2671 1528
rect 3894 1458 3958 1522
rect 5736 1458 5800 1522
rect 930 1277 994 1341
rect 3943 1277 4007 1341
rect 5418 1142 5482 1206
rect -3193 932 -3137 988
rect 9503 929 9567 993
rect 4731 833 4795 897
rect 6700 429 6764 493
rect 1423 285 1487 349
rect -2879 124 -2823 180
rect 9198 115 9210 175
rect 9210 115 9262 175
rect 9198 111 9262 115
rect 160 -282 224 -218
rect -3200 -865 -3136 -801
rect -364 -1138 -300 -1074
rect 9503 -875 9567 -811
rect 6817 -1363 6881 -1299
rect -2885 -1684 -2824 -1620
rect -2824 -1684 -2821 -1620
rect 9197 -1683 9209 -1622
rect 9209 -1683 9261 -1622
rect 9197 -1686 9261 -1683
<< metal3 >>
rect -3782 9961 -3718 9967
rect -3782 8192 -3718 9897
rect 10120 9961 10184 9969
rect -3490 9563 -3426 9569
rect -3783 8187 -3717 8192
rect -3783 8131 -3778 8187
rect -3722 8131 -3717 8187
rect -3783 8126 -3717 8131
rect -3782 6391 -3718 8126
rect -3490 7382 -3426 9499
rect 9786 9497 9796 9561
rect 9860 9497 9870 9561
rect -3199 9160 -3135 9166
rect 9496 9097 9506 9161
rect 9570 9097 9580 9161
rect -3494 7377 -3418 7382
rect -3494 7321 -3484 7377
rect -3428 7321 -3418 7377
rect -3494 7316 -3418 7321
rect -3790 6386 -3714 6391
rect -3790 6330 -3780 6386
rect -3724 6330 -3714 6386
rect -3790 6325 -3714 6330
rect -3782 4592 -3718 6325
rect -3490 5583 -3426 7316
rect -3492 5578 -3416 5583
rect -3492 5522 -3482 5578
rect -3426 5522 -3416 5578
rect -3492 5517 -3416 5522
rect -3790 4587 -3714 4592
rect -3790 4531 -3780 4587
rect -3724 4531 -3714 4587
rect -3790 4526 -3714 4531
rect -3782 4524 -3718 4526
rect -3490 3784 -3426 5517
rect -3497 3779 -3421 3784
rect -3497 3723 -3487 3779
rect -3431 3723 -3421 3779
rect -3497 3718 -3421 3723
rect -3490 3715 -3426 3718
rect -3199 2792 -3135 9096
rect -2889 8762 -2825 8768
rect -3202 2787 -3126 2792
rect -3202 2731 -3192 2787
rect -3136 2731 -3126 2787
rect -3202 2726 -3126 2731
rect -3199 993 -3135 2726
rect -2889 1984 -2825 8698
rect 9188 8697 9198 8761
rect 9262 8697 9272 8761
rect 6851 7697 6935 7702
rect 6851 7633 6861 7697
rect 6925 7633 6935 7697
rect 6851 7628 6935 7633
rect 6861 6879 6925 7628
rect 6191 6815 6925 6879
rect 1975 6756 2080 6780
rect 1975 6692 1996 6756
rect 2060 6692 2080 6756
rect 1975 6669 2080 6692
rect 6191 6515 6255 6815
rect 2896 6448 3638 6512
rect 1752 6398 1826 6403
rect 1752 6334 1757 6398
rect 1821 6334 1826 6398
rect 1752 6329 1826 6334
rect 4719 6361 4793 6366
rect 4719 6297 4724 6361
rect 4788 6297 4793 6361
rect 4719 6292 4793 6297
rect -497 5893 -391 5915
rect -497 5829 -477 5893
rect -413 5829 -391 5893
rect -497 5808 -391 5829
rect 6686 5895 6784 5914
rect 6686 5831 6704 5895
rect 6768 5831 6784 5895
rect 6686 5814 6784 5831
rect 3400 5781 3484 5810
rect 3400 5717 3410 5781
rect 3474 5717 3484 5781
rect 3400 5693 3484 5717
rect 1152 5612 1236 5617
rect 1150 5548 1162 5612
rect 1226 5548 1236 5612
rect 1152 5543 1236 5548
rect 1616 5613 1708 5646
rect 1616 5549 1630 5613
rect 1694 5549 1708 5613
rect 1616 5524 1708 5549
rect -238 5170 -98 5201
rect -238 5106 -197 5170
rect -133 5106 -98 5170
rect -238 5072 -98 5106
rect 3379 5169 3508 5177
rect 3379 5105 3410 5169
rect 3474 5105 3508 5169
rect 5418 5111 5482 5460
rect 3379 5097 3508 5105
rect 4648 5106 4732 5111
rect 4648 5042 4658 5106
rect 4722 5042 4732 5106
rect 4648 5037 4732 5042
rect 5408 5106 5492 5111
rect 5408 5042 5418 5106
rect 5482 5042 5492 5106
rect 5408 5037 5492 5042
rect 4061 4928 4171 4944
rect 4061 4864 4084 4928
rect 4148 4864 4171 4928
rect 4061 4850 4171 4864
rect 526 4777 600 4782
rect 526 4713 531 4777
rect 595 4713 600 4777
rect 526 4708 600 4713
rect 4658 4712 4722 5037
rect 5683 4928 5793 4943
rect 5683 4864 5706 4928
rect 5770 4864 5793 4928
rect 5683 4849 5793 4864
rect 6428 4764 6502 4769
rect 6428 4700 6433 4764
rect 6497 4700 6502 4764
rect 6428 4695 6502 4700
rect 3081 4563 3190 4586
rect 3081 4499 3106 4563
rect 3170 4499 3190 4563
rect 3081 4479 3190 4499
rect 1424 4219 1498 4224
rect 1424 4155 1429 4219
rect 1493 4155 1905 4219
rect 3249 4212 3333 4217
rect 1424 4150 1498 4155
rect 3249 4148 3259 4212
rect 3323 4148 3698 4212
rect 3249 4143 3333 4148
rect 4862 3980 4953 4019
rect 4862 3916 4876 3980
rect 4940 3916 4953 3980
rect 3234 3862 3340 3885
rect 4862 3879 4953 3916
rect 5193 3980 5284 4018
rect 5193 3916 5206 3980
rect 5270 3916 5284 3980
rect 5193 3878 5284 3916
rect 3234 3798 3257 3862
rect 3321 3798 3340 3862
rect 3234 3778 3340 3798
rect 333 3672 397 3761
rect 321 3483 410 3672
rect 321 3419 333 3483
rect 397 3419 410 3483
rect 321 3327 410 3419
rect 743 3483 849 3501
rect 743 3419 765 3483
rect 829 3419 849 3483
rect 743 3404 849 3419
rect 1397 3483 1484 3517
rect 1397 3419 1408 3483
rect 1472 3419 1484 3483
rect 1397 3388 1484 3419
rect 321 3263 333 3327
rect 397 3263 410 3327
rect 2348 3339 2412 3740
rect 4479 3462 4604 3492
rect 4479 3398 4510 3462
rect 4574 3398 4604 3462
rect 4479 3371 4604 3398
rect 2348 3275 3912 3339
rect 321 2948 410 3263
rect 745 3158 837 3183
rect 745 3153 838 3158
rect 745 3089 764 3153
rect 828 3089 838 3153
rect 745 3084 838 3089
rect 745 3061 837 3084
rect 333 2812 397 2948
rect 3848 2819 3912 3275
rect 4486 3151 4590 3171
rect 4486 3087 4508 3151
rect 4572 3087 4590 3151
rect 4486 3071 4590 3087
rect 6468 2920 6542 3631
rect 3235 2623 3341 2645
rect 3235 2559 3257 2623
rect 3321 2559 3341 2623
rect 3235 2538 3341 2559
rect 3249 2223 3333 2228
rect 2887 2159 3259 2223
rect 3323 2159 3333 2223
rect 3249 2154 3333 2159
rect 9199 1987 9263 8697
rect 9506 2797 9570 9097
rect 9796 7392 9860 9497
rect 10120 8201 10184 9897
rect 10111 8196 10195 8201
rect 10111 8132 10121 8196
rect 10185 8132 10195 8196
rect 10111 8127 10195 8132
rect 9786 7387 9870 7392
rect 9786 7323 9796 7387
rect 9860 7323 9870 7387
rect 9786 7318 9870 7323
rect 9796 5587 9860 7318
rect 10120 6397 10184 8127
rect 10110 6392 10194 6397
rect 10110 6328 10120 6392
rect 10184 6328 10194 6392
rect 10110 6323 10194 6328
rect 9782 5582 9866 5587
rect 9782 5518 9792 5582
rect 9856 5518 9866 5582
rect 9782 5513 9866 5518
rect 9796 3788 9860 5513
rect 10120 4602 10184 6323
rect 10110 4597 10194 4602
rect 10110 4533 10120 4597
rect 10184 4533 10194 4597
rect 10110 4528 10194 4533
rect 10120 4526 10184 4528
rect 9783 3783 9867 3788
rect 9783 3719 9793 3783
rect 9857 3719 9867 3783
rect 9783 3714 9867 3719
rect 9494 2792 9578 2797
rect 9494 2728 9504 2792
rect 9568 2728 9578 2792
rect 9494 2723 9578 2728
rect -2894 1979 -2818 1984
rect -2894 1923 -2884 1979
rect -2828 1923 -2818 1979
rect -2894 1918 -2818 1923
rect 9183 1982 9267 1987
rect 9183 1918 9193 1982
rect 9257 1918 9267 1982
rect -3203 988 -3127 993
rect -3203 932 -3193 988
rect -3137 932 -3127 988
rect -3203 927 -3127 932
rect -3199 -796 -3135 927
rect -2889 185 -2825 1918
rect 9183 1913 9267 1918
rect 1830 1866 1894 1868
rect 157 1518 221 1827
rect 1818 1674 1905 1866
rect 6468 1822 6542 1827
rect 4654 1811 4728 1816
rect 4654 1747 4659 1811
rect 4723 1747 4728 1811
rect 6468 1758 6473 1822
rect 6537 1758 6542 1822
rect 6468 1753 6542 1758
rect 4654 1742 4728 1747
rect 1818 1610 1830 1674
rect 1894 1610 1905 1674
rect 1818 1601 1905 1610
rect 2307 1640 2415 1666
rect 2307 1576 2330 1640
rect 2394 1576 2415 1640
rect 2307 1553 2415 1576
rect 2602 1528 2676 1533
rect 152 1513 226 1518
rect 152 1449 157 1513
rect 221 1449 226 1513
rect 539 1513 605 1518
rect 539 1457 544 1513
rect 600 1457 605 1513
rect 2602 1464 2607 1528
rect 2671 1464 2676 1528
rect 2602 1459 2676 1464
rect 3873 1522 3978 1546
rect 539 1452 605 1457
rect 152 1444 226 1449
rect 540 1112 604 1452
rect 910 1341 1011 1357
rect 910 1277 930 1341
rect 994 1277 1011 1341
rect 910 1259 1011 1277
rect 1733 1042 1807 1116
rect 2607 1115 2671 1459
rect 3873 1458 3894 1522
rect 3958 1458 3978 1522
rect 3873 1437 3978 1458
rect 5715 1522 5820 1544
rect 5715 1458 5736 1522
rect 5800 1458 5820 1522
rect 5715 1435 5820 1458
rect 3923 1341 4024 1360
rect 3923 1277 3943 1341
rect 4007 1277 4024 1341
rect 3923 1262 4024 1277
rect 5413 1206 5487 1211
rect 5413 1142 5418 1206
rect 5482 1142 5487 1206
rect 5413 1137 5487 1142
rect 4726 897 4800 902
rect 4726 833 4731 897
rect 4795 833 4800 897
rect 4726 828 4800 833
rect 5547 552 5566 616
rect 6683 493 6785 514
rect 6683 429 6700 493
rect 6764 429 6785 493
rect 6683 411 6785 429
rect 1405 349 1503 380
rect 1405 285 1423 349
rect 1487 285 1503 349
rect 2812 299 3629 363
rect 1405 260 1503 285
rect -2889 180 -2813 185
rect 9199 180 9263 1913
rect 9506 998 9570 2723
rect 9493 993 9577 998
rect 9493 929 9503 993
rect 9567 929 9577 993
rect 9493 924 9577 929
rect -2889 124 -2879 180
rect -2823 124 -2813 180
rect -2889 119 -2813 124
rect 9188 175 9272 180
rect -3210 -801 -3126 -796
rect -3210 -865 -3200 -801
rect -3136 -865 -3126 -801
rect -3210 -870 -3126 -865
rect -3199 -877 -3135 -870
rect -2889 -1615 -2825 119
rect 139 -218 245 -195
rect 139 -282 160 -218
rect 224 -282 245 -218
rect 139 -299 245 -282
rect 6179 -303 6243 116
rect 9188 111 9198 175
rect 9262 111 9272 175
rect 9188 106 9272 111
rect 6179 -367 6881 -303
rect -378 -1074 -280 -1056
rect -378 -1138 -364 -1074
rect -300 -1138 -280 -1074
rect -378 -1159 -280 -1138
rect 6817 -1294 6881 -367
rect 6807 -1299 6891 -1294
rect 6807 -1363 6817 -1299
rect 6881 -1363 6891 -1299
rect 6807 -1368 6891 -1363
rect 6817 -1372 6881 -1368
rect -2895 -1620 -2811 -1615
rect 9199 -1617 9263 106
rect 9506 -806 9570 924
rect 9493 -811 9577 -806
rect 9493 -875 9503 -811
rect 9567 -875 9577 -811
rect 9493 -880 9577 -875
rect 9506 -889 9570 -880
rect -2895 -1684 -2885 -1620
rect -2821 -1684 -2811 -1620
rect -2895 -1689 -2811 -1684
rect 9187 -1622 9271 -1617
rect 9187 -1686 9197 -1622
rect 9261 -1686 9271 -1622
rect 9187 -1691 9271 -1686
rect 9199 -1692 9263 -1691
<< via3 >>
rect -3782 9897 -3718 9961
rect 10120 9897 10184 9961
rect -3490 9499 -3426 9563
rect 9796 9497 9860 9561
rect -3199 9096 -3135 9160
rect 9506 9097 9570 9161
rect -2889 8698 -2825 8762
rect 9198 8697 9262 8761
rect 1996 6692 2060 6756
rect -477 5829 -413 5893
rect 6704 5831 6768 5895
rect 3410 5717 3474 5781
rect 1630 5549 1694 5613
rect -197 5106 -133 5170
rect 3410 5105 3474 5169
rect 4084 4864 4148 4928
rect 5706 4864 5770 4928
rect 3106 4499 3170 4563
rect 4876 3916 4940 3980
rect 5206 3916 5270 3980
rect 3257 3798 3321 3862
rect 765 3419 829 3483
rect 1408 3419 1472 3483
rect 4510 3398 4574 3462
rect 764 3089 828 3153
rect 4508 3087 4572 3151
rect 3257 2559 3321 2623
rect 2330 1576 2394 1640
rect 930 1277 994 1341
rect 3894 1458 3958 1522
rect 5736 1458 5800 1522
rect 3943 1277 4007 1341
rect 6700 429 6764 493
rect 1423 285 1487 349
rect 160 -282 224 -218
rect -364 -1138 -300 -1074
<< metal4 >>
rect -3783 9961 -3717 9962
rect 10119 9961 10185 9962
rect -3799 9897 -3782 9961
rect -3718 9897 10120 9961
rect 10184 9897 10185 9961
rect -3783 9896 -3717 9897
rect 10119 9896 10185 9897
rect -3491 9563 -3425 9564
rect -3491 9561 -3490 9563
rect -3799 9499 -3490 9561
rect -3426 9561 -3425 9563
rect 9795 9561 9861 9562
rect -3426 9499 9796 9561
rect -3799 9497 9796 9499
rect 9860 9497 10184 9561
rect 9795 9496 9861 9497
rect 9505 9161 9571 9162
rect -3799 9160 9506 9161
rect -3799 9097 -3199 9160
rect -3200 9096 -3199 9097
rect -3135 9097 9506 9160
rect 9570 9097 10184 9161
rect -3135 9096 -3134 9097
rect 9505 9096 9571 9097
rect -3200 9095 -3134 9096
rect -2890 8762 -2824 8763
rect -2890 8761 -2889 8762
rect -3799 8698 -2889 8761
rect -2825 8761 -2824 8762
rect 9197 8761 9263 8762
rect -2825 8698 9198 8761
rect -3799 8697 9198 8698
rect 9262 8697 10184 8761
rect 9197 8696 9263 8697
rect 1995 6756 2061 6757
rect 1995 6692 1996 6756
rect 2060 6692 2061 6756
rect 1995 6691 2061 6692
rect 1996 6377 2060 6691
rect 6703 5895 6769 5896
rect -478 5893 -412 5894
rect -478 5829 -477 5893
rect -413 5829 155 5893
rect 6322 5831 6704 5895
rect 6768 5831 6769 5895
rect 6703 5830 6769 5831
rect -478 5828 -412 5829
rect 3409 5781 3475 5782
rect 3409 5717 3410 5781
rect 3474 5717 3744 5781
rect 3409 5716 3475 5717
rect 1629 5613 1695 5614
rect 544 5311 608 5551
rect 1629 5549 1630 5613
rect 1694 5549 1949 5613
rect 1629 5548 1695 5549
rect 544 5247 5105 5311
rect -198 5170 -132 5171
rect -198 5106 -197 5170
rect -133 5169 -132 5170
rect 3409 5169 3475 5170
rect -133 5106 3410 5169
rect -198 5105 3410 5106
rect 3474 5105 3475 5169
rect 320 4612 384 5105
rect 3409 5104 3475 5105
rect 4083 4928 4149 4929
rect 1242 4864 4084 4928
rect 4148 4864 4150 4928
rect 765 3484 829 3761
rect 764 3483 830 3484
rect 764 3419 765 3483
rect 829 3419 830 3483
rect 764 3418 830 3419
rect 763 3153 829 3154
rect 763 3089 764 3153
rect 828 3089 829 3153
rect 763 3088 829 3089
rect 764 2811 828 3088
rect -364 1985 213 2049
rect -364 -1073 -300 1985
rect 930 1342 994 1946
rect 929 1341 995 1342
rect 929 1277 930 1341
rect 994 1277 995 1341
rect 929 1276 995 1277
rect 1242 859 1306 4864
rect 4083 4863 4149 4864
rect 3105 4563 3171 4564
rect 2808 4499 3106 4563
rect 3170 4499 3171 4563
rect 3105 4498 3171 4499
rect 4875 3980 4941 3981
rect 4875 3916 4876 3980
rect 4940 3916 4941 3980
rect 4875 3915 4941 3916
rect 3256 3862 3322 3863
rect 3256 3798 3257 3862
rect 3321 3798 3746 3862
rect 3256 3797 3322 3798
rect 1407 3483 1473 3484
rect 1407 3419 1408 3483
rect 1472 3419 1473 3483
rect 1407 3418 1473 3419
rect 998 795 1306 859
rect 1408 813 1472 3418
rect 2348 3339 2412 3740
rect 4510 3463 4574 3790
rect 4509 3462 4575 3463
rect 4509 3398 4510 3462
rect 4574 3398 4575 3462
rect 4509 3397 4575 3398
rect 2348 3275 3912 3339
rect 3848 2820 3912 3275
rect 4507 3151 4573 3152
rect 4507 3087 4508 3151
rect 4572 3087 4573 3151
rect 4507 3086 4573 3087
rect 4508 2788 4572 3086
rect 3256 2623 3322 2624
rect 2816 2559 3257 2623
rect 3321 2559 3322 2623
rect 3256 2558 3322 2559
rect 2330 1641 2394 1961
rect 2329 1640 2395 1641
rect 2329 1576 2330 1640
rect 2394 1576 2395 1640
rect 2329 1575 2395 1576
rect 3893 1522 3959 1523
rect 3224 1458 3894 1522
rect 3958 1458 3959 1522
rect 1408 749 1954 813
rect 3224 812 3288 1458
rect 3893 1457 3959 1458
rect 3943 1342 4007 1345
rect 3942 1341 4008 1342
rect 3942 1277 3943 1341
rect 4007 1277 4008 1341
rect 3942 1276 4008 1277
rect 3943 1007 4007 1276
rect 4876 844 4940 3915
rect 2812 748 3288 812
rect 4609 780 4940 844
rect 5041 616 5105 5247
rect 5706 4929 5770 5552
rect 5705 4928 5771 4929
rect 5705 4864 5706 4928
rect 5770 4864 5771 4928
rect 5705 4863 5771 4864
rect 5205 3980 5271 3981
rect 5205 3916 5206 3980
rect 5270 3916 5546 3980
rect 5205 3915 5271 3916
rect 5736 1523 5800 1953
rect 5735 1522 5801 1523
rect 5735 1458 5736 1522
rect 5800 1458 5801 1522
rect 5735 1457 5801 1458
rect 5041 552 5566 616
rect 6699 493 6765 494
rect 6384 429 6700 493
rect 6764 429 6766 493
rect 6699 428 6765 429
rect 1422 349 1488 350
rect 1420 285 1423 349
rect 1487 285 1953 349
rect 1422 284 1488 285
rect 160 -217 224 179
rect 159 -218 225 -217
rect 159 -282 160 -218
rect 224 -282 225 -218
rect 159 -283 225 -282
rect -365 -1074 -299 -1073
rect -365 -1138 -364 -1074
rect -300 -1138 -299 -1074
rect -365 -1139 -299 -1138
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1654898484
transform -1 0 10253 0 1 51
box -53 -49 1241 1063
use transmission_gate  transmission_gate_1
timestamp 1654898484
transform -1 0 10253 0 1 1851
box -53 -49 1241 1063
use transmission_gate  transmission_gate_2
timestamp 1654898484
transform -1 0 10253 0 1 -1749
box -53 -49 1241 1063
use transmission_gate  transmission_gate_3
timestamp 1654898484
transform -1 0 10253 0 1 3651
box -53 -49 1241 1063
use transmission_gate  transmission_gate_4
timestamp 1654898484
transform -1 0 10253 0 1 5451
box -53 -49 1241 1063
use transmission_gate  transmission_gate_5
timestamp 1654898484
transform -1 0 10253 0 1 7251
box -53 -49 1241 1063
use transmission_gate  transmission_gate_6
timestamp 1654898484
transform -1 0 -2677 0 1 7251
box -53 -49 1241 1063
use transmission_gate  transmission_gate_7
timestamp 1654898484
transform -1 0 -2677 0 1 5451
box -53 -49 1241 1063
use transmission_gate  transmission_gate_8
timestamp 1654898484
transform -1 0 -2677 0 1 3651
box -53 -49 1241 1063
use transmission_gate  transmission_gate_9
timestamp 1654898484
transform -1 0 -2677 0 1 1851
box -53 -49 1241 1063
use transmission_gate  transmission_gate_10
timestamp 1654898484
transform -1 0 -2677 0 1 51
box -53 -49 1241 1063
use transmission_gate  transmission_gate_11
timestamp 1654898484
transform -1 0 -2677 0 1 -1749
box -53 -49 1241 1063
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_0
timestamp 1654898484
transform 1 0 630 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_1
timestamp 1654898484
transform 1 0 2430 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_2
timestamp 1654898484
transform 1 0 4230 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_3
timestamp 1654898484
transform 1 0 6030 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_4
timestamp 1654898484
transform 1 0 6030 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_5
timestamp 1654898484
transform 1 0 4230 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_6
timestamp 1654898484
transform 1 0 2430 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_7
timestamp 1654898484
transform 1 0 630 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_8
timestamp 1654898484
transform 1 0 6030 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_9
timestamp 1654898484
transform 1 0 4230 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_10
timestamp 1654898484
transform 1 0 2430 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_11
timestamp 1654898484
transform 1 0 630 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_12
timestamp 1654898484
transform 1 0 6030 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_13
timestamp 1654898484
transform 1 0 4230 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_14
timestamp 1654898484
transform 1 0 2430 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_15
timestamp 1654898484
transform 1 0 630 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_16
timestamp 1654898484
transform 1 0 7830 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_17
timestamp 1654898484
transform 1 0 7830 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_18
timestamp 1654898484
transform 1 0 7830 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_19
timestamp 1654898484
transform 1 0 7830 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_20
timestamp 1654898484
transform 1 0 -1170 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_21
timestamp 1654898484
transform 1 0 -1170 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_22
timestamp 1654898484
transform 1 0 -1170 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_23
timestamp 1654898484
transform 1 0 -1170 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_24
timestamp 1654898484
transform 1 0 7830 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_25
timestamp 1654898484
transform 1 0 6030 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_26
timestamp 1654898484
transform 1 0 4230 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_27
timestamp 1654898484
transform 1 0 2430 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_28
timestamp 1654898484
transform 1 0 630 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_29
timestamp 1654898484
transform 1 0 -1170 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_30
timestamp 1654898484
transform 1 0 -1170 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_31
timestamp 1654898484
transform 1 0 630 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_32
timestamp 1654898484
transform 1 0 2430 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_33
timestamp 1654898484
transform 1 0 4230 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_34
timestamp 1654898484
transform 1 0 6030 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_35
timestamp 1654898484
transform 1 0 7830 0 1 -1220
box -630 -580 528 580
<< labels >>
flabel metal1 -5304 3369 -5304 3369 1 FreeSans 400 0 0 0 op
port 4 n
flabel metal1 -4692 3368 -4692 3368 1 FreeSans 400 0 0 0 on
port 1 n
flabel metal1 -4232 3371 -4232 3371 1 FreeSans 400 0 0 0 cmc
port 5 n
flabel metal1 10900 3295 10900 3295 1 FreeSans 400 0 0 0 cm
port 2 n
flabel metal1 11402 3298 11402 3298 1 FreeSans 400 0 0 0 bias_a
port 3 n
flabel locali -1902 9423 -1902 9423 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel locali -1884 8465 -1884 8465 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal4 -3651 9926 -3651 9926 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal4 -3653 9530 -3653 9530 1 FreeSans 400 0 0 0 p2
port 7 n
flabel metal4 -3652 9123 -3652 9123 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal4 -3653 8733 -3653 8733 1 FreeSans 400 0 0 0 p1
port 9 n
<< end >>
