magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -4124 181 -4066 187
rect -3704 181 -3646 187
rect -3284 181 -3226 187
rect -2864 181 -2806 187
rect -2444 181 -2386 187
rect -2024 181 -1966 187
rect -1604 181 -1546 187
rect -1184 181 -1126 187
rect -764 181 -706 187
rect -344 181 -286 187
rect 76 181 134 187
rect 496 181 554 187
rect 916 181 974 187
rect 1336 181 1394 187
rect 1756 181 1814 187
rect 2176 181 2234 187
rect 2596 181 2654 187
rect 3016 181 3074 187
rect 3436 181 3494 187
rect 3856 181 3914 187
rect -4124 147 -4112 181
rect -3704 147 -3692 181
rect -3284 147 -3272 181
rect -2864 147 -2852 181
rect -2444 147 -2432 181
rect -2024 147 -2012 181
rect -1604 147 -1592 181
rect -1184 147 -1172 181
rect -764 147 -752 181
rect -344 147 -332 181
rect 76 147 88 181
rect 496 147 508 181
rect 916 147 928 181
rect 1336 147 1348 181
rect 1756 147 1768 181
rect 2176 147 2188 181
rect 2596 147 2608 181
rect 3016 147 3028 181
rect 3436 147 3448 181
rect 3856 147 3868 181
rect -4124 141 -4066 147
rect -3704 141 -3646 147
rect -3284 141 -3226 147
rect -2864 141 -2806 147
rect -2444 141 -2386 147
rect -2024 141 -1966 147
rect -1604 141 -1546 147
rect -1184 141 -1126 147
rect -764 141 -706 147
rect -344 141 -286 147
rect 76 141 134 147
rect 496 141 554 147
rect 916 141 974 147
rect 1336 141 1394 147
rect 1756 141 1814 147
rect 2176 141 2234 147
rect 2596 141 2654 147
rect 3016 141 3074 147
rect 3436 141 3494 147
rect 3856 141 3914 147
rect -3914 -147 -3856 -141
rect -3494 -147 -3436 -141
rect -3074 -147 -3016 -141
rect -2654 -147 -2596 -141
rect -2234 -147 -2176 -141
rect -1814 -147 -1756 -141
rect -1394 -147 -1336 -141
rect -974 -147 -916 -141
rect -554 -147 -496 -141
rect -134 -147 -76 -141
rect 286 -147 344 -141
rect 706 -147 764 -141
rect 1126 -147 1184 -141
rect 1546 -147 1604 -141
rect 1966 -147 2024 -141
rect 2386 -147 2444 -141
rect 2806 -147 2864 -141
rect 3226 -147 3284 -141
rect 3646 -147 3704 -141
rect 4066 -147 4124 -141
rect -3914 -181 -3902 -147
rect -3494 -181 -3482 -147
rect -3074 -181 -3062 -147
rect -2654 -181 -2642 -147
rect -2234 -181 -2222 -147
rect -1814 -181 -1802 -147
rect -1394 -181 -1382 -147
rect -974 -181 -962 -147
rect -554 -181 -542 -147
rect -134 -181 -122 -147
rect 286 -181 298 -147
rect 706 -181 718 -147
rect 1126 -181 1138 -147
rect 1546 -181 1558 -147
rect 1966 -181 1978 -147
rect 2386 -181 2398 -147
rect 2806 -181 2818 -147
rect 3226 -181 3238 -147
rect 3646 -181 3658 -147
rect 4066 -181 4078 -147
rect -3914 -187 -3856 -181
rect -3494 -187 -3436 -181
rect -3074 -187 -3016 -181
rect -2654 -187 -2596 -181
rect -2234 -187 -2176 -181
rect -1814 -187 -1756 -181
rect -1394 -187 -1336 -181
rect -974 -187 -916 -181
rect -554 -187 -496 -181
rect -134 -187 -76 -181
rect 286 -187 344 -181
rect 706 -187 764 -181
rect 1126 -187 1184 -181
rect 1546 -187 1604 -181
rect 1966 -187 2024 -181
rect 2386 -187 2444 -181
rect 2806 -187 2864 -181
rect 3226 -187 3284 -181
rect 3646 -187 3704 -181
rect 4066 -187 4124 -181
rect -4122 -351 -4064 -345
rect -3702 -351 -3644 -345
rect -3282 -351 -3224 -345
rect -2862 -351 -2804 -345
rect -2442 -351 -2384 -345
rect -2022 -351 -1964 -345
rect -1602 -351 -1544 -345
rect -1182 -351 -1124 -345
rect -762 -351 -704 -345
rect -342 -351 -284 -345
rect 78 -351 136 -345
rect 498 -351 556 -345
rect 918 -351 976 -345
rect 1338 -351 1396 -345
rect 1758 -351 1816 -345
rect 2178 -351 2236 -345
rect 2598 -351 2656 -345
rect 3018 -351 3076 -345
rect 3438 -351 3496 -345
rect 3858 -351 3916 -345
rect -4122 -385 -4110 -351
rect -3702 -385 -3690 -351
rect -3282 -385 -3270 -351
rect -2862 -385 -2850 -351
rect -2442 -385 -2430 -351
rect -2022 -385 -2010 -351
rect -1602 -385 -1590 -351
rect -1182 -385 -1170 -351
rect -762 -385 -750 -351
rect -342 -385 -330 -351
rect 78 -385 90 -351
rect 498 -385 510 -351
rect 918 -385 930 -351
rect 1338 -385 1350 -351
rect 1758 -385 1770 -351
rect 2178 -385 2190 -351
rect 2598 -385 2610 -351
rect 3018 -385 3030 -351
rect 3438 -385 3450 -351
rect 3858 -385 3870 -351
rect -4122 -391 -4064 -385
rect -3702 -391 -3644 -385
rect -3282 -391 -3224 -385
rect -2862 -391 -2804 -385
rect -2442 -391 -2384 -385
rect -2022 -391 -1964 -385
rect -1602 -391 -1544 -385
rect -1182 -391 -1124 -385
rect -762 -391 -704 -385
rect -342 -391 -284 -385
rect 78 -391 136 -385
rect 498 -391 556 -385
rect 918 -391 976 -385
rect 1338 -391 1396 -385
rect 1758 -391 1816 -385
rect 2178 -391 2236 -385
rect 2598 -391 2656 -385
rect 3018 -391 3076 -385
rect 3438 -391 3496 -385
rect 3858 -391 3916 -385
rect -3912 -679 -3854 -673
rect -3492 -679 -3434 -673
rect -3072 -679 -3014 -673
rect -2652 -679 -2594 -673
rect -2232 -679 -2174 -673
rect -1812 -679 -1754 -673
rect -1392 -679 -1334 -673
rect -972 -679 -914 -673
rect -552 -679 -494 -673
rect -132 -679 -74 -673
rect 288 -679 346 -673
rect 708 -679 766 -673
rect 1128 -679 1186 -673
rect 1548 -679 1606 -673
rect 1968 -679 2026 -673
rect 2388 -679 2446 -673
rect 2808 -679 2866 -673
rect 3228 -679 3286 -673
rect 3648 -679 3706 -673
rect 4068 -679 4126 -673
rect -3912 -713 -3900 -679
rect -3492 -713 -3480 -679
rect -3072 -713 -3060 -679
rect -2652 -713 -2640 -679
rect -2232 -713 -2220 -679
rect -1812 -713 -1800 -679
rect -1392 -713 -1380 -679
rect -972 -713 -960 -679
rect -552 -713 -540 -679
rect -132 -713 -120 -679
rect 288 -713 300 -679
rect 708 -713 720 -679
rect 1128 -713 1140 -679
rect 1548 -713 1560 -679
rect 1968 -713 1980 -679
rect 2388 -713 2400 -679
rect 2808 -713 2820 -679
rect 3228 -713 3240 -679
rect 3648 -713 3660 -679
rect 4068 -713 4080 -679
rect -3912 -719 -3854 -713
rect -3492 -719 -3434 -713
rect -3072 -719 -3014 -713
rect -2652 -719 -2594 -713
rect -2232 -719 -2174 -713
rect -1812 -719 -1754 -713
rect -1392 -719 -1334 -713
rect -972 -719 -914 -713
rect -552 -719 -494 -713
rect -132 -719 -74 -713
rect 288 -719 346 -713
rect 708 -719 766 -713
rect 1128 -719 1186 -713
rect 1548 -719 1606 -713
rect 1968 -719 2026 -713
rect 2388 -719 2446 -713
rect 2808 -719 2866 -713
rect 3228 -719 3286 -713
rect 3648 -719 3706 -713
rect 4068 -719 4126 -713
<< nwell >>
rect -4520 -851 4520 319
<< pmos >>
rect -4320 -100 -4290 100
rect -4110 -100 -4080 100
rect -3900 -100 -3870 100
rect -3690 -100 -3660 100
rect -3480 -100 -3450 100
rect -3270 -100 -3240 100
rect -3060 -100 -3030 100
rect -2850 -100 -2820 100
rect -2640 -100 -2610 100
rect -2430 -100 -2400 100
rect -2220 -100 -2190 100
rect -2010 -100 -1980 100
rect -1800 -100 -1770 100
rect -1590 -100 -1560 100
rect -1380 -100 -1350 100
rect -1170 -100 -1140 100
rect -960 -100 -930 100
rect -750 -100 -720 100
rect -540 -100 -510 100
rect -330 -100 -300 100
rect -120 -100 -90 100
rect 90 -100 120 100
rect 300 -100 330 100
rect 510 -100 540 100
rect 720 -100 750 100
rect 930 -100 960 100
rect 1140 -100 1170 100
rect 1350 -100 1380 100
rect 1560 -100 1590 100
rect 1770 -100 1800 100
rect 1980 -100 2010 100
rect 2190 -100 2220 100
rect 2400 -100 2430 100
rect 2610 -100 2640 100
rect 2820 -100 2850 100
rect 3030 -100 3060 100
rect 3240 -100 3270 100
rect 3450 -100 3480 100
rect 3660 -100 3690 100
rect 3870 -100 3900 100
rect 4080 -100 4110 100
rect 4290 -100 4320 100
rect -4318 -632 -4288 -432
rect -4108 -632 -4078 -432
rect -3898 -632 -3868 -432
rect -3688 -632 -3658 -432
rect -3478 -632 -3448 -432
rect -3268 -632 -3238 -432
rect -3058 -632 -3028 -432
rect -2848 -632 -2818 -432
rect -2638 -632 -2608 -432
rect -2428 -632 -2398 -432
rect -2218 -632 -2188 -432
rect -2008 -632 -1978 -432
rect -1798 -632 -1768 -432
rect -1588 -632 -1558 -432
rect -1378 -632 -1348 -432
rect -1168 -632 -1138 -432
rect -958 -632 -928 -432
rect -748 -632 -718 -432
rect -538 -632 -508 -432
rect -328 -632 -298 -432
rect -118 -632 -88 -432
rect 92 -632 122 -432
rect 302 -632 332 -432
rect 512 -632 542 -432
rect 722 -632 752 -432
rect 932 -632 962 -432
rect 1142 -632 1172 -432
rect 1352 -632 1382 -432
rect 1562 -632 1592 -432
rect 1772 -632 1802 -432
rect 1982 -632 2012 -432
rect 2192 -632 2222 -432
rect 2402 -632 2432 -432
rect 2612 -632 2642 -432
rect 2822 -632 2852 -432
rect 3032 -632 3062 -432
rect 3242 -632 3272 -432
rect 3452 -632 3482 -432
rect 3662 -632 3692 -432
rect 3872 -632 3902 -432
rect 4082 -632 4112 -432
rect 4292 -632 4322 -432
<< pdiff >>
rect -4382 85 -4320 100
rect -4382 51 -4370 85
rect -4336 51 -4320 85
rect -4382 17 -4320 51
rect -4382 -17 -4370 17
rect -4336 -17 -4320 17
rect -4382 -51 -4320 -17
rect -4382 -85 -4370 -51
rect -4336 -85 -4320 -51
rect -4382 -100 -4320 -85
rect -4290 85 -4228 100
rect -4290 51 -4274 85
rect -4240 51 -4228 85
rect -4290 17 -4228 51
rect -4290 -17 -4274 17
rect -4240 -17 -4228 17
rect -4290 -51 -4228 -17
rect -4290 -85 -4274 -51
rect -4240 -85 -4228 -51
rect -4290 -100 -4228 -85
rect -4172 85 -4110 100
rect -4172 51 -4160 85
rect -4126 51 -4110 85
rect -4172 17 -4110 51
rect -4172 -17 -4160 17
rect -4126 -17 -4110 17
rect -4172 -51 -4110 -17
rect -4172 -85 -4160 -51
rect -4126 -85 -4110 -51
rect -4172 -100 -4110 -85
rect -4080 85 -4018 100
rect -4080 51 -4064 85
rect -4030 51 -4018 85
rect -4080 17 -4018 51
rect -4080 -17 -4064 17
rect -4030 -17 -4018 17
rect -4080 -51 -4018 -17
rect -4080 -85 -4064 -51
rect -4030 -85 -4018 -51
rect -4080 -100 -4018 -85
rect -3962 85 -3900 100
rect -3962 51 -3950 85
rect -3916 51 -3900 85
rect -3962 17 -3900 51
rect -3962 -17 -3950 17
rect -3916 -17 -3900 17
rect -3962 -51 -3900 -17
rect -3962 -85 -3950 -51
rect -3916 -85 -3900 -51
rect -3962 -100 -3900 -85
rect -3870 85 -3808 100
rect -3870 51 -3854 85
rect -3820 51 -3808 85
rect -3870 17 -3808 51
rect -3870 -17 -3854 17
rect -3820 -17 -3808 17
rect -3870 -51 -3808 -17
rect -3870 -85 -3854 -51
rect -3820 -85 -3808 -51
rect -3870 -100 -3808 -85
rect -3752 85 -3690 100
rect -3752 51 -3740 85
rect -3706 51 -3690 85
rect -3752 17 -3690 51
rect -3752 -17 -3740 17
rect -3706 -17 -3690 17
rect -3752 -51 -3690 -17
rect -3752 -85 -3740 -51
rect -3706 -85 -3690 -51
rect -3752 -100 -3690 -85
rect -3660 85 -3598 100
rect -3660 51 -3644 85
rect -3610 51 -3598 85
rect -3660 17 -3598 51
rect -3660 -17 -3644 17
rect -3610 -17 -3598 17
rect -3660 -51 -3598 -17
rect -3660 -85 -3644 -51
rect -3610 -85 -3598 -51
rect -3660 -100 -3598 -85
rect -3542 85 -3480 100
rect -3542 51 -3530 85
rect -3496 51 -3480 85
rect -3542 17 -3480 51
rect -3542 -17 -3530 17
rect -3496 -17 -3480 17
rect -3542 -51 -3480 -17
rect -3542 -85 -3530 -51
rect -3496 -85 -3480 -51
rect -3542 -100 -3480 -85
rect -3450 85 -3388 100
rect -3450 51 -3434 85
rect -3400 51 -3388 85
rect -3450 17 -3388 51
rect -3450 -17 -3434 17
rect -3400 -17 -3388 17
rect -3450 -51 -3388 -17
rect -3450 -85 -3434 -51
rect -3400 -85 -3388 -51
rect -3450 -100 -3388 -85
rect -3332 85 -3270 100
rect -3332 51 -3320 85
rect -3286 51 -3270 85
rect -3332 17 -3270 51
rect -3332 -17 -3320 17
rect -3286 -17 -3270 17
rect -3332 -51 -3270 -17
rect -3332 -85 -3320 -51
rect -3286 -85 -3270 -51
rect -3332 -100 -3270 -85
rect -3240 85 -3178 100
rect -3240 51 -3224 85
rect -3190 51 -3178 85
rect -3240 17 -3178 51
rect -3240 -17 -3224 17
rect -3190 -17 -3178 17
rect -3240 -51 -3178 -17
rect -3240 -85 -3224 -51
rect -3190 -85 -3178 -51
rect -3240 -100 -3178 -85
rect -3122 85 -3060 100
rect -3122 51 -3110 85
rect -3076 51 -3060 85
rect -3122 17 -3060 51
rect -3122 -17 -3110 17
rect -3076 -17 -3060 17
rect -3122 -51 -3060 -17
rect -3122 -85 -3110 -51
rect -3076 -85 -3060 -51
rect -3122 -100 -3060 -85
rect -3030 85 -2968 100
rect -3030 51 -3014 85
rect -2980 51 -2968 85
rect -3030 17 -2968 51
rect -3030 -17 -3014 17
rect -2980 -17 -2968 17
rect -3030 -51 -2968 -17
rect -3030 -85 -3014 -51
rect -2980 -85 -2968 -51
rect -3030 -100 -2968 -85
rect -2912 85 -2850 100
rect -2912 51 -2900 85
rect -2866 51 -2850 85
rect -2912 17 -2850 51
rect -2912 -17 -2900 17
rect -2866 -17 -2850 17
rect -2912 -51 -2850 -17
rect -2912 -85 -2900 -51
rect -2866 -85 -2850 -51
rect -2912 -100 -2850 -85
rect -2820 85 -2758 100
rect -2820 51 -2804 85
rect -2770 51 -2758 85
rect -2820 17 -2758 51
rect -2820 -17 -2804 17
rect -2770 -17 -2758 17
rect -2820 -51 -2758 -17
rect -2820 -85 -2804 -51
rect -2770 -85 -2758 -51
rect -2820 -100 -2758 -85
rect -2702 85 -2640 100
rect -2702 51 -2690 85
rect -2656 51 -2640 85
rect -2702 17 -2640 51
rect -2702 -17 -2690 17
rect -2656 -17 -2640 17
rect -2702 -51 -2640 -17
rect -2702 -85 -2690 -51
rect -2656 -85 -2640 -51
rect -2702 -100 -2640 -85
rect -2610 85 -2548 100
rect -2610 51 -2594 85
rect -2560 51 -2548 85
rect -2610 17 -2548 51
rect -2610 -17 -2594 17
rect -2560 -17 -2548 17
rect -2610 -51 -2548 -17
rect -2610 -85 -2594 -51
rect -2560 -85 -2548 -51
rect -2610 -100 -2548 -85
rect -2492 85 -2430 100
rect -2492 51 -2480 85
rect -2446 51 -2430 85
rect -2492 17 -2430 51
rect -2492 -17 -2480 17
rect -2446 -17 -2430 17
rect -2492 -51 -2430 -17
rect -2492 -85 -2480 -51
rect -2446 -85 -2430 -51
rect -2492 -100 -2430 -85
rect -2400 85 -2338 100
rect -2400 51 -2384 85
rect -2350 51 -2338 85
rect -2400 17 -2338 51
rect -2400 -17 -2384 17
rect -2350 -17 -2338 17
rect -2400 -51 -2338 -17
rect -2400 -85 -2384 -51
rect -2350 -85 -2338 -51
rect -2400 -100 -2338 -85
rect -2282 85 -2220 100
rect -2282 51 -2270 85
rect -2236 51 -2220 85
rect -2282 17 -2220 51
rect -2282 -17 -2270 17
rect -2236 -17 -2220 17
rect -2282 -51 -2220 -17
rect -2282 -85 -2270 -51
rect -2236 -85 -2220 -51
rect -2282 -100 -2220 -85
rect -2190 85 -2128 100
rect -2190 51 -2174 85
rect -2140 51 -2128 85
rect -2190 17 -2128 51
rect -2190 -17 -2174 17
rect -2140 -17 -2128 17
rect -2190 -51 -2128 -17
rect -2190 -85 -2174 -51
rect -2140 -85 -2128 -51
rect -2190 -100 -2128 -85
rect -2072 85 -2010 100
rect -2072 51 -2060 85
rect -2026 51 -2010 85
rect -2072 17 -2010 51
rect -2072 -17 -2060 17
rect -2026 -17 -2010 17
rect -2072 -51 -2010 -17
rect -2072 -85 -2060 -51
rect -2026 -85 -2010 -51
rect -2072 -100 -2010 -85
rect -1980 85 -1918 100
rect -1980 51 -1964 85
rect -1930 51 -1918 85
rect -1980 17 -1918 51
rect -1980 -17 -1964 17
rect -1930 -17 -1918 17
rect -1980 -51 -1918 -17
rect -1980 -85 -1964 -51
rect -1930 -85 -1918 -51
rect -1980 -100 -1918 -85
rect -1862 85 -1800 100
rect -1862 51 -1850 85
rect -1816 51 -1800 85
rect -1862 17 -1800 51
rect -1862 -17 -1850 17
rect -1816 -17 -1800 17
rect -1862 -51 -1800 -17
rect -1862 -85 -1850 -51
rect -1816 -85 -1800 -51
rect -1862 -100 -1800 -85
rect -1770 85 -1708 100
rect -1770 51 -1754 85
rect -1720 51 -1708 85
rect -1770 17 -1708 51
rect -1770 -17 -1754 17
rect -1720 -17 -1708 17
rect -1770 -51 -1708 -17
rect -1770 -85 -1754 -51
rect -1720 -85 -1708 -51
rect -1770 -100 -1708 -85
rect -1652 85 -1590 100
rect -1652 51 -1640 85
rect -1606 51 -1590 85
rect -1652 17 -1590 51
rect -1652 -17 -1640 17
rect -1606 -17 -1590 17
rect -1652 -51 -1590 -17
rect -1652 -85 -1640 -51
rect -1606 -85 -1590 -51
rect -1652 -100 -1590 -85
rect -1560 85 -1498 100
rect -1560 51 -1544 85
rect -1510 51 -1498 85
rect -1560 17 -1498 51
rect -1560 -17 -1544 17
rect -1510 -17 -1498 17
rect -1560 -51 -1498 -17
rect -1560 -85 -1544 -51
rect -1510 -85 -1498 -51
rect -1560 -100 -1498 -85
rect -1442 85 -1380 100
rect -1442 51 -1430 85
rect -1396 51 -1380 85
rect -1442 17 -1380 51
rect -1442 -17 -1430 17
rect -1396 -17 -1380 17
rect -1442 -51 -1380 -17
rect -1442 -85 -1430 -51
rect -1396 -85 -1380 -51
rect -1442 -100 -1380 -85
rect -1350 85 -1288 100
rect -1350 51 -1334 85
rect -1300 51 -1288 85
rect -1350 17 -1288 51
rect -1350 -17 -1334 17
rect -1300 -17 -1288 17
rect -1350 -51 -1288 -17
rect -1350 -85 -1334 -51
rect -1300 -85 -1288 -51
rect -1350 -100 -1288 -85
rect -1232 85 -1170 100
rect -1232 51 -1220 85
rect -1186 51 -1170 85
rect -1232 17 -1170 51
rect -1232 -17 -1220 17
rect -1186 -17 -1170 17
rect -1232 -51 -1170 -17
rect -1232 -85 -1220 -51
rect -1186 -85 -1170 -51
rect -1232 -100 -1170 -85
rect -1140 85 -1078 100
rect -1140 51 -1124 85
rect -1090 51 -1078 85
rect -1140 17 -1078 51
rect -1140 -17 -1124 17
rect -1090 -17 -1078 17
rect -1140 -51 -1078 -17
rect -1140 -85 -1124 -51
rect -1090 -85 -1078 -51
rect -1140 -100 -1078 -85
rect -1022 85 -960 100
rect -1022 51 -1010 85
rect -976 51 -960 85
rect -1022 17 -960 51
rect -1022 -17 -1010 17
rect -976 -17 -960 17
rect -1022 -51 -960 -17
rect -1022 -85 -1010 -51
rect -976 -85 -960 -51
rect -1022 -100 -960 -85
rect -930 85 -868 100
rect -930 51 -914 85
rect -880 51 -868 85
rect -930 17 -868 51
rect -930 -17 -914 17
rect -880 -17 -868 17
rect -930 -51 -868 -17
rect -930 -85 -914 -51
rect -880 -85 -868 -51
rect -930 -100 -868 -85
rect -812 85 -750 100
rect -812 51 -800 85
rect -766 51 -750 85
rect -812 17 -750 51
rect -812 -17 -800 17
rect -766 -17 -750 17
rect -812 -51 -750 -17
rect -812 -85 -800 -51
rect -766 -85 -750 -51
rect -812 -100 -750 -85
rect -720 85 -658 100
rect -720 51 -704 85
rect -670 51 -658 85
rect -720 17 -658 51
rect -720 -17 -704 17
rect -670 -17 -658 17
rect -720 -51 -658 -17
rect -720 -85 -704 -51
rect -670 -85 -658 -51
rect -720 -100 -658 -85
rect -602 85 -540 100
rect -602 51 -590 85
rect -556 51 -540 85
rect -602 17 -540 51
rect -602 -17 -590 17
rect -556 -17 -540 17
rect -602 -51 -540 -17
rect -602 -85 -590 -51
rect -556 -85 -540 -51
rect -602 -100 -540 -85
rect -510 85 -448 100
rect -510 51 -494 85
rect -460 51 -448 85
rect -510 17 -448 51
rect -510 -17 -494 17
rect -460 -17 -448 17
rect -510 -51 -448 -17
rect -510 -85 -494 -51
rect -460 -85 -448 -51
rect -510 -100 -448 -85
rect -392 85 -330 100
rect -392 51 -380 85
rect -346 51 -330 85
rect -392 17 -330 51
rect -392 -17 -380 17
rect -346 -17 -330 17
rect -392 -51 -330 -17
rect -392 -85 -380 -51
rect -346 -85 -330 -51
rect -392 -100 -330 -85
rect -300 85 -238 100
rect -300 51 -284 85
rect -250 51 -238 85
rect -300 17 -238 51
rect -300 -17 -284 17
rect -250 -17 -238 17
rect -300 -51 -238 -17
rect -300 -85 -284 -51
rect -250 -85 -238 -51
rect -300 -100 -238 -85
rect -182 85 -120 100
rect -182 51 -170 85
rect -136 51 -120 85
rect -182 17 -120 51
rect -182 -17 -170 17
rect -136 -17 -120 17
rect -182 -51 -120 -17
rect -182 -85 -170 -51
rect -136 -85 -120 -51
rect -182 -100 -120 -85
rect -90 85 -28 100
rect -90 51 -74 85
rect -40 51 -28 85
rect -90 17 -28 51
rect -90 -17 -74 17
rect -40 -17 -28 17
rect -90 -51 -28 -17
rect -90 -85 -74 -51
rect -40 -85 -28 -51
rect -90 -100 -28 -85
rect 28 85 90 100
rect 28 51 40 85
rect 74 51 90 85
rect 28 17 90 51
rect 28 -17 40 17
rect 74 -17 90 17
rect 28 -51 90 -17
rect 28 -85 40 -51
rect 74 -85 90 -51
rect 28 -100 90 -85
rect 120 85 182 100
rect 120 51 136 85
rect 170 51 182 85
rect 120 17 182 51
rect 120 -17 136 17
rect 170 -17 182 17
rect 120 -51 182 -17
rect 120 -85 136 -51
rect 170 -85 182 -51
rect 120 -100 182 -85
rect 238 85 300 100
rect 238 51 250 85
rect 284 51 300 85
rect 238 17 300 51
rect 238 -17 250 17
rect 284 -17 300 17
rect 238 -51 300 -17
rect 238 -85 250 -51
rect 284 -85 300 -51
rect 238 -100 300 -85
rect 330 85 392 100
rect 330 51 346 85
rect 380 51 392 85
rect 330 17 392 51
rect 330 -17 346 17
rect 380 -17 392 17
rect 330 -51 392 -17
rect 330 -85 346 -51
rect 380 -85 392 -51
rect 330 -100 392 -85
rect 448 85 510 100
rect 448 51 460 85
rect 494 51 510 85
rect 448 17 510 51
rect 448 -17 460 17
rect 494 -17 510 17
rect 448 -51 510 -17
rect 448 -85 460 -51
rect 494 -85 510 -51
rect 448 -100 510 -85
rect 540 85 602 100
rect 540 51 556 85
rect 590 51 602 85
rect 540 17 602 51
rect 540 -17 556 17
rect 590 -17 602 17
rect 540 -51 602 -17
rect 540 -85 556 -51
rect 590 -85 602 -51
rect 540 -100 602 -85
rect 658 85 720 100
rect 658 51 670 85
rect 704 51 720 85
rect 658 17 720 51
rect 658 -17 670 17
rect 704 -17 720 17
rect 658 -51 720 -17
rect 658 -85 670 -51
rect 704 -85 720 -51
rect 658 -100 720 -85
rect 750 85 812 100
rect 750 51 766 85
rect 800 51 812 85
rect 750 17 812 51
rect 750 -17 766 17
rect 800 -17 812 17
rect 750 -51 812 -17
rect 750 -85 766 -51
rect 800 -85 812 -51
rect 750 -100 812 -85
rect 868 85 930 100
rect 868 51 880 85
rect 914 51 930 85
rect 868 17 930 51
rect 868 -17 880 17
rect 914 -17 930 17
rect 868 -51 930 -17
rect 868 -85 880 -51
rect 914 -85 930 -51
rect 868 -100 930 -85
rect 960 85 1022 100
rect 960 51 976 85
rect 1010 51 1022 85
rect 960 17 1022 51
rect 960 -17 976 17
rect 1010 -17 1022 17
rect 960 -51 1022 -17
rect 960 -85 976 -51
rect 1010 -85 1022 -51
rect 960 -100 1022 -85
rect 1078 85 1140 100
rect 1078 51 1090 85
rect 1124 51 1140 85
rect 1078 17 1140 51
rect 1078 -17 1090 17
rect 1124 -17 1140 17
rect 1078 -51 1140 -17
rect 1078 -85 1090 -51
rect 1124 -85 1140 -51
rect 1078 -100 1140 -85
rect 1170 85 1232 100
rect 1170 51 1186 85
rect 1220 51 1232 85
rect 1170 17 1232 51
rect 1170 -17 1186 17
rect 1220 -17 1232 17
rect 1170 -51 1232 -17
rect 1170 -85 1186 -51
rect 1220 -85 1232 -51
rect 1170 -100 1232 -85
rect 1288 85 1350 100
rect 1288 51 1300 85
rect 1334 51 1350 85
rect 1288 17 1350 51
rect 1288 -17 1300 17
rect 1334 -17 1350 17
rect 1288 -51 1350 -17
rect 1288 -85 1300 -51
rect 1334 -85 1350 -51
rect 1288 -100 1350 -85
rect 1380 85 1442 100
rect 1380 51 1396 85
rect 1430 51 1442 85
rect 1380 17 1442 51
rect 1380 -17 1396 17
rect 1430 -17 1442 17
rect 1380 -51 1442 -17
rect 1380 -85 1396 -51
rect 1430 -85 1442 -51
rect 1380 -100 1442 -85
rect 1498 85 1560 100
rect 1498 51 1510 85
rect 1544 51 1560 85
rect 1498 17 1560 51
rect 1498 -17 1510 17
rect 1544 -17 1560 17
rect 1498 -51 1560 -17
rect 1498 -85 1510 -51
rect 1544 -85 1560 -51
rect 1498 -100 1560 -85
rect 1590 85 1652 100
rect 1590 51 1606 85
rect 1640 51 1652 85
rect 1590 17 1652 51
rect 1590 -17 1606 17
rect 1640 -17 1652 17
rect 1590 -51 1652 -17
rect 1590 -85 1606 -51
rect 1640 -85 1652 -51
rect 1590 -100 1652 -85
rect 1708 85 1770 100
rect 1708 51 1720 85
rect 1754 51 1770 85
rect 1708 17 1770 51
rect 1708 -17 1720 17
rect 1754 -17 1770 17
rect 1708 -51 1770 -17
rect 1708 -85 1720 -51
rect 1754 -85 1770 -51
rect 1708 -100 1770 -85
rect 1800 85 1862 100
rect 1800 51 1816 85
rect 1850 51 1862 85
rect 1800 17 1862 51
rect 1800 -17 1816 17
rect 1850 -17 1862 17
rect 1800 -51 1862 -17
rect 1800 -85 1816 -51
rect 1850 -85 1862 -51
rect 1800 -100 1862 -85
rect 1918 85 1980 100
rect 1918 51 1930 85
rect 1964 51 1980 85
rect 1918 17 1980 51
rect 1918 -17 1930 17
rect 1964 -17 1980 17
rect 1918 -51 1980 -17
rect 1918 -85 1930 -51
rect 1964 -85 1980 -51
rect 1918 -100 1980 -85
rect 2010 85 2072 100
rect 2010 51 2026 85
rect 2060 51 2072 85
rect 2010 17 2072 51
rect 2010 -17 2026 17
rect 2060 -17 2072 17
rect 2010 -51 2072 -17
rect 2010 -85 2026 -51
rect 2060 -85 2072 -51
rect 2010 -100 2072 -85
rect 2128 85 2190 100
rect 2128 51 2140 85
rect 2174 51 2190 85
rect 2128 17 2190 51
rect 2128 -17 2140 17
rect 2174 -17 2190 17
rect 2128 -51 2190 -17
rect 2128 -85 2140 -51
rect 2174 -85 2190 -51
rect 2128 -100 2190 -85
rect 2220 85 2282 100
rect 2220 51 2236 85
rect 2270 51 2282 85
rect 2220 17 2282 51
rect 2220 -17 2236 17
rect 2270 -17 2282 17
rect 2220 -51 2282 -17
rect 2220 -85 2236 -51
rect 2270 -85 2282 -51
rect 2220 -100 2282 -85
rect 2338 85 2400 100
rect 2338 51 2350 85
rect 2384 51 2400 85
rect 2338 17 2400 51
rect 2338 -17 2350 17
rect 2384 -17 2400 17
rect 2338 -51 2400 -17
rect 2338 -85 2350 -51
rect 2384 -85 2400 -51
rect 2338 -100 2400 -85
rect 2430 85 2492 100
rect 2430 51 2446 85
rect 2480 51 2492 85
rect 2430 17 2492 51
rect 2430 -17 2446 17
rect 2480 -17 2492 17
rect 2430 -51 2492 -17
rect 2430 -85 2446 -51
rect 2480 -85 2492 -51
rect 2430 -100 2492 -85
rect 2548 85 2610 100
rect 2548 51 2560 85
rect 2594 51 2610 85
rect 2548 17 2610 51
rect 2548 -17 2560 17
rect 2594 -17 2610 17
rect 2548 -51 2610 -17
rect 2548 -85 2560 -51
rect 2594 -85 2610 -51
rect 2548 -100 2610 -85
rect 2640 85 2702 100
rect 2640 51 2656 85
rect 2690 51 2702 85
rect 2640 17 2702 51
rect 2640 -17 2656 17
rect 2690 -17 2702 17
rect 2640 -51 2702 -17
rect 2640 -85 2656 -51
rect 2690 -85 2702 -51
rect 2640 -100 2702 -85
rect 2758 85 2820 100
rect 2758 51 2770 85
rect 2804 51 2820 85
rect 2758 17 2820 51
rect 2758 -17 2770 17
rect 2804 -17 2820 17
rect 2758 -51 2820 -17
rect 2758 -85 2770 -51
rect 2804 -85 2820 -51
rect 2758 -100 2820 -85
rect 2850 85 2912 100
rect 2850 51 2866 85
rect 2900 51 2912 85
rect 2850 17 2912 51
rect 2850 -17 2866 17
rect 2900 -17 2912 17
rect 2850 -51 2912 -17
rect 2850 -85 2866 -51
rect 2900 -85 2912 -51
rect 2850 -100 2912 -85
rect 2968 85 3030 100
rect 2968 51 2980 85
rect 3014 51 3030 85
rect 2968 17 3030 51
rect 2968 -17 2980 17
rect 3014 -17 3030 17
rect 2968 -51 3030 -17
rect 2968 -85 2980 -51
rect 3014 -85 3030 -51
rect 2968 -100 3030 -85
rect 3060 85 3122 100
rect 3060 51 3076 85
rect 3110 51 3122 85
rect 3060 17 3122 51
rect 3060 -17 3076 17
rect 3110 -17 3122 17
rect 3060 -51 3122 -17
rect 3060 -85 3076 -51
rect 3110 -85 3122 -51
rect 3060 -100 3122 -85
rect 3178 85 3240 100
rect 3178 51 3190 85
rect 3224 51 3240 85
rect 3178 17 3240 51
rect 3178 -17 3190 17
rect 3224 -17 3240 17
rect 3178 -51 3240 -17
rect 3178 -85 3190 -51
rect 3224 -85 3240 -51
rect 3178 -100 3240 -85
rect 3270 85 3332 100
rect 3270 51 3286 85
rect 3320 51 3332 85
rect 3270 17 3332 51
rect 3270 -17 3286 17
rect 3320 -17 3332 17
rect 3270 -51 3332 -17
rect 3270 -85 3286 -51
rect 3320 -85 3332 -51
rect 3270 -100 3332 -85
rect 3388 85 3450 100
rect 3388 51 3400 85
rect 3434 51 3450 85
rect 3388 17 3450 51
rect 3388 -17 3400 17
rect 3434 -17 3450 17
rect 3388 -51 3450 -17
rect 3388 -85 3400 -51
rect 3434 -85 3450 -51
rect 3388 -100 3450 -85
rect 3480 85 3542 100
rect 3480 51 3496 85
rect 3530 51 3542 85
rect 3480 17 3542 51
rect 3480 -17 3496 17
rect 3530 -17 3542 17
rect 3480 -51 3542 -17
rect 3480 -85 3496 -51
rect 3530 -85 3542 -51
rect 3480 -100 3542 -85
rect 3598 85 3660 100
rect 3598 51 3610 85
rect 3644 51 3660 85
rect 3598 17 3660 51
rect 3598 -17 3610 17
rect 3644 -17 3660 17
rect 3598 -51 3660 -17
rect 3598 -85 3610 -51
rect 3644 -85 3660 -51
rect 3598 -100 3660 -85
rect 3690 85 3752 100
rect 3690 51 3706 85
rect 3740 51 3752 85
rect 3690 17 3752 51
rect 3690 -17 3706 17
rect 3740 -17 3752 17
rect 3690 -51 3752 -17
rect 3690 -85 3706 -51
rect 3740 -85 3752 -51
rect 3690 -100 3752 -85
rect 3808 85 3870 100
rect 3808 51 3820 85
rect 3854 51 3870 85
rect 3808 17 3870 51
rect 3808 -17 3820 17
rect 3854 -17 3870 17
rect 3808 -51 3870 -17
rect 3808 -85 3820 -51
rect 3854 -85 3870 -51
rect 3808 -100 3870 -85
rect 3900 85 3962 100
rect 3900 51 3916 85
rect 3950 51 3962 85
rect 3900 17 3962 51
rect 3900 -17 3916 17
rect 3950 -17 3962 17
rect 3900 -51 3962 -17
rect 3900 -85 3916 -51
rect 3950 -85 3962 -51
rect 3900 -100 3962 -85
rect 4018 85 4080 100
rect 4018 51 4030 85
rect 4064 51 4080 85
rect 4018 17 4080 51
rect 4018 -17 4030 17
rect 4064 -17 4080 17
rect 4018 -51 4080 -17
rect 4018 -85 4030 -51
rect 4064 -85 4080 -51
rect 4018 -100 4080 -85
rect 4110 85 4172 100
rect 4110 51 4126 85
rect 4160 51 4172 85
rect 4110 17 4172 51
rect 4110 -17 4126 17
rect 4160 -17 4172 17
rect 4110 -51 4172 -17
rect 4110 -85 4126 -51
rect 4160 -85 4172 -51
rect 4110 -100 4172 -85
rect 4228 85 4290 100
rect 4228 51 4240 85
rect 4274 51 4290 85
rect 4228 17 4290 51
rect 4228 -17 4240 17
rect 4274 -17 4290 17
rect 4228 -51 4290 -17
rect 4228 -85 4240 -51
rect 4274 -85 4290 -51
rect 4228 -100 4290 -85
rect 4320 85 4382 100
rect 4320 51 4336 85
rect 4370 51 4382 85
rect 4320 17 4382 51
rect 4320 -17 4336 17
rect 4370 -17 4382 17
rect 4320 -51 4382 -17
rect 4320 -85 4336 -51
rect 4370 -85 4382 -51
rect 4320 -100 4382 -85
rect -4380 -447 -4318 -432
rect -4380 -481 -4368 -447
rect -4334 -481 -4318 -447
rect -4380 -515 -4318 -481
rect -4380 -549 -4368 -515
rect -4334 -549 -4318 -515
rect -4380 -583 -4318 -549
rect -4380 -617 -4368 -583
rect -4334 -617 -4318 -583
rect -4380 -632 -4318 -617
rect -4288 -447 -4226 -432
rect -4288 -481 -4272 -447
rect -4238 -481 -4226 -447
rect -4288 -515 -4226 -481
rect -4288 -549 -4272 -515
rect -4238 -549 -4226 -515
rect -4288 -583 -4226 -549
rect -4288 -617 -4272 -583
rect -4238 -617 -4226 -583
rect -4288 -632 -4226 -617
rect -4170 -447 -4108 -432
rect -4170 -481 -4158 -447
rect -4124 -481 -4108 -447
rect -4170 -515 -4108 -481
rect -4170 -549 -4158 -515
rect -4124 -549 -4108 -515
rect -4170 -583 -4108 -549
rect -4170 -617 -4158 -583
rect -4124 -617 -4108 -583
rect -4170 -632 -4108 -617
rect -4078 -447 -4016 -432
rect -4078 -481 -4062 -447
rect -4028 -481 -4016 -447
rect -4078 -515 -4016 -481
rect -4078 -549 -4062 -515
rect -4028 -549 -4016 -515
rect -4078 -583 -4016 -549
rect -4078 -617 -4062 -583
rect -4028 -617 -4016 -583
rect -4078 -632 -4016 -617
rect -3960 -447 -3898 -432
rect -3960 -481 -3948 -447
rect -3914 -481 -3898 -447
rect -3960 -515 -3898 -481
rect -3960 -549 -3948 -515
rect -3914 -549 -3898 -515
rect -3960 -583 -3898 -549
rect -3960 -617 -3948 -583
rect -3914 -617 -3898 -583
rect -3960 -632 -3898 -617
rect -3868 -447 -3806 -432
rect -3868 -481 -3852 -447
rect -3818 -481 -3806 -447
rect -3868 -515 -3806 -481
rect -3868 -549 -3852 -515
rect -3818 -549 -3806 -515
rect -3868 -583 -3806 -549
rect -3868 -617 -3852 -583
rect -3818 -617 -3806 -583
rect -3868 -632 -3806 -617
rect -3750 -447 -3688 -432
rect -3750 -481 -3738 -447
rect -3704 -481 -3688 -447
rect -3750 -515 -3688 -481
rect -3750 -549 -3738 -515
rect -3704 -549 -3688 -515
rect -3750 -583 -3688 -549
rect -3750 -617 -3738 -583
rect -3704 -617 -3688 -583
rect -3750 -632 -3688 -617
rect -3658 -447 -3596 -432
rect -3658 -481 -3642 -447
rect -3608 -481 -3596 -447
rect -3658 -515 -3596 -481
rect -3658 -549 -3642 -515
rect -3608 -549 -3596 -515
rect -3658 -583 -3596 -549
rect -3658 -617 -3642 -583
rect -3608 -617 -3596 -583
rect -3658 -632 -3596 -617
rect -3540 -447 -3478 -432
rect -3540 -481 -3528 -447
rect -3494 -481 -3478 -447
rect -3540 -515 -3478 -481
rect -3540 -549 -3528 -515
rect -3494 -549 -3478 -515
rect -3540 -583 -3478 -549
rect -3540 -617 -3528 -583
rect -3494 -617 -3478 -583
rect -3540 -632 -3478 -617
rect -3448 -447 -3386 -432
rect -3448 -481 -3432 -447
rect -3398 -481 -3386 -447
rect -3448 -515 -3386 -481
rect -3448 -549 -3432 -515
rect -3398 -549 -3386 -515
rect -3448 -583 -3386 -549
rect -3448 -617 -3432 -583
rect -3398 -617 -3386 -583
rect -3448 -632 -3386 -617
rect -3330 -447 -3268 -432
rect -3330 -481 -3318 -447
rect -3284 -481 -3268 -447
rect -3330 -515 -3268 -481
rect -3330 -549 -3318 -515
rect -3284 -549 -3268 -515
rect -3330 -583 -3268 -549
rect -3330 -617 -3318 -583
rect -3284 -617 -3268 -583
rect -3330 -632 -3268 -617
rect -3238 -447 -3176 -432
rect -3238 -481 -3222 -447
rect -3188 -481 -3176 -447
rect -3238 -515 -3176 -481
rect -3238 -549 -3222 -515
rect -3188 -549 -3176 -515
rect -3238 -583 -3176 -549
rect -3238 -617 -3222 -583
rect -3188 -617 -3176 -583
rect -3238 -632 -3176 -617
rect -3120 -447 -3058 -432
rect -3120 -481 -3108 -447
rect -3074 -481 -3058 -447
rect -3120 -515 -3058 -481
rect -3120 -549 -3108 -515
rect -3074 -549 -3058 -515
rect -3120 -583 -3058 -549
rect -3120 -617 -3108 -583
rect -3074 -617 -3058 -583
rect -3120 -632 -3058 -617
rect -3028 -447 -2966 -432
rect -3028 -481 -3012 -447
rect -2978 -481 -2966 -447
rect -3028 -515 -2966 -481
rect -3028 -549 -3012 -515
rect -2978 -549 -2966 -515
rect -3028 -583 -2966 -549
rect -3028 -617 -3012 -583
rect -2978 -617 -2966 -583
rect -3028 -632 -2966 -617
rect -2910 -447 -2848 -432
rect -2910 -481 -2898 -447
rect -2864 -481 -2848 -447
rect -2910 -515 -2848 -481
rect -2910 -549 -2898 -515
rect -2864 -549 -2848 -515
rect -2910 -583 -2848 -549
rect -2910 -617 -2898 -583
rect -2864 -617 -2848 -583
rect -2910 -632 -2848 -617
rect -2818 -447 -2756 -432
rect -2818 -481 -2802 -447
rect -2768 -481 -2756 -447
rect -2818 -515 -2756 -481
rect -2818 -549 -2802 -515
rect -2768 -549 -2756 -515
rect -2818 -583 -2756 -549
rect -2818 -617 -2802 -583
rect -2768 -617 -2756 -583
rect -2818 -632 -2756 -617
rect -2700 -447 -2638 -432
rect -2700 -481 -2688 -447
rect -2654 -481 -2638 -447
rect -2700 -515 -2638 -481
rect -2700 -549 -2688 -515
rect -2654 -549 -2638 -515
rect -2700 -583 -2638 -549
rect -2700 -617 -2688 -583
rect -2654 -617 -2638 -583
rect -2700 -632 -2638 -617
rect -2608 -447 -2546 -432
rect -2608 -481 -2592 -447
rect -2558 -481 -2546 -447
rect -2608 -515 -2546 -481
rect -2608 -549 -2592 -515
rect -2558 -549 -2546 -515
rect -2608 -583 -2546 -549
rect -2608 -617 -2592 -583
rect -2558 -617 -2546 -583
rect -2608 -632 -2546 -617
rect -2490 -447 -2428 -432
rect -2490 -481 -2478 -447
rect -2444 -481 -2428 -447
rect -2490 -515 -2428 -481
rect -2490 -549 -2478 -515
rect -2444 -549 -2428 -515
rect -2490 -583 -2428 -549
rect -2490 -617 -2478 -583
rect -2444 -617 -2428 -583
rect -2490 -632 -2428 -617
rect -2398 -447 -2336 -432
rect -2398 -481 -2382 -447
rect -2348 -481 -2336 -447
rect -2398 -515 -2336 -481
rect -2398 -549 -2382 -515
rect -2348 -549 -2336 -515
rect -2398 -583 -2336 -549
rect -2398 -617 -2382 -583
rect -2348 -617 -2336 -583
rect -2398 -632 -2336 -617
rect -2280 -447 -2218 -432
rect -2280 -481 -2268 -447
rect -2234 -481 -2218 -447
rect -2280 -515 -2218 -481
rect -2280 -549 -2268 -515
rect -2234 -549 -2218 -515
rect -2280 -583 -2218 -549
rect -2280 -617 -2268 -583
rect -2234 -617 -2218 -583
rect -2280 -632 -2218 -617
rect -2188 -447 -2126 -432
rect -2188 -481 -2172 -447
rect -2138 -481 -2126 -447
rect -2188 -515 -2126 -481
rect -2188 -549 -2172 -515
rect -2138 -549 -2126 -515
rect -2188 -583 -2126 -549
rect -2188 -617 -2172 -583
rect -2138 -617 -2126 -583
rect -2188 -632 -2126 -617
rect -2070 -447 -2008 -432
rect -2070 -481 -2058 -447
rect -2024 -481 -2008 -447
rect -2070 -515 -2008 -481
rect -2070 -549 -2058 -515
rect -2024 -549 -2008 -515
rect -2070 -583 -2008 -549
rect -2070 -617 -2058 -583
rect -2024 -617 -2008 -583
rect -2070 -632 -2008 -617
rect -1978 -447 -1916 -432
rect -1978 -481 -1962 -447
rect -1928 -481 -1916 -447
rect -1978 -515 -1916 -481
rect -1978 -549 -1962 -515
rect -1928 -549 -1916 -515
rect -1978 -583 -1916 -549
rect -1978 -617 -1962 -583
rect -1928 -617 -1916 -583
rect -1978 -632 -1916 -617
rect -1860 -447 -1798 -432
rect -1860 -481 -1848 -447
rect -1814 -481 -1798 -447
rect -1860 -515 -1798 -481
rect -1860 -549 -1848 -515
rect -1814 -549 -1798 -515
rect -1860 -583 -1798 -549
rect -1860 -617 -1848 -583
rect -1814 -617 -1798 -583
rect -1860 -632 -1798 -617
rect -1768 -447 -1706 -432
rect -1768 -481 -1752 -447
rect -1718 -481 -1706 -447
rect -1768 -515 -1706 -481
rect -1768 -549 -1752 -515
rect -1718 -549 -1706 -515
rect -1768 -583 -1706 -549
rect -1768 -617 -1752 -583
rect -1718 -617 -1706 -583
rect -1768 -632 -1706 -617
rect -1650 -447 -1588 -432
rect -1650 -481 -1638 -447
rect -1604 -481 -1588 -447
rect -1650 -515 -1588 -481
rect -1650 -549 -1638 -515
rect -1604 -549 -1588 -515
rect -1650 -583 -1588 -549
rect -1650 -617 -1638 -583
rect -1604 -617 -1588 -583
rect -1650 -632 -1588 -617
rect -1558 -447 -1496 -432
rect -1558 -481 -1542 -447
rect -1508 -481 -1496 -447
rect -1558 -515 -1496 -481
rect -1558 -549 -1542 -515
rect -1508 -549 -1496 -515
rect -1558 -583 -1496 -549
rect -1558 -617 -1542 -583
rect -1508 -617 -1496 -583
rect -1558 -632 -1496 -617
rect -1440 -447 -1378 -432
rect -1440 -481 -1428 -447
rect -1394 -481 -1378 -447
rect -1440 -515 -1378 -481
rect -1440 -549 -1428 -515
rect -1394 -549 -1378 -515
rect -1440 -583 -1378 -549
rect -1440 -617 -1428 -583
rect -1394 -617 -1378 -583
rect -1440 -632 -1378 -617
rect -1348 -447 -1286 -432
rect -1348 -481 -1332 -447
rect -1298 -481 -1286 -447
rect -1348 -515 -1286 -481
rect -1348 -549 -1332 -515
rect -1298 -549 -1286 -515
rect -1348 -583 -1286 -549
rect -1348 -617 -1332 -583
rect -1298 -617 -1286 -583
rect -1348 -632 -1286 -617
rect -1230 -447 -1168 -432
rect -1230 -481 -1218 -447
rect -1184 -481 -1168 -447
rect -1230 -515 -1168 -481
rect -1230 -549 -1218 -515
rect -1184 -549 -1168 -515
rect -1230 -583 -1168 -549
rect -1230 -617 -1218 -583
rect -1184 -617 -1168 -583
rect -1230 -632 -1168 -617
rect -1138 -447 -1076 -432
rect -1138 -481 -1122 -447
rect -1088 -481 -1076 -447
rect -1138 -515 -1076 -481
rect -1138 -549 -1122 -515
rect -1088 -549 -1076 -515
rect -1138 -583 -1076 -549
rect -1138 -617 -1122 -583
rect -1088 -617 -1076 -583
rect -1138 -632 -1076 -617
rect -1020 -447 -958 -432
rect -1020 -481 -1008 -447
rect -974 -481 -958 -447
rect -1020 -515 -958 -481
rect -1020 -549 -1008 -515
rect -974 -549 -958 -515
rect -1020 -583 -958 -549
rect -1020 -617 -1008 -583
rect -974 -617 -958 -583
rect -1020 -632 -958 -617
rect -928 -447 -866 -432
rect -928 -481 -912 -447
rect -878 -481 -866 -447
rect -928 -515 -866 -481
rect -928 -549 -912 -515
rect -878 -549 -866 -515
rect -928 -583 -866 -549
rect -928 -617 -912 -583
rect -878 -617 -866 -583
rect -928 -632 -866 -617
rect -810 -447 -748 -432
rect -810 -481 -798 -447
rect -764 -481 -748 -447
rect -810 -515 -748 -481
rect -810 -549 -798 -515
rect -764 -549 -748 -515
rect -810 -583 -748 -549
rect -810 -617 -798 -583
rect -764 -617 -748 -583
rect -810 -632 -748 -617
rect -718 -447 -656 -432
rect -718 -481 -702 -447
rect -668 -481 -656 -447
rect -718 -515 -656 -481
rect -718 -549 -702 -515
rect -668 -549 -656 -515
rect -718 -583 -656 -549
rect -718 -617 -702 -583
rect -668 -617 -656 -583
rect -718 -632 -656 -617
rect -600 -447 -538 -432
rect -600 -481 -588 -447
rect -554 -481 -538 -447
rect -600 -515 -538 -481
rect -600 -549 -588 -515
rect -554 -549 -538 -515
rect -600 -583 -538 -549
rect -600 -617 -588 -583
rect -554 -617 -538 -583
rect -600 -632 -538 -617
rect -508 -447 -446 -432
rect -508 -481 -492 -447
rect -458 -481 -446 -447
rect -508 -515 -446 -481
rect -508 -549 -492 -515
rect -458 -549 -446 -515
rect -508 -583 -446 -549
rect -508 -617 -492 -583
rect -458 -617 -446 -583
rect -508 -632 -446 -617
rect -390 -447 -328 -432
rect -390 -481 -378 -447
rect -344 -481 -328 -447
rect -390 -515 -328 -481
rect -390 -549 -378 -515
rect -344 -549 -328 -515
rect -390 -583 -328 -549
rect -390 -617 -378 -583
rect -344 -617 -328 -583
rect -390 -632 -328 -617
rect -298 -447 -236 -432
rect -298 -481 -282 -447
rect -248 -481 -236 -447
rect -298 -515 -236 -481
rect -298 -549 -282 -515
rect -248 -549 -236 -515
rect -298 -583 -236 -549
rect -298 -617 -282 -583
rect -248 -617 -236 -583
rect -298 -632 -236 -617
rect -180 -447 -118 -432
rect -180 -481 -168 -447
rect -134 -481 -118 -447
rect -180 -515 -118 -481
rect -180 -549 -168 -515
rect -134 -549 -118 -515
rect -180 -583 -118 -549
rect -180 -617 -168 -583
rect -134 -617 -118 -583
rect -180 -632 -118 -617
rect -88 -447 -26 -432
rect -88 -481 -72 -447
rect -38 -481 -26 -447
rect -88 -515 -26 -481
rect -88 -549 -72 -515
rect -38 -549 -26 -515
rect -88 -583 -26 -549
rect -88 -617 -72 -583
rect -38 -617 -26 -583
rect -88 -632 -26 -617
rect 30 -447 92 -432
rect 30 -481 42 -447
rect 76 -481 92 -447
rect 30 -515 92 -481
rect 30 -549 42 -515
rect 76 -549 92 -515
rect 30 -583 92 -549
rect 30 -617 42 -583
rect 76 -617 92 -583
rect 30 -632 92 -617
rect 122 -447 184 -432
rect 122 -481 138 -447
rect 172 -481 184 -447
rect 122 -515 184 -481
rect 122 -549 138 -515
rect 172 -549 184 -515
rect 122 -583 184 -549
rect 122 -617 138 -583
rect 172 -617 184 -583
rect 122 -632 184 -617
rect 240 -447 302 -432
rect 240 -481 252 -447
rect 286 -481 302 -447
rect 240 -515 302 -481
rect 240 -549 252 -515
rect 286 -549 302 -515
rect 240 -583 302 -549
rect 240 -617 252 -583
rect 286 -617 302 -583
rect 240 -632 302 -617
rect 332 -447 394 -432
rect 332 -481 348 -447
rect 382 -481 394 -447
rect 332 -515 394 -481
rect 332 -549 348 -515
rect 382 -549 394 -515
rect 332 -583 394 -549
rect 332 -617 348 -583
rect 382 -617 394 -583
rect 332 -632 394 -617
rect 450 -447 512 -432
rect 450 -481 462 -447
rect 496 -481 512 -447
rect 450 -515 512 -481
rect 450 -549 462 -515
rect 496 -549 512 -515
rect 450 -583 512 -549
rect 450 -617 462 -583
rect 496 -617 512 -583
rect 450 -632 512 -617
rect 542 -447 604 -432
rect 542 -481 558 -447
rect 592 -481 604 -447
rect 542 -515 604 -481
rect 542 -549 558 -515
rect 592 -549 604 -515
rect 542 -583 604 -549
rect 542 -617 558 -583
rect 592 -617 604 -583
rect 542 -632 604 -617
rect 660 -447 722 -432
rect 660 -481 672 -447
rect 706 -481 722 -447
rect 660 -515 722 -481
rect 660 -549 672 -515
rect 706 -549 722 -515
rect 660 -583 722 -549
rect 660 -617 672 -583
rect 706 -617 722 -583
rect 660 -632 722 -617
rect 752 -447 814 -432
rect 752 -481 768 -447
rect 802 -481 814 -447
rect 752 -515 814 -481
rect 752 -549 768 -515
rect 802 -549 814 -515
rect 752 -583 814 -549
rect 752 -617 768 -583
rect 802 -617 814 -583
rect 752 -632 814 -617
rect 870 -447 932 -432
rect 870 -481 882 -447
rect 916 -481 932 -447
rect 870 -515 932 -481
rect 870 -549 882 -515
rect 916 -549 932 -515
rect 870 -583 932 -549
rect 870 -617 882 -583
rect 916 -617 932 -583
rect 870 -632 932 -617
rect 962 -447 1024 -432
rect 962 -481 978 -447
rect 1012 -481 1024 -447
rect 962 -515 1024 -481
rect 962 -549 978 -515
rect 1012 -549 1024 -515
rect 962 -583 1024 -549
rect 962 -617 978 -583
rect 1012 -617 1024 -583
rect 962 -632 1024 -617
rect 1080 -447 1142 -432
rect 1080 -481 1092 -447
rect 1126 -481 1142 -447
rect 1080 -515 1142 -481
rect 1080 -549 1092 -515
rect 1126 -549 1142 -515
rect 1080 -583 1142 -549
rect 1080 -617 1092 -583
rect 1126 -617 1142 -583
rect 1080 -632 1142 -617
rect 1172 -447 1234 -432
rect 1172 -481 1188 -447
rect 1222 -481 1234 -447
rect 1172 -515 1234 -481
rect 1172 -549 1188 -515
rect 1222 -549 1234 -515
rect 1172 -583 1234 -549
rect 1172 -617 1188 -583
rect 1222 -617 1234 -583
rect 1172 -632 1234 -617
rect 1290 -447 1352 -432
rect 1290 -481 1302 -447
rect 1336 -481 1352 -447
rect 1290 -515 1352 -481
rect 1290 -549 1302 -515
rect 1336 -549 1352 -515
rect 1290 -583 1352 -549
rect 1290 -617 1302 -583
rect 1336 -617 1352 -583
rect 1290 -632 1352 -617
rect 1382 -447 1444 -432
rect 1382 -481 1398 -447
rect 1432 -481 1444 -447
rect 1382 -515 1444 -481
rect 1382 -549 1398 -515
rect 1432 -549 1444 -515
rect 1382 -583 1444 -549
rect 1382 -617 1398 -583
rect 1432 -617 1444 -583
rect 1382 -632 1444 -617
rect 1500 -447 1562 -432
rect 1500 -481 1512 -447
rect 1546 -481 1562 -447
rect 1500 -515 1562 -481
rect 1500 -549 1512 -515
rect 1546 -549 1562 -515
rect 1500 -583 1562 -549
rect 1500 -617 1512 -583
rect 1546 -617 1562 -583
rect 1500 -632 1562 -617
rect 1592 -447 1654 -432
rect 1592 -481 1608 -447
rect 1642 -481 1654 -447
rect 1592 -515 1654 -481
rect 1592 -549 1608 -515
rect 1642 -549 1654 -515
rect 1592 -583 1654 -549
rect 1592 -617 1608 -583
rect 1642 -617 1654 -583
rect 1592 -632 1654 -617
rect 1710 -447 1772 -432
rect 1710 -481 1722 -447
rect 1756 -481 1772 -447
rect 1710 -515 1772 -481
rect 1710 -549 1722 -515
rect 1756 -549 1772 -515
rect 1710 -583 1772 -549
rect 1710 -617 1722 -583
rect 1756 -617 1772 -583
rect 1710 -632 1772 -617
rect 1802 -447 1864 -432
rect 1802 -481 1818 -447
rect 1852 -481 1864 -447
rect 1802 -515 1864 -481
rect 1802 -549 1818 -515
rect 1852 -549 1864 -515
rect 1802 -583 1864 -549
rect 1802 -617 1818 -583
rect 1852 -617 1864 -583
rect 1802 -632 1864 -617
rect 1920 -447 1982 -432
rect 1920 -481 1932 -447
rect 1966 -481 1982 -447
rect 1920 -515 1982 -481
rect 1920 -549 1932 -515
rect 1966 -549 1982 -515
rect 1920 -583 1982 -549
rect 1920 -617 1932 -583
rect 1966 -617 1982 -583
rect 1920 -632 1982 -617
rect 2012 -447 2074 -432
rect 2012 -481 2028 -447
rect 2062 -481 2074 -447
rect 2012 -515 2074 -481
rect 2012 -549 2028 -515
rect 2062 -549 2074 -515
rect 2012 -583 2074 -549
rect 2012 -617 2028 -583
rect 2062 -617 2074 -583
rect 2012 -632 2074 -617
rect 2130 -447 2192 -432
rect 2130 -481 2142 -447
rect 2176 -481 2192 -447
rect 2130 -515 2192 -481
rect 2130 -549 2142 -515
rect 2176 -549 2192 -515
rect 2130 -583 2192 -549
rect 2130 -617 2142 -583
rect 2176 -617 2192 -583
rect 2130 -632 2192 -617
rect 2222 -447 2284 -432
rect 2222 -481 2238 -447
rect 2272 -481 2284 -447
rect 2222 -515 2284 -481
rect 2222 -549 2238 -515
rect 2272 -549 2284 -515
rect 2222 -583 2284 -549
rect 2222 -617 2238 -583
rect 2272 -617 2284 -583
rect 2222 -632 2284 -617
rect 2340 -447 2402 -432
rect 2340 -481 2352 -447
rect 2386 -481 2402 -447
rect 2340 -515 2402 -481
rect 2340 -549 2352 -515
rect 2386 -549 2402 -515
rect 2340 -583 2402 -549
rect 2340 -617 2352 -583
rect 2386 -617 2402 -583
rect 2340 -632 2402 -617
rect 2432 -447 2494 -432
rect 2432 -481 2448 -447
rect 2482 -481 2494 -447
rect 2432 -515 2494 -481
rect 2432 -549 2448 -515
rect 2482 -549 2494 -515
rect 2432 -583 2494 -549
rect 2432 -617 2448 -583
rect 2482 -617 2494 -583
rect 2432 -632 2494 -617
rect 2550 -447 2612 -432
rect 2550 -481 2562 -447
rect 2596 -481 2612 -447
rect 2550 -515 2612 -481
rect 2550 -549 2562 -515
rect 2596 -549 2612 -515
rect 2550 -583 2612 -549
rect 2550 -617 2562 -583
rect 2596 -617 2612 -583
rect 2550 -632 2612 -617
rect 2642 -447 2704 -432
rect 2642 -481 2658 -447
rect 2692 -481 2704 -447
rect 2642 -515 2704 -481
rect 2642 -549 2658 -515
rect 2692 -549 2704 -515
rect 2642 -583 2704 -549
rect 2642 -617 2658 -583
rect 2692 -617 2704 -583
rect 2642 -632 2704 -617
rect 2760 -447 2822 -432
rect 2760 -481 2772 -447
rect 2806 -481 2822 -447
rect 2760 -515 2822 -481
rect 2760 -549 2772 -515
rect 2806 -549 2822 -515
rect 2760 -583 2822 -549
rect 2760 -617 2772 -583
rect 2806 -617 2822 -583
rect 2760 -632 2822 -617
rect 2852 -447 2914 -432
rect 2852 -481 2868 -447
rect 2902 -481 2914 -447
rect 2852 -515 2914 -481
rect 2852 -549 2868 -515
rect 2902 -549 2914 -515
rect 2852 -583 2914 -549
rect 2852 -617 2868 -583
rect 2902 -617 2914 -583
rect 2852 -632 2914 -617
rect 2970 -447 3032 -432
rect 2970 -481 2982 -447
rect 3016 -481 3032 -447
rect 2970 -515 3032 -481
rect 2970 -549 2982 -515
rect 3016 -549 3032 -515
rect 2970 -583 3032 -549
rect 2970 -617 2982 -583
rect 3016 -617 3032 -583
rect 2970 -632 3032 -617
rect 3062 -447 3124 -432
rect 3062 -481 3078 -447
rect 3112 -481 3124 -447
rect 3062 -515 3124 -481
rect 3062 -549 3078 -515
rect 3112 -549 3124 -515
rect 3062 -583 3124 -549
rect 3062 -617 3078 -583
rect 3112 -617 3124 -583
rect 3062 -632 3124 -617
rect 3180 -447 3242 -432
rect 3180 -481 3192 -447
rect 3226 -481 3242 -447
rect 3180 -515 3242 -481
rect 3180 -549 3192 -515
rect 3226 -549 3242 -515
rect 3180 -583 3242 -549
rect 3180 -617 3192 -583
rect 3226 -617 3242 -583
rect 3180 -632 3242 -617
rect 3272 -447 3334 -432
rect 3272 -481 3288 -447
rect 3322 -481 3334 -447
rect 3272 -515 3334 -481
rect 3272 -549 3288 -515
rect 3322 -549 3334 -515
rect 3272 -583 3334 -549
rect 3272 -617 3288 -583
rect 3322 -617 3334 -583
rect 3272 -632 3334 -617
rect 3390 -447 3452 -432
rect 3390 -481 3402 -447
rect 3436 -481 3452 -447
rect 3390 -515 3452 -481
rect 3390 -549 3402 -515
rect 3436 -549 3452 -515
rect 3390 -583 3452 -549
rect 3390 -617 3402 -583
rect 3436 -617 3452 -583
rect 3390 -632 3452 -617
rect 3482 -447 3544 -432
rect 3482 -481 3498 -447
rect 3532 -481 3544 -447
rect 3482 -515 3544 -481
rect 3482 -549 3498 -515
rect 3532 -549 3544 -515
rect 3482 -583 3544 -549
rect 3482 -617 3498 -583
rect 3532 -617 3544 -583
rect 3482 -632 3544 -617
rect 3600 -447 3662 -432
rect 3600 -481 3612 -447
rect 3646 -481 3662 -447
rect 3600 -515 3662 -481
rect 3600 -549 3612 -515
rect 3646 -549 3662 -515
rect 3600 -583 3662 -549
rect 3600 -617 3612 -583
rect 3646 -617 3662 -583
rect 3600 -632 3662 -617
rect 3692 -447 3754 -432
rect 3692 -481 3708 -447
rect 3742 -481 3754 -447
rect 3692 -515 3754 -481
rect 3692 -549 3708 -515
rect 3742 -549 3754 -515
rect 3692 -583 3754 -549
rect 3692 -617 3708 -583
rect 3742 -617 3754 -583
rect 3692 -632 3754 -617
rect 3810 -447 3872 -432
rect 3810 -481 3822 -447
rect 3856 -481 3872 -447
rect 3810 -515 3872 -481
rect 3810 -549 3822 -515
rect 3856 -549 3872 -515
rect 3810 -583 3872 -549
rect 3810 -617 3822 -583
rect 3856 -617 3872 -583
rect 3810 -632 3872 -617
rect 3902 -447 3964 -432
rect 3902 -481 3918 -447
rect 3952 -481 3964 -447
rect 3902 -515 3964 -481
rect 3902 -549 3918 -515
rect 3952 -549 3964 -515
rect 3902 -583 3964 -549
rect 3902 -617 3918 -583
rect 3952 -617 3964 -583
rect 3902 -632 3964 -617
rect 4020 -447 4082 -432
rect 4020 -481 4032 -447
rect 4066 -481 4082 -447
rect 4020 -515 4082 -481
rect 4020 -549 4032 -515
rect 4066 -549 4082 -515
rect 4020 -583 4082 -549
rect 4020 -617 4032 -583
rect 4066 -617 4082 -583
rect 4020 -632 4082 -617
rect 4112 -447 4174 -432
rect 4112 -481 4128 -447
rect 4162 -481 4174 -447
rect 4112 -515 4174 -481
rect 4112 -549 4128 -515
rect 4162 -549 4174 -515
rect 4112 -583 4174 -549
rect 4112 -617 4128 -583
rect 4162 -617 4174 -583
rect 4112 -632 4174 -617
rect 4230 -447 4292 -432
rect 4230 -481 4242 -447
rect 4276 -481 4292 -447
rect 4230 -515 4292 -481
rect 4230 -549 4242 -515
rect 4276 -549 4292 -515
rect 4230 -583 4292 -549
rect 4230 -617 4242 -583
rect 4276 -617 4292 -583
rect 4230 -632 4292 -617
rect 4322 -447 4384 -432
rect 4322 -481 4338 -447
rect 4372 -481 4384 -447
rect 4322 -515 4384 -481
rect 4322 -549 4338 -515
rect 4372 -549 4384 -515
rect 4322 -583 4384 -549
rect 4322 -617 4338 -583
rect 4372 -617 4384 -583
rect 4322 -632 4384 -617
<< pdiffc >>
rect -4370 51 -4336 85
rect -4370 -17 -4336 17
rect -4370 -85 -4336 -51
rect -4274 51 -4240 85
rect -4274 -17 -4240 17
rect -4274 -85 -4240 -51
rect -4160 51 -4126 85
rect -4160 -17 -4126 17
rect -4160 -85 -4126 -51
rect -4064 51 -4030 85
rect -4064 -17 -4030 17
rect -4064 -85 -4030 -51
rect -3950 51 -3916 85
rect -3950 -17 -3916 17
rect -3950 -85 -3916 -51
rect -3854 51 -3820 85
rect -3854 -17 -3820 17
rect -3854 -85 -3820 -51
rect -3740 51 -3706 85
rect -3740 -17 -3706 17
rect -3740 -85 -3706 -51
rect -3644 51 -3610 85
rect -3644 -17 -3610 17
rect -3644 -85 -3610 -51
rect -3530 51 -3496 85
rect -3530 -17 -3496 17
rect -3530 -85 -3496 -51
rect -3434 51 -3400 85
rect -3434 -17 -3400 17
rect -3434 -85 -3400 -51
rect -3320 51 -3286 85
rect -3320 -17 -3286 17
rect -3320 -85 -3286 -51
rect -3224 51 -3190 85
rect -3224 -17 -3190 17
rect -3224 -85 -3190 -51
rect -3110 51 -3076 85
rect -3110 -17 -3076 17
rect -3110 -85 -3076 -51
rect -3014 51 -2980 85
rect -3014 -17 -2980 17
rect -3014 -85 -2980 -51
rect -2900 51 -2866 85
rect -2900 -17 -2866 17
rect -2900 -85 -2866 -51
rect -2804 51 -2770 85
rect -2804 -17 -2770 17
rect -2804 -85 -2770 -51
rect -2690 51 -2656 85
rect -2690 -17 -2656 17
rect -2690 -85 -2656 -51
rect -2594 51 -2560 85
rect -2594 -17 -2560 17
rect -2594 -85 -2560 -51
rect -2480 51 -2446 85
rect -2480 -17 -2446 17
rect -2480 -85 -2446 -51
rect -2384 51 -2350 85
rect -2384 -17 -2350 17
rect -2384 -85 -2350 -51
rect -2270 51 -2236 85
rect -2270 -17 -2236 17
rect -2270 -85 -2236 -51
rect -2174 51 -2140 85
rect -2174 -17 -2140 17
rect -2174 -85 -2140 -51
rect -2060 51 -2026 85
rect -2060 -17 -2026 17
rect -2060 -85 -2026 -51
rect -1964 51 -1930 85
rect -1964 -17 -1930 17
rect -1964 -85 -1930 -51
rect -1850 51 -1816 85
rect -1850 -17 -1816 17
rect -1850 -85 -1816 -51
rect -1754 51 -1720 85
rect -1754 -17 -1720 17
rect -1754 -85 -1720 -51
rect -1640 51 -1606 85
rect -1640 -17 -1606 17
rect -1640 -85 -1606 -51
rect -1544 51 -1510 85
rect -1544 -17 -1510 17
rect -1544 -85 -1510 -51
rect -1430 51 -1396 85
rect -1430 -17 -1396 17
rect -1430 -85 -1396 -51
rect -1334 51 -1300 85
rect -1334 -17 -1300 17
rect -1334 -85 -1300 -51
rect -1220 51 -1186 85
rect -1220 -17 -1186 17
rect -1220 -85 -1186 -51
rect -1124 51 -1090 85
rect -1124 -17 -1090 17
rect -1124 -85 -1090 -51
rect -1010 51 -976 85
rect -1010 -17 -976 17
rect -1010 -85 -976 -51
rect -914 51 -880 85
rect -914 -17 -880 17
rect -914 -85 -880 -51
rect -800 51 -766 85
rect -800 -17 -766 17
rect -800 -85 -766 -51
rect -704 51 -670 85
rect -704 -17 -670 17
rect -704 -85 -670 -51
rect -590 51 -556 85
rect -590 -17 -556 17
rect -590 -85 -556 -51
rect -494 51 -460 85
rect -494 -17 -460 17
rect -494 -85 -460 -51
rect -380 51 -346 85
rect -380 -17 -346 17
rect -380 -85 -346 -51
rect -284 51 -250 85
rect -284 -17 -250 17
rect -284 -85 -250 -51
rect -170 51 -136 85
rect -170 -17 -136 17
rect -170 -85 -136 -51
rect -74 51 -40 85
rect -74 -17 -40 17
rect -74 -85 -40 -51
rect 40 51 74 85
rect 40 -17 74 17
rect 40 -85 74 -51
rect 136 51 170 85
rect 136 -17 170 17
rect 136 -85 170 -51
rect 250 51 284 85
rect 250 -17 284 17
rect 250 -85 284 -51
rect 346 51 380 85
rect 346 -17 380 17
rect 346 -85 380 -51
rect 460 51 494 85
rect 460 -17 494 17
rect 460 -85 494 -51
rect 556 51 590 85
rect 556 -17 590 17
rect 556 -85 590 -51
rect 670 51 704 85
rect 670 -17 704 17
rect 670 -85 704 -51
rect 766 51 800 85
rect 766 -17 800 17
rect 766 -85 800 -51
rect 880 51 914 85
rect 880 -17 914 17
rect 880 -85 914 -51
rect 976 51 1010 85
rect 976 -17 1010 17
rect 976 -85 1010 -51
rect 1090 51 1124 85
rect 1090 -17 1124 17
rect 1090 -85 1124 -51
rect 1186 51 1220 85
rect 1186 -17 1220 17
rect 1186 -85 1220 -51
rect 1300 51 1334 85
rect 1300 -17 1334 17
rect 1300 -85 1334 -51
rect 1396 51 1430 85
rect 1396 -17 1430 17
rect 1396 -85 1430 -51
rect 1510 51 1544 85
rect 1510 -17 1544 17
rect 1510 -85 1544 -51
rect 1606 51 1640 85
rect 1606 -17 1640 17
rect 1606 -85 1640 -51
rect 1720 51 1754 85
rect 1720 -17 1754 17
rect 1720 -85 1754 -51
rect 1816 51 1850 85
rect 1816 -17 1850 17
rect 1816 -85 1850 -51
rect 1930 51 1964 85
rect 1930 -17 1964 17
rect 1930 -85 1964 -51
rect 2026 51 2060 85
rect 2026 -17 2060 17
rect 2026 -85 2060 -51
rect 2140 51 2174 85
rect 2140 -17 2174 17
rect 2140 -85 2174 -51
rect 2236 51 2270 85
rect 2236 -17 2270 17
rect 2236 -85 2270 -51
rect 2350 51 2384 85
rect 2350 -17 2384 17
rect 2350 -85 2384 -51
rect 2446 51 2480 85
rect 2446 -17 2480 17
rect 2446 -85 2480 -51
rect 2560 51 2594 85
rect 2560 -17 2594 17
rect 2560 -85 2594 -51
rect 2656 51 2690 85
rect 2656 -17 2690 17
rect 2656 -85 2690 -51
rect 2770 51 2804 85
rect 2770 -17 2804 17
rect 2770 -85 2804 -51
rect 2866 51 2900 85
rect 2866 -17 2900 17
rect 2866 -85 2900 -51
rect 2980 51 3014 85
rect 2980 -17 3014 17
rect 2980 -85 3014 -51
rect 3076 51 3110 85
rect 3076 -17 3110 17
rect 3076 -85 3110 -51
rect 3190 51 3224 85
rect 3190 -17 3224 17
rect 3190 -85 3224 -51
rect 3286 51 3320 85
rect 3286 -17 3320 17
rect 3286 -85 3320 -51
rect 3400 51 3434 85
rect 3400 -17 3434 17
rect 3400 -85 3434 -51
rect 3496 51 3530 85
rect 3496 -17 3530 17
rect 3496 -85 3530 -51
rect 3610 51 3644 85
rect 3610 -17 3644 17
rect 3610 -85 3644 -51
rect 3706 51 3740 85
rect 3706 -17 3740 17
rect 3706 -85 3740 -51
rect 3820 51 3854 85
rect 3820 -17 3854 17
rect 3820 -85 3854 -51
rect 3916 51 3950 85
rect 3916 -17 3950 17
rect 3916 -85 3950 -51
rect 4030 51 4064 85
rect 4030 -17 4064 17
rect 4030 -85 4064 -51
rect 4126 51 4160 85
rect 4126 -17 4160 17
rect 4126 -85 4160 -51
rect 4240 51 4274 85
rect 4240 -17 4274 17
rect 4240 -85 4274 -51
rect 4336 51 4370 85
rect 4336 -17 4370 17
rect 4336 -85 4370 -51
rect -4368 -481 -4334 -447
rect -4368 -549 -4334 -515
rect -4368 -617 -4334 -583
rect -4272 -481 -4238 -447
rect -4272 -549 -4238 -515
rect -4272 -617 -4238 -583
rect -4158 -481 -4124 -447
rect -4158 -549 -4124 -515
rect -4158 -617 -4124 -583
rect -4062 -481 -4028 -447
rect -4062 -549 -4028 -515
rect -4062 -617 -4028 -583
rect -3948 -481 -3914 -447
rect -3948 -549 -3914 -515
rect -3948 -617 -3914 -583
rect -3852 -481 -3818 -447
rect -3852 -549 -3818 -515
rect -3852 -617 -3818 -583
rect -3738 -481 -3704 -447
rect -3738 -549 -3704 -515
rect -3738 -617 -3704 -583
rect -3642 -481 -3608 -447
rect -3642 -549 -3608 -515
rect -3642 -617 -3608 -583
rect -3528 -481 -3494 -447
rect -3528 -549 -3494 -515
rect -3528 -617 -3494 -583
rect -3432 -481 -3398 -447
rect -3432 -549 -3398 -515
rect -3432 -617 -3398 -583
rect -3318 -481 -3284 -447
rect -3318 -549 -3284 -515
rect -3318 -617 -3284 -583
rect -3222 -481 -3188 -447
rect -3222 -549 -3188 -515
rect -3222 -617 -3188 -583
rect -3108 -481 -3074 -447
rect -3108 -549 -3074 -515
rect -3108 -617 -3074 -583
rect -3012 -481 -2978 -447
rect -3012 -549 -2978 -515
rect -3012 -617 -2978 -583
rect -2898 -481 -2864 -447
rect -2898 -549 -2864 -515
rect -2898 -617 -2864 -583
rect -2802 -481 -2768 -447
rect -2802 -549 -2768 -515
rect -2802 -617 -2768 -583
rect -2688 -481 -2654 -447
rect -2688 -549 -2654 -515
rect -2688 -617 -2654 -583
rect -2592 -481 -2558 -447
rect -2592 -549 -2558 -515
rect -2592 -617 -2558 -583
rect -2478 -481 -2444 -447
rect -2478 -549 -2444 -515
rect -2478 -617 -2444 -583
rect -2382 -481 -2348 -447
rect -2382 -549 -2348 -515
rect -2382 -617 -2348 -583
rect -2268 -481 -2234 -447
rect -2268 -549 -2234 -515
rect -2268 -617 -2234 -583
rect -2172 -481 -2138 -447
rect -2172 -549 -2138 -515
rect -2172 -617 -2138 -583
rect -2058 -481 -2024 -447
rect -2058 -549 -2024 -515
rect -2058 -617 -2024 -583
rect -1962 -481 -1928 -447
rect -1962 -549 -1928 -515
rect -1962 -617 -1928 -583
rect -1848 -481 -1814 -447
rect -1848 -549 -1814 -515
rect -1848 -617 -1814 -583
rect -1752 -481 -1718 -447
rect -1752 -549 -1718 -515
rect -1752 -617 -1718 -583
rect -1638 -481 -1604 -447
rect -1638 -549 -1604 -515
rect -1638 -617 -1604 -583
rect -1542 -481 -1508 -447
rect -1542 -549 -1508 -515
rect -1542 -617 -1508 -583
rect -1428 -481 -1394 -447
rect -1428 -549 -1394 -515
rect -1428 -617 -1394 -583
rect -1332 -481 -1298 -447
rect -1332 -549 -1298 -515
rect -1332 -617 -1298 -583
rect -1218 -481 -1184 -447
rect -1218 -549 -1184 -515
rect -1218 -617 -1184 -583
rect -1122 -481 -1088 -447
rect -1122 -549 -1088 -515
rect -1122 -617 -1088 -583
rect -1008 -481 -974 -447
rect -1008 -549 -974 -515
rect -1008 -617 -974 -583
rect -912 -481 -878 -447
rect -912 -549 -878 -515
rect -912 -617 -878 -583
rect -798 -481 -764 -447
rect -798 -549 -764 -515
rect -798 -617 -764 -583
rect -702 -481 -668 -447
rect -702 -549 -668 -515
rect -702 -617 -668 -583
rect -588 -481 -554 -447
rect -588 -549 -554 -515
rect -588 -617 -554 -583
rect -492 -481 -458 -447
rect -492 -549 -458 -515
rect -492 -617 -458 -583
rect -378 -481 -344 -447
rect -378 -549 -344 -515
rect -378 -617 -344 -583
rect -282 -481 -248 -447
rect -282 -549 -248 -515
rect -282 -617 -248 -583
rect -168 -481 -134 -447
rect -168 -549 -134 -515
rect -168 -617 -134 -583
rect -72 -481 -38 -447
rect -72 -549 -38 -515
rect -72 -617 -38 -583
rect 42 -481 76 -447
rect 42 -549 76 -515
rect 42 -617 76 -583
rect 138 -481 172 -447
rect 138 -549 172 -515
rect 138 -617 172 -583
rect 252 -481 286 -447
rect 252 -549 286 -515
rect 252 -617 286 -583
rect 348 -481 382 -447
rect 348 -549 382 -515
rect 348 -617 382 -583
rect 462 -481 496 -447
rect 462 -549 496 -515
rect 462 -617 496 -583
rect 558 -481 592 -447
rect 558 -549 592 -515
rect 558 -617 592 -583
rect 672 -481 706 -447
rect 672 -549 706 -515
rect 672 -617 706 -583
rect 768 -481 802 -447
rect 768 -549 802 -515
rect 768 -617 802 -583
rect 882 -481 916 -447
rect 882 -549 916 -515
rect 882 -617 916 -583
rect 978 -481 1012 -447
rect 978 -549 1012 -515
rect 978 -617 1012 -583
rect 1092 -481 1126 -447
rect 1092 -549 1126 -515
rect 1092 -617 1126 -583
rect 1188 -481 1222 -447
rect 1188 -549 1222 -515
rect 1188 -617 1222 -583
rect 1302 -481 1336 -447
rect 1302 -549 1336 -515
rect 1302 -617 1336 -583
rect 1398 -481 1432 -447
rect 1398 -549 1432 -515
rect 1398 -617 1432 -583
rect 1512 -481 1546 -447
rect 1512 -549 1546 -515
rect 1512 -617 1546 -583
rect 1608 -481 1642 -447
rect 1608 -549 1642 -515
rect 1608 -617 1642 -583
rect 1722 -481 1756 -447
rect 1722 -549 1756 -515
rect 1722 -617 1756 -583
rect 1818 -481 1852 -447
rect 1818 -549 1852 -515
rect 1818 -617 1852 -583
rect 1932 -481 1966 -447
rect 1932 -549 1966 -515
rect 1932 -617 1966 -583
rect 2028 -481 2062 -447
rect 2028 -549 2062 -515
rect 2028 -617 2062 -583
rect 2142 -481 2176 -447
rect 2142 -549 2176 -515
rect 2142 -617 2176 -583
rect 2238 -481 2272 -447
rect 2238 -549 2272 -515
rect 2238 -617 2272 -583
rect 2352 -481 2386 -447
rect 2352 -549 2386 -515
rect 2352 -617 2386 -583
rect 2448 -481 2482 -447
rect 2448 -549 2482 -515
rect 2448 -617 2482 -583
rect 2562 -481 2596 -447
rect 2562 -549 2596 -515
rect 2562 -617 2596 -583
rect 2658 -481 2692 -447
rect 2658 -549 2692 -515
rect 2658 -617 2692 -583
rect 2772 -481 2806 -447
rect 2772 -549 2806 -515
rect 2772 -617 2806 -583
rect 2868 -481 2902 -447
rect 2868 -549 2902 -515
rect 2868 -617 2902 -583
rect 2982 -481 3016 -447
rect 2982 -549 3016 -515
rect 2982 -617 3016 -583
rect 3078 -481 3112 -447
rect 3078 -549 3112 -515
rect 3078 -617 3112 -583
rect 3192 -481 3226 -447
rect 3192 -549 3226 -515
rect 3192 -617 3226 -583
rect 3288 -481 3322 -447
rect 3288 -549 3322 -515
rect 3288 -617 3322 -583
rect 3402 -481 3436 -447
rect 3402 -549 3436 -515
rect 3402 -617 3436 -583
rect 3498 -481 3532 -447
rect 3498 -549 3532 -515
rect 3498 -617 3532 -583
rect 3612 -481 3646 -447
rect 3612 -549 3646 -515
rect 3612 -617 3646 -583
rect 3708 -481 3742 -447
rect 3708 -549 3742 -515
rect 3708 -617 3742 -583
rect 3822 -481 3856 -447
rect 3822 -549 3856 -515
rect 3822 -617 3856 -583
rect 3918 -481 3952 -447
rect 3918 -549 3952 -515
rect 3918 -617 3952 -583
rect 4032 -481 4066 -447
rect 4032 -549 4066 -515
rect 4032 -617 4066 -583
rect 4128 -481 4162 -447
rect 4128 -549 4162 -515
rect 4128 -617 4162 -583
rect 4242 -481 4276 -447
rect 4242 -549 4276 -515
rect 4242 -617 4276 -583
rect 4338 -481 4372 -447
rect 4338 -549 4372 -515
rect 4338 -617 4372 -583
<< nsubdiff >>
rect -4484 249 -4369 283
rect -4335 249 -4301 283
rect -4267 249 -4233 283
rect -4199 249 -4165 283
rect -4131 249 -4097 283
rect -4063 249 -4029 283
rect -3995 249 -3961 283
rect -3927 249 -3893 283
rect -3859 249 -3825 283
rect -3791 249 -3757 283
rect -3723 249 -3689 283
rect -3655 249 -3621 283
rect -3587 249 -3553 283
rect -3519 249 -3485 283
rect -3451 249 -3417 283
rect -3383 249 -3349 283
rect -3315 249 -3281 283
rect -3247 249 -3213 283
rect -3179 249 -3145 283
rect -3111 249 -3077 283
rect -3043 249 -3009 283
rect -2975 249 -2941 283
rect -2907 249 -2873 283
rect -2839 249 -2805 283
rect -2771 249 -2737 283
rect -2703 249 -2669 283
rect -2635 249 -2601 283
rect -2567 249 -2533 283
rect -2499 249 -2465 283
rect -2431 249 -2397 283
rect -2363 249 -2329 283
rect -2295 249 -2261 283
rect -2227 249 -2193 283
rect -2159 249 -2125 283
rect -2091 249 -2057 283
rect -2023 249 -1989 283
rect -1955 249 -1921 283
rect -1887 249 -1853 283
rect -1819 249 -1785 283
rect -1751 249 -1717 283
rect -1683 249 -1649 283
rect -1615 249 -1581 283
rect -1547 249 -1513 283
rect -1479 249 -1445 283
rect -1411 249 -1377 283
rect -1343 249 -1309 283
rect -1275 249 -1241 283
rect -1207 249 -1173 283
rect -1139 249 -1105 283
rect -1071 249 -1037 283
rect -1003 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1003 283
rect 1037 249 1071 283
rect 1105 249 1139 283
rect 1173 249 1207 283
rect 1241 249 1275 283
rect 1309 249 1343 283
rect 1377 249 1411 283
rect 1445 249 1479 283
rect 1513 249 1547 283
rect 1581 249 1615 283
rect 1649 249 1683 283
rect 1717 249 1751 283
rect 1785 249 1819 283
rect 1853 249 1887 283
rect 1921 249 1955 283
rect 1989 249 2023 283
rect 2057 249 2091 283
rect 2125 249 2159 283
rect 2193 249 2227 283
rect 2261 249 2295 283
rect 2329 249 2363 283
rect 2397 249 2431 283
rect 2465 249 2499 283
rect 2533 249 2567 283
rect 2601 249 2635 283
rect 2669 249 2703 283
rect 2737 249 2771 283
rect 2805 249 2839 283
rect 2873 249 2907 283
rect 2941 249 2975 283
rect 3009 249 3043 283
rect 3077 249 3111 283
rect 3145 249 3179 283
rect 3213 249 3247 283
rect 3281 249 3315 283
rect 3349 249 3383 283
rect 3417 249 3451 283
rect 3485 249 3519 283
rect 3553 249 3587 283
rect 3621 249 3655 283
rect 3689 249 3723 283
rect 3757 249 3791 283
rect 3825 249 3859 283
rect 3893 249 3927 283
rect 3961 249 3995 283
rect 4029 249 4063 283
rect 4097 249 4131 283
rect 4165 249 4199 283
rect 4233 249 4267 283
rect 4301 249 4335 283
rect 4369 249 4484 283
rect -4484 187 -4450 249
rect -4484 119 -4450 153
rect 4450 187 4484 249
rect 4450 119 4484 153
rect -4484 51 -4450 85
rect -4484 -17 -4450 17
rect -4484 -85 -4450 -51
rect 4450 51 4484 85
rect 4450 -17 4484 17
rect 4450 -85 4484 -51
rect -4484 -153 -4450 -119
rect -4484 -345 -4450 -187
rect 4450 -153 4484 -119
rect -4484 -413 -4450 -379
rect 4450 -345 4484 -187
rect 4450 -413 4484 -379
rect -4484 -481 -4450 -447
rect -4484 -549 -4450 -515
rect -4484 -617 -4450 -583
rect 4450 -481 4484 -447
rect 4450 -549 4484 -515
rect 4450 -617 4484 -583
rect -4484 -685 -4450 -651
rect -4484 -781 -4450 -719
rect 4450 -685 4484 -651
rect 4450 -781 4484 -719
rect -4484 -815 -4369 -781
rect -4335 -815 -4301 -781
rect -4267 -815 -4233 -781
rect -4199 -815 -4165 -781
rect -4131 -815 -4097 -781
rect -4063 -815 -4029 -781
rect -3995 -815 -3961 -781
rect -3927 -815 -3893 -781
rect -3859 -815 -3825 -781
rect -3791 -815 -3757 -781
rect -3723 -815 -3689 -781
rect -3655 -815 -3621 -781
rect -3587 -815 -3553 -781
rect -3519 -815 -3485 -781
rect -3451 -815 -3417 -781
rect -3383 -815 -3349 -781
rect -3315 -815 -3281 -781
rect -3247 -815 -3213 -781
rect -3179 -815 -3145 -781
rect -3111 -815 -3077 -781
rect -3043 -815 -3009 -781
rect -2975 -815 -2941 -781
rect -2907 -815 -2873 -781
rect -2839 -815 -2805 -781
rect -2771 -815 -2737 -781
rect -2703 -815 -2669 -781
rect -2635 -815 -2601 -781
rect -2567 -815 -2533 -781
rect -2499 -815 -2465 -781
rect -2431 -815 -2397 -781
rect -2363 -815 -2329 -781
rect -2295 -815 -2261 -781
rect -2227 -815 -2193 -781
rect -2159 -815 -2125 -781
rect -2091 -815 -2057 -781
rect -2023 -815 -1989 -781
rect -1955 -815 -1921 -781
rect -1887 -815 -1853 -781
rect -1819 -815 -1785 -781
rect -1751 -815 -1717 -781
rect -1683 -815 -1649 -781
rect -1615 -815 -1581 -781
rect -1547 -815 -1513 -781
rect -1479 -815 -1445 -781
rect -1411 -815 -1377 -781
rect -1343 -815 -1309 -781
rect -1275 -815 -1241 -781
rect -1207 -815 -1173 -781
rect -1139 -815 -1105 -781
rect -1071 -815 -1037 -781
rect -1003 -815 -969 -781
rect -935 -815 -901 -781
rect -867 -815 -833 -781
rect -799 -815 -765 -781
rect -731 -815 -697 -781
rect -663 -815 -629 -781
rect -595 -815 -561 -781
rect -527 -815 -493 -781
rect -459 -815 -425 -781
rect -391 -815 -357 -781
rect -323 -815 -289 -781
rect -255 -815 -221 -781
rect -187 -815 -153 -781
rect -119 -815 -85 -781
rect -51 -815 -17 -781
rect 17 -815 51 -781
rect 85 -815 119 -781
rect 153 -815 187 -781
rect 221 -815 255 -781
rect 289 -815 323 -781
rect 357 -815 391 -781
rect 425 -815 459 -781
rect 493 -815 527 -781
rect 561 -815 595 -781
rect 629 -815 663 -781
rect 697 -815 731 -781
rect 765 -815 799 -781
rect 833 -815 867 -781
rect 901 -815 935 -781
rect 969 -815 1003 -781
rect 1037 -815 1071 -781
rect 1105 -815 1139 -781
rect 1173 -815 1207 -781
rect 1241 -815 1275 -781
rect 1309 -815 1343 -781
rect 1377 -815 1411 -781
rect 1445 -815 1479 -781
rect 1513 -815 1547 -781
rect 1581 -815 1615 -781
rect 1649 -815 1683 -781
rect 1717 -815 1751 -781
rect 1785 -815 1819 -781
rect 1853 -815 1887 -781
rect 1921 -815 1955 -781
rect 1989 -815 2023 -781
rect 2057 -815 2091 -781
rect 2125 -815 2159 -781
rect 2193 -815 2227 -781
rect 2261 -815 2295 -781
rect 2329 -815 2363 -781
rect 2397 -815 2431 -781
rect 2465 -815 2499 -781
rect 2533 -815 2567 -781
rect 2601 -815 2635 -781
rect 2669 -815 2703 -781
rect 2737 -815 2771 -781
rect 2805 -815 2839 -781
rect 2873 -815 2907 -781
rect 2941 -815 2975 -781
rect 3009 -815 3043 -781
rect 3077 -815 3111 -781
rect 3145 -815 3179 -781
rect 3213 -815 3247 -781
rect 3281 -815 3315 -781
rect 3349 -815 3383 -781
rect 3417 -815 3451 -781
rect 3485 -815 3519 -781
rect 3553 -815 3587 -781
rect 3621 -815 3655 -781
rect 3689 -815 3723 -781
rect 3757 -815 3791 -781
rect 3825 -815 3859 -781
rect 3893 -815 3927 -781
rect 3961 -815 3995 -781
rect 4029 -815 4063 -781
rect 4097 -815 4131 -781
rect 4165 -815 4199 -781
rect 4233 -815 4267 -781
rect 4301 -815 4335 -781
rect 4369 -815 4484 -781
<< nsubdiffcont >>
rect -4369 249 -4335 283
rect -4301 249 -4267 283
rect -4233 249 -4199 283
rect -4165 249 -4131 283
rect -4097 249 -4063 283
rect -4029 249 -3995 283
rect -3961 249 -3927 283
rect -3893 249 -3859 283
rect -3825 249 -3791 283
rect -3757 249 -3723 283
rect -3689 249 -3655 283
rect -3621 249 -3587 283
rect -3553 249 -3519 283
rect -3485 249 -3451 283
rect -3417 249 -3383 283
rect -3349 249 -3315 283
rect -3281 249 -3247 283
rect -3213 249 -3179 283
rect -3145 249 -3111 283
rect -3077 249 -3043 283
rect -3009 249 -2975 283
rect -2941 249 -2907 283
rect -2873 249 -2839 283
rect -2805 249 -2771 283
rect -2737 249 -2703 283
rect -2669 249 -2635 283
rect -2601 249 -2567 283
rect -2533 249 -2499 283
rect -2465 249 -2431 283
rect -2397 249 -2363 283
rect -2329 249 -2295 283
rect -2261 249 -2227 283
rect -2193 249 -2159 283
rect -2125 249 -2091 283
rect -2057 249 -2023 283
rect -1989 249 -1955 283
rect -1921 249 -1887 283
rect -1853 249 -1819 283
rect -1785 249 -1751 283
rect -1717 249 -1683 283
rect -1649 249 -1615 283
rect -1581 249 -1547 283
rect -1513 249 -1479 283
rect -1445 249 -1411 283
rect -1377 249 -1343 283
rect -1309 249 -1275 283
rect -1241 249 -1207 283
rect -1173 249 -1139 283
rect -1105 249 -1071 283
rect -1037 249 -1003 283
rect -969 249 -935 283
rect -901 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 901 283
rect 935 249 969 283
rect 1003 249 1037 283
rect 1071 249 1105 283
rect 1139 249 1173 283
rect 1207 249 1241 283
rect 1275 249 1309 283
rect 1343 249 1377 283
rect 1411 249 1445 283
rect 1479 249 1513 283
rect 1547 249 1581 283
rect 1615 249 1649 283
rect 1683 249 1717 283
rect 1751 249 1785 283
rect 1819 249 1853 283
rect 1887 249 1921 283
rect 1955 249 1989 283
rect 2023 249 2057 283
rect 2091 249 2125 283
rect 2159 249 2193 283
rect 2227 249 2261 283
rect 2295 249 2329 283
rect 2363 249 2397 283
rect 2431 249 2465 283
rect 2499 249 2533 283
rect 2567 249 2601 283
rect 2635 249 2669 283
rect 2703 249 2737 283
rect 2771 249 2805 283
rect 2839 249 2873 283
rect 2907 249 2941 283
rect 2975 249 3009 283
rect 3043 249 3077 283
rect 3111 249 3145 283
rect 3179 249 3213 283
rect 3247 249 3281 283
rect 3315 249 3349 283
rect 3383 249 3417 283
rect 3451 249 3485 283
rect 3519 249 3553 283
rect 3587 249 3621 283
rect 3655 249 3689 283
rect 3723 249 3757 283
rect 3791 249 3825 283
rect 3859 249 3893 283
rect 3927 249 3961 283
rect 3995 249 4029 283
rect 4063 249 4097 283
rect 4131 249 4165 283
rect 4199 249 4233 283
rect 4267 249 4301 283
rect 4335 249 4369 283
rect -4484 153 -4450 187
rect 4450 153 4484 187
rect -4484 85 -4450 119
rect -4484 17 -4450 51
rect -4484 -51 -4450 -17
rect -4484 -119 -4450 -85
rect 4450 85 4484 119
rect 4450 17 4484 51
rect 4450 -51 4484 -17
rect 4450 -119 4484 -85
rect -4484 -187 -4450 -153
rect 4450 -187 4484 -153
rect -4484 -379 -4450 -345
rect 4450 -379 4484 -345
rect -4484 -447 -4450 -413
rect -4484 -515 -4450 -481
rect -4484 -583 -4450 -549
rect -4484 -651 -4450 -617
rect 4450 -447 4484 -413
rect 4450 -515 4484 -481
rect 4450 -583 4484 -549
rect 4450 -651 4484 -617
rect -4484 -719 -4450 -685
rect 4450 -719 4484 -685
rect -4369 -815 -4335 -781
rect -4301 -815 -4267 -781
rect -4233 -815 -4199 -781
rect -4165 -815 -4131 -781
rect -4097 -815 -4063 -781
rect -4029 -815 -3995 -781
rect -3961 -815 -3927 -781
rect -3893 -815 -3859 -781
rect -3825 -815 -3791 -781
rect -3757 -815 -3723 -781
rect -3689 -815 -3655 -781
rect -3621 -815 -3587 -781
rect -3553 -815 -3519 -781
rect -3485 -815 -3451 -781
rect -3417 -815 -3383 -781
rect -3349 -815 -3315 -781
rect -3281 -815 -3247 -781
rect -3213 -815 -3179 -781
rect -3145 -815 -3111 -781
rect -3077 -815 -3043 -781
rect -3009 -815 -2975 -781
rect -2941 -815 -2907 -781
rect -2873 -815 -2839 -781
rect -2805 -815 -2771 -781
rect -2737 -815 -2703 -781
rect -2669 -815 -2635 -781
rect -2601 -815 -2567 -781
rect -2533 -815 -2499 -781
rect -2465 -815 -2431 -781
rect -2397 -815 -2363 -781
rect -2329 -815 -2295 -781
rect -2261 -815 -2227 -781
rect -2193 -815 -2159 -781
rect -2125 -815 -2091 -781
rect -2057 -815 -2023 -781
rect -1989 -815 -1955 -781
rect -1921 -815 -1887 -781
rect -1853 -815 -1819 -781
rect -1785 -815 -1751 -781
rect -1717 -815 -1683 -781
rect -1649 -815 -1615 -781
rect -1581 -815 -1547 -781
rect -1513 -815 -1479 -781
rect -1445 -815 -1411 -781
rect -1377 -815 -1343 -781
rect -1309 -815 -1275 -781
rect -1241 -815 -1207 -781
rect -1173 -815 -1139 -781
rect -1105 -815 -1071 -781
rect -1037 -815 -1003 -781
rect -969 -815 -935 -781
rect -901 -815 -867 -781
rect -833 -815 -799 -781
rect -765 -815 -731 -781
rect -697 -815 -663 -781
rect -629 -815 -595 -781
rect -561 -815 -527 -781
rect -493 -815 -459 -781
rect -425 -815 -391 -781
rect -357 -815 -323 -781
rect -289 -815 -255 -781
rect -221 -815 -187 -781
rect -153 -815 -119 -781
rect -85 -815 -51 -781
rect -17 -815 17 -781
rect 51 -815 85 -781
rect 119 -815 153 -781
rect 187 -815 221 -781
rect 255 -815 289 -781
rect 323 -815 357 -781
rect 391 -815 425 -781
rect 459 -815 493 -781
rect 527 -815 561 -781
rect 595 -815 629 -781
rect 663 -815 697 -781
rect 731 -815 765 -781
rect 799 -815 833 -781
rect 867 -815 901 -781
rect 935 -815 969 -781
rect 1003 -815 1037 -781
rect 1071 -815 1105 -781
rect 1139 -815 1173 -781
rect 1207 -815 1241 -781
rect 1275 -815 1309 -781
rect 1343 -815 1377 -781
rect 1411 -815 1445 -781
rect 1479 -815 1513 -781
rect 1547 -815 1581 -781
rect 1615 -815 1649 -781
rect 1683 -815 1717 -781
rect 1751 -815 1785 -781
rect 1819 -815 1853 -781
rect 1887 -815 1921 -781
rect 1955 -815 1989 -781
rect 2023 -815 2057 -781
rect 2091 -815 2125 -781
rect 2159 -815 2193 -781
rect 2227 -815 2261 -781
rect 2295 -815 2329 -781
rect 2363 -815 2397 -781
rect 2431 -815 2465 -781
rect 2499 -815 2533 -781
rect 2567 -815 2601 -781
rect 2635 -815 2669 -781
rect 2703 -815 2737 -781
rect 2771 -815 2805 -781
rect 2839 -815 2873 -781
rect 2907 -815 2941 -781
rect 2975 -815 3009 -781
rect 3043 -815 3077 -781
rect 3111 -815 3145 -781
rect 3179 -815 3213 -781
rect 3247 -815 3281 -781
rect 3315 -815 3349 -781
rect 3383 -815 3417 -781
rect 3451 -815 3485 -781
rect 3519 -815 3553 -781
rect 3587 -815 3621 -781
rect 3655 -815 3689 -781
rect 3723 -815 3757 -781
rect 3791 -815 3825 -781
rect 3859 -815 3893 -781
rect 3927 -815 3961 -781
rect 3995 -815 4029 -781
rect 4063 -815 4097 -781
rect 4131 -815 4165 -781
rect 4199 -815 4233 -781
rect 4267 -815 4301 -781
rect 4335 -815 4369 -781
<< poly >>
rect -4128 181 -4062 197
rect -4128 147 -4112 181
rect -4078 147 -4062 181
rect -4128 131 -4062 147
rect -3708 181 -3642 197
rect -3708 147 -3692 181
rect -3658 147 -3642 181
rect -3708 131 -3642 147
rect -3288 181 -3222 197
rect -3288 147 -3272 181
rect -3238 147 -3222 181
rect -3288 131 -3222 147
rect -2868 181 -2802 197
rect -2868 147 -2852 181
rect -2818 147 -2802 181
rect -2868 131 -2802 147
rect -2448 181 -2382 197
rect -2448 147 -2432 181
rect -2398 147 -2382 181
rect -2448 131 -2382 147
rect -2028 181 -1962 197
rect -2028 147 -2012 181
rect -1978 147 -1962 181
rect -2028 131 -1962 147
rect -1608 181 -1542 197
rect -1608 147 -1592 181
rect -1558 147 -1542 181
rect -1608 131 -1542 147
rect -1188 181 -1122 197
rect -1188 147 -1172 181
rect -1138 147 -1122 181
rect -1188 131 -1122 147
rect -768 181 -702 197
rect -768 147 -752 181
rect -718 147 -702 181
rect -768 131 -702 147
rect -348 181 -282 197
rect -348 147 -332 181
rect -298 147 -282 181
rect -348 131 -282 147
rect 72 181 138 197
rect 72 147 88 181
rect 122 147 138 181
rect 72 131 138 147
rect 492 181 558 197
rect 492 147 508 181
rect 542 147 558 181
rect 492 131 558 147
rect 912 181 978 197
rect 912 147 928 181
rect 962 147 978 181
rect 912 131 978 147
rect 1332 181 1398 197
rect 1332 147 1348 181
rect 1382 147 1398 181
rect 1332 131 1398 147
rect 1752 181 1818 197
rect 1752 147 1768 181
rect 1802 147 1818 181
rect 1752 131 1818 147
rect 2172 181 2238 197
rect 2172 147 2188 181
rect 2222 147 2238 181
rect 2172 131 2238 147
rect 2592 181 2658 197
rect 2592 147 2608 181
rect 2642 147 2658 181
rect 2592 131 2658 147
rect 3012 181 3078 197
rect 3012 147 3028 181
rect 3062 147 3078 181
rect 3012 131 3078 147
rect 3432 181 3498 197
rect 3432 147 3448 181
rect 3482 147 3498 181
rect 3432 131 3498 147
rect 3852 181 3918 197
rect 3852 147 3868 181
rect 3902 147 3918 181
rect 3852 131 3918 147
rect 4272 181 4338 197
rect 4272 147 4288 181
rect 4322 147 4338 181
rect 4272 131 4338 147
rect -4320 100 -4290 126
rect -4110 100 -4080 131
rect -3900 100 -3870 126
rect -3690 100 -3660 131
rect -3480 100 -3450 126
rect -3270 100 -3240 131
rect -3060 100 -3030 126
rect -2850 100 -2820 131
rect -2640 100 -2610 126
rect -2430 100 -2400 131
rect -2220 100 -2190 126
rect -2010 100 -1980 131
rect -1800 100 -1770 126
rect -1590 100 -1560 131
rect -1380 100 -1350 126
rect -1170 100 -1140 131
rect -960 100 -930 126
rect -750 100 -720 131
rect -540 100 -510 126
rect -330 100 -300 131
rect -120 100 -90 126
rect 90 100 120 131
rect 300 100 330 126
rect 510 100 540 131
rect 720 100 750 126
rect 930 100 960 131
rect 1140 100 1170 126
rect 1350 100 1380 131
rect 1560 100 1590 126
rect 1770 100 1800 131
rect 1980 100 2010 126
rect 2190 100 2220 131
rect 2400 100 2430 126
rect 2610 100 2640 131
rect 2820 100 2850 126
rect 3030 100 3060 131
rect 3240 100 3270 126
rect 3450 100 3480 131
rect 3660 100 3690 126
rect 3870 100 3900 131
rect 4080 100 4110 126
rect 4290 100 4320 131
rect -4320 -131 -4290 -100
rect -4110 -126 -4080 -100
rect -3900 -131 -3870 -100
rect -3690 -126 -3660 -100
rect -3480 -131 -3450 -100
rect -3270 -126 -3240 -100
rect -3060 -131 -3030 -100
rect -2850 -126 -2820 -100
rect -2640 -131 -2610 -100
rect -2430 -126 -2400 -100
rect -2220 -131 -2190 -100
rect -2010 -126 -1980 -100
rect -1800 -131 -1770 -100
rect -1590 -126 -1560 -100
rect -1380 -131 -1350 -100
rect -1170 -126 -1140 -100
rect -960 -131 -930 -100
rect -750 -126 -720 -100
rect -540 -131 -510 -100
rect -330 -126 -300 -100
rect -120 -131 -90 -100
rect 90 -126 120 -100
rect 300 -131 330 -100
rect 510 -126 540 -100
rect 720 -131 750 -100
rect 930 -126 960 -100
rect 1140 -131 1170 -100
rect 1350 -126 1380 -100
rect 1560 -131 1590 -100
rect 1770 -126 1800 -100
rect 1980 -131 2010 -100
rect 2190 -126 2220 -100
rect 2400 -131 2430 -100
rect 2610 -126 2640 -100
rect 2820 -131 2850 -100
rect 3030 -126 3060 -100
rect 3240 -131 3270 -100
rect 3450 -126 3480 -100
rect 3660 -131 3690 -100
rect 3870 -126 3900 -100
rect 4080 -131 4110 -100
rect 4290 -126 4320 -100
rect -4338 -147 -4272 -131
rect -4338 -181 -4322 -147
rect -4288 -181 -4272 -147
rect -4338 -197 -4272 -181
rect -3918 -147 -3852 -131
rect -3918 -181 -3902 -147
rect -3868 -181 -3852 -147
rect -3918 -197 -3852 -181
rect -3498 -147 -3432 -131
rect -3498 -181 -3482 -147
rect -3448 -181 -3432 -147
rect -3498 -197 -3432 -181
rect -3078 -147 -3012 -131
rect -3078 -181 -3062 -147
rect -3028 -181 -3012 -147
rect -3078 -197 -3012 -181
rect -2658 -147 -2592 -131
rect -2658 -181 -2642 -147
rect -2608 -181 -2592 -147
rect -2658 -197 -2592 -181
rect -2238 -147 -2172 -131
rect -2238 -181 -2222 -147
rect -2188 -181 -2172 -147
rect -2238 -197 -2172 -181
rect -1818 -147 -1752 -131
rect -1818 -181 -1802 -147
rect -1768 -181 -1752 -147
rect -1818 -197 -1752 -181
rect -1398 -147 -1332 -131
rect -1398 -181 -1382 -147
rect -1348 -181 -1332 -147
rect -1398 -197 -1332 -181
rect -978 -147 -912 -131
rect -978 -181 -962 -147
rect -928 -181 -912 -147
rect -978 -197 -912 -181
rect -558 -147 -492 -131
rect -558 -181 -542 -147
rect -508 -181 -492 -147
rect -558 -197 -492 -181
rect -138 -147 -72 -131
rect -138 -181 -122 -147
rect -88 -181 -72 -147
rect -138 -197 -72 -181
rect 282 -147 348 -131
rect 282 -181 298 -147
rect 332 -181 348 -147
rect 282 -197 348 -181
rect 702 -147 768 -131
rect 702 -181 718 -147
rect 752 -181 768 -147
rect 702 -197 768 -181
rect 1122 -147 1188 -131
rect 1122 -181 1138 -147
rect 1172 -181 1188 -147
rect 1122 -197 1188 -181
rect 1542 -147 1608 -131
rect 1542 -181 1558 -147
rect 1592 -181 1608 -147
rect 1542 -197 1608 -181
rect 1962 -147 2028 -131
rect 1962 -181 1978 -147
rect 2012 -181 2028 -147
rect 1962 -197 2028 -181
rect 2382 -147 2448 -131
rect 2382 -181 2398 -147
rect 2432 -181 2448 -147
rect 2382 -197 2448 -181
rect 2802 -147 2868 -131
rect 2802 -181 2818 -147
rect 2852 -181 2868 -147
rect 2802 -197 2868 -181
rect 3222 -147 3288 -131
rect 3222 -181 3238 -147
rect 3272 -181 3288 -147
rect 3222 -197 3288 -181
rect 3642 -147 3708 -131
rect 3642 -181 3658 -147
rect 3692 -181 3708 -147
rect 3642 -197 3708 -181
rect 4062 -147 4128 -131
rect 4062 -181 4078 -147
rect 4112 -181 4128 -147
rect 4062 -197 4128 -181
rect -4126 -351 -4060 -335
rect -4126 -385 -4110 -351
rect -4076 -385 -4060 -351
rect -4126 -401 -4060 -385
rect -3706 -351 -3640 -335
rect -3706 -385 -3690 -351
rect -3656 -385 -3640 -351
rect -3706 -401 -3640 -385
rect -3286 -351 -3220 -335
rect -3286 -385 -3270 -351
rect -3236 -385 -3220 -351
rect -3286 -401 -3220 -385
rect -2866 -351 -2800 -335
rect -2866 -385 -2850 -351
rect -2816 -385 -2800 -351
rect -2866 -401 -2800 -385
rect -2446 -351 -2380 -335
rect -2446 -385 -2430 -351
rect -2396 -385 -2380 -351
rect -2446 -401 -2380 -385
rect -2026 -351 -1960 -335
rect -2026 -385 -2010 -351
rect -1976 -385 -1960 -351
rect -2026 -401 -1960 -385
rect -1606 -351 -1540 -335
rect -1606 -385 -1590 -351
rect -1556 -385 -1540 -351
rect -1606 -401 -1540 -385
rect -1186 -351 -1120 -335
rect -1186 -385 -1170 -351
rect -1136 -385 -1120 -351
rect -1186 -401 -1120 -385
rect -766 -351 -700 -335
rect -766 -385 -750 -351
rect -716 -385 -700 -351
rect -766 -401 -700 -385
rect -346 -351 -280 -335
rect -346 -385 -330 -351
rect -296 -385 -280 -351
rect -346 -401 -280 -385
rect 74 -351 140 -335
rect 74 -385 90 -351
rect 124 -385 140 -351
rect 74 -401 140 -385
rect 494 -351 560 -335
rect 494 -385 510 -351
rect 544 -385 560 -351
rect 494 -401 560 -385
rect 914 -351 980 -335
rect 914 -385 930 -351
rect 964 -385 980 -351
rect 914 -401 980 -385
rect 1334 -351 1400 -335
rect 1334 -385 1350 -351
rect 1384 -385 1400 -351
rect 1334 -401 1400 -385
rect 1754 -351 1820 -335
rect 1754 -385 1770 -351
rect 1804 -385 1820 -351
rect 1754 -401 1820 -385
rect 2174 -351 2240 -335
rect 2174 -385 2190 -351
rect 2224 -385 2240 -351
rect 2174 -401 2240 -385
rect 2594 -351 2660 -335
rect 2594 -385 2610 -351
rect 2644 -385 2660 -351
rect 2594 -401 2660 -385
rect 3014 -351 3080 -335
rect 3014 -385 3030 -351
rect 3064 -385 3080 -351
rect 3014 -401 3080 -385
rect 3434 -351 3500 -335
rect 3434 -385 3450 -351
rect 3484 -385 3500 -351
rect 3434 -401 3500 -385
rect 3854 -351 3920 -335
rect 3854 -385 3870 -351
rect 3904 -385 3920 -351
rect 3854 -401 3920 -385
rect 4274 -351 4340 -335
rect 4274 -385 4290 -351
rect 4324 -385 4340 -351
rect 4274 -401 4340 -385
rect -4318 -432 -4288 -406
rect -4108 -432 -4078 -401
rect -3898 -432 -3868 -406
rect -3688 -432 -3658 -401
rect -3478 -432 -3448 -406
rect -3268 -432 -3238 -401
rect -3058 -432 -3028 -406
rect -2848 -432 -2818 -401
rect -2638 -432 -2608 -406
rect -2428 -432 -2398 -401
rect -2218 -432 -2188 -406
rect -2008 -432 -1978 -401
rect -1798 -432 -1768 -406
rect -1588 -432 -1558 -401
rect -1378 -432 -1348 -406
rect -1168 -432 -1138 -401
rect -958 -432 -928 -406
rect -748 -432 -718 -401
rect -538 -432 -508 -406
rect -328 -432 -298 -401
rect -118 -432 -88 -406
rect 92 -432 122 -401
rect 302 -432 332 -406
rect 512 -432 542 -401
rect 722 -432 752 -406
rect 932 -432 962 -401
rect 1142 -432 1172 -406
rect 1352 -432 1382 -401
rect 1562 -432 1592 -406
rect 1772 -432 1802 -401
rect 1982 -432 2012 -406
rect 2192 -432 2222 -401
rect 2402 -432 2432 -406
rect 2612 -432 2642 -401
rect 2822 -432 2852 -406
rect 3032 -432 3062 -401
rect 3242 -432 3272 -406
rect 3452 -432 3482 -401
rect 3662 -432 3692 -406
rect 3872 -432 3902 -401
rect 4082 -432 4112 -406
rect 4292 -432 4322 -401
rect -4318 -663 -4288 -632
rect -4108 -658 -4078 -632
rect -3898 -663 -3868 -632
rect -3688 -658 -3658 -632
rect -3478 -663 -3448 -632
rect -3268 -658 -3238 -632
rect -3058 -663 -3028 -632
rect -2848 -658 -2818 -632
rect -2638 -663 -2608 -632
rect -2428 -658 -2398 -632
rect -2218 -663 -2188 -632
rect -2008 -658 -1978 -632
rect -1798 -663 -1768 -632
rect -1588 -658 -1558 -632
rect -1378 -663 -1348 -632
rect -1168 -658 -1138 -632
rect -958 -663 -928 -632
rect -748 -658 -718 -632
rect -538 -663 -508 -632
rect -328 -658 -298 -632
rect -118 -663 -88 -632
rect 92 -658 122 -632
rect 302 -663 332 -632
rect 512 -658 542 -632
rect 722 -663 752 -632
rect 932 -658 962 -632
rect 1142 -663 1172 -632
rect 1352 -658 1382 -632
rect 1562 -663 1592 -632
rect 1772 -658 1802 -632
rect 1982 -663 2012 -632
rect 2192 -658 2222 -632
rect 2402 -663 2432 -632
rect 2612 -658 2642 -632
rect 2822 -663 2852 -632
rect 3032 -658 3062 -632
rect 3242 -663 3272 -632
rect 3452 -658 3482 -632
rect 3662 -663 3692 -632
rect 3872 -658 3902 -632
rect 4082 -663 4112 -632
rect 4292 -658 4322 -632
rect -4336 -679 -4270 -663
rect -4336 -713 -4320 -679
rect -4286 -713 -4270 -679
rect -4336 -729 -4270 -713
rect -3916 -679 -3850 -663
rect -3916 -713 -3900 -679
rect -3866 -713 -3850 -679
rect -3916 -729 -3850 -713
rect -3496 -679 -3430 -663
rect -3496 -713 -3480 -679
rect -3446 -713 -3430 -679
rect -3496 -729 -3430 -713
rect -3076 -679 -3010 -663
rect -3076 -713 -3060 -679
rect -3026 -713 -3010 -679
rect -3076 -729 -3010 -713
rect -2656 -679 -2590 -663
rect -2656 -713 -2640 -679
rect -2606 -713 -2590 -679
rect -2656 -729 -2590 -713
rect -2236 -679 -2170 -663
rect -2236 -713 -2220 -679
rect -2186 -713 -2170 -679
rect -2236 -729 -2170 -713
rect -1816 -679 -1750 -663
rect -1816 -713 -1800 -679
rect -1766 -713 -1750 -679
rect -1816 -729 -1750 -713
rect -1396 -679 -1330 -663
rect -1396 -713 -1380 -679
rect -1346 -713 -1330 -679
rect -1396 -729 -1330 -713
rect -976 -679 -910 -663
rect -976 -713 -960 -679
rect -926 -713 -910 -679
rect -976 -729 -910 -713
rect -556 -679 -490 -663
rect -556 -713 -540 -679
rect -506 -713 -490 -679
rect -556 -729 -490 -713
rect -136 -679 -70 -663
rect -136 -713 -120 -679
rect -86 -713 -70 -679
rect -136 -729 -70 -713
rect 284 -679 350 -663
rect 284 -713 300 -679
rect 334 -713 350 -679
rect 284 -729 350 -713
rect 704 -679 770 -663
rect 704 -713 720 -679
rect 754 -713 770 -679
rect 704 -729 770 -713
rect 1124 -679 1190 -663
rect 1124 -713 1140 -679
rect 1174 -713 1190 -679
rect 1124 -729 1190 -713
rect 1544 -679 1610 -663
rect 1544 -713 1560 -679
rect 1594 -713 1610 -679
rect 1544 -729 1610 -713
rect 1964 -679 2030 -663
rect 1964 -713 1980 -679
rect 2014 -713 2030 -679
rect 1964 -729 2030 -713
rect 2384 -679 2450 -663
rect 2384 -713 2400 -679
rect 2434 -713 2450 -679
rect 2384 -729 2450 -713
rect 2804 -679 2870 -663
rect 2804 -713 2820 -679
rect 2854 -713 2870 -679
rect 2804 -729 2870 -713
rect 3224 -679 3290 -663
rect 3224 -713 3240 -679
rect 3274 -713 3290 -679
rect 3224 -729 3290 -713
rect 3644 -679 3710 -663
rect 3644 -713 3660 -679
rect 3694 -713 3710 -679
rect 3644 -729 3710 -713
rect 4064 -679 4130 -663
rect 4064 -713 4080 -679
rect 4114 -713 4130 -679
rect 4064 -729 4130 -713
<< polycont >>
rect -4112 147 -4078 181
rect -3692 147 -3658 181
rect -3272 147 -3238 181
rect -2852 147 -2818 181
rect -2432 147 -2398 181
rect -2012 147 -1978 181
rect -1592 147 -1558 181
rect -1172 147 -1138 181
rect -752 147 -718 181
rect -332 147 -298 181
rect 88 147 122 181
rect 508 147 542 181
rect 928 147 962 181
rect 1348 147 1382 181
rect 1768 147 1802 181
rect 2188 147 2222 181
rect 2608 147 2642 181
rect 3028 147 3062 181
rect 3448 147 3482 181
rect 3868 147 3902 181
rect 4288 147 4322 181
rect -4322 -181 -4288 -147
rect -3902 -181 -3868 -147
rect -3482 -181 -3448 -147
rect -3062 -181 -3028 -147
rect -2642 -181 -2608 -147
rect -2222 -181 -2188 -147
rect -1802 -181 -1768 -147
rect -1382 -181 -1348 -147
rect -962 -181 -928 -147
rect -542 -181 -508 -147
rect -122 -181 -88 -147
rect 298 -181 332 -147
rect 718 -181 752 -147
rect 1138 -181 1172 -147
rect 1558 -181 1592 -147
rect 1978 -181 2012 -147
rect 2398 -181 2432 -147
rect 2818 -181 2852 -147
rect 3238 -181 3272 -147
rect 3658 -181 3692 -147
rect 4078 -181 4112 -147
rect -4110 -385 -4076 -351
rect -3690 -385 -3656 -351
rect -3270 -385 -3236 -351
rect -2850 -385 -2816 -351
rect -2430 -385 -2396 -351
rect -2010 -385 -1976 -351
rect -1590 -385 -1556 -351
rect -1170 -385 -1136 -351
rect -750 -385 -716 -351
rect -330 -385 -296 -351
rect 90 -385 124 -351
rect 510 -385 544 -351
rect 930 -385 964 -351
rect 1350 -385 1384 -351
rect 1770 -385 1804 -351
rect 2190 -385 2224 -351
rect 2610 -385 2644 -351
rect 3030 -385 3064 -351
rect 3450 -385 3484 -351
rect 3870 -385 3904 -351
rect 4290 -385 4324 -351
rect -4320 -713 -4286 -679
rect -3900 -713 -3866 -679
rect -3480 -713 -3446 -679
rect -3060 -713 -3026 -679
rect -2640 -713 -2606 -679
rect -2220 -713 -2186 -679
rect -1800 -713 -1766 -679
rect -1380 -713 -1346 -679
rect -960 -713 -926 -679
rect -540 -713 -506 -679
rect -120 -713 -86 -679
rect 300 -713 334 -679
rect 720 -713 754 -679
rect 1140 -713 1174 -679
rect 1560 -713 1594 -679
rect 1980 -713 2014 -679
rect 2400 -713 2434 -679
rect 2820 -713 2854 -679
rect 3240 -713 3274 -679
rect 3660 -713 3694 -679
rect 4080 -713 4114 -679
<< locali >>
rect -4484 249 -4369 283
rect -4335 249 -4301 283
rect -4267 249 -4233 283
rect -4199 249 -4165 283
rect -4131 249 -4097 283
rect -4063 249 -4029 283
rect -3995 249 -3961 283
rect -3927 249 -3893 283
rect -3859 249 -3825 283
rect -3791 249 -3757 283
rect -3723 249 -3689 283
rect -3655 249 -3621 283
rect -3587 249 -3553 283
rect -3519 249 -3485 283
rect -3451 249 -3417 283
rect -3383 249 -3349 283
rect -3315 249 -3281 283
rect -3247 249 -3213 283
rect -3179 249 -3145 283
rect -3111 249 -3077 283
rect -3043 249 -3009 283
rect -2975 249 -2941 283
rect -2907 249 -2873 283
rect -2839 249 -2805 283
rect -2771 249 -2737 283
rect -2703 249 -2669 283
rect -2635 249 -2601 283
rect -2567 249 -2533 283
rect -2499 249 -2465 283
rect -2431 249 -2397 283
rect -2363 249 -2329 283
rect -2295 249 -2261 283
rect -2227 249 -2193 283
rect -2159 249 -2125 283
rect -2091 249 -2057 283
rect -2023 249 -1989 283
rect -1955 249 -1921 283
rect -1887 249 -1853 283
rect -1819 249 -1785 283
rect -1751 249 -1717 283
rect -1683 249 -1649 283
rect -1615 249 -1581 283
rect -1547 249 -1513 283
rect -1479 249 -1445 283
rect -1411 249 -1377 283
rect -1343 249 -1309 283
rect -1275 249 -1241 283
rect -1207 249 -1173 283
rect -1139 249 -1105 283
rect -1071 249 -1037 283
rect -1003 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1003 283
rect 1037 249 1071 283
rect 1105 249 1139 283
rect 1173 249 1207 283
rect 1241 249 1275 283
rect 1309 249 1343 283
rect 1377 249 1411 283
rect 1445 249 1479 283
rect 1513 249 1547 283
rect 1581 249 1615 283
rect 1649 249 1683 283
rect 1717 249 1751 283
rect 1785 249 1819 283
rect 1853 249 1887 283
rect 1921 249 1955 283
rect 1989 249 2023 283
rect 2057 249 2091 283
rect 2125 249 2159 283
rect 2193 249 2227 283
rect 2261 249 2295 283
rect 2329 249 2363 283
rect 2397 249 2431 283
rect 2465 249 2499 283
rect 2533 249 2567 283
rect 2601 249 2635 283
rect 2669 249 2703 283
rect 2737 249 2771 283
rect 2805 249 2839 283
rect 2873 249 2907 283
rect 2941 249 2975 283
rect 3009 249 3043 283
rect 3077 249 3111 283
rect 3145 249 3179 283
rect 3213 249 3247 283
rect 3281 249 3315 283
rect 3349 249 3383 283
rect 3417 249 3451 283
rect 3485 249 3519 283
rect 3553 249 3587 283
rect 3621 249 3655 283
rect 3689 249 3723 283
rect 3757 249 3791 283
rect 3825 249 3859 283
rect 3893 249 3927 283
rect 3961 249 3995 283
rect 4029 249 4063 283
rect 4097 249 4131 283
rect 4165 249 4199 283
rect 4233 249 4267 283
rect 4301 249 4335 283
rect 4369 249 4484 283
rect -4484 187 -4450 249
rect 4450 187 4484 249
rect -4484 119 -4450 153
rect -4128 147 -4112 181
rect -4078 147 -4062 181
rect -3708 147 -3692 181
rect -3658 147 -3642 181
rect -3288 147 -3272 181
rect -3238 147 -3222 181
rect -2868 147 -2852 181
rect -2818 147 -2802 181
rect -2448 147 -2432 181
rect -2398 147 -2382 181
rect -2028 147 -2012 181
rect -1978 147 -1962 181
rect -1608 147 -1592 181
rect -1558 147 -1542 181
rect -1188 147 -1172 181
rect -1138 147 -1122 181
rect -768 147 -752 181
rect -718 147 -702 181
rect -348 147 -332 181
rect -298 147 -282 181
rect 72 147 88 181
rect 122 147 138 181
rect 492 147 508 181
rect 542 147 558 181
rect 912 147 928 181
rect 962 147 978 181
rect 1332 147 1348 181
rect 1382 147 1398 181
rect 1752 147 1768 181
rect 1802 147 1818 181
rect 2172 147 2188 181
rect 2222 147 2238 181
rect 2592 147 2608 181
rect 2642 147 2658 181
rect 3012 147 3028 181
rect 3062 147 3078 181
rect 3432 147 3448 181
rect 3482 147 3498 181
rect 3852 147 3868 181
rect 3902 147 3918 181
rect 4240 147 4288 181
rect 4322 153 4450 181
rect 4322 147 4484 153
rect -4484 51 -4450 85
rect -4484 -17 -4450 17
rect -4484 -85 -4450 -51
rect -4484 -147 -4450 -119
rect -4370 85 -4336 104
rect -4370 17 -4336 51
rect -4370 -51 -4336 -17
rect -4370 -147 -4336 -85
rect -4274 85 -4240 104
rect -4274 17 -4240 51
rect -4274 -51 -4240 -17
rect -4274 -147 -4240 -85
rect -4160 85 -4126 104
rect -4160 17 -4126 51
rect -4160 -51 -4126 -17
rect -4160 -104 -4126 -85
rect -4064 85 -4030 104
rect -4064 17 -4030 51
rect -4064 -51 -4030 -17
rect -4064 -104 -4030 -85
rect -3950 85 -3916 104
rect -3950 17 -3916 51
rect -3950 -51 -3916 -17
rect -3950 -104 -3916 -85
rect -3854 85 -3820 104
rect -3854 17 -3820 51
rect -3854 -51 -3820 -17
rect -3854 -104 -3820 -85
rect -3740 85 -3706 104
rect -3740 17 -3706 51
rect -3740 -51 -3706 -17
rect -3740 -104 -3706 -85
rect -3644 85 -3610 104
rect -3644 17 -3610 51
rect -3644 -51 -3610 -17
rect -3644 -104 -3610 -85
rect -3530 85 -3496 104
rect -3530 17 -3496 51
rect -3530 -51 -3496 -17
rect -3530 -104 -3496 -85
rect -3434 85 -3400 104
rect -3434 17 -3400 51
rect -3434 -51 -3400 -17
rect -3434 -104 -3400 -85
rect -3320 85 -3286 104
rect -3320 17 -3286 51
rect -3320 -51 -3286 -17
rect -3320 -104 -3286 -85
rect -3224 85 -3190 104
rect -3224 17 -3190 51
rect -3224 -51 -3190 -17
rect -3224 -104 -3190 -85
rect -3110 85 -3076 104
rect -3110 17 -3076 51
rect -3110 -51 -3076 -17
rect -3110 -104 -3076 -85
rect -3014 85 -2980 104
rect -3014 17 -2980 51
rect -3014 -51 -2980 -17
rect -3014 -104 -2980 -85
rect -2900 85 -2866 104
rect -2900 17 -2866 51
rect -2900 -51 -2866 -17
rect -2900 -104 -2866 -85
rect -2804 85 -2770 104
rect -2804 17 -2770 51
rect -2804 -51 -2770 -17
rect -2804 -104 -2770 -85
rect -2690 85 -2656 104
rect -2690 17 -2656 51
rect -2690 -51 -2656 -17
rect -2690 -104 -2656 -85
rect -2594 85 -2560 104
rect -2594 17 -2560 51
rect -2594 -51 -2560 -17
rect -2594 -104 -2560 -85
rect -2480 85 -2446 104
rect -2480 17 -2446 51
rect -2480 -51 -2446 -17
rect -2480 -104 -2446 -85
rect -2384 85 -2350 104
rect -2384 17 -2350 51
rect -2384 -51 -2350 -17
rect -2384 -104 -2350 -85
rect -2270 85 -2236 104
rect -2270 17 -2236 51
rect -2270 -51 -2236 -17
rect -2270 -104 -2236 -85
rect -2174 85 -2140 104
rect -2174 17 -2140 51
rect -2174 -51 -2140 -17
rect -2174 -104 -2140 -85
rect -2060 85 -2026 104
rect -2060 17 -2026 51
rect -2060 -51 -2026 -17
rect -2060 -104 -2026 -85
rect -1964 85 -1930 104
rect -1964 17 -1930 51
rect -1964 -51 -1930 -17
rect -1964 -104 -1930 -85
rect -1850 85 -1816 104
rect -1850 17 -1816 51
rect -1850 -51 -1816 -17
rect -1850 -104 -1816 -85
rect -1754 85 -1720 104
rect -1754 17 -1720 51
rect -1754 -51 -1720 -17
rect -1754 -104 -1720 -85
rect -1640 85 -1606 104
rect -1640 17 -1606 51
rect -1640 -51 -1606 -17
rect -1640 -104 -1606 -85
rect -1544 85 -1510 104
rect -1544 17 -1510 51
rect -1544 -51 -1510 -17
rect -1544 -104 -1510 -85
rect -1430 85 -1396 104
rect -1430 17 -1396 51
rect -1430 -51 -1396 -17
rect -1430 -104 -1396 -85
rect -1334 85 -1300 104
rect -1334 17 -1300 51
rect -1334 -51 -1300 -17
rect -1334 -104 -1300 -85
rect -1220 85 -1186 104
rect -1220 17 -1186 51
rect -1220 -51 -1186 -17
rect -1220 -104 -1186 -85
rect -1124 85 -1090 104
rect -1124 17 -1090 51
rect -1124 -51 -1090 -17
rect -1124 -104 -1090 -85
rect -1010 85 -976 104
rect -1010 17 -976 51
rect -1010 -51 -976 -17
rect -1010 -104 -976 -85
rect -914 85 -880 104
rect -914 17 -880 51
rect -914 -51 -880 -17
rect -914 -104 -880 -85
rect -800 85 -766 104
rect -800 17 -766 51
rect -800 -51 -766 -17
rect -800 -104 -766 -85
rect -704 85 -670 104
rect -704 17 -670 51
rect -704 -51 -670 -17
rect -704 -104 -670 -85
rect -590 85 -556 104
rect -590 17 -556 51
rect -590 -51 -556 -17
rect -590 -104 -556 -85
rect -494 85 -460 104
rect -494 17 -460 51
rect -494 -51 -460 -17
rect -494 -104 -460 -85
rect -380 85 -346 104
rect -380 17 -346 51
rect -380 -51 -346 -17
rect -380 -104 -346 -85
rect -284 85 -250 104
rect -284 17 -250 51
rect -284 -51 -250 -17
rect -284 -104 -250 -85
rect -170 85 -136 104
rect -170 17 -136 51
rect -170 -51 -136 -17
rect -170 -104 -136 -85
rect -74 85 -40 104
rect -74 17 -40 51
rect -74 -51 -40 -17
rect -74 -104 -40 -85
rect 40 85 74 104
rect 40 17 74 51
rect 40 -51 74 -17
rect 40 -104 74 -85
rect 136 85 170 104
rect 136 17 170 51
rect 136 -51 170 -17
rect 136 -104 170 -85
rect 250 85 284 104
rect 250 17 284 51
rect 250 -51 284 -17
rect 250 -104 284 -85
rect 346 85 380 104
rect 346 17 380 51
rect 346 -51 380 -17
rect 346 -104 380 -85
rect 460 85 494 104
rect 460 17 494 51
rect 460 -51 494 -17
rect 460 -104 494 -85
rect 556 85 590 104
rect 556 17 590 51
rect 556 -51 590 -17
rect 556 -104 590 -85
rect 670 85 704 104
rect 670 17 704 51
rect 670 -51 704 -17
rect 670 -104 704 -85
rect 766 85 800 104
rect 766 17 800 51
rect 766 -51 800 -17
rect 766 -104 800 -85
rect 880 85 914 104
rect 880 17 914 51
rect 880 -51 914 -17
rect 880 -104 914 -85
rect 976 85 1010 104
rect 976 17 1010 51
rect 976 -51 1010 -17
rect 976 -104 1010 -85
rect 1090 85 1124 104
rect 1090 17 1124 51
rect 1090 -51 1124 -17
rect 1090 -104 1124 -85
rect 1186 85 1220 104
rect 1186 17 1220 51
rect 1186 -51 1220 -17
rect 1186 -104 1220 -85
rect 1300 85 1334 104
rect 1300 17 1334 51
rect 1300 -51 1334 -17
rect 1300 -104 1334 -85
rect 1396 85 1430 104
rect 1396 17 1430 51
rect 1396 -51 1430 -17
rect 1396 -104 1430 -85
rect 1510 85 1544 104
rect 1510 17 1544 51
rect 1510 -51 1544 -17
rect 1510 -104 1544 -85
rect 1606 85 1640 104
rect 1606 17 1640 51
rect 1606 -51 1640 -17
rect 1606 -104 1640 -85
rect 1720 85 1754 104
rect 1720 17 1754 51
rect 1720 -51 1754 -17
rect 1720 -104 1754 -85
rect 1816 85 1850 104
rect 1816 17 1850 51
rect 1816 -51 1850 -17
rect 1816 -104 1850 -85
rect 1930 85 1964 104
rect 1930 17 1964 51
rect 1930 -51 1964 -17
rect 1930 -104 1964 -85
rect 2026 85 2060 104
rect 2026 17 2060 51
rect 2026 -51 2060 -17
rect 2026 -104 2060 -85
rect 2140 85 2174 104
rect 2140 17 2174 51
rect 2140 -51 2174 -17
rect 2140 -104 2174 -85
rect 2236 85 2270 104
rect 2236 17 2270 51
rect 2236 -51 2270 -17
rect 2236 -104 2270 -85
rect 2350 85 2384 104
rect 2350 17 2384 51
rect 2350 -51 2384 -17
rect 2350 -104 2384 -85
rect 2446 85 2480 104
rect 2446 17 2480 51
rect 2446 -51 2480 -17
rect 2446 -104 2480 -85
rect 2560 85 2594 104
rect 2560 17 2594 51
rect 2560 -51 2594 -17
rect 2560 -104 2594 -85
rect 2656 85 2690 104
rect 2656 17 2690 51
rect 2656 -51 2690 -17
rect 2656 -104 2690 -85
rect 2770 85 2804 104
rect 2770 17 2804 51
rect 2770 -51 2804 -17
rect 2770 -104 2804 -85
rect 2866 85 2900 104
rect 2866 17 2900 51
rect 2866 -51 2900 -17
rect 2866 -104 2900 -85
rect 2980 85 3014 104
rect 2980 17 3014 51
rect 2980 -51 3014 -17
rect 2980 -104 3014 -85
rect 3076 85 3110 104
rect 3076 17 3110 51
rect 3076 -51 3110 -17
rect 3076 -104 3110 -85
rect 3190 85 3224 104
rect 3190 17 3224 51
rect 3190 -51 3224 -17
rect 3190 -104 3224 -85
rect 3286 85 3320 104
rect 3286 17 3320 51
rect 3286 -51 3320 -17
rect 3286 -104 3320 -85
rect 3400 85 3434 104
rect 3400 17 3434 51
rect 3400 -51 3434 -17
rect 3400 -104 3434 -85
rect 3496 85 3530 104
rect 3496 17 3530 51
rect 3496 -51 3530 -17
rect 3496 -104 3530 -85
rect 3610 85 3644 104
rect 3610 17 3644 51
rect 3610 -51 3644 -17
rect 3610 -104 3644 -85
rect 3706 85 3740 104
rect 3706 17 3740 51
rect 3706 -51 3740 -17
rect 3706 -104 3740 -85
rect 3820 85 3854 104
rect 3820 17 3854 51
rect 3820 -51 3854 -17
rect 3820 -104 3854 -85
rect 3916 85 3950 104
rect 3916 17 3950 51
rect 3916 -51 3950 -17
rect 3916 -104 3950 -85
rect 4030 85 4064 104
rect 4030 17 4064 51
rect 4030 -51 4064 -17
rect 4030 -104 4064 -85
rect 4126 85 4160 104
rect 4126 17 4160 51
rect 4126 -51 4160 -17
rect 4126 -104 4160 -85
rect 4240 85 4274 147
rect 4240 17 4274 51
rect 4240 -51 4274 -17
rect 4240 -104 4274 -85
rect 4336 85 4370 147
rect 4336 17 4370 51
rect 4336 -51 4370 -17
rect 4336 -104 4370 -85
rect 4450 119 4484 147
rect 4450 51 4484 85
rect 4450 -17 4484 17
rect 4450 -85 4484 -51
rect -4484 -153 -4322 -147
rect -4450 -181 -4322 -153
rect -4288 -181 -4240 -147
rect -3918 -181 -3902 -147
rect -3868 -181 -3852 -147
rect -3498 -181 -3482 -147
rect -3448 -181 -3432 -147
rect -3078 -181 -3062 -147
rect -3028 -181 -3012 -147
rect -2658 -181 -2642 -147
rect -2608 -181 -2592 -147
rect -2238 -181 -2222 -147
rect -2188 -181 -2172 -147
rect -1818 -181 -1802 -147
rect -1768 -181 -1752 -147
rect -1398 -181 -1382 -147
rect -1348 -181 -1332 -147
rect -978 -181 -962 -147
rect -928 -181 -912 -147
rect -558 -181 -542 -147
rect -508 -181 -492 -147
rect -138 -181 -122 -147
rect -88 -181 -72 -147
rect 282 -181 298 -147
rect 332 -181 348 -147
rect 702 -181 718 -147
rect 752 -181 768 -147
rect 1122 -181 1138 -147
rect 1172 -181 1188 -147
rect 1542 -181 1558 -147
rect 1592 -181 1608 -147
rect 1962 -181 1978 -147
rect 2012 -181 2028 -147
rect 2382 -181 2398 -147
rect 2432 -181 2448 -147
rect 2802 -181 2818 -147
rect 2852 -181 2868 -147
rect 3222 -181 3238 -147
rect 3272 -181 3288 -147
rect 3642 -181 3658 -147
rect 3692 -181 3708 -147
rect 4062 -181 4078 -147
rect 4112 -181 4128 -147
rect 4450 -153 4484 -119
rect -4484 -345 -4450 -187
rect 4450 -345 4484 -187
rect -4484 -413 -4450 -379
rect -4126 -385 -4110 -351
rect -4076 -385 -4060 -351
rect -3706 -385 -3690 -351
rect -3656 -385 -3640 -351
rect -3286 -385 -3270 -351
rect -3236 -385 -3220 -351
rect -2866 -385 -2850 -351
rect -2816 -385 -2800 -351
rect -2446 -385 -2430 -351
rect -2396 -385 -2380 -351
rect -2026 -385 -2010 -351
rect -1976 -385 -1960 -351
rect -1606 -385 -1590 -351
rect -1556 -385 -1540 -351
rect -1186 -385 -1170 -351
rect -1136 -385 -1120 -351
rect -766 -385 -750 -351
rect -716 -385 -700 -351
rect -346 -385 -330 -351
rect -296 -385 -280 -351
rect 74 -385 90 -351
rect 124 -385 140 -351
rect 494 -385 510 -351
rect 544 -385 560 -351
rect 914 -385 930 -351
rect 964 -385 980 -351
rect 1334 -385 1350 -351
rect 1384 -385 1400 -351
rect 1754 -385 1770 -351
rect 1804 -385 1820 -351
rect 2174 -385 2190 -351
rect 2224 -385 2240 -351
rect 2594 -385 2610 -351
rect 2644 -385 2660 -351
rect 3014 -385 3030 -351
rect 3064 -385 3080 -351
rect 3434 -385 3450 -351
rect 3484 -385 3500 -351
rect 3854 -385 3870 -351
rect 3904 -385 3920 -351
rect 4242 -385 4290 -351
rect 4324 -379 4450 -351
rect 4324 -385 4484 -379
rect -4484 -481 -4450 -447
rect -4484 -549 -4450 -515
rect -4484 -617 -4450 -583
rect -4484 -679 -4450 -651
rect -4368 -447 -4334 -428
rect -4368 -515 -4334 -481
rect -4368 -583 -4334 -549
rect -4368 -679 -4334 -617
rect -4272 -447 -4238 -428
rect -4272 -515 -4238 -481
rect -4272 -583 -4238 -549
rect -4272 -679 -4238 -617
rect -4158 -447 -4124 -428
rect -4158 -515 -4124 -481
rect -4158 -583 -4124 -549
rect -4158 -636 -4124 -617
rect -4062 -447 -4028 -428
rect -4062 -515 -4028 -481
rect -4062 -583 -4028 -549
rect -4062 -636 -4028 -617
rect -3948 -447 -3914 -428
rect -3948 -515 -3914 -481
rect -3948 -583 -3914 -549
rect -3948 -636 -3914 -617
rect -3852 -447 -3818 -428
rect -3852 -515 -3818 -481
rect -3852 -583 -3818 -549
rect -3852 -636 -3818 -617
rect -3738 -447 -3704 -428
rect -3738 -515 -3704 -481
rect -3738 -583 -3704 -549
rect -3738 -636 -3704 -617
rect -3642 -447 -3608 -428
rect -3642 -515 -3608 -481
rect -3642 -583 -3608 -549
rect -3642 -636 -3608 -617
rect -3528 -447 -3494 -428
rect -3528 -515 -3494 -481
rect -3528 -583 -3494 -549
rect -3528 -636 -3494 -617
rect -3432 -447 -3398 -428
rect -3432 -515 -3398 -481
rect -3432 -583 -3398 -549
rect -3432 -636 -3398 -617
rect -3318 -447 -3284 -428
rect -3318 -515 -3284 -481
rect -3318 -583 -3284 -549
rect -3318 -636 -3284 -617
rect -3222 -447 -3188 -428
rect -3222 -515 -3188 -481
rect -3222 -583 -3188 -549
rect -3222 -636 -3188 -617
rect -3108 -447 -3074 -428
rect -3108 -515 -3074 -481
rect -3108 -583 -3074 -549
rect -3108 -636 -3074 -617
rect -3012 -447 -2978 -428
rect -3012 -515 -2978 -481
rect -3012 -583 -2978 -549
rect -3012 -636 -2978 -617
rect -2898 -447 -2864 -428
rect -2898 -515 -2864 -481
rect -2898 -583 -2864 -549
rect -2898 -636 -2864 -617
rect -2802 -447 -2768 -428
rect -2802 -515 -2768 -481
rect -2802 -583 -2768 -549
rect -2802 -636 -2768 -617
rect -2688 -447 -2654 -428
rect -2688 -515 -2654 -481
rect -2688 -583 -2654 -549
rect -2688 -636 -2654 -617
rect -2592 -447 -2558 -428
rect -2592 -515 -2558 -481
rect -2592 -583 -2558 -549
rect -2592 -636 -2558 -617
rect -2478 -447 -2444 -428
rect -2478 -515 -2444 -481
rect -2478 -583 -2444 -549
rect -2478 -636 -2444 -617
rect -2382 -447 -2348 -428
rect -2382 -515 -2348 -481
rect -2382 -583 -2348 -549
rect -2382 -636 -2348 -617
rect -2268 -447 -2234 -428
rect -2268 -515 -2234 -481
rect -2268 -583 -2234 -549
rect -2268 -636 -2234 -617
rect -2172 -447 -2138 -428
rect -2172 -515 -2138 -481
rect -2172 -583 -2138 -549
rect -2172 -636 -2138 -617
rect -2058 -447 -2024 -428
rect -2058 -515 -2024 -481
rect -2058 -583 -2024 -549
rect -2058 -636 -2024 -617
rect -1962 -447 -1928 -428
rect -1962 -515 -1928 -481
rect -1962 -583 -1928 -549
rect -1962 -636 -1928 -617
rect -1848 -447 -1814 -428
rect -1848 -515 -1814 -481
rect -1848 -583 -1814 -549
rect -1848 -636 -1814 -617
rect -1752 -447 -1718 -428
rect -1752 -515 -1718 -481
rect -1752 -583 -1718 -549
rect -1752 -636 -1718 -617
rect -1638 -447 -1604 -428
rect -1638 -515 -1604 -481
rect -1638 -583 -1604 -549
rect -1638 -636 -1604 -617
rect -1542 -447 -1508 -428
rect -1542 -515 -1508 -481
rect -1542 -583 -1508 -549
rect -1542 -636 -1508 -617
rect -1428 -447 -1394 -428
rect -1428 -515 -1394 -481
rect -1428 -583 -1394 -549
rect -1428 -636 -1394 -617
rect -1332 -447 -1298 -428
rect -1332 -515 -1298 -481
rect -1332 -583 -1298 -549
rect -1332 -636 -1298 -617
rect -1218 -447 -1184 -428
rect -1218 -515 -1184 -481
rect -1218 -583 -1184 -549
rect -1218 -636 -1184 -617
rect -1122 -447 -1088 -428
rect -1122 -515 -1088 -481
rect -1122 -583 -1088 -549
rect -1122 -636 -1088 -617
rect -1008 -447 -974 -428
rect -1008 -515 -974 -481
rect -1008 -583 -974 -549
rect -1008 -636 -974 -617
rect -912 -447 -878 -428
rect -912 -515 -878 -481
rect -912 -583 -878 -549
rect -912 -636 -878 -617
rect -798 -447 -764 -428
rect -798 -515 -764 -481
rect -798 -583 -764 -549
rect -798 -636 -764 -617
rect -702 -447 -668 -428
rect -702 -515 -668 -481
rect -702 -583 -668 -549
rect -702 -636 -668 -617
rect -588 -447 -554 -428
rect -588 -515 -554 -481
rect -588 -583 -554 -549
rect -588 -636 -554 -617
rect -492 -447 -458 -428
rect -492 -515 -458 -481
rect -492 -583 -458 -549
rect -492 -636 -458 -617
rect -378 -447 -344 -428
rect -378 -515 -344 -481
rect -378 -583 -344 -549
rect -378 -636 -344 -617
rect -282 -447 -248 -428
rect -282 -515 -248 -481
rect -282 -583 -248 -549
rect -282 -636 -248 -617
rect -168 -447 -134 -428
rect -168 -515 -134 -481
rect -168 -583 -134 -549
rect -168 -636 -134 -617
rect -72 -447 -38 -428
rect -72 -515 -38 -481
rect -72 -583 -38 -549
rect -72 -636 -38 -617
rect 42 -447 76 -428
rect 42 -515 76 -481
rect 42 -583 76 -549
rect 42 -636 76 -617
rect 138 -447 172 -428
rect 138 -515 172 -481
rect 138 -583 172 -549
rect 138 -636 172 -617
rect 252 -447 286 -428
rect 252 -515 286 -481
rect 252 -583 286 -549
rect 252 -636 286 -617
rect 348 -447 382 -428
rect 348 -515 382 -481
rect 348 -583 382 -549
rect 348 -636 382 -617
rect 462 -447 496 -428
rect 462 -515 496 -481
rect 462 -583 496 -549
rect 462 -636 496 -617
rect 558 -447 592 -428
rect 558 -515 592 -481
rect 558 -583 592 -549
rect 558 -636 592 -617
rect 672 -447 706 -428
rect 672 -515 706 -481
rect 672 -583 706 -549
rect 672 -636 706 -617
rect 768 -447 802 -428
rect 768 -515 802 -481
rect 768 -583 802 -549
rect 768 -636 802 -617
rect 882 -447 916 -428
rect 882 -515 916 -481
rect 882 -583 916 -549
rect 882 -636 916 -617
rect 978 -447 1012 -428
rect 978 -515 1012 -481
rect 978 -583 1012 -549
rect 978 -636 1012 -617
rect 1092 -447 1126 -428
rect 1092 -515 1126 -481
rect 1092 -583 1126 -549
rect 1092 -636 1126 -617
rect 1188 -447 1222 -428
rect 1188 -515 1222 -481
rect 1188 -583 1222 -549
rect 1188 -636 1222 -617
rect 1302 -447 1336 -428
rect 1302 -515 1336 -481
rect 1302 -583 1336 -549
rect 1302 -636 1336 -617
rect 1398 -447 1432 -428
rect 1398 -515 1432 -481
rect 1398 -583 1432 -549
rect 1398 -636 1432 -617
rect 1512 -447 1546 -428
rect 1512 -515 1546 -481
rect 1512 -583 1546 -549
rect 1512 -636 1546 -617
rect 1608 -447 1642 -428
rect 1608 -515 1642 -481
rect 1608 -583 1642 -549
rect 1608 -636 1642 -617
rect 1722 -447 1756 -428
rect 1722 -515 1756 -481
rect 1722 -583 1756 -549
rect 1722 -636 1756 -617
rect 1818 -447 1852 -428
rect 1818 -515 1852 -481
rect 1818 -583 1852 -549
rect 1818 -636 1852 -617
rect 1932 -447 1966 -428
rect 1932 -515 1966 -481
rect 1932 -583 1966 -549
rect 1932 -636 1966 -617
rect 2028 -447 2062 -428
rect 2028 -515 2062 -481
rect 2028 -583 2062 -549
rect 2028 -636 2062 -617
rect 2142 -447 2176 -428
rect 2142 -515 2176 -481
rect 2142 -583 2176 -549
rect 2142 -636 2176 -617
rect 2238 -447 2272 -428
rect 2238 -515 2272 -481
rect 2238 -583 2272 -549
rect 2238 -636 2272 -617
rect 2352 -447 2386 -428
rect 2352 -515 2386 -481
rect 2352 -583 2386 -549
rect 2352 -636 2386 -617
rect 2448 -447 2482 -428
rect 2448 -515 2482 -481
rect 2448 -583 2482 -549
rect 2448 -636 2482 -617
rect 2562 -447 2596 -428
rect 2562 -515 2596 -481
rect 2562 -583 2596 -549
rect 2562 -636 2596 -617
rect 2658 -447 2692 -428
rect 2658 -515 2692 -481
rect 2658 -583 2692 -549
rect 2658 -636 2692 -617
rect 2772 -447 2806 -428
rect 2772 -515 2806 -481
rect 2772 -583 2806 -549
rect 2772 -636 2806 -617
rect 2868 -447 2902 -428
rect 2868 -515 2902 -481
rect 2868 -583 2902 -549
rect 2868 -636 2902 -617
rect 2982 -447 3016 -428
rect 2982 -515 3016 -481
rect 2982 -583 3016 -549
rect 2982 -636 3016 -617
rect 3078 -447 3112 -428
rect 3078 -515 3112 -481
rect 3078 -583 3112 -549
rect 3078 -636 3112 -617
rect 3192 -447 3226 -428
rect 3192 -515 3226 -481
rect 3192 -583 3226 -549
rect 3192 -636 3226 -617
rect 3288 -447 3322 -428
rect 3288 -515 3322 -481
rect 3288 -583 3322 -549
rect 3288 -636 3322 -617
rect 3402 -447 3436 -428
rect 3402 -515 3436 -481
rect 3402 -583 3436 -549
rect 3402 -636 3436 -617
rect 3498 -447 3532 -428
rect 3498 -515 3532 -481
rect 3498 -583 3532 -549
rect 3498 -636 3532 -617
rect 3612 -447 3646 -428
rect 3612 -515 3646 -481
rect 3612 -583 3646 -549
rect 3612 -636 3646 -617
rect 3708 -447 3742 -428
rect 3708 -515 3742 -481
rect 3708 -583 3742 -549
rect 3708 -636 3742 -617
rect 3822 -447 3856 -428
rect 3822 -515 3856 -481
rect 3822 -583 3856 -549
rect 3822 -636 3856 -617
rect 3918 -447 3952 -428
rect 3918 -515 3952 -481
rect 3918 -583 3952 -549
rect 3918 -636 3952 -617
rect 4032 -447 4066 -428
rect 4032 -515 4066 -481
rect 4032 -583 4066 -549
rect 4032 -636 4066 -617
rect 4128 -447 4162 -428
rect 4128 -515 4162 -481
rect 4128 -583 4162 -549
rect 4128 -636 4162 -617
rect 4242 -447 4276 -385
rect 4242 -515 4276 -481
rect 4242 -583 4276 -549
rect 4242 -636 4276 -617
rect 4338 -447 4372 -385
rect 4338 -515 4372 -481
rect 4338 -583 4372 -549
rect 4338 -636 4372 -617
rect 4450 -413 4484 -385
rect 4450 -481 4484 -447
rect 4450 -549 4484 -515
rect 4450 -617 4484 -583
rect -4484 -685 -4320 -679
rect -4450 -713 -4320 -685
rect -4286 -713 -4238 -679
rect -3916 -713 -3900 -679
rect -3866 -713 -3850 -679
rect -3496 -713 -3480 -679
rect -3446 -713 -3430 -679
rect -3076 -713 -3060 -679
rect -3026 -713 -3010 -679
rect -2656 -713 -2640 -679
rect -2606 -713 -2590 -679
rect -2236 -713 -2220 -679
rect -2186 -713 -2170 -679
rect -1816 -713 -1800 -679
rect -1766 -713 -1750 -679
rect -1396 -713 -1380 -679
rect -1346 -713 -1330 -679
rect -976 -713 -960 -679
rect -926 -713 -910 -679
rect -556 -713 -540 -679
rect -506 -713 -490 -679
rect -136 -713 -120 -679
rect -86 -713 -70 -679
rect 284 -713 300 -679
rect 334 -713 350 -679
rect 704 -713 720 -679
rect 754 -713 770 -679
rect 1124 -713 1140 -679
rect 1174 -713 1190 -679
rect 1544 -713 1560 -679
rect 1594 -713 1610 -679
rect 1964 -713 1980 -679
rect 2014 -713 2030 -679
rect 2384 -713 2400 -679
rect 2434 -713 2450 -679
rect 2804 -713 2820 -679
rect 2854 -713 2870 -679
rect 3224 -713 3240 -679
rect 3274 -713 3290 -679
rect 3644 -713 3660 -679
rect 3694 -713 3710 -679
rect 4064 -713 4080 -679
rect 4114 -713 4130 -679
rect 4450 -685 4484 -651
rect -4484 -781 -4450 -719
rect 4450 -781 4484 -719
rect -4484 -815 -4369 -781
rect -4335 -815 -4301 -781
rect -4267 -815 -4233 -781
rect -4199 -815 -4165 -781
rect -4131 -815 -4097 -781
rect -4063 -815 -4029 -781
rect -3995 -815 -3961 -781
rect -3927 -815 -3893 -781
rect -3859 -815 -3825 -781
rect -3791 -815 -3757 -781
rect -3723 -815 -3689 -781
rect -3655 -815 -3621 -781
rect -3587 -815 -3553 -781
rect -3519 -815 -3485 -781
rect -3451 -815 -3417 -781
rect -3383 -815 -3349 -781
rect -3315 -815 -3281 -781
rect -3247 -815 -3213 -781
rect -3179 -815 -3145 -781
rect -3111 -815 -3077 -781
rect -3043 -815 -3009 -781
rect -2975 -815 -2941 -781
rect -2907 -815 -2873 -781
rect -2839 -815 -2805 -781
rect -2771 -815 -2737 -781
rect -2703 -815 -2669 -781
rect -2635 -815 -2601 -781
rect -2567 -815 -2533 -781
rect -2499 -815 -2465 -781
rect -2431 -815 -2397 -781
rect -2363 -815 -2329 -781
rect -2295 -815 -2261 -781
rect -2227 -815 -2193 -781
rect -2159 -815 -2125 -781
rect -2091 -815 -2057 -781
rect -2023 -815 -1989 -781
rect -1955 -815 -1921 -781
rect -1887 -815 -1853 -781
rect -1819 -815 -1785 -781
rect -1751 -815 -1717 -781
rect -1683 -815 -1649 -781
rect -1615 -815 -1581 -781
rect -1547 -815 -1513 -781
rect -1479 -815 -1445 -781
rect -1411 -815 -1377 -781
rect -1343 -815 -1309 -781
rect -1275 -815 -1241 -781
rect -1207 -815 -1173 -781
rect -1139 -815 -1105 -781
rect -1071 -815 -1037 -781
rect -1003 -815 -969 -781
rect -935 -815 -901 -781
rect -867 -815 -833 -781
rect -799 -815 -765 -781
rect -731 -815 -697 -781
rect -663 -815 -629 -781
rect -595 -815 -561 -781
rect -527 -815 -493 -781
rect -459 -815 -425 -781
rect -391 -815 -357 -781
rect -323 -815 -289 -781
rect -255 -815 -221 -781
rect -187 -815 -153 -781
rect -119 -815 -85 -781
rect -51 -815 -17 -781
rect 17 -815 51 -781
rect 85 -815 119 -781
rect 153 -815 187 -781
rect 221 -815 255 -781
rect 289 -815 323 -781
rect 357 -815 391 -781
rect 425 -815 459 -781
rect 493 -815 527 -781
rect 561 -815 595 -781
rect 629 -815 663 -781
rect 697 -815 731 -781
rect 765 -815 799 -781
rect 833 -815 867 -781
rect 901 -815 935 -781
rect 969 -815 1003 -781
rect 1037 -815 1071 -781
rect 1105 -815 1139 -781
rect 1173 -815 1207 -781
rect 1241 -815 1275 -781
rect 1309 -815 1343 -781
rect 1377 -815 1411 -781
rect 1445 -815 1479 -781
rect 1513 -815 1547 -781
rect 1581 -815 1615 -781
rect 1649 -815 1683 -781
rect 1717 -815 1751 -781
rect 1785 -815 1819 -781
rect 1853 -815 1887 -781
rect 1921 -815 1955 -781
rect 1989 -815 2023 -781
rect 2057 -815 2091 -781
rect 2125 -815 2159 -781
rect 2193 -815 2227 -781
rect 2261 -815 2295 -781
rect 2329 -815 2363 -781
rect 2397 -815 2431 -781
rect 2465 -815 2499 -781
rect 2533 -815 2567 -781
rect 2601 -815 2635 -781
rect 2669 -815 2703 -781
rect 2737 -815 2771 -781
rect 2805 -815 2839 -781
rect 2873 -815 2907 -781
rect 2941 -815 2975 -781
rect 3009 -815 3043 -781
rect 3077 -815 3111 -781
rect 3145 -815 3179 -781
rect 3213 -815 3247 -781
rect 3281 -815 3315 -781
rect 3349 -815 3383 -781
rect 3417 -815 3451 -781
rect 3485 -815 3519 -781
rect 3553 -815 3587 -781
rect 3621 -815 3655 -781
rect 3689 -815 3723 -781
rect 3757 -815 3791 -781
rect 3825 -815 3859 -781
rect 3893 -815 3927 -781
rect 3961 -815 3995 -781
rect 4029 -815 4063 -781
rect 4097 -815 4131 -781
rect 4165 -815 4199 -781
rect 4233 -815 4267 -781
rect 4301 -815 4335 -781
rect 4369 -815 4484 -781
<< viali >>
rect -4112 147 -4078 181
rect -3692 147 -3658 181
rect -3272 147 -3238 181
rect -2852 147 -2818 181
rect -2432 147 -2398 181
rect -2012 147 -1978 181
rect -1592 147 -1558 181
rect -1172 147 -1138 181
rect -752 147 -718 181
rect -332 147 -298 181
rect 88 147 122 181
rect 508 147 542 181
rect 928 147 962 181
rect 1348 147 1382 181
rect 1768 147 1802 181
rect 2188 147 2222 181
rect 2608 147 2642 181
rect 3028 147 3062 181
rect 3448 147 3482 181
rect 3868 147 3902 181
rect -3902 -181 -3868 -147
rect -3482 -181 -3448 -147
rect -3062 -181 -3028 -147
rect -2642 -181 -2608 -147
rect -2222 -181 -2188 -147
rect -1802 -181 -1768 -147
rect -1382 -181 -1348 -147
rect -962 -181 -928 -147
rect -542 -181 -508 -147
rect -122 -181 -88 -147
rect 298 -181 332 -147
rect 718 -181 752 -147
rect 1138 -181 1172 -147
rect 1558 -181 1592 -147
rect 1978 -181 2012 -147
rect 2398 -181 2432 -147
rect 2818 -181 2852 -147
rect 3238 -181 3272 -147
rect 3658 -181 3692 -147
rect 4078 -181 4112 -147
rect -4110 -385 -4076 -351
rect -3690 -385 -3656 -351
rect -3270 -385 -3236 -351
rect -2850 -385 -2816 -351
rect -2430 -385 -2396 -351
rect -2010 -385 -1976 -351
rect -1590 -385 -1556 -351
rect -1170 -385 -1136 -351
rect -750 -385 -716 -351
rect -330 -385 -296 -351
rect 90 -385 124 -351
rect 510 -385 544 -351
rect 930 -385 964 -351
rect 1350 -385 1384 -351
rect 1770 -385 1804 -351
rect 2190 -385 2224 -351
rect 2610 -385 2644 -351
rect 3030 -385 3064 -351
rect 3450 -385 3484 -351
rect 3870 -385 3904 -351
rect -3900 -713 -3866 -679
rect -3480 -713 -3446 -679
rect -3060 -713 -3026 -679
rect -2640 -713 -2606 -679
rect -2220 -713 -2186 -679
rect -1800 -713 -1766 -679
rect -1380 -713 -1346 -679
rect -960 -713 -926 -679
rect -540 -713 -506 -679
rect -120 -713 -86 -679
rect 300 -713 334 -679
rect 720 -713 754 -679
rect 1140 -713 1174 -679
rect 1560 -713 1594 -679
rect 1980 -713 2014 -679
rect 2400 -713 2434 -679
rect 2820 -713 2854 -679
rect 3240 -713 3274 -679
rect 3660 -713 3694 -679
rect 4080 -713 4114 -679
<< metal1 >>
rect -4124 181 -4066 187
rect -4124 147 -4112 181
rect -4078 147 -4066 181
rect -4124 141 -4066 147
rect -3704 181 -3646 187
rect -3704 147 -3692 181
rect -3658 147 -3646 181
rect -3704 141 -3646 147
rect -3284 181 -3226 187
rect -3284 147 -3272 181
rect -3238 147 -3226 181
rect -3284 141 -3226 147
rect -2864 181 -2806 187
rect -2864 147 -2852 181
rect -2818 147 -2806 181
rect -2864 141 -2806 147
rect -2444 181 -2386 187
rect -2444 147 -2432 181
rect -2398 147 -2386 181
rect -2444 141 -2386 147
rect -2024 181 -1966 187
rect -2024 147 -2012 181
rect -1978 147 -1966 181
rect -2024 141 -1966 147
rect -1604 181 -1546 187
rect -1604 147 -1592 181
rect -1558 147 -1546 181
rect -1604 141 -1546 147
rect -1184 181 -1126 187
rect -1184 147 -1172 181
rect -1138 147 -1126 181
rect -1184 141 -1126 147
rect -764 181 -706 187
rect -764 147 -752 181
rect -718 147 -706 181
rect -764 141 -706 147
rect -344 181 -286 187
rect -344 147 -332 181
rect -298 147 -286 181
rect -344 141 -286 147
rect 76 181 134 187
rect 76 147 88 181
rect 122 147 134 181
rect 76 141 134 147
rect 496 181 554 187
rect 496 147 508 181
rect 542 147 554 181
rect 496 141 554 147
rect 916 181 974 187
rect 916 147 928 181
rect 962 147 974 181
rect 916 141 974 147
rect 1336 181 1394 187
rect 1336 147 1348 181
rect 1382 147 1394 181
rect 1336 141 1394 147
rect 1756 181 1814 187
rect 1756 147 1768 181
rect 1802 147 1814 181
rect 1756 141 1814 147
rect 2176 181 2234 187
rect 2176 147 2188 181
rect 2222 147 2234 181
rect 2176 141 2234 147
rect 2596 181 2654 187
rect 2596 147 2608 181
rect 2642 147 2654 181
rect 2596 141 2654 147
rect 3016 181 3074 187
rect 3016 147 3028 181
rect 3062 147 3074 181
rect 3016 141 3074 147
rect 3436 181 3494 187
rect 3436 147 3448 181
rect 3482 147 3494 181
rect 3436 141 3494 147
rect 3856 181 3914 187
rect 3856 147 3868 181
rect 3902 147 3914 181
rect 3856 141 3914 147
rect -3914 -147 -3856 -141
rect -3914 -181 -3902 -147
rect -3868 -181 -3856 -147
rect -3914 -187 -3856 -181
rect -3494 -147 -3436 -141
rect -3494 -181 -3482 -147
rect -3448 -181 -3436 -147
rect -3494 -187 -3436 -181
rect -3074 -147 -3016 -141
rect -3074 -181 -3062 -147
rect -3028 -181 -3016 -147
rect -3074 -187 -3016 -181
rect -2654 -147 -2596 -141
rect -2654 -181 -2642 -147
rect -2608 -181 -2596 -147
rect -2654 -187 -2596 -181
rect -2234 -147 -2176 -141
rect -2234 -181 -2222 -147
rect -2188 -181 -2176 -147
rect -2234 -187 -2176 -181
rect -1814 -147 -1756 -141
rect -1814 -181 -1802 -147
rect -1768 -181 -1756 -147
rect -1814 -187 -1756 -181
rect -1394 -147 -1336 -141
rect -1394 -181 -1382 -147
rect -1348 -181 -1336 -147
rect -1394 -187 -1336 -181
rect -974 -147 -916 -141
rect -974 -181 -962 -147
rect -928 -181 -916 -147
rect -974 -187 -916 -181
rect -554 -147 -496 -141
rect -554 -181 -542 -147
rect -508 -181 -496 -147
rect -554 -187 -496 -181
rect -134 -147 -76 -141
rect -134 -181 -122 -147
rect -88 -181 -76 -147
rect -134 -187 -76 -181
rect 286 -147 344 -141
rect 286 -181 298 -147
rect 332 -181 344 -147
rect 286 -187 344 -181
rect 706 -147 764 -141
rect 706 -181 718 -147
rect 752 -181 764 -147
rect 706 -187 764 -181
rect 1126 -147 1184 -141
rect 1126 -181 1138 -147
rect 1172 -181 1184 -147
rect 1126 -187 1184 -181
rect 1546 -147 1604 -141
rect 1546 -181 1558 -147
rect 1592 -181 1604 -147
rect 1546 -187 1604 -181
rect 1966 -147 2024 -141
rect 1966 -181 1978 -147
rect 2012 -181 2024 -147
rect 1966 -187 2024 -181
rect 2386 -147 2444 -141
rect 2386 -181 2398 -147
rect 2432 -181 2444 -147
rect 2386 -187 2444 -181
rect 2806 -147 2864 -141
rect 2806 -181 2818 -147
rect 2852 -181 2864 -147
rect 2806 -187 2864 -181
rect 3226 -147 3284 -141
rect 3226 -181 3238 -147
rect 3272 -181 3284 -147
rect 3226 -187 3284 -181
rect 3646 -147 3704 -141
rect 3646 -181 3658 -147
rect 3692 -181 3704 -147
rect 3646 -187 3704 -181
rect 4066 -147 4124 -141
rect 4066 -181 4078 -147
rect 4112 -181 4124 -147
rect 4066 -187 4124 -181
rect -4122 -351 -4064 -345
rect -4122 -385 -4110 -351
rect -4076 -385 -4064 -351
rect -4122 -391 -4064 -385
rect -3702 -351 -3644 -345
rect -3702 -385 -3690 -351
rect -3656 -385 -3644 -351
rect -3702 -391 -3644 -385
rect -3282 -351 -3224 -345
rect -3282 -385 -3270 -351
rect -3236 -385 -3224 -351
rect -3282 -391 -3224 -385
rect -2862 -351 -2804 -345
rect -2862 -385 -2850 -351
rect -2816 -385 -2804 -351
rect -2862 -391 -2804 -385
rect -2442 -351 -2384 -345
rect -2442 -385 -2430 -351
rect -2396 -385 -2384 -351
rect -2442 -391 -2384 -385
rect -2022 -351 -1964 -345
rect -2022 -385 -2010 -351
rect -1976 -385 -1964 -351
rect -2022 -391 -1964 -385
rect -1602 -351 -1544 -345
rect -1602 -385 -1590 -351
rect -1556 -385 -1544 -351
rect -1602 -391 -1544 -385
rect -1182 -351 -1124 -345
rect -1182 -385 -1170 -351
rect -1136 -385 -1124 -351
rect -1182 -391 -1124 -385
rect -762 -351 -704 -345
rect -762 -385 -750 -351
rect -716 -385 -704 -351
rect -762 -391 -704 -385
rect -342 -351 -284 -345
rect -342 -385 -330 -351
rect -296 -385 -284 -351
rect -342 -391 -284 -385
rect 78 -351 136 -345
rect 78 -385 90 -351
rect 124 -385 136 -351
rect 78 -391 136 -385
rect 498 -351 556 -345
rect 498 -385 510 -351
rect 544 -385 556 -351
rect 498 -391 556 -385
rect 918 -351 976 -345
rect 918 -385 930 -351
rect 964 -385 976 -351
rect 918 -391 976 -385
rect 1338 -351 1396 -345
rect 1338 -385 1350 -351
rect 1384 -385 1396 -351
rect 1338 -391 1396 -385
rect 1758 -351 1816 -345
rect 1758 -385 1770 -351
rect 1804 -385 1816 -351
rect 1758 -391 1816 -385
rect 2178 -351 2236 -345
rect 2178 -385 2190 -351
rect 2224 -385 2236 -351
rect 2178 -391 2236 -385
rect 2598 -351 2656 -345
rect 2598 -385 2610 -351
rect 2644 -385 2656 -351
rect 2598 -391 2656 -385
rect 3018 -351 3076 -345
rect 3018 -385 3030 -351
rect 3064 -385 3076 -351
rect 3018 -391 3076 -385
rect 3438 -351 3496 -345
rect 3438 -385 3450 -351
rect 3484 -385 3496 -351
rect 3438 -391 3496 -385
rect 3858 -351 3916 -345
rect 3858 -385 3870 -351
rect 3904 -385 3916 -351
rect 3858 -391 3916 -385
rect -3912 -679 -3854 -673
rect -3912 -713 -3900 -679
rect -3866 -713 -3854 -679
rect -3912 -719 -3854 -713
rect -3492 -679 -3434 -673
rect -3492 -713 -3480 -679
rect -3446 -713 -3434 -679
rect -3492 -719 -3434 -713
rect -3072 -679 -3014 -673
rect -3072 -713 -3060 -679
rect -3026 -713 -3014 -679
rect -3072 -719 -3014 -713
rect -2652 -679 -2594 -673
rect -2652 -713 -2640 -679
rect -2606 -713 -2594 -679
rect -2652 -719 -2594 -713
rect -2232 -679 -2174 -673
rect -2232 -713 -2220 -679
rect -2186 -713 -2174 -679
rect -2232 -719 -2174 -713
rect -1812 -679 -1754 -673
rect -1812 -713 -1800 -679
rect -1766 -713 -1754 -679
rect -1812 -719 -1754 -713
rect -1392 -679 -1334 -673
rect -1392 -713 -1380 -679
rect -1346 -713 -1334 -679
rect -1392 -719 -1334 -713
rect -972 -679 -914 -673
rect -972 -713 -960 -679
rect -926 -713 -914 -679
rect -972 -719 -914 -713
rect -552 -679 -494 -673
rect -552 -713 -540 -679
rect -506 -713 -494 -679
rect -552 -719 -494 -713
rect -132 -679 -74 -673
rect -132 -713 -120 -679
rect -86 -713 -74 -679
rect -132 -719 -74 -713
rect 288 -679 346 -673
rect 288 -713 300 -679
rect 334 -713 346 -679
rect 288 -719 346 -713
rect 708 -679 766 -673
rect 708 -713 720 -679
rect 754 -713 766 -679
rect 708 -719 766 -713
rect 1128 -679 1186 -673
rect 1128 -713 1140 -679
rect 1174 -713 1186 -679
rect 1128 -719 1186 -713
rect 1548 -679 1606 -673
rect 1548 -713 1560 -679
rect 1594 -713 1606 -679
rect 1548 -719 1606 -713
rect 1968 -679 2026 -673
rect 1968 -713 1980 -679
rect 2014 -713 2026 -679
rect 1968 -719 2026 -713
rect 2388 -679 2446 -673
rect 2388 -713 2400 -679
rect 2434 -713 2446 -679
rect 2388 -719 2446 -713
rect 2808 -679 2866 -673
rect 2808 -713 2820 -679
rect 2854 -713 2866 -679
rect 2808 -719 2866 -713
rect 3228 -679 3286 -673
rect 3228 -713 3240 -679
rect 3274 -713 3286 -679
rect 3228 -719 3286 -713
rect 3648 -679 3706 -673
rect 3648 -713 3660 -679
rect 3694 -713 3706 -679
rect 3648 -719 3706 -713
rect 4068 -679 4126 -673
rect 4068 -713 4080 -679
rect 4114 -713 4126 -679
rect 4068 -719 4126 -713
<< properties >>
string FIXED_BBOX -4467 -266 4467 266
<< end >>
