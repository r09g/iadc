magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< nwell >>
rect -455 -558 455 338
<< pmos >>
rect -255 -49 -225 51
rect -159 -49 -129 51
rect -63 -49 -33 51
rect 33 -49 63 51
rect 129 -49 159 51
rect 225 -49 255 51
rect -255 -271 -225 -171
rect -159 -271 -129 -171
rect -63 -271 -33 -171
rect 33 -271 63 -171
rect 129 -271 159 -171
rect 225 -271 255 -171
<< pdiff >>
rect -317 39 -255 51
rect -317 -37 -305 39
rect -271 -37 -255 39
rect -317 -49 -255 -37
rect -225 39 -159 51
rect -225 -37 -209 39
rect -175 -37 -159 39
rect -225 -49 -159 -37
rect -129 39 -63 51
rect -129 -37 -113 39
rect -79 -37 -63 39
rect -129 -49 -63 -37
rect -33 39 33 51
rect -33 -37 -17 39
rect 17 -37 33 39
rect -33 -49 33 -37
rect 63 39 129 51
rect 63 -37 79 39
rect 113 -37 129 39
rect 63 -49 129 -37
rect 159 39 225 51
rect 159 -37 175 39
rect 209 -37 225 39
rect 159 -49 225 -37
rect 255 39 317 51
rect 255 -37 271 39
rect 305 -37 317 39
rect 255 -49 317 -37
rect -317 -183 -255 -171
rect -317 -259 -305 -183
rect -271 -259 -255 -183
rect -317 -271 -255 -259
rect -225 -183 -159 -171
rect -225 -259 -209 -183
rect -175 -259 -159 -183
rect -225 -271 -159 -259
rect -129 -183 -63 -171
rect -129 -259 -113 -183
rect -79 -259 -63 -183
rect -129 -271 -63 -259
rect -33 -183 33 -171
rect -33 -259 -17 -183
rect 17 -259 33 -183
rect -33 -271 33 -259
rect 63 -183 129 -171
rect 63 -259 79 -183
rect 113 -259 129 -183
rect 63 -271 129 -259
rect 159 -183 225 -171
rect 159 -259 175 -183
rect 209 -259 225 -183
rect 159 -271 225 -259
rect 255 -183 317 -171
rect 255 -259 271 -183
rect 305 -259 317 -183
rect 255 -271 317 -259
<< pdiffc >>
rect -305 -37 -271 39
rect -209 -37 -175 39
rect -113 -37 -79 39
rect -17 -37 17 39
rect 79 -37 113 39
rect 175 -37 209 39
rect 271 -37 305 39
rect -305 -259 -271 -183
rect -209 -259 -175 -183
rect -113 -259 -79 -183
rect -17 -259 17 -183
rect 79 -259 113 -183
rect 175 -259 209 -183
rect 271 -259 305 -183
<< nsubdiff >>
rect -419 268 -323 302
rect 323 268 419 302
rect -419 206 -385 268
rect 385 206 419 268
rect -419 -488 -385 -426
rect 385 -488 419 -426
rect -419 -522 -323 -488
rect 323 -522 419 -488
<< nsubdiffcont >>
rect -323 268 323 302
rect -419 -426 -385 206
rect 385 -426 419 206
rect -323 -522 323 -488
<< poly >>
rect -63 200 63 216
rect -63 166 -17 200
rect 17 166 63 200
rect -63 150 63 166
rect -291 132 -225 148
rect -291 98 -275 132
rect -241 98 -225 132
rect -291 82 -225 98
rect -177 132 -111 148
rect -177 98 -161 132
rect -127 98 -111 132
rect -177 82 -111 98
rect -255 51 -225 82
rect -159 51 -129 82
rect -63 51 -33 150
rect 33 51 63 150
rect 111 132 177 148
rect 111 98 127 132
rect 161 98 177 132
rect 111 82 177 98
rect 225 132 291 148
rect 225 98 241 132
rect 275 98 291 132
rect 225 82 291 98
rect 129 51 159 82
rect 225 51 255 82
rect -255 -75 -225 -49
rect -159 -75 -129 -49
rect -63 -75 -33 -49
rect 33 -75 63 -49
rect 129 -75 159 -49
rect 225 -75 255 -49
rect -255 -171 -225 -145
rect -159 -171 -129 -145
rect -63 -171 -33 -145
rect 33 -171 63 -145
rect 129 -171 159 -145
rect 225 -171 255 -145
rect -255 -302 -225 -271
rect -159 -302 -129 -271
rect -291 -318 -225 -302
rect -291 -352 -275 -318
rect -241 -352 -225 -318
rect -291 -368 -225 -352
rect -177 -318 -111 -302
rect -177 -352 -161 -318
rect -127 -352 -111 -318
rect -177 -368 -111 -352
rect -63 -370 -33 -271
rect 33 -370 63 -271
rect 129 -302 159 -271
rect 225 -302 255 -271
rect 111 -318 177 -302
rect 111 -352 127 -318
rect 161 -352 177 -318
rect 111 -368 177 -352
rect 225 -318 291 -302
rect 225 -352 241 -318
rect 275 -352 291 -318
rect 225 -368 291 -352
rect -63 -386 63 -370
rect -63 -420 -17 -386
rect 17 -420 63 -386
rect -63 -436 63 -420
<< polycont >>
rect -17 166 17 200
rect -275 98 -241 132
rect -161 98 -127 132
rect 127 98 161 132
rect 241 98 275 132
rect -275 -352 -241 -318
rect -161 -352 -127 -318
rect 127 -352 161 -318
rect 241 -352 275 -318
rect -17 -420 17 -386
<< locali >>
rect -419 268 -323 302
rect 323 268 419 302
rect -419 206 -385 268
rect 385 206 419 268
rect -33 166 -17 200
rect 17 166 33 200
rect -385 98 -275 132
rect -241 98 -225 132
rect -177 98 -161 132
rect -127 98 -111 132
rect 111 98 127 132
rect 161 98 177 132
rect 225 98 241 132
rect 275 98 385 132
rect -305 39 -271 98
rect -305 -53 -271 -37
rect -209 47 -175 55
rect -209 -53 -175 -37
rect -113 39 -79 55
rect -113 -93 -79 -37
rect -17 39 17 55
rect 79 39 113 55
rect -305 -183 -271 -167
rect -305 -318 -271 -259
rect -209 -183 -175 -167
rect -209 -275 -175 -267
rect -113 -183 -79 -127
rect 79 -93 113 -37
rect 175 47 209 55
rect 175 -53 209 -37
rect 271 39 305 98
rect 271 -53 305 -37
rect -113 -275 -79 -259
rect -17 -275 17 -259
rect 79 -183 113 -127
rect 79 -275 113 -259
rect 175 -183 209 -167
rect 175 -275 209 -267
rect 271 -183 305 -167
rect 271 -318 305 -259
rect -385 -352 -275 -318
rect -241 -352 -225 -318
rect -177 -352 -161 -318
rect -127 -352 -111 -318
rect 111 -352 127 -318
rect 161 -352 177 -318
rect 225 -352 241 -318
rect 275 -352 385 -318
rect -33 -420 -17 -386
rect 17 -420 33 -386
rect -419 -488 -385 -426
rect 385 -488 419 -426
rect -419 -522 -323 -488
rect 323 -522 419 -488
<< viali >>
rect -17 268 17 302
rect -17 166 17 200
rect -161 98 -127 132
rect 127 98 161 132
rect -209 39 -175 47
rect -209 13 -175 39
rect -17 -37 17 -21
rect -17 -55 17 -37
rect -113 -127 -79 -93
rect -209 -259 -175 -233
rect -209 -267 -175 -259
rect 175 39 209 47
rect 175 13 209 39
rect 79 -127 113 -93
rect -17 -183 17 -165
rect -17 -199 17 -183
rect 175 -259 209 -233
rect 175 -267 209 -259
rect -161 -352 -127 -318
rect 127 -352 161 -318
rect -17 -420 17 -386
<< metal1 >>
rect -37 258 -27 310
rect 27 258 37 310
rect -303 200 -293 218
rect -455 166 -293 200
rect -241 200 -231 218
rect -29 200 29 206
rect -241 166 -17 200
rect 17 166 63 200
rect -29 160 29 166
rect -173 132 -115 138
rect 115 132 173 138
rect 231 132 241 150
rect -177 98 -161 132
rect -127 98 127 132
rect 161 98 241 132
rect 293 132 303 150
rect 293 98 455 132
rect -173 92 -115 98
rect 115 92 173 98
rect -221 47 -163 53
rect 163 47 221 53
rect -221 13 -209 47
rect -175 13 175 47
rect 209 13 455 47
rect -221 7 -163 13
rect 163 7 221 13
rect -29 -21 29 -15
rect -455 -55 -17 -21
rect 17 -55 29 -21
rect -305 -233 -271 -55
rect -29 -61 29 -55
rect -133 -135 -123 -83
rect -71 -93 -61 -83
rect 61 -93 71 -83
rect -71 -127 71 -93
rect -71 -135 -61 -127
rect 61 -135 71 -127
rect 123 -135 133 -83
rect -29 -165 29 -159
rect 271 -165 305 13
rect -29 -199 -17 -165
rect 17 -199 305 -165
rect -29 -205 29 -199
rect -221 -233 -163 -227
rect 163 -233 221 -227
rect -305 -267 -209 -233
rect -175 -267 175 -233
rect 209 -267 221 -233
rect -221 -273 -163 -267
rect 163 -273 221 -267
rect -173 -318 -115 -312
rect 115 -318 173 -312
rect -303 -370 -293 -318
rect -241 -352 -161 -318
rect -127 -352 127 -318
rect 161 -352 177 -318
rect -241 -370 -231 -352
rect -173 -358 -115 -352
rect 115 -358 173 -352
rect -29 -386 29 -380
rect -63 -420 -17 -386
rect 17 -420 241 -386
rect -29 -426 29 -420
rect 231 -438 241 -420
rect 293 -438 303 -386
<< via1 >>
rect -27 302 27 310
rect -27 268 -17 302
rect -17 268 17 302
rect 17 268 27 302
rect -27 258 27 268
rect -293 166 -241 218
rect 241 98 293 150
rect -123 -93 -71 -83
rect 71 -93 123 -83
rect -123 -127 -113 -93
rect -113 -127 -79 -93
rect -79 -127 -71 -93
rect 71 -127 79 -93
rect 79 -127 113 -93
rect 113 -127 123 -93
rect -123 -135 -71 -127
rect 71 -135 123 -127
rect -293 -370 -241 -318
rect 241 -438 293 -386
<< metal2 >>
rect -27 310 27 320
rect -293 218 -241 228
rect -293 -318 -241 166
rect -27 -83 27 258
rect 241 150 293 160
rect -129 -135 -123 -83
rect -71 -135 71 -83
rect 123 -135 129 -83
rect -293 -380 -241 -370
rect 241 -386 293 98
rect 241 -448 293 -438
<< properties >>
string FIXED_BBOX -402 -206 402 206
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
