magic
tech sky130A
magscale 1 2
timestamp 1653437277
<< nwell >>
rect -51 2940 246 3012
rect 417 3000 983 3284
rect 866 2991 983 3000
rect 1136 2940 1501 3012
rect -51 2936 1501 2940
rect -51 2117 246 2936
rect 1136 2192 1501 2936
rect 1154 2117 1501 2192
<< pwell >>
rect 204 3077 339 4732
rect 1061 3077 1196 4732
rect -40 1884 36 1997
rect -128 1831 36 1884
rect -40 1717 36 1831
rect 1364 1883 1440 1997
rect 1364 1827 1585 1883
rect 1364 1717 1440 1827
rect 293 749 389 795
<< viali >>
rect 378 3957 412 3991
rect 987 3958 1021 3992
rect 445 3841 479 3875
rect 921 3841 955 3875
rect 377 3514 411 3548
rect 989 3529 1023 3563
rect 377 3306 411 3340
rect 987 3306 1021 3340
rect 371 3114 405 3148
rect 995 3114 1029 3148
rect 377 2943 1023 2977
rect -4 1729 30 1985
rect 1370 1729 1404 1985
rect 377 1527 1023 1561
rect 377 755 1023 789
rect 184 235 1214 269
<< metal1 >>
rect 108 4036 204 4870
rect 266 3881 300 4870
rect 652 4018 748 4870
rect 359 3947 369 3999
rect 421 3947 431 3999
rect 853 3947 863 3999
rect 915 3947 925 3999
rect 967 3949 977 4001
rect 1029 3949 1039 4001
rect 517 3881 527 3884
rect 266 3875 527 3881
rect 266 3841 445 3875
rect 479 3841 527 3875
rect 266 3835 527 3841
rect 517 3832 527 3835
rect 579 3832 589 3884
rect 867 3881 911 3947
rect 1100 3881 1134 4870
rect 1196 3976 1292 4870
rect 867 3875 1134 3881
rect 867 3841 921 3875
rect 955 3841 1134 3875
rect 867 3835 1134 3841
rect 977 3563 1035 3569
rect 365 3548 423 3556
rect 365 3514 377 3548
rect 411 3514 423 3548
rect 365 3340 423 3514
rect 977 3529 989 3563
rect 1023 3529 1035 3563
rect 977 3523 1035 3529
rect 977 3346 1033 3523
rect 365 3306 377 3340
rect 411 3306 423 3340
rect 365 3300 423 3306
rect 975 3340 1033 3346
rect 975 3306 987 3340
rect 1021 3306 1033 3340
rect 975 3300 1033 3306
rect 350 3105 360 3157
rect 412 3105 422 3157
rect 974 3106 984 3158
rect 1036 3106 1046 3158
rect 652 2983 748 3088
rect 245 2979 1155 2983
rect 245 2977 1365 2979
rect 85 2943 377 2977
rect 1023 2945 1365 2977
rect 1023 2943 1155 2945
rect -31 2578 -21 2630
rect 31 2578 41 2630
rect 85 2560 119 2943
rect 245 2936 1155 2943
rect 1149 2670 1159 2722
rect 1211 2670 1221 2722
rect 167 2602 245 2654
rect 297 2602 307 2654
rect -171 2473 161 2507
rect 1149 2357 1159 2366
rect 788 2323 1159 2357
rect 1149 2314 1159 2323
rect 1211 2357 1269 2366
rect 1211 2323 1277 2357
rect 1211 2314 1269 2323
rect 235 2255 245 2264
rect 158 2221 245 2255
rect -40 1985 36 1997
rect -40 1884 -4 1985
rect -128 1831 -4 1884
rect -40 1729 -4 1831
rect 30 1729 36 1985
rect 158 1769 192 2221
rect 235 2212 245 2221
rect 297 2255 307 2264
rect 523 2255 820 2288
rect 1331 2287 1365 2945
rect 1409 2303 1419 2355
rect 1471 2303 1481 2355
rect 297 2221 557 2255
rect 297 2212 307 2221
rect 1289 2198 1571 2232
rect 1364 1985 1440 1997
rect 352 1945 1278 1979
rect 158 1735 838 1769
rect -40 1717 36 1729
rect 1364 1729 1370 1985
rect 1404 1883 1440 1985
rect 1404 1827 1585 1883
rect 1404 1729 1440 1827
rect 1364 1717 1440 1729
rect -171 1561 1571 1567
rect -171 1527 377 1561
rect 1023 1527 1571 1561
rect -171 1521 1571 1527
rect -171 1425 386 1459
rect 1121 1357 1571 1391
rect 235 1213 245 1265
rect 297 1213 307 1265
rect 1093 1263 1103 1315
rect 1155 1263 1165 1315
rect -171 789 1571 795
rect -171 755 377 789
rect 1023 755 1571 789
rect -171 749 1571 755
rect 664 433 674 485
rect 726 433 736 485
rect -171 337 1050 371
rect -147 269 1571 275
rect -147 235 184 269
rect 1214 235 1571 269
rect -147 229 1571 235
<< via1 >>
rect 369 3991 421 3999
rect 369 3957 378 3991
rect 378 3957 412 3991
rect 412 3957 421 3991
rect 369 3947 421 3957
rect 863 3947 915 3999
rect 977 3992 1029 4001
rect 977 3958 987 3992
rect 987 3958 1021 3992
rect 1021 3958 1029 3992
rect 977 3949 1029 3958
rect 527 3832 579 3884
rect 360 3148 412 3157
rect 360 3114 371 3148
rect 371 3114 405 3148
rect 405 3114 412 3148
rect 360 3105 412 3114
rect 984 3148 1036 3158
rect 984 3114 995 3148
rect 995 3114 1029 3148
rect 1029 3114 1036 3148
rect 984 3106 1036 3114
rect -21 2578 31 2630
rect 1159 2670 1211 2722
rect 245 2602 297 2654
rect 1159 2314 1211 2366
rect 245 2212 297 2264
rect 1419 2303 1471 2355
rect 245 1213 297 1265
rect 1103 1263 1155 1315
rect 674 433 726 485
<< metal2 >>
rect 369 3999 421 4009
rect 863 3999 915 4009
rect 421 3947 863 3999
rect 369 3937 421 3947
rect 863 3937 915 3947
rect 977 4001 1029 4011
rect 527 3884 579 3894
rect 977 3884 1029 3949
rect 579 3832 1029 3884
rect 527 3822 579 3832
rect 360 3157 412 3167
rect 245 3105 360 3151
rect 984 3158 1036 3168
rect 412 3105 428 3151
rect 245 3099 428 3105
rect 973 3106 984 3154
rect 1036 3106 1211 3154
rect 973 3102 1211 3106
rect 245 2654 297 3099
rect 360 3095 412 3099
rect 984 3096 1036 3102
rect -21 2630 31 2640
rect -21 1769 31 2578
rect 245 2264 297 2602
rect 245 2007 297 2212
rect 1159 2722 1211 3102
rect 1159 2366 1211 2670
rect 245 1973 479 2007
rect 1159 1945 1211 2314
rect 1419 2355 1471 2365
rect -21 1735 297 1769
rect -21 1726 31 1735
rect 245 1265 297 1735
rect 1419 1711 1471 2303
rect 1103 1315 1155 1711
rect 1253 1677 1471 1711
rect 1419 1667 1471 1677
rect 1103 1253 1155 1263
rect 245 1203 297 1213
rect 674 485 726 816
rect 674 423 726 433
use input_diff_pair  input_diff_pair_0
timestamp 1653369986
transform 1 0 700 0 1 1267
box -455 -548 455 330
use latch_nmos_pair  latch_nmos_pair_0
timestamp 1653369027
transform 1 0 700 0 1 1857
box -740 -260 740 260
use latch_pmos_pair  latch_pmos_pair_0
timestamp 1653369027
transform 1 0 700 0 1 2675
box -455 -558 455 338
use nfet_tail_current_source  nfet_tail_current_source_0
timestamp 1653369027
transform -1 0 699 0 -1 459
box -647 -261 647 261
use sky130_fd_pr__pfet_01v8_8EMFFC  sky130_fd_pr__pfet_01v8_8EMFFC_0
timestamp 1653369027
transform -1 0 1392 0 -1 2329
box -108 -88 196 150
use sky130_fd_pr__pfet_01v8_8EMFFC  sky130_fd_pr__pfet_01v8_8EMFFC_1
timestamp 1653369027
transform -1 0 144 0 -1 2604
box -108 -88 196 150
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 -1 1244 1 0 3077
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1650294714
transform 0 1 156 1 0 3077
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 1 156 -1 0 4733
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1650294714
transform 0 -1 1244 1 0 4365
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 1 156 -1 0 4273
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_1
timestamp 1650294714
transform 0 -1 1244 -1 0 4273
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 1 156 -1 0 4365
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform 0 -1 1244 1 0 4273
box -38 -48 130 592
<< labels >>
flabel metal1 283 4868 283 4868 5 FreeSans 400 0 0 0 outp
flabel metal1 1117 4868 1117 4868 5 FreeSans 400 0 0 0 outn
flabel metal1 -166 2489 -166 2489 3 FreeSans 400 0 0 0 clk
flabel metal1 1564 2214 1564 2214 1 FreeSans 400 0 0 0 clk
flabel metal1 -123 1858 -123 1858 1 FreeSans 400 0 0 0 VSS
flabel metal1 1582 1855 1582 1855 7 FreeSans 400 0 0 0 VSS
flabel metal1 -166 1544 -166 1544 3 FreeSans 400 0 0 0 VSS
flabel metal1 -164 771 -164 771 1 FreeSans 400 0 0 0 VSS
flabel metal1 -134 250 -134 250 1 FreeSans 400 0 0 0 VSS
flabel metal1 -165 1442 -165 1442 1 FreeSans 400 0 0 0 ip
flabel metal1 1563 1373 1563 1373 1 FreeSans 400 0 0 0 in
flabel metal1 -160 353 -160 353 1 FreeSans 400 0 0 0 clk
flabel metal1 156 4865 156 4865 5 FreeSans 400 0 0 0 VSS
flabel metal1 1243 4868 1243 4868 5 FreeSans 400 0 0 0 VSS
flabel metal1 700 4864 700 4864 1 FreeSans 800 0 0 0 VDD
<< end >>
