magic
tech sky130A
timestamp 1653475914
<< pwell >>
rect -323 -131 324 100
<< nmos >>
rect -223 -26 -208 26
rect -175 -26 -160 26
rect -127 -26 -112 26
rect -79 -26 -64 26
rect -31 -26 -16 26
rect 17 -26 32 26
rect 65 -26 80 26
rect 113 -26 128 26
rect 161 -26 176 26
rect 209 -26 224 26
<< ndiff >>
rect -254 20 -223 26
rect -254 -20 -248 20
rect -231 -20 -223 20
rect -254 -26 -223 -20
rect -208 20 -175 26
rect -208 -20 -200 20
rect -183 -20 -175 20
rect -208 -26 -175 -20
rect -160 20 -127 26
rect -160 -20 -152 20
rect -135 -20 -127 20
rect -160 -26 -127 -20
rect -112 20 -79 26
rect -112 -20 -104 20
rect -87 -20 -79 20
rect -112 -26 -79 -20
rect -64 20 -31 26
rect -64 -20 -56 20
rect -39 -20 -31 20
rect -64 -26 -31 -20
rect -16 20 17 26
rect -16 -20 -8 20
rect 9 -20 17 20
rect -16 -26 17 -20
rect 32 20 65 26
rect 32 -20 40 20
rect 57 -20 65 20
rect 32 -26 65 -20
rect 80 20 113 26
rect 80 -20 88 20
rect 105 -20 113 20
rect 80 -26 113 -20
rect 128 20 161 26
rect 128 -20 136 20
rect 153 -20 161 20
rect 128 -26 161 -20
rect 176 20 209 26
rect 176 -20 184 20
rect 201 -20 209 20
rect 176 -26 209 -20
rect 224 20 255 26
rect 224 -20 232 20
rect 249 -20 255 20
rect 224 -26 255 -20
<< ndiffc >>
rect -248 -20 -231 20
rect -200 -20 -183 20
rect -152 -20 -135 20
rect -104 -20 -87 20
rect -56 -20 -39 20
rect -8 -20 9 20
rect 40 -20 57 20
rect 88 -20 105 20
rect 136 -20 153 20
rect 184 -20 201 20
rect 232 -20 249 20
<< psubdiff >>
rect -305 65 -257 82
rect 258 65 306 82
rect -305 34 -288 65
rect 289 34 306 65
rect -305 -96 -288 -65
rect 289 -96 306 -65
rect -305 -113 -257 -96
rect 258 -113 306 -96
<< psubdiffcont >>
rect -257 65 258 82
rect -305 -65 -288 34
rect 289 -65 306 34
rect -257 -113 258 -96
<< poly >>
rect -223 26 -208 39
rect -175 26 -160 39
rect -127 26 -112 39
rect -79 26 -64 39
rect -31 26 -16 39
rect 17 26 32 39
rect 65 26 80 39
rect 113 26 128 39
rect 161 26 176 39
rect 209 26 224 39
rect -223 -37 -208 -26
rect -175 -37 -160 -26
rect -127 -37 -112 -26
rect -79 -37 -64 -26
rect -31 -37 -16 -26
rect 17 -37 32 -26
rect 65 -37 80 -26
rect 113 -37 128 -26
rect 161 -37 176 -26
rect 209 -37 224 -26
rect -256 -47 257 -37
rect -256 -64 -248 -47
rect -231 -64 -152 -47
rect -135 -64 -56 -47
rect -39 -64 40 -47
rect 57 -64 136 -47
rect 153 -64 232 -47
rect 249 -64 257 -47
rect -256 -70 257 -64
<< polycont >>
rect -248 -64 -231 -47
rect -152 -64 -135 -47
rect -56 -64 -39 -47
rect 40 -64 57 -47
rect 136 -64 153 -47
rect 232 -64 249 -47
<< locali >>
rect -305 65 -257 82
rect 258 65 306 82
rect -305 34 -288 65
rect 289 34 306 65
rect -248 20 -231 28
rect -248 -28 -231 -20
rect -200 20 -183 28
rect -200 -28 -183 -20
rect -152 20 -135 28
rect -152 -28 -135 -20
rect -104 20 -87 28
rect -104 -28 -87 -20
rect -56 20 -39 28
rect -56 -28 -39 -20
rect -8 20 9 28
rect -8 -28 9 -20
rect 40 20 57 28
rect 40 -28 57 -20
rect 88 20 105 28
rect 88 -28 105 -20
rect 136 20 153 28
rect 136 -28 153 -20
rect 184 20 201 28
rect 184 -28 201 -20
rect 232 20 249 28
rect 232 -28 249 -20
rect -256 -64 -248 -47
rect -231 -64 -223 -47
rect -160 -64 -152 -47
rect -135 -64 -127 -47
rect -64 -64 -56 -47
rect -39 -64 -31 -47
rect 32 -64 40 -47
rect 57 -64 65 -47
rect 128 -64 136 -47
rect 153 -64 161 -47
rect 224 -64 232 -47
rect 249 -64 257 -47
rect -305 -96 -288 -65
rect 289 -96 306 -65
rect -305 -113 -257 -96
rect 258 -113 306 -96
<< viali >>
rect -248 -20 -231 20
rect -200 -20 -183 20
rect -152 -20 -135 20
rect -104 -20 -87 20
rect -56 -20 -39 20
rect -8 -20 9 20
rect 40 -20 57 20
rect 88 -20 105 20
rect 136 -20 153 20
rect 184 -20 201 20
rect 232 -20 249 20
rect -248 -64 -231 -47
rect -152 -64 -135 -47
rect -56 -64 -39 -47
rect 40 -64 57 -47
rect 136 -64 153 -47
rect 232 -64 249 -47
<< metal1 >>
rect -251 20 -228 26
rect -251 -20 -248 20
rect -231 -20 -228 20
rect -251 -26 -228 -20
rect -203 20 -180 26
rect -203 -20 -200 20
rect -183 -20 -180 20
rect -203 -26 -180 -20
rect -155 20 -132 26
rect -155 -20 -152 20
rect -135 -20 -132 20
rect -155 -26 -132 -20
rect -107 20 -84 26
rect -107 -20 -104 20
rect -87 -20 -84 20
rect -107 -26 -84 -20
rect -59 20 -36 26
rect -59 -20 -56 20
rect -39 -20 -36 20
rect -59 -26 -36 -20
rect -11 20 12 26
rect -11 -20 -8 20
rect 9 -20 12 20
rect -11 -26 12 -20
rect 37 20 60 26
rect 37 -20 40 20
rect 57 -20 60 20
rect 37 -26 60 -20
rect 85 20 108 26
rect 85 -20 88 20
rect 105 -20 108 20
rect 85 -26 108 -20
rect 133 20 156 26
rect 133 -20 136 20
rect 153 -20 156 20
rect 133 -26 156 -20
rect 181 20 204 26
rect 181 -20 184 20
rect 201 -20 204 20
rect 181 -26 204 -20
rect 229 20 252 26
rect 229 -20 232 20
rect 249 -20 252 20
rect 229 -26 252 -20
rect -256 -47 -223 -40
rect -256 -64 -248 -47
rect -231 -64 -223 -47
rect -256 -70 -223 -64
rect -160 -47 -127 -40
rect -160 -64 -152 -47
rect -135 -64 -127 -47
rect -160 -70 -127 -64
rect -64 -47 -31 -40
rect -64 -64 -56 -47
rect -39 -64 -31 -47
rect -64 -70 -31 -64
rect 32 -47 65 -40
rect 32 -64 40 -47
rect 57 -64 65 -47
rect 32 -70 65 -64
rect 128 -47 161 -40
rect 128 -64 136 -47
rect 153 -64 161 -47
rect 128 -70 161 -64
rect 224 -47 257 -40
rect 224 -64 232 -47
rect 249 -64 257 -47
rect 224 -70 257 -64
<< properties >>
string FIXED_BBOX -297 -105 297 105
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.53 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
