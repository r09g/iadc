magic
tech sky130A
magscale 1 2
timestamp 1653437290
<< nwell >>
rect 417 3013 983 4771
rect 245 3012 1155 3013
rect -51 2692 1501 3012
rect -52 2454 1501 2692
rect -51 2117 1501 2454
<< pwell >>
rect 177 4704 339 4732
rect 139 4670 339 4704
rect 177 4366 339 4670
rect 204 4362 339 4366
rect 194 4276 351 4362
rect 204 4272 339 4276
rect 177 4243 359 4272
rect 139 4209 359 4243
rect 177 3498 359 4209
rect 204 3444 339 3498
rect 177 3175 359 3444
rect 177 3140 339 3175
rect 139 3106 339 3140
rect 177 3078 339 3106
rect 204 3077 339 3078
rect 1061 4428 1223 4732
rect 1061 4394 1261 4428
rect 1061 4366 1223 4394
rect 1061 4362 1196 4366
rect 1049 4276 1206 4362
rect 1061 4272 1196 4276
rect 1041 4243 1223 4272
rect 1041 4209 1261 4243
rect 1041 3498 1223 4209
rect 1061 3444 1196 3498
rect 1041 3175 1223 3444
rect 1061 3140 1223 3175
rect 1061 3106 1261 3140
rect 1061 3078 1223 3106
rect 1061 3077 1196 3078
rect -40 1884 1440 2117
rect -128 1883 1440 1884
rect -128 1831 1585 1883
rect -40 1827 1585 1831
rect -40 1597 1440 1827
rect 245 720 1155 1597
rect 52 199 1346 720
rect 52 198 1345 199
<< nmos >>
rect 160 1807 190 1907
rect 370 1807 400 1907
rect 580 1807 610 1907
rect 790 1807 820 1907
rect 1000 1807 1030 1907
rect 1210 1807 1240 1907
rect 445 1219 475 1319
rect 541 1219 571 1319
rect 637 1219 667 1319
rect 733 1219 763 1319
rect 829 1219 859 1319
rect 925 1219 955 1319
rect 445 997 475 1097
rect 541 997 571 1097
rect 637 997 667 1097
rect 733 997 763 1097
rect 829 997 859 1097
rect 925 997 955 1097
rect 252 408 282 510
rect 348 408 378 510
rect 444 408 474 510
rect 540 408 570 510
rect 636 408 666 510
rect 732 408 762 510
rect 828 408 858 510
rect 924 408 954 510
rect 1020 408 1050 510
rect 1116 408 1146 510
<< scnmos >>
rect 203 4444 313 4654
rect 1087 4444 1197 4654
rect 203 4164 333 4194
rect 1067 4164 1197 4194
rect 203 4080 333 4110
rect 1067 4080 1197 4110
rect 203 3996 333 4026
rect 1067 3996 1197 4026
rect 203 3912 333 3942
rect 1067 3912 1197 3942
rect 203 3828 333 3858
rect 1067 3828 1197 3858
rect 203 3744 333 3774
rect 1067 3744 1197 3774
rect 203 3660 333 3690
rect 1067 3660 1197 3690
rect 203 3576 333 3606
rect 1067 3576 1197 3606
rect 203 3335 333 3365
rect 1067 3335 1197 3365
rect 203 3251 333 3281
rect 1067 3251 1197 3281
rect 203 3156 287 3186
rect 1113 3156 1197 3186
<< pmos >>
rect 42 2554 72 2654
rect 129 2554 159 2654
rect 445 2626 475 2726
rect 541 2626 571 2726
rect 637 2626 667 2726
rect 733 2626 763 2726
rect 829 2626 859 2726
rect 925 2626 955 2726
rect 445 2404 475 2504
rect 541 2404 571 2504
rect 637 2404 667 2504
rect 733 2404 763 2504
rect 829 2404 859 2504
rect 925 2404 955 2504
rect 1290 2279 1320 2379
rect 1377 2279 1407 2379
<< scpmoshvt >>
rect 479 4444 653 4654
rect 747 4444 921 4654
rect 453 4164 653 4194
rect 747 4164 947 4194
rect 453 4080 653 4110
rect 747 4080 947 4110
rect 453 3996 653 4026
rect 747 3996 947 4026
rect 453 3912 653 3942
rect 747 3912 947 3942
rect 453 3828 653 3858
rect 747 3828 947 3858
rect 453 3744 653 3774
rect 747 3744 947 3774
rect 453 3660 653 3690
rect 747 3660 947 3690
rect 453 3576 653 3606
rect 747 3576 947 3606
rect 453 3335 653 3365
rect 747 3335 947 3365
rect 453 3251 653 3281
rect 747 3251 947 3281
rect 517 3156 645 3186
rect 755 3156 883 3186
<< ndiff >>
rect 203 4698 313 4706
rect 203 4664 241 4698
rect 275 4664 313 4698
rect 203 4654 313 4664
rect 1087 4698 1197 4706
rect 1087 4664 1125 4698
rect 1159 4664 1197 4698
rect 1087 4654 1197 4664
rect 203 4434 313 4444
rect 203 4400 241 4434
rect 275 4400 313 4434
rect 203 4392 313 4400
rect 1087 4434 1197 4444
rect 1087 4400 1125 4434
rect 1159 4400 1197 4434
rect 1087 4392 1197 4400
rect 203 4238 333 4246
rect 203 4204 215 4238
rect 249 4204 283 4238
rect 317 4204 333 4238
rect 203 4194 333 4204
rect 1067 4238 1197 4246
rect 1067 4204 1083 4238
rect 1117 4204 1151 4238
rect 1185 4204 1197 4238
rect 1067 4194 1197 4204
rect 203 4154 333 4164
rect 203 4120 215 4154
rect 249 4120 333 4154
rect 203 4110 333 4120
rect 1067 4154 1197 4164
rect 1067 4120 1151 4154
rect 1185 4120 1197 4154
rect 1067 4110 1197 4120
rect 203 4070 333 4080
rect 203 4036 215 4070
rect 249 4036 283 4070
rect 317 4036 333 4070
rect 203 4026 333 4036
rect 1067 4070 1197 4080
rect 1067 4036 1083 4070
rect 1117 4036 1151 4070
rect 1185 4036 1197 4070
rect 1067 4026 1197 4036
rect 203 3986 333 3996
rect 203 3952 215 3986
rect 249 3952 333 3986
rect 203 3942 333 3952
rect 1067 3986 1197 3996
rect 1067 3952 1151 3986
rect 1185 3952 1197 3986
rect 1067 3942 1197 3952
rect 203 3902 333 3912
rect 203 3868 215 3902
rect 249 3868 283 3902
rect 317 3868 333 3902
rect 203 3858 333 3868
rect 1067 3902 1197 3912
rect 1067 3868 1083 3902
rect 1117 3868 1151 3902
rect 1185 3868 1197 3902
rect 1067 3858 1197 3868
rect 203 3818 333 3828
rect 203 3784 283 3818
rect 317 3784 333 3818
rect 203 3774 333 3784
rect 1067 3818 1197 3828
rect 1067 3784 1083 3818
rect 1117 3784 1197 3818
rect 1067 3774 1197 3784
rect 203 3734 333 3744
rect 203 3700 215 3734
rect 249 3700 333 3734
rect 203 3690 333 3700
rect 1067 3734 1197 3744
rect 1067 3700 1151 3734
rect 1185 3700 1197 3734
rect 1067 3690 1197 3700
rect 203 3650 333 3660
rect 203 3616 283 3650
rect 317 3616 333 3650
rect 203 3606 333 3616
rect 1067 3650 1197 3660
rect 1067 3616 1083 3650
rect 1117 3616 1197 3650
rect 1067 3606 1197 3616
rect 203 3566 333 3576
rect 203 3532 215 3566
rect 249 3532 283 3566
rect 317 3532 333 3566
rect 203 3524 333 3532
rect 1067 3566 1197 3576
rect 1067 3532 1083 3566
rect 1117 3532 1151 3566
rect 1185 3532 1197 3566
rect 1067 3524 1197 3532
rect 203 3409 333 3418
rect 203 3375 219 3409
rect 253 3375 287 3409
rect 321 3375 333 3409
rect 203 3365 333 3375
rect 1067 3409 1197 3418
rect 1067 3375 1079 3409
rect 1113 3375 1147 3409
rect 1181 3375 1197 3409
rect 1067 3365 1197 3375
rect 203 3325 333 3335
rect 203 3291 245 3325
rect 279 3291 333 3325
rect 203 3281 333 3291
rect 1067 3325 1197 3335
rect 1067 3291 1121 3325
rect 1155 3291 1197 3325
rect 1067 3281 1197 3291
rect 203 3239 333 3251
rect 203 3205 215 3239
rect 249 3205 333 3239
rect 203 3201 333 3205
rect 1067 3239 1197 3251
rect 1067 3205 1151 3239
rect 1185 3205 1197 3239
rect 1067 3201 1197 3205
rect 203 3186 287 3201
rect 1113 3186 1197 3201
rect 203 3146 287 3156
rect 203 3112 228 3146
rect 262 3112 287 3146
rect 203 3104 287 3112
rect 1113 3146 1197 3156
rect 1113 3112 1138 3146
rect 1172 3112 1197 3146
rect 1113 3104 1197 3112
rect 98 1895 160 1907
rect 98 1819 110 1895
rect 144 1819 160 1895
rect 98 1807 160 1819
rect 190 1895 252 1907
rect 190 1819 206 1895
rect 240 1819 252 1895
rect 190 1807 252 1819
rect 308 1895 370 1907
rect 308 1819 320 1895
rect 354 1819 370 1895
rect 308 1807 370 1819
rect 400 1895 462 1907
rect 400 1819 416 1895
rect 450 1819 462 1895
rect 400 1807 462 1819
rect 518 1895 580 1907
rect 518 1819 530 1895
rect 564 1819 580 1895
rect 518 1807 580 1819
rect 610 1895 672 1907
rect 610 1819 626 1895
rect 660 1819 672 1895
rect 610 1807 672 1819
rect 728 1895 790 1907
rect 728 1819 740 1895
rect 774 1819 790 1895
rect 728 1807 790 1819
rect 820 1895 882 1907
rect 820 1819 836 1895
rect 870 1819 882 1895
rect 820 1807 882 1819
rect 938 1895 1000 1907
rect 938 1819 950 1895
rect 984 1819 1000 1895
rect 938 1807 1000 1819
rect 1030 1895 1092 1907
rect 1030 1819 1046 1895
rect 1080 1819 1092 1895
rect 1030 1807 1092 1819
rect 1148 1895 1210 1907
rect 1148 1819 1160 1895
rect 1194 1819 1210 1895
rect 1148 1807 1210 1819
rect 1240 1895 1302 1907
rect 1240 1819 1256 1895
rect 1290 1819 1302 1895
rect 1240 1807 1302 1819
rect 383 1307 445 1319
rect 383 1231 395 1307
rect 429 1231 445 1307
rect 383 1219 445 1231
rect 475 1307 541 1319
rect 475 1231 491 1307
rect 525 1231 541 1307
rect 475 1219 541 1231
rect 571 1307 637 1319
rect 571 1231 587 1307
rect 621 1231 637 1307
rect 571 1219 637 1231
rect 667 1307 733 1319
rect 667 1231 683 1307
rect 717 1231 733 1307
rect 667 1219 733 1231
rect 763 1307 829 1319
rect 763 1231 779 1307
rect 813 1231 829 1307
rect 763 1219 829 1231
rect 859 1307 925 1319
rect 859 1231 875 1307
rect 909 1231 925 1307
rect 859 1219 925 1231
rect 955 1307 1017 1319
rect 955 1231 971 1307
rect 1005 1231 1017 1307
rect 955 1219 1017 1231
rect 383 1085 445 1097
rect 383 1009 395 1085
rect 429 1009 445 1085
rect 383 997 445 1009
rect 475 1085 541 1097
rect 475 1009 491 1085
rect 525 1009 541 1085
rect 475 997 541 1009
rect 571 1085 637 1097
rect 571 1009 587 1085
rect 621 1009 637 1085
rect 571 997 637 1009
rect 667 1085 733 1097
rect 667 1009 683 1085
rect 717 1009 733 1085
rect 667 997 733 1009
rect 763 1085 829 1097
rect 763 1009 779 1085
rect 813 1009 829 1085
rect 763 997 829 1009
rect 859 1085 925 1097
rect 859 1009 875 1085
rect 909 1009 925 1085
rect 859 997 925 1009
rect 955 1085 1017 1097
rect 955 1009 971 1085
rect 1005 1009 1017 1085
rect 955 997 1017 1009
rect 190 498 252 510
rect 190 420 202 498
rect 236 420 252 498
rect 190 408 252 420
rect 282 498 348 510
rect 282 420 298 498
rect 332 420 348 498
rect 282 408 348 420
rect 378 498 444 510
rect 378 420 394 498
rect 428 420 444 498
rect 378 408 444 420
rect 474 498 540 510
rect 474 420 490 498
rect 524 420 540 498
rect 474 408 540 420
rect 570 498 636 510
rect 570 420 586 498
rect 620 420 636 498
rect 570 408 636 420
rect 666 498 732 510
rect 666 420 682 498
rect 716 420 732 498
rect 666 408 732 420
rect 762 498 828 510
rect 762 420 778 498
rect 812 420 828 498
rect 762 408 828 420
rect 858 498 924 510
rect 858 420 874 498
rect 908 420 924 498
rect 858 408 924 420
rect 954 498 1020 510
rect 954 420 970 498
rect 1004 420 1020 498
rect 954 408 1020 420
rect 1050 498 1116 510
rect 1050 420 1066 498
rect 1100 420 1116 498
rect 1050 408 1116 420
rect 1146 498 1208 510
rect 1146 420 1162 498
rect 1196 420 1208 498
rect 1146 408 1208 420
<< pdiff >>
rect 479 4698 653 4706
rect 479 4664 505 4698
rect 539 4664 607 4698
rect 641 4664 653 4698
rect 479 4654 653 4664
rect 747 4698 921 4706
rect 747 4664 759 4698
rect 793 4664 861 4698
rect 895 4664 921 4698
rect 747 4654 921 4664
rect 479 4434 653 4444
rect 479 4400 505 4434
rect 539 4400 607 4434
rect 641 4400 653 4434
rect 479 4392 653 4400
rect 747 4434 921 4444
rect 747 4400 759 4434
rect 793 4400 861 4434
rect 895 4400 921 4434
rect 747 4392 921 4400
rect 453 4238 653 4246
rect 453 4204 471 4238
rect 505 4204 539 4238
rect 573 4204 607 4238
rect 641 4204 653 4238
rect 453 4194 653 4204
rect 747 4238 947 4246
rect 747 4204 759 4238
rect 793 4204 827 4238
rect 861 4204 895 4238
rect 929 4204 947 4238
rect 747 4194 947 4204
rect 453 4154 653 4164
rect 453 4120 471 4154
rect 505 4120 539 4154
rect 573 4120 607 4154
rect 641 4120 653 4154
rect 453 4110 653 4120
rect 747 4154 947 4164
rect 747 4120 759 4154
rect 793 4120 827 4154
rect 861 4120 895 4154
rect 929 4120 947 4154
rect 747 4110 947 4120
rect 453 4070 653 4080
rect 453 4036 539 4070
rect 573 4036 607 4070
rect 641 4036 653 4070
rect 453 4026 653 4036
rect 747 4070 947 4080
rect 747 4036 759 4070
rect 793 4036 827 4070
rect 861 4036 947 4070
rect 747 4026 947 4036
rect 453 3986 653 3996
rect 453 3952 471 3986
rect 505 3952 539 3986
rect 573 3952 607 3986
rect 641 3952 653 3986
rect 453 3942 653 3952
rect 747 3986 947 3996
rect 747 3952 759 3986
rect 793 3952 827 3986
rect 861 3952 895 3986
rect 929 3952 947 3986
rect 747 3942 947 3952
rect 453 3902 653 3912
rect 453 3868 539 3902
rect 573 3868 607 3902
rect 641 3868 653 3902
rect 453 3858 653 3868
rect 747 3902 947 3912
rect 747 3868 759 3902
rect 793 3868 827 3902
rect 861 3868 947 3902
rect 747 3858 947 3868
rect 453 3818 653 3828
rect 453 3784 471 3818
rect 505 3784 539 3818
rect 573 3784 607 3818
rect 641 3784 653 3818
rect 453 3774 653 3784
rect 747 3818 947 3828
rect 747 3784 759 3818
rect 793 3784 827 3818
rect 861 3784 895 3818
rect 929 3784 947 3818
rect 747 3774 947 3784
rect 453 3734 653 3744
rect 453 3700 539 3734
rect 573 3700 607 3734
rect 641 3700 653 3734
rect 453 3690 653 3700
rect 747 3734 947 3744
rect 747 3700 759 3734
rect 793 3700 827 3734
rect 861 3700 947 3734
rect 747 3690 947 3700
rect 453 3650 653 3660
rect 453 3616 471 3650
rect 505 3616 539 3650
rect 573 3616 607 3650
rect 641 3616 653 3650
rect 453 3606 653 3616
rect 747 3650 947 3660
rect 747 3616 759 3650
rect 793 3616 827 3650
rect 861 3616 895 3650
rect 929 3616 947 3650
rect 747 3606 947 3616
rect 453 3566 653 3576
rect 453 3532 539 3566
rect 573 3532 607 3566
rect 641 3532 653 3566
rect 453 3524 653 3532
rect 747 3566 947 3576
rect 747 3532 759 3566
rect 793 3532 827 3566
rect 861 3532 947 3566
rect 747 3524 947 3532
rect 453 3409 653 3418
rect 453 3375 471 3409
rect 505 3375 539 3409
rect 573 3375 607 3409
rect 641 3375 653 3409
rect 453 3365 653 3375
rect 747 3409 947 3418
rect 747 3375 759 3409
rect 793 3375 827 3409
rect 861 3375 895 3409
rect 929 3375 947 3409
rect 747 3365 947 3375
rect 453 3325 653 3335
rect 453 3291 502 3325
rect 536 3291 583 3325
rect 617 3291 653 3325
rect 453 3281 653 3291
rect 747 3325 947 3335
rect 747 3291 783 3325
rect 817 3291 864 3325
rect 898 3291 947 3325
rect 747 3281 947 3291
rect 453 3239 653 3251
rect 453 3205 531 3239
rect 565 3205 599 3239
rect 633 3205 653 3239
rect 453 3201 653 3205
rect 747 3239 947 3251
rect 747 3205 767 3239
rect 801 3205 835 3239
rect 869 3205 947 3239
rect 747 3201 947 3205
rect 517 3186 645 3201
rect 755 3186 883 3201
rect 517 3146 645 3156
rect 517 3112 531 3146
rect 565 3112 599 3146
rect 633 3112 645 3146
rect 517 3104 645 3112
rect 755 3146 883 3156
rect 755 3112 767 3146
rect 801 3112 835 3146
rect 869 3112 883 3146
rect 755 3104 883 3112
rect -16 2642 42 2654
rect -16 2566 -4 2642
rect 30 2566 42 2642
rect -16 2554 42 2566
rect 72 2642 129 2654
rect 72 2566 84 2642
rect 118 2566 129 2642
rect 72 2554 129 2566
rect 159 2642 216 2654
rect 159 2566 170 2642
rect 204 2566 216 2642
rect 159 2554 216 2566
rect 383 2714 445 2726
rect 383 2638 395 2714
rect 429 2638 445 2714
rect 383 2626 445 2638
rect 475 2714 541 2726
rect 475 2638 491 2714
rect 525 2638 541 2714
rect 475 2626 541 2638
rect 571 2714 637 2726
rect 571 2638 587 2714
rect 621 2638 637 2714
rect 571 2626 637 2638
rect 667 2714 733 2726
rect 667 2638 683 2714
rect 717 2638 733 2714
rect 667 2626 733 2638
rect 763 2714 829 2726
rect 763 2638 779 2714
rect 813 2638 829 2714
rect 763 2626 829 2638
rect 859 2714 925 2726
rect 859 2638 875 2714
rect 909 2638 925 2714
rect 859 2626 925 2638
rect 955 2714 1017 2726
rect 955 2638 971 2714
rect 1005 2638 1017 2714
rect 955 2626 1017 2638
rect 383 2492 445 2504
rect 383 2416 395 2492
rect 429 2416 445 2492
rect 383 2404 445 2416
rect 475 2492 541 2504
rect 475 2416 491 2492
rect 525 2416 541 2492
rect 475 2404 541 2416
rect 571 2492 637 2504
rect 571 2416 587 2492
rect 621 2416 637 2492
rect 571 2404 637 2416
rect 667 2492 733 2504
rect 667 2416 683 2492
rect 717 2416 733 2492
rect 667 2404 733 2416
rect 763 2492 829 2504
rect 763 2416 779 2492
rect 813 2416 829 2492
rect 763 2404 829 2416
rect 859 2492 925 2504
rect 859 2416 875 2492
rect 909 2416 925 2492
rect 859 2404 925 2416
rect 955 2492 1017 2504
rect 955 2416 971 2492
rect 1005 2416 1017 2492
rect 955 2404 1017 2416
rect 1232 2367 1290 2379
rect 1232 2291 1244 2367
rect 1278 2291 1290 2367
rect 1232 2279 1290 2291
rect 1320 2367 1377 2379
rect 1320 2291 1332 2367
rect 1366 2291 1377 2367
rect 1320 2279 1377 2291
rect 1407 2367 1464 2379
rect 1407 2291 1418 2367
rect 1452 2291 1464 2367
rect 1407 2279 1464 2291
<< ndiffc >>
rect 241 4664 275 4698
rect 1125 4664 1159 4698
rect 241 4400 275 4434
rect 1125 4400 1159 4434
rect 215 4204 249 4238
rect 283 4204 317 4238
rect 1083 4204 1117 4238
rect 1151 4204 1185 4238
rect 215 4120 249 4154
rect 1151 4120 1185 4154
rect 215 4036 249 4070
rect 283 4036 317 4070
rect 1083 4036 1117 4070
rect 1151 4036 1185 4070
rect 215 3952 249 3986
rect 1151 3952 1185 3986
rect 215 3868 249 3902
rect 283 3868 317 3902
rect 1083 3868 1117 3902
rect 1151 3868 1185 3902
rect 283 3784 317 3818
rect 1083 3784 1117 3818
rect 215 3700 249 3734
rect 1151 3700 1185 3734
rect 283 3616 317 3650
rect 1083 3616 1117 3650
rect 215 3532 249 3566
rect 283 3532 317 3566
rect 1083 3532 1117 3566
rect 1151 3532 1185 3566
rect 219 3375 253 3409
rect 287 3375 321 3409
rect 1079 3375 1113 3409
rect 1147 3375 1181 3409
rect 245 3291 279 3325
rect 1121 3291 1155 3325
rect 215 3205 249 3239
rect 1151 3205 1185 3239
rect 228 3112 262 3146
rect 1138 3112 1172 3146
rect 110 1819 144 1895
rect 206 1819 240 1895
rect 320 1819 354 1895
rect 416 1819 450 1895
rect 530 1819 564 1895
rect 626 1819 660 1895
rect 740 1819 774 1895
rect 836 1819 870 1895
rect 950 1819 984 1895
rect 1046 1819 1080 1895
rect 1160 1819 1194 1895
rect 1256 1819 1290 1895
rect 395 1231 429 1307
rect 491 1231 525 1307
rect 587 1231 621 1307
rect 683 1231 717 1307
rect 779 1231 813 1307
rect 875 1231 909 1307
rect 971 1231 1005 1307
rect 395 1009 429 1085
rect 491 1009 525 1085
rect 587 1009 621 1085
rect 683 1009 717 1085
rect 779 1009 813 1085
rect 875 1009 909 1085
rect 971 1009 1005 1085
rect 202 420 236 498
rect 298 420 332 498
rect 394 420 428 498
rect 490 420 524 498
rect 586 420 620 498
rect 682 420 716 498
rect 778 420 812 498
rect 874 420 908 498
rect 970 420 1004 498
rect 1066 420 1100 498
rect 1162 420 1196 498
<< pdiffc >>
rect 505 4664 539 4698
rect 607 4664 641 4698
rect 759 4664 793 4698
rect 861 4664 895 4698
rect 505 4400 539 4434
rect 607 4400 641 4434
rect 759 4400 793 4434
rect 861 4400 895 4434
rect 471 4204 505 4238
rect 539 4204 573 4238
rect 607 4204 641 4238
rect 759 4204 793 4238
rect 827 4204 861 4238
rect 895 4204 929 4238
rect 471 4120 505 4154
rect 539 4120 573 4154
rect 607 4120 641 4154
rect 759 4120 793 4154
rect 827 4120 861 4154
rect 895 4120 929 4154
rect 539 4036 573 4070
rect 607 4036 641 4070
rect 759 4036 793 4070
rect 827 4036 861 4070
rect 471 3952 505 3986
rect 539 3952 573 3986
rect 607 3952 641 3986
rect 759 3952 793 3986
rect 827 3952 861 3986
rect 895 3952 929 3986
rect 539 3868 573 3902
rect 607 3868 641 3902
rect 759 3868 793 3902
rect 827 3868 861 3902
rect 471 3784 505 3818
rect 539 3784 573 3818
rect 607 3784 641 3818
rect 759 3784 793 3818
rect 827 3784 861 3818
rect 895 3784 929 3818
rect 539 3700 573 3734
rect 607 3700 641 3734
rect 759 3700 793 3734
rect 827 3700 861 3734
rect 471 3616 505 3650
rect 539 3616 573 3650
rect 607 3616 641 3650
rect 759 3616 793 3650
rect 827 3616 861 3650
rect 895 3616 929 3650
rect 539 3532 573 3566
rect 607 3532 641 3566
rect 759 3532 793 3566
rect 827 3532 861 3566
rect 471 3375 505 3409
rect 539 3375 573 3409
rect 607 3375 641 3409
rect 759 3375 793 3409
rect 827 3375 861 3409
rect 895 3375 929 3409
rect 502 3291 536 3325
rect 583 3291 617 3325
rect 783 3291 817 3325
rect 864 3291 898 3325
rect 531 3205 565 3239
rect 599 3205 633 3239
rect 767 3205 801 3239
rect 835 3205 869 3239
rect 531 3112 565 3146
rect 599 3112 633 3146
rect 767 3112 801 3146
rect 835 3112 869 3146
rect -4 2566 30 2642
rect 84 2566 118 2642
rect 170 2566 204 2642
rect 395 2638 429 2714
rect 491 2638 525 2714
rect 587 2638 621 2714
rect 683 2638 717 2714
rect 779 2638 813 2714
rect 875 2638 909 2714
rect 971 2638 1005 2714
rect 395 2416 429 2492
rect 491 2416 525 2492
rect 587 2416 621 2492
rect 683 2416 717 2492
rect 779 2416 813 2492
rect 875 2416 909 2492
rect 971 2416 1005 2492
rect 1244 2291 1278 2367
rect 1332 2291 1366 2367
rect 1418 2291 1452 2367
<< psubdiff >>
rect 220 4302 267 4336
rect 301 4302 325 4336
rect 1075 4302 1099 4336
rect 1133 4302 1180 4336
rect -4 2047 92 2081
rect 1308 2047 1404 2081
rect -4 1985 30 2047
rect 1370 1985 1404 2047
rect -4 1667 30 1729
rect 1370 1667 1404 1729
rect -4 1633 92 1667
rect 1308 1633 1404 1667
rect 281 1527 377 1561
rect 1023 1527 1119 1561
rect 281 1465 315 1527
rect 1085 1465 1119 1527
rect 281 789 315 851
rect 1085 789 1119 851
rect 281 755 377 789
rect 1023 755 1119 789
rect 88 650 184 684
rect 1214 650 1310 684
rect 88 588 122 650
rect 1276 588 1310 650
rect 88 268 122 330
rect 1276 268 1310 330
rect 88 234 184 268
rect 1214 234 1310 268
<< nsubdiff >>
rect 461 4302 485 4336
rect 519 4302 578 4336
rect 612 4302 636 4336
rect 764 4302 788 4336
rect 822 4302 881 4336
rect 915 4302 939 4336
rect 281 2943 377 2977
rect 1023 2943 1119 2977
rect 281 2881 315 2943
rect 1085 2881 1119 2943
rect 281 2187 315 2249
rect 1085 2187 1119 2249
rect 281 2153 377 2187
rect 1023 2153 1119 2187
<< psubdiffcont >>
rect 267 4302 301 4336
rect 1099 4302 1133 4336
rect 92 2047 1308 2081
rect -4 1729 30 1985
rect 1370 1729 1404 1985
rect 92 1633 1308 1667
rect 377 1527 1023 1561
rect 281 851 315 1465
rect 1085 851 1119 1465
rect 377 755 1023 789
rect 184 650 1214 684
rect 88 330 122 588
rect 1276 330 1310 588
rect 184 234 1214 268
<< nsubdiffcont >>
rect 485 4302 519 4336
rect 578 4302 612 4336
rect 788 4302 822 4336
rect 881 4302 915 4336
rect 377 2943 1023 2977
rect 281 2249 315 2881
rect 1085 2249 1119 2881
rect 377 2153 1023 2187
<< poly >>
rect 381 4696 447 4712
rect 381 4662 397 4696
rect 431 4662 447 4696
rect 381 4654 447 4662
rect 989 4696 1055 4712
rect 989 4662 1005 4696
rect 1039 4662 1055 4696
rect 989 4654 1055 4662
rect 177 4444 203 4654
rect 313 4528 339 4654
rect 381 4570 479 4654
rect 313 4444 411 4528
rect 453 4444 479 4570
rect 653 4444 679 4654
rect 721 4444 747 4654
rect 921 4528 947 4654
rect 989 4570 1087 4654
rect 921 4444 1019 4528
rect 1061 4444 1087 4570
rect 1197 4444 1223 4654
rect 345 4436 411 4444
rect 345 4402 361 4436
rect 395 4402 411 4436
rect 345 4386 411 4402
rect 953 4436 1019 4444
rect 953 4402 969 4436
rect 1003 4402 1019 4436
rect 953 4386 1019 4402
rect 355 4235 421 4251
rect 355 4201 371 4235
rect 405 4201 421 4235
rect 355 4194 421 4201
rect 979 4235 1045 4251
rect 979 4201 995 4235
rect 1029 4201 1045 4235
rect 979 4194 1045 4201
rect 177 4164 203 4194
rect 333 4164 453 4194
rect 653 4164 679 4194
rect 721 4164 747 4194
rect 947 4164 1067 4194
rect 1197 4164 1223 4194
rect 355 4154 421 4164
rect 355 4120 371 4154
rect 405 4120 421 4154
rect 355 4110 421 4120
rect 979 4154 1045 4164
rect 979 4120 995 4154
rect 1029 4120 1045 4154
rect 979 4110 1045 4120
rect 177 4080 203 4110
rect 333 4080 453 4110
rect 653 4080 679 4110
rect 721 4080 747 4110
rect 947 4080 1067 4110
rect 1197 4080 1223 4110
rect 355 4070 421 4080
rect 355 4036 371 4070
rect 405 4036 421 4070
rect 355 4026 421 4036
rect 979 4070 1045 4080
rect 979 4036 995 4070
rect 1029 4036 1045 4070
rect 979 4026 1045 4036
rect 177 3996 203 4026
rect 333 3996 453 4026
rect 653 3996 679 4026
rect 721 3996 747 4026
rect 947 3996 1067 4026
rect 1197 3996 1223 4026
rect 355 3986 421 3996
rect 355 3952 371 3986
rect 405 3952 421 3986
rect 355 3942 421 3952
rect 979 3986 1045 3996
rect 979 3952 995 3986
rect 1029 3952 1045 3986
rect 979 3942 1045 3952
rect 177 3912 203 3942
rect 333 3912 453 3942
rect 653 3912 679 3942
rect 721 3912 747 3942
rect 947 3912 1067 3942
rect 1197 3912 1223 3942
rect 177 3828 203 3858
rect 333 3828 453 3858
rect 653 3828 679 3858
rect 721 3828 747 3858
rect 947 3828 1067 3858
rect 1197 3828 1223 3858
rect 355 3774 421 3828
rect 979 3774 1045 3828
rect 177 3744 203 3774
rect 333 3744 453 3774
rect 653 3744 679 3774
rect 721 3744 747 3774
rect 947 3744 1067 3774
rect 1197 3744 1223 3774
rect 355 3734 421 3744
rect 355 3700 371 3734
rect 405 3700 421 3734
rect 355 3690 421 3700
rect 979 3734 1045 3744
rect 979 3700 995 3734
rect 1029 3700 1045 3734
rect 979 3690 1045 3700
rect 177 3660 203 3690
rect 333 3660 453 3690
rect 653 3660 679 3690
rect 721 3660 747 3690
rect 947 3660 1067 3690
rect 1197 3660 1223 3690
rect 355 3650 421 3660
rect 355 3616 371 3650
rect 405 3616 421 3650
rect 355 3606 421 3616
rect 979 3650 1045 3660
rect 979 3616 995 3650
rect 1029 3616 1045 3650
rect 979 3606 1045 3616
rect 177 3576 203 3606
rect 333 3576 453 3606
rect 653 3576 679 3606
rect 721 3576 747 3606
rect 947 3576 1067 3606
rect 1197 3576 1223 3606
rect 177 3335 203 3365
rect 333 3335 453 3365
rect 653 3335 679 3365
rect 721 3335 747 3365
rect 947 3335 1067 3365
rect 1197 3335 1223 3365
rect 355 3281 421 3335
rect 979 3281 1045 3335
rect 177 3251 203 3281
rect 333 3272 453 3281
rect 333 3251 371 3272
rect 355 3238 371 3251
rect 405 3251 453 3272
rect 653 3251 679 3281
rect 721 3251 747 3281
rect 947 3272 1067 3281
rect 947 3251 995 3272
rect 405 3238 421 3251
rect 355 3228 421 3238
rect 979 3238 995 3251
rect 1029 3251 1067 3272
rect 1197 3251 1223 3281
rect 1029 3238 1045 3251
rect 979 3228 1045 3238
rect 177 3156 203 3186
rect 287 3156 517 3186
rect 645 3156 671 3186
rect 729 3156 755 3186
rect 883 3156 1113 3186
rect 1197 3156 1223 3186
rect 355 3148 421 3156
rect 355 3114 371 3148
rect 405 3114 421 3148
rect 355 3104 421 3114
rect 979 3148 1045 3156
rect 979 3114 995 3148
rect 1029 3114 1045 3148
rect 979 3104 1045 3114
rect 42 2654 72 2684
rect 129 2654 159 2684
rect 42 2524 72 2554
rect 129 2524 159 2554
rect 42 2507 159 2524
rect 42 2473 84 2507
rect 118 2473 159 2507
rect 42 2458 159 2473
rect 637 2875 763 2891
rect 637 2841 683 2875
rect 717 2841 763 2875
rect 637 2825 763 2841
rect 409 2807 475 2823
rect 409 2773 425 2807
rect 459 2773 475 2807
rect 409 2757 475 2773
rect 523 2807 589 2823
rect 523 2773 539 2807
rect 573 2773 589 2807
rect 523 2757 589 2773
rect 445 2726 475 2757
rect 541 2726 571 2757
rect 637 2726 667 2825
rect 733 2726 763 2825
rect 811 2807 877 2823
rect 811 2773 827 2807
rect 861 2773 877 2807
rect 811 2757 877 2773
rect 925 2807 991 2823
rect 925 2773 941 2807
rect 975 2773 991 2807
rect 925 2757 991 2773
rect 829 2726 859 2757
rect 925 2726 955 2757
rect 445 2600 475 2626
rect 541 2600 571 2626
rect 637 2600 667 2626
rect 733 2600 763 2626
rect 829 2600 859 2626
rect 925 2600 955 2626
rect 445 2504 475 2530
rect 541 2504 571 2530
rect 637 2504 667 2530
rect 733 2504 763 2530
rect 829 2504 859 2530
rect 925 2504 955 2530
rect 445 2373 475 2404
rect 541 2373 571 2404
rect 409 2357 475 2373
rect 409 2323 425 2357
rect 459 2323 475 2357
rect 409 2307 475 2323
rect 523 2357 589 2373
rect 523 2323 539 2357
rect 573 2323 589 2357
rect 523 2307 589 2323
rect 637 2305 667 2404
rect 733 2305 763 2404
rect 829 2373 859 2404
rect 925 2373 955 2404
rect 811 2357 877 2373
rect 811 2323 827 2357
rect 861 2323 877 2357
rect 811 2307 877 2323
rect 925 2357 991 2373
rect 925 2323 941 2357
rect 975 2323 991 2357
rect 925 2307 991 2323
rect 637 2289 763 2305
rect 637 2255 683 2289
rect 717 2255 763 2289
rect 637 2239 763 2255
rect 1290 2379 1320 2409
rect 1377 2379 1407 2409
rect 1290 2249 1320 2279
rect 1377 2249 1407 2279
rect 1290 2232 1407 2249
rect 1290 2198 1332 2232
rect 1366 2198 1407 2232
rect 1290 2183 1407 2198
rect 142 1979 208 1995
rect 142 1945 158 1979
rect 192 1945 208 1979
rect 142 1929 208 1945
rect 352 1979 418 1995
rect 352 1945 368 1979
rect 402 1945 418 1979
rect 352 1929 418 1945
rect 982 1979 1048 1995
rect 982 1945 998 1979
rect 1032 1945 1048 1979
rect 160 1907 190 1929
rect 370 1907 400 1929
rect 580 1907 610 1933
rect 790 1907 820 1933
rect 982 1929 1048 1945
rect 1192 1979 1258 1995
rect 1192 1945 1208 1979
rect 1242 1945 1258 1979
rect 1192 1929 1258 1945
rect 1000 1907 1030 1929
rect 1210 1907 1240 1929
rect 160 1785 190 1807
rect 142 1769 208 1785
rect 370 1781 400 1807
rect 580 1785 610 1807
rect 790 1785 820 1807
rect 142 1735 158 1769
rect 192 1735 208 1769
rect 142 1719 208 1735
rect 562 1769 628 1785
rect 562 1735 578 1769
rect 612 1735 628 1769
rect 562 1719 628 1735
rect 772 1769 838 1785
rect 1000 1781 1030 1807
rect 1210 1785 1240 1807
rect 772 1735 788 1769
rect 822 1735 838 1769
rect 772 1719 838 1735
rect 1192 1769 1258 1785
rect 1192 1735 1208 1769
rect 1242 1735 1258 1769
rect 1192 1719 1258 1735
rect 637 1459 763 1475
rect 637 1425 683 1459
rect 717 1425 763 1459
rect 637 1409 763 1425
rect 409 1391 475 1407
rect 409 1357 425 1391
rect 459 1357 475 1391
rect 409 1341 475 1357
rect 523 1391 589 1407
rect 523 1357 539 1391
rect 573 1357 589 1391
rect 523 1341 589 1357
rect 445 1319 475 1341
rect 541 1319 571 1341
rect 637 1319 667 1409
rect 733 1319 763 1409
rect 811 1391 877 1407
rect 811 1357 827 1391
rect 861 1357 877 1391
rect 811 1341 877 1357
rect 925 1391 991 1407
rect 925 1357 941 1391
rect 975 1357 991 1391
rect 925 1341 991 1357
rect 829 1319 859 1341
rect 925 1319 955 1341
rect 445 1193 475 1219
rect 541 1193 571 1219
rect 637 1193 667 1219
rect 733 1193 763 1219
rect 829 1193 859 1219
rect 925 1193 955 1219
rect 445 1097 475 1123
rect 541 1097 571 1123
rect 637 1097 667 1123
rect 733 1097 763 1123
rect 829 1097 859 1123
rect 925 1097 955 1123
rect 445 975 475 997
rect 541 975 571 997
rect 409 959 475 975
rect 409 925 425 959
rect 459 925 475 959
rect 409 909 475 925
rect 523 959 589 975
rect 523 925 539 959
rect 573 925 589 959
rect 523 909 589 925
rect 637 907 667 997
rect 733 907 763 997
rect 829 975 859 997
rect 925 975 955 997
rect 811 959 877 975
rect 811 925 827 959
rect 861 925 877 959
rect 811 909 877 925
rect 925 959 991 975
rect 925 925 941 959
rect 975 925 991 959
rect 925 909 991 925
rect 637 891 763 907
rect 637 857 683 891
rect 717 857 763 891
rect 637 841 763 857
rect 216 582 282 598
rect 216 548 232 582
rect 266 548 282 582
rect 216 532 282 548
rect 1116 582 1182 598
rect 1116 548 1132 582
rect 1166 548 1182 582
rect 252 510 282 532
rect 348 510 378 536
rect 444 510 474 536
rect 540 510 570 536
rect 636 510 666 536
rect 732 510 762 536
rect 828 510 858 536
rect 924 510 954 536
rect 1020 510 1050 536
rect 1116 532 1182 548
rect 1116 510 1146 532
rect 252 386 282 408
rect 216 370 282 386
rect 216 336 232 370
rect 266 336 282 370
rect 216 320 282 336
rect 348 386 378 408
rect 444 386 474 408
rect 540 386 570 408
rect 636 386 666 408
rect 732 386 762 408
rect 828 386 858 408
rect 924 386 954 408
rect 1020 386 1050 408
rect 348 370 1050 386
rect 348 336 394 370
rect 428 336 586 370
rect 620 336 778 370
rect 812 336 952 370
rect 986 336 1050 370
rect 348 320 1050 336
rect 1116 386 1146 408
rect 1116 370 1182 386
rect 1116 336 1132 370
rect 1166 336 1182 370
rect 1116 320 1182 336
<< polycont >>
rect 397 4662 431 4696
rect 1005 4662 1039 4696
rect 361 4402 395 4436
rect 969 4402 1003 4436
rect 371 4201 405 4235
rect 995 4201 1029 4235
rect 371 4120 405 4154
rect 995 4120 1029 4154
rect 371 4036 405 4070
rect 995 4036 1029 4070
rect 371 3952 405 3986
rect 995 3952 1029 3986
rect 371 3700 405 3734
rect 995 3700 1029 3734
rect 371 3616 405 3650
rect 995 3616 1029 3650
rect 371 3238 405 3272
rect 995 3238 1029 3272
rect 371 3114 405 3148
rect 995 3114 1029 3148
rect 84 2473 118 2507
rect 683 2841 717 2875
rect 425 2773 459 2807
rect 539 2773 573 2807
rect 827 2773 861 2807
rect 941 2773 975 2807
rect 425 2323 459 2357
rect 539 2323 573 2357
rect 827 2323 861 2357
rect 941 2323 975 2357
rect 683 2255 717 2289
rect 1332 2198 1366 2232
rect 158 1945 192 1979
rect 368 1945 402 1979
rect 998 1945 1032 1979
rect 1208 1945 1242 1979
rect 158 1735 192 1769
rect 578 1735 612 1769
rect 788 1735 822 1769
rect 1208 1735 1242 1769
rect 683 1425 717 1459
rect 425 1357 459 1391
rect 539 1357 573 1391
rect 827 1357 861 1391
rect 941 1357 975 1391
rect 425 925 459 959
rect 539 925 573 959
rect 827 925 861 959
rect 941 925 975 959
rect 683 857 717 891
rect 232 548 266 582
rect 1132 548 1166 582
rect 232 336 266 370
rect 394 336 428 370
rect 586 336 620 370
rect 778 336 812 370
rect 952 336 986 370
rect 1132 336 1166 370
<< locali >>
rect 139 4716 173 4733
rect 683 4716 717 4733
rect 1227 4716 1261 4733
rect 139 4704 431 4716
rect 173 4698 431 4704
rect 173 4670 241 4698
rect 139 4664 241 4670
rect 275 4696 431 4698
rect 275 4664 397 4696
rect 139 4662 397 4664
rect 139 4612 431 4662
rect 173 4578 431 4612
rect 139 4566 431 4578
rect 465 4704 1039 4716
rect 465 4698 683 4704
rect 465 4664 505 4698
rect 539 4664 607 4698
rect 641 4670 683 4698
rect 717 4698 1039 4704
rect 717 4670 759 4698
rect 641 4664 759 4670
rect 793 4664 861 4698
rect 895 4696 1039 4698
rect 895 4664 1005 4696
rect 465 4662 1005 4664
rect 465 4612 1039 4662
rect 465 4578 683 4612
rect 717 4578 1039 4612
rect 465 4566 1039 4578
rect 1073 4704 1261 4716
rect 1073 4698 1227 4704
rect 1073 4664 1125 4698
rect 1159 4670 1227 4698
rect 1159 4664 1261 4670
rect 1073 4612 1261 4664
rect 1073 4578 1227 4612
rect 139 4520 327 4566
rect 465 4532 935 4566
rect 1073 4532 1261 4578
rect 173 4486 327 4520
rect 139 4434 327 4486
rect 139 4428 241 4434
rect 173 4400 241 4428
rect 275 4400 327 4434
rect 173 4394 327 4400
rect 139 4382 327 4394
rect 361 4520 935 4532
rect 361 4486 683 4520
rect 717 4486 935 4520
rect 361 4436 935 4486
rect 395 4434 935 4436
rect 395 4402 505 4434
rect 361 4400 505 4402
rect 539 4400 607 4434
rect 641 4428 759 4434
rect 641 4400 683 4428
rect 361 4394 683 4400
rect 717 4400 759 4428
rect 793 4400 861 4434
rect 895 4400 935 4434
rect 717 4394 935 4400
rect 361 4382 935 4394
rect 969 4520 1261 4532
rect 969 4486 1227 4520
rect 969 4436 1261 4486
rect 1003 4434 1261 4436
rect 1003 4402 1125 4434
rect 969 4400 1125 4402
rect 1159 4428 1261 4434
rect 1159 4400 1227 4428
rect 969 4394 1227 4400
rect 969 4382 1261 4394
rect 139 4348 173 4382
rect 683 4348 717 4382
rect 1227 4348 1261 4382
rect 139 4336 318 4348
rect 173 4302 267 4336
rect 301 4302 318 4336
rect 139 4290 318 4302
rect 450 4336 950 4348
rect 450 4302 485 4336
rect 519 4302 578 4336
rect 612 4302 683 4336
rect 717 4302 788 4336
rect 822 4302 881 4336
rect 915 4302 950 4336
rect 450 4290 950 4302
rect 1082 4336 1261 4348
rect 1082 4302 1099 4336
rect 1133 4302 1227 4336
rect 1082 4290 1261 4302
rect 139 4244 173 4290
rect 683 4255 717 4290
rect 139 4154 173 4210
rect 207 4238 337 4255
rect 207 4204 215 4238
rect 249 4204 283 4238
rect 317 4204 337 4238
rect 207 4188 337 4204
rect 139 4152 215 4154
rect 173 4120 215 4152
rect 249 4120 265 4154
rect 139 4060 173 4118
rect 299 4086 337 4188
rect 139 3986 173 4026
rect 207 4070 337 4086
rect 207 4036 215 4070
rect 249 4036 283 4070
rect 317 4036 337 4070
rect 207 4020 337 4036
rect 139 3968 215 3986
rect 173 3952 215 3968
rect 249 3952 265 3986
rect 139 3876 173 3934
rect 299 3918 337 4020
rect 371 4235 421 4251
rect 405 4201 421 4235
rect 455 4244 945 4255
rect 455 4238 683 4244
rect 455 4204 471 4238
rect 505 4204 539 4238
rect 573 4204 607 4238
rect 641 4210 683 4238
rect 717 4238 945 4244
rect 717 4210 759 4238
rect 641 4204 759 4210
rect 793 4204 827 4238
rect 861 4204 895 4238
rect 929 4204 945 4238
rect 979 4235 1029 4251
rect 371 4154 421 4201
rect 405 4120 421 4154
rect 371 4070 421 4120
rect 405 4036 421 4070
rect 371 3991 421 4036
rect 371 3986 378 3991
rect 412 3957 421 3991
rect 405 3952 421 3957
rect 371 3927 421 3952
rect 455 4154 649 4170
rect 455 4120 471 4154
rect 505 4120 539 4154
rect 573 4120 607 4154
rect 641 4120 649 4154
rect 455 4104 649 4120
rect 683 4152 717 4204
rect 979 4201 995 4235
rect 455 4002 489 4104
rect 683 4070 717 4118
rect 751 4154 945 4170
rect 751 4120 759 4154
rect 793 4120 827 4154
rect 861 4120 895 4154
rect 929 4120 945 4154
rect 751 4104 945 4120
rect 523 4036 539 4070
rect 573 4036 607 4070
rect 641 4060 759 4070
rect 641 4036 683 4060
rect 717 4036 759 4060
rect 793 4036 827 4070
rect 861 4036 877 4070
rect 455 3986 649 4002
rect 455 3952 471 3986
rect 505 3952 539 3986
rect 573 3952 607 3986
rect 641 3952 649 3986
rect 455 3936 649 3952
rect 683 3968 717 4026
rect 911 4002 945 4104
rect 139 3784 173 3842
rect 139 3692 173 3750
rect 139 3600 173 3658
rect 139 3508 173 3566
rect 207 3902 337 3918
rect 207 3868 215 3902
rect 249 3868 283 3902
rect 317 3868 337 3902
rect 455 3891 489 3936
rect 751 3986 945 4002
rect 751 3952 759 3986
rect 793 3952 827 3986
rect 861 3952 895 3986
rect 929 3952 945 3986
rect 751 3936 945 3952
rect 683 3902 717 3934
rect 371 3875 489 3891
rect 207 3734 249 3868
rect 371 3841 445 3875
rect 479 3841 489 3875
rect 523 3868 539 3902
rect 573 3868 607 3902
rect 641 3876 759 3902
rect 641 3868 683 3876
rect 371 3834 489 3841
rect 717 3868 759 3876
rect 793 3868 827 3902
rect 861 3868 877 3902
rect 911 3891 945 3936
rect 979 4154 1029 4201
rect 979 4120 995 4154
rect 979 4070 1029 4120
rect 979 4036 995 4070
rect 979 3992 1029 4036
rect 979 3958 987 3992
rect 1021 3986 1029 3992
rect 979 3952 995 3958
rect 979 3927 1029 3952
rect 1063 4238 1193 4255
rect 1063 4204 1083 4238
rect 1117 4204 1151 4238
rect 1185 4204 1193 4238
rect 1063 4188 1193 4204
rect 1227 4244 1261 4290
rect 1063 4086 1101 4188
rect 1227 4154 1261 4210
rect 1135 4120 1151 4154
rect 1185 4152 1261 4154
rect 1185 4120 1227 4152
rect 1063 4070 1193 4086
rect 1063 4036 1083 4070
rect 1117 4036 1151 4070
rect 1185 4036 1193 4070
rect 1063 4020 1193 4036
rect 1227 4060 1261 4118
rect 1063 3918 1101 4020
rect 1227 3986 1261 4026
rect 1135 3952 1151 3986
rect 1185 3968 1261 3986
rect 1185 3952 1227 3968
rect 1063 3902 1193 3918
rect 911 3875 1029 3891
rect 207 3700 215 3734
rect 207 3566 249 3700
rect 283 3818 649 3834
rect 317 3784 471 3818
rect 505 3784 539 3818
rect 573 3784 607 3818
rect 641 3784 649 3818
rect 283 3650 317 3784
rect 455 3768 649 3784
rect 683 3784 717 3842
rect 911 3841 921 3875
rect 955 3841 1029 3875
rect 1063 3868 1083 3902
rect 1117 3868 1151 3902
rect 1185 3868 1193 3902
rect 911 3834 1029 3841
rect 283 3600 317 3616
rect 371 3734 421 3750
rect 405 3700 421 3734
rect 371 3650 421 3700
rect 405 3616 421 3650
rect 207 3532 215 3566
rect 249 3532 283 3566
rect 317 3532 333 3566
rect 207 3516 333 3532
rect 371 3548 421 3616
rect 455 3666 489 3768
rect 751 3818 1117 3834
rect 751 3784 759 3818
rect 793 3784 827 3818
rect 861 3784 895 3818
rect 929 3784 1083 3818
rect 751 3768 945 3784
rect 683 3734 717 3750
rect 523 3700 539 3734
rect 573 3700 607 3734
rect 641 3700 759 3734
rect 793 3700 827 3734
rect 861 3700 877 3734
rect 683 3692 717 3700
rect 455 3650 649 3666
rect 455 3616 471 3650
rect 505 3616 539 3650
rect 573 3616 607 3650
rect 641 3616 649 3650
rect 455 3600 649 3616
rect 911 3666 945 3768
rect 683 3600 717 3658
rect 751 3650 945 3666
rect 751 3616 759 3650
rect 793 3616 827 3650
rect 861 3616 895 3650
rect 929 3616 945 3650
rect 751 3600 945 3616
rect 979 3734 1029 3750
rect 979 3700 995 3734
rect 979 3650 1029 3700
rect 979 3616 995 3650
rect 139 3427 173 3474
rect 371 3514 377 3548
rect 411 3514 421 3548
rect 523 3532 539 3566
rect 573 3532 607 3566
rect 641 3532 759 3566
rect 793 3532 827 3566
rect 861 3532 877 3566
rect 523 3516 877 3532
rect 979 3563 1029 3616
rect 1083 3650 1117 3784
rect 1083 3600 1117 3616
rect 1151 3734 1193 3868
rect 1185 3700 1193 3734
rect 1151 3566 1193 3700
rect 979 3529 989 3563
rect 1023 3529 1029 3563
rect 371 3462 421 3514
rect 683 3508 717 3516
rect 683 3427 717 3474
rect 979 3462 1029 3529
rect 1067 3532 1083 3566
rect 1117 3532 1151 3566
rect 1185 3532 1193 3566
rect 1067 3516 1193 3532
rect 1227 3876 1261 3934
rect 1227 3784 1261 3842
rect 1227 3692 1261 3750
rect 1227 3600 1261 3658
rect 1227 3508 1261 3566
rect 1227 3427 1261 3474
rect 139 3416 341 3427
rect 173 3409 341 3416
rect 173 3382 219 3409
rect 139 3375 219 3382
rect 253 3375 287 3409
rect 321 3375 341 3409
rect 453 3416 947 3427
rect 453 3409 683 3416
rect 453 3375 471 3409
rect 505 3375 539 3409
rect 573 3375 607 3409
rect 641 3382 683 3409
rect 717 3409 947 3416
rect 717 3382 759 3409
rect 641 3375 759 3382
rect 793 3375 827 3409
rect 861 3375 895 3409
rect 929 3375 947 3409
rect 1059 3416 1261 3427
rect 1059 3409 1227 3416
rect 1059 3375 1079 3409
rect 1113 3375 1147 3409
rect 1181 3382 1227 3409
rect 1181 3375 1261 3382
rect 139 3324 173 3375
rect 139 3255 173 3290
rect 207 3325 377 3340
rect 207 3291 245 3325
rect 279 3306 377 3325
rect 411 3325 649 3340
rect 411 3306 502 3325
rect 279 3291 322 3306
rect 207 3289 322 3291
rect 468 3291 502 3306
rect 536 3291 583 3325
rect 617 3291 649 3325
rect 468 3289 649 3291
rect 683 3324 717 3375
rect 355 3255 371 3272
rect 139 3239 249 3255
rect 139 3232 215 3239
rect 173 3205 215 3232
rect 173 3198 249 3205
rect 139 3189 249 3198
rect 283 3238 371 3255
rect 405 3255 421 3272
rect 683 3255 717 3290
rect 751 3325 987 3340
rect 751 3291 783 3325
rect 817 3291 864 3325
rect 898 3306 987 3325
rect 1021 3325 1193 3340
rect 1021 3306 1121 3325
rect 898 3291 932 3306
rect 751 3289 932 3291
rect 1078 3291 1121 3306
rect 1155 3291 1193 3325
rect 1078 3289 1193 3291
rect 1227 3324 1261 3375
rect 979 3255 995 3272
rect 405 3238 497 3255
rect 283 3221 497 3238
rect 139 3140 173 3189
rect 283 3146 317 3221
rect 207 3112 228 3146
rect 262 3112 317 3146
rect 353 3148 427 3165
rect 353 3114 371 3148
rect 405 3114 427 3148
rect 139 3077 173 3106
rect 353 3094 427 3114
rect 463 3146 497 3221
rect 531 3239 869 3255
rect 565 3205 599 3239
rect 633 3232 767 3239
rect 633 3205 683 3232
rect 531 3198 683 3205
rect 717 3205 767 3232
rect 801 3205 835 3239
rect 717 3198 869 3205
rect 531 3189 869 3198
rect 903 3238 995 3255
rect 1029 3255 1045 3272
rect 1227 3255 1261 3290
rect 1029 3238 1117 3255
rect 903 3221 1117 3238
rect 463 3112 531 3146
rect 565 3112 599 3146
rect 633 3112 649 3146
rect 683 3140 717 3189
rect 903 3146 937 3221
rect 751 3112 767 3146
rect 801 3112 835 3146
rect 869 3112 937 3146
rect 973 3148 1047 3165
rect 973 3114 995 3148
rect 1029 3114 1047 3148
rect 683 3077 717 3106
rect 973 3094 1047 3114
rect 1083 3146 1117 3221
rect 1151 3239 1261 3255
rect 1185 3232 1261 3239
rect 1185 3205 1227 3232
rect 1151 3198 1227 3205
rect 1151 3189 1261 3198
rect 1083 3112 1138 3146
rect 1172 3112 1193 3146
rect 1227 3140 1261 3189
rect 1227 3077 1261 3106
rect 281 2943 377 2977
rect 1023 2943 1119 2977
rect 281 2881 315 2943
rect -4 2642 30 2658
rect -4 2550 30 2566
rect 84 2642 118 2658
rect 84 2550 118 2566
rect 170 2642 204 2658
rect 170 2550 204 2566
rect 42 2473 84 2507
rect 118 2473 159 2507
rect 1085 2881 1119 2943
rect 667 2841 683 2875
rect 717 2841 733 2875
rect 315 2773 425 2807
rect 459 2773 475 2807
rect 523 2773 539 2807
rect 573 2773 589 2807
rect 811 2773 827 2807
rect 861 2773 877 2807
rect 925 2773 941 2807
rect 975 2773 1085 2807
rect 395 2714 429 2773
rect 395 2622 429 2638
rect 491 2722 525 2730
rect 491 2622 525 2638
rect 587 2714 621 2730
rect 587 2582 621 2638
rect 683 2714 717 2730
rect 779 2714 813 2730
rect 395 2492 429 2508
rect 395 2357 429 2416
rect 491 2492 525 2508
rect 491 2400 525 2408
rect 587 2492 621 2548
rect 779 2582 813 2638
rect 875 2722 909 2730
rect 875 2622 909 2638
rect 971 2714 1005 2773
rect 971 2622 1005 2638
rect 587 2400 621 2416
rect 683 2400 717 2416
rect 779 2492 813 2548
rect 779 2400 813 2416
rect 875 2492 909 2508
rect 875 2400 909 2408
rect 971 2492 1005 2508
rect 971 2357 1005 2416
rect 315 2323 425 2357
rect 459 2323 475 2357
rect 523 2323 539 2357
rect 573 2323 589 2357
rect 811 2323 827 2357
rect 861 2323 877 2357
rect 925 2323 941 2357
rect 975 2323 1085 2357
rect 667 2255 683 2289
rect 717 2255 733 2289
rect 281 2187 315 2249
rect 1244 2367 1278 2383
rect 1244 2275 1278 2291
rect 1332 2367 1366 2383
rect 1332 2275 1366 2291
rect 1418 2367 1452 2383
rect 1418 2275 1452 2291
rect 1085 2187 1119 2249
rect 1290 2198 1332 2232
rect 1366 2198 1407 2232
rect 281 2153 377 2187
rect 1023 2153 1119 2187
rect -4 2047 92 2081
rect 1308 2047 1404 2081
rect -4 1985 30 2047
rect 158 1979 192 2047
rect 1208 1979 1242 2047
rect 1370 1985 1404 2047
rect 110 1945 158 1979
rect 192 1945 240 1979
rect 352 1945 368 1979
rect 402 1945 998 1979
rect 1032 1945 1048 1979
rect 1160 1945 1208 1979
rect 1242 1945 1290 1979
rect 110 1895 144 1945
rect 110 1769 144 1819
rect 206 1895 240 1945
rect 206 1769 240 1819
rect 320 1905 354 1911
rect 320 1803 354 1819
rect 416 1905 450 1911
rect 416 1803 450 1819
rect 530 1909 564 1911
rect 530 1803 564 1819
rect 626 1895 660 1911
rect 626 1803 660 1809
rect 740 1895 774 1911
rect 740 1803 774 1809
rect 836 1909 870 1911
rect 836 1803 870 1819
rect 950 1905 984 1911
rect 950 1803 984 1819
rect 1046 1905 1080 1911
rect 1046 1803 1080 1819
rect 1160 1895 1194 1945
rect 1160 1769 1194 1819
rect 1256 1895 1290 1945
rect 1256 1769 1290 1819
rect 110 1735 158 1769
rect 192 1735 240 1769
rect 562 1735 578 1769
rect 612 1735 788 1769
rect 822 1735 838 1769
rect 1160 1735 1208 1769
rect 1242 1735 1290 1769
rect -4 1667 30 1729
rect 158 1667 192 1735
rect 1208 1667 1242 1735
rect 1370 1667 1404 1729
rect -4 1633 92 1667
rect 1308 1633 1404 1667
rect 281 1527 377 1561
rect 1023 1527 1119 1561
rect 281 1465 315 1527
rect 1085 1465 1119 1527
rect 667 1425 683 1459
rect 717 1425 733 1459
rect 315 1357 425 1391
rect 459 1357 475 1391
rect 523 1357 539 1391
rect 573 1357 589 1391
rect 811 1357 827 1391
rect 861 1357 877 1391
rect 925 1357 941 1391
rect 975 1357 1085 1391
rect 395 1307 429 1357
rect 395 1215 429 1231
rect 491 1315 525 1323
rect 491 1215 525 1231
rect 587 1307 621 1323
rect 587 1175 621 1231
rect 683 1307 717 1323
rect 779 1307 813 1323
rect 779 1175 813 1231
rect 875 1315 909 1323
rect 875 1215 909 1231
rect 971 1307 1005 1357
rect 971 1215 1005 1231
rect 621 1141 779 1175
rect 395 1085 429 1101
rect 395 959 429 1009
rect 491 1085 525 1101
rect 491 993 525 1001
rect 587 1085 621 1141
rect 587 993 621 1009
rect 683 993 717 1009
rect 779 1085 813 1141
rect 779 993 813 1009
rect 875 1085 909 1101
rect 875 993 909 1001
rect 971 1085 1005 1101
rect 971 959 1005 1009
rect 315 925 425 959
rect 459 925 475 959
rect 523 925 539 959
rect 573 925 589 959
rect 811 925 827 959
rect 861 925 877 959
rect 925 925 941 959
rect 975 925 1085 959
rect 667 857 683 891
rect 717 857 733 891
rect 281 789 315 851
rect 1085 789 1119 851
rect 281 755 377 789
rect 1023 755 1119 789
rect 88 650 184 684
rect 1214 650 1310 684
rect 88 588 122 650
rect 88 268 122 330
rect 202 582 236 650
rect 202 548 232 582
rect 266 548 282 582
rect 202 498 236 548
rect 202 370 236 420
rect 298 498 332 514
rect 298 404 332 420
rect 394 498 428 650
rect 394 404 428 420
rect 490 498 524 514
rect 490 404 524 420
rect 586 498 620 650
rect 586 404 620 420
rect 682 498 716 514
rect 682 404 716 420
rect 778 498 812 650
rect 778 404 812 420
rect 874 498 908 514
rect 874 404 908 420
rect 970 498 1004 650
rect 1162 582 1196 650
rect 1116 548 1132 582
rect 1166 548 1196 582
rect 970 404 1004 420
rect 1066 498 1100 514
rect 1066 404 1100 420
rect 1162 498 1196 548
rect 1162 370 1196 420
rect 202 336 232 370
rect 266 336 282 370
rect 378 336 394 370
rect 428 336 444 370
rect 570 336 586 370
rect 620 336 636 370
rect 762 336 778 370
rect 812 336 828 370
rect 936 336 952 370
rect 986 336 1002 370
rect 1116 336 1132 370
rect 1166 336 1196 370
rect 202 269 236 336
rect 1162 269 1196 336
rect 1276 588 1310 650
rect 1276 268 1310 330
rect 88 234 184 268
rect 1214 234 1310 268
<< viali >>
rect 139 4670 173 4704
rect 139 4578 173 4612
rect 683 4670 717 4704
rect 683 4578 717 4612
rect 1227 4670 1261 4704
rect 1227 4578 1261 4612
rect 139 4486 173 4520
rect 139 4394 173 4428
rect 683 4486 717 4520
rect 683 4394 717 4428
rect 1227 4486 1261 4520
rect 1227 4394 1261 4428
rect 139 4302 173 4336
rect 683 4302 717 4336
rect 1227 4302 1261 4336
rect 139 4210 173 4244
rect 139 4118 173 4152
rect 139 4026 173 4060
rect 139 3934 173 3968
rect 683 4210 717 4244
rect 378 3986 412 3991
rect 378 3957 405 3986
rect 405 3957 412 3986
rect 683 4118 717 4152
rect 683 4026 717 4060
rect 139 3842 173 3876
rect 139 3750 173 3784
rect 139 3658 173 3692
rect 139 3566 173 3600
rect 683 3934 717 3968
rect 445 3841 479 3875
rect 683 3842 717 3876
rect 987 3986 1021 3992
rect 987 3958 995 3986
rect 995 3958 1021 3986
rect 1227 4210 1261 4244
rect 1227 4118 1261 4152
rect 1227 4026 1261 4060
rect 1227 3934 1261 3968
rect 921 3841 955 3875
rect 683 3750 717 3784
rect 683 3658 717 3692
rect 683 3566 717 3600
rect 139 3474 173 3508
rect 377 3514 411 3548
rect 989 3529 1023 3563
rect 683 3474 717 3508
rect 1227 3842 1261 3876
rect 1227 3750 1261 3784
rect 1227 3658 1261 3692
rect 1227 3566 1261 3600
rect 1227 3474 1261 3508
rect 139 3382 173 3416
rect 683 3382 717 3416
rect 1227 3382 1261 3416
rect 139 3290 173 3324
rect 377 3306 411 3340
rect 683 3290 717 3324
rect 139 3198 173 3232
rect 987 3306 1021 3340
rect 1227 3290 1261 3324
rect 139 3106 173 3140
rect 371 3114 405 3148
rect 683 3198 717 3232
rect 683 3106 717 3140
rect 995 3114 1029 3148
rect 1227 3198 1261 3232
rect 1227 3106 1261 3140
rect 377 2943 1023 2977
rect -4 2566 30 2642
rect 84 2566 118 2642
rect 170 2566 204 2642
rect 84 2473 118 2507
rect 683 2841 717 2875
rect 539 2773 573 2807
rect 827 2773 861 2807
rect 491 2714 525 2722
rect 491 2688 525 2714
rect 683 2638 717 2654
rect 683 2620 717 2638
rect 587 2548 621 2582
rect 491 2416 525 2442
rect 491 2408 525 2416
rect 875 2714 909 2722
rect 875 2688 909 2714
rect 779 2548 813 2582
rect 683 2492 717 2510
rect 683 2476 717 2492
rect 875 2416 909 2442
rect 875 2408 909 2416
rect 539 2323 573 2357
rect 827 2323 861 2357
rect 683 2255 717 2289
rect 1244 2291 1278 2367
rect 1332 2291 1366 2367
rect 1418 2291 1452 2367
rect 1332 2198 1366 2232
rect -4 1729 30 1985
rect 368 1945 402 1979
rect 998 1945 1032 1979
rect 320 1895 354 1905
rect 320 1871 354 1895
rect 416 1895 450 1905
rect 416 1871 450 1895
rect 530 1895 564 1909
rect 530 1875 564 1895
rect 626 1819 660 1843
rect 626 1809 660 1819
rect 740 1819 774 1843
rect 740 1809 774 1819
rect 836 1895 870 1909
rect 836 1875 870 1895
rect 950 1895 984 1905
rect 950 1871 984 1895
rect 1046 1895 1080 1905
rect 1046 1871 1080 1895
rect 578 1735 612 1769
rect 788 1735 822 1769
rect 1370 1729 1404 1985
rect 377 1527 1023 1561
rect 683 1425 717 1459
rect 539 1357 573 1391
rect 827 1357 861 1391
rect 491 1307 525 1315
rect 491 1281 525 1307
rect 683 1231 717 1247
rect 683 1213 717 1231
rect 875 1307 909 1315
rect 875 1281 909 1307
rect 587 1141 621 1175
rect 779 1141 813 1175
rect 491 1009 525 1035
rect 491 1001 525 1009
rect 683 1085 717 1103
rect 683 1069 717 1085
rect 875 1009 909 1035
rect 875 1001 909 1009
rect 539 925 573 959
rect 827 925 861 959
rect 683 857 717 891
rect 377 755 1023 789
rect 298 442 332 476
rect 490 442 524 476
rect 682 442 716 476
rect 874 442 908 476
rect 1066 442 1100 476
rect 394 336 428 370
rect 586 336 620 370
rect 778 336 812 370
rect 952 336 986 370
rect 184 268 1214 269
rect 184 235 1214 268
<< metal1 >>
rect 108 4704 204 4870
rect 108 4670 139 4704
rect 173 4670 204 4704
rect 108 4612 204 4670
rect 108 4578 139 4612
rect 173 4578 204 4612
rect 108 4520 204 4578
rect 108 4486 139 4520
rect 173 4486 204 4520
rect 108 4428 204 4486
rect 108 4394 139 4428
rect 173 4394 204 4428
rect 108 4336 204 4394
rect 108 4302 139 4336
rect 173 4302 204 4336
rect 108 4244 204 4302
rect 108 4210 139 4244
rect 173 4210 204 4244
rect 108 4152 204 4210
rect 108 4118 139 4152
rect 173 4118 204 4152
rect 108 4060 204 4118
rect 108 4026 139 4060
rect 173 4026 204 4060
rect 108 3968 204 4026
rect 108 3934 139 3968
rect 173 3934 204 3968
rect 108 3876 204 3934
rect 108 3842 139 3876
rect 173 3842 204 3876
rect 108 3784 204 3842
rect 266 3881 300 4870
rect 652 4704 748 4870
rect 652 4670 683 4704
rect 717 4670 748 4704
rect 652 4612 748 4670
rect 652 4578 683 4612
rect 717 4578 748 4612
rect 652 4520 748 4578
rect 652 4486 683 4520
rect 717 4486 748 4520
rect 652 4428 748 4486
rect 652 4394 683 4428
rect 717 4394 748 4428
rect 652 4336 748 4394
rect 652 4302 683 4336
rect 717 4302 748 4336
rect 652 4244 748 4302
rect 652 4210 683 4244
rect 717 4210 748 4244
rect 652 4152 748 4210
rect 652 4118 683 4152
rect 717 4118 748 4152
rect 652 4060 748 4118
rect 652 4026 683 4060
rect 717 4026 748 4060
rect 359 3947 369 3999
rect 421 3947 431 3999
rect 652 3968 748 4026
rect 652 3934 683 3968
rect 717 3934 748 3968
rect 853 3947 863 3999
rect 915 3947 925 3999
rect 967 3949 977 4001
rect 1029 3949 1039 4001
rect 517 3881 527 3884
rect 266 3875 527 3881
rect 266 3841 445 3875
rect 479 3841 527 3875
rect 266 3835 527 3841
rect 517 3832 527 3835
rect 579 3832 589 3884
rect 652 3876 748 3934
rect 652 3842 683 3876
rect 717 3842 748 3876
rect 108 3750 139 3784
rect 173 3750 204 3784
rect 108 3692 204 3750
rect 108 3658 139 3692
rect 173 3658 204 3692
rect 108 3600 204 3658
rect 108 3566 139 3600
rect 173 3566 204 3600
rect 108 3508 204 3566
rect 652 3784 748 3842
rect 867 3881 911 3947
rect 1100 3881 1134 4870
rect 867 3875 1134 3881
rect 867 3841 921 3875
rect 955 3841 1134 3875
rect 867 3835 1134 3841
rect 1196 4704 1292 4870
rect 1196 4670 1227 4704
rect 1261 4670 1292 4704
rect 1196 4612 1292 4670
rect 1196 4578 1227 4612
rect 1261 4578 1292 4612
rect 1196 4520 1292 4578
rect 1196 4486 1227 4520
rect 1261 4486 1292 4520
rect 1196 4428 1292 4486
rect 1196 4394 1227 4428
rect 1261 4394 1292 4428
rect 1196 4336 1292 4394
rect 1196 4302 1227 4336
rect 1261 4302 1292 4336
rect 1196 4244 1292 4302
rect 1196 4210 1227 4244
rect 1261 4210 1292 4244
rect 1196 4152 1292 4210
rect 1196 4118 1227 4152
rect 1261 4118 1292 4152
rect 1196 4060 1292 4118
rect 1196 4026 1227 4060
rect 1261 4026 1292 4060
rect 1196 3968 1292 4026
rect 1196 3934 1227 3968
rect 1261 3934 1292 3968
rect 1196 3876 1292 3934
rect 1196 3842 1227 3876
rect 1261 3842 1292 3876
rect 652 3750 683 3784
rect 717 3750 748 3784
rect 652 3692 748 3750
rect 652 3658 683 3692
rect 717 3658 748 3692
rect 652 3600 748 3658
rect 652 3566 683 3600
rect 717 3566 748 3600
rect 1196 3784 1292 3842
rect 1196 3750 1227 3784
rect 1261 3750 1292 3784
rect 1196 3692 1292 3750
rect 1196 3658 1227 3692
rect 1261 3658 1292 3692
rect 1196 3600 1292 3658
rect 108 3474 139 3508
rect 173 3474 204 3508
rect 108 3416 204 3474
rect 108 3382 139 3416
rect 173 3382 204 3416
rect 108 3324 204 3382
rect 108 3290 139 3324
rect 173 3290 204 3324
rect 365 3548 423 3556
rect 365 3514 377 3548
rect 411 3514 423 3548
rect 365 3340 423 3514
rect 365 3306 377 3340
rect 411 3306 423 3340
rect 365 3300 423 3306
rect 652 3508 748 3566
rect 652 3474 683 3508
rect 717 3474 748 3508
rect 652 3416 748 3474
rect 652 3382 683 3416
rect 717 3382 748 3416
rect 652 3324 748 3382
rect 977 3563 1035 3569
rect 977 3529 989 3563
rect 1023 3529 1035 3563
rect 977 3523 1035 3529
rect 1196 3566 1227 3600
rect 1261 3566 1292 3600
rect 977 3346 1033 3523
rect 108 3232 204 3290
rect 108 3198 139 3232
rect 173 3198 204 3232
rect 108 3140 204 3198
rect 652 3290 683 3324
rect 717 3290 748 3324
rect 975 3340 1033 3346
rect 975 3306 987 3340
rect 1021 3306 1033 3340
rect 975 3300 1033 3306
rect 1196 3508 1292 3566
rect 1196 3474 1227 3508
rect 1261 3474 1292 3508
rect 1196 3416 1292 3474
rect 1196 3382 1227 3416
rect 1261 3382 1292 3416
rect 1196 3324 1292 3382
rect 652 3232 748 3290
rect 652 3198 683 3232
rect 717 3198 748 3232
rect 108 3106 139 3140
rect 173 3106 204 3140
rect 108 3077 204 3106
rect 350 3105 360 3157
rect 412 3105 422 3157
rect 652 3140 748 3198
rect 1196 3290 1227 3324
rect 1261 3290 1292 3324
rect 1196 3232 1292 3290
rect 1196 3198 1227 3232
rect 1261 3198 1292 3232
rect 652 3106 683 3140
rect 717 3106 748 3140
rect 974 3106 984 3158
rect 1036 3106 1046 3158
rect 1196 3140 1292 3198
rect 1196 3106 1227 3140
rect 1261 3106 1292 3140
rect 652 2985 748 3106
rect 1196 3077 1292 3106
rect 652 2983 673 2985
rect 245 2977 673 2983
rect 727 2983 748 2985
rect 727 2979 1155 2983
rect 727 2977 1365 2979
rect 85 2943 377 2977
rect 1023 2945 1365 2977
rect 1023 2943 1155 2945
rect 85 2654 119 2943
rect 245 2936 673 2943
rect 663 2933 673 2936
rect 727 2936 1155 2943
rect 727 2933 737 2936
rect 397 2875 407 2893
rect 245 2841 407 2875
rect 459 2875 469 2893
rect 671 2875 729 2881
rect 459 2841 683 2875
rect 717 2841 763 2875
rect 671 2835 729 2841
rect 527 2807 585 2813
rect 815 2807 873 2813
rect 931 2807 941 2825
rect 523 2773 539 2807
rect 573 2773 827 2807
rect 861 2773 941 2807
rect 993 2807 1003 2825
rect 993 2773 1155 2807
rect 527 2767 585 2773
rect 815 2767 873 2773
rect 479 2722 537 2728
rect 863 2722 921 2728
rect 479 2688 491 2722
rect 525 2688 875 2722
rect 909 2688 1159 2722
rect 479 2682 537 2688
rect 863 2682 921 2688
rect 671 2654 729 2660
rect -10 2642 36 2654
rect -10 2630 -4 2642
rect 30 2630 36 2642
rect 78 2642 124 2654
rect -31 2578 -21 2630
rect 31 2578 41 2630
rect -10 2566 -4 2578
rect 30 2566 36 2578
rect -10 2554 36 2566
rect 78 2566 84 2642
rect 118 2566 124 2642
rect 78 2554 124 2566
rect 164 2642 245 2654
rect 164 2566 170 2642
rect 204 2602 245 2642
rect 297 2620 683 2654
rect 717 2620 729 2654
rect 297 2602 307 2620
rect 204 2566 210 2602
rect 164 2554 210 2566
rect 72 2507 130 2513
rect -171 2473 84 2507
rect 118 2473 161 2507
rect 72 2467 130 2473
rect 395 2442 429 2620
rect 671 2614 729 2620
rect 567 2540 577 2592
rect 629 2582 639 2592
rect 761 2582 771 2592
rect 629 2548 771 2582
rect 629 2540 639 2548
rect 761 2540 771 2548
rect 823 2540 833 2592
rect 671 2510 729 2516
rect 971 2510 1005 2688
rect 1149 2670 1159 2688
rect 1211 2670 1221 2722
rect 671 2476 683 2510
rect 717 2476 1005 2510
rect 671 2470 729 2476
rect 479 2442 537 2448
rect 863 2442 921 2448
rect 395 2408 491 2442
rect 525 2408 875 2442
rect 909 2408 921 2442
rect 479 2402 537 2408
rect 863 2402 921 2408
rect 1331 2379 1365 2945
rect 1238 2367 1284 2379
rect 1238 2366 1244 2367
rect 527 2357 585 2363
rect 815 2357 873 2363
rect 1149 2357 1159 2366
rect 397 2305 407 2357
rect 459 2323 539 2357
rect 573 2323 827 2357
rect 861 2323 1159 2357
rect 459 2305 469 2323
rect 527 2317 585 2323
rect 815 2317 873 2323
rect 1149 2314 1159 2323
rect 1211 2314 1244 2366
rect 671 2289 729 2295
rect 1238 2291 1244 2314
rect 1278 2291 1284 2367
rect 637 2288 683 2289
rect 235 2255 245 2264
rect 158 2221 245 2255
rect -40 1985 36 1997
rect -40 1884 -4 1985
rect -128 1831 -4 1884
rect -40 1729 -4 1831
rect 30 1729 36 1985
rect 158 1769 192 2221
rect 235 2212 245 2221
rect 297 2255 307 2264
rect 523 2255 683 2288
rect 717 2255 941 2289
rect 297 2221 557 2255
rect 671 2249 729 2255
rect 931 2237 941 2255
rect 993 2237 1003 2289
rect 1238 2279 1284 2291
rect 1326 2367 1372 2379
rect 1326 2291 1332 2367
rect 1366 2291 1372 2367
rect 1412 2367 1458 2379
rect 1412 2355 1418 2367
rect 1452 2355 1458 2367
rect 1409 2303 1418 2355
rect 1471 2303 1481 2355
rect 1326 2279 1372 2291
rect 1412 2291 1418 2303
rect 1452 2291 1458 2303
rect 1412 2279 1458 2291
rect 1320 2232 1378 2238
rect 297 2212 307 2221
rect 1289 2198 1332 2232
rect 1366 2198 1571 2232
rect 1320 2192 1378 2198
rect 356 1979 414 1985
rect 986 1979 1044 1985
rect 1148 1979 1158 1997
rect 352 1945 368 1979
rect 402 1945 998 1979
rect 1032 1945 1158 1979
rect 1210 1979 1218 1997
rect 1364 1985 1440 1997
rect 1210 1945 1278 1979
rect 356 1939 414 1945
rect 986 1939 1044 1945
rect 308 1905 366 1911
rect 292 1853 302 1905
rect 354 1865 366 1905
rect 404 1905 462 1911
rect 518 1909 576 1915
rect 824 1909 882 1915
rect 404 1865 416 1905
rect 354 1853 364 1865
rect 406 1853 416 1865
rect 468 1853 478 1905
rect 518 1875 530 1909
rect 564 1877 836 1909
rect 564 1875 576 1877
rect 518 1869 576 1875
rect 824 1875 836 1877
rect 870 1875 882 1909
rect 938 1905 996 1911
rect 824 1859 882 1875
rect 614 1843 674 1849
rect 614 1809 626 1843
rect 660 1809 674 1843
rect 614 1803 674 1809
rect 664 1797 674 1803
rect 726 1843 786 1849
rect 726 1809 740 1843
rect 774 1809 786 1843
rect 726 1803 786 1809
rect 824 1807 836 1859
rect 888 1807 894 1859
rect 926 1853 932 1905
rect 984 1865 996 1905
rect 1034 1905 1092 1911
rect 1034 1865 1046 1905
rect 984 1853 994 1865
rect 1036 1853 1046 1865
rect 1098 1853 1108 1905
rect 726 1797 736 1803
rect 566 1769 624 1775
rect 776 1773 834 1775
rect 770 1769 834 1773
rect 158 1735 578 1769
rect 612 1735 788 1769
rect 822 1735 838 1769
rect 566 1729 624 1735
rect 776 1729 834 1735
rect 1364 1729 1370 1985
rect 1404 1883 1440 1985
rect 1404 1827 1585 1883
rect 1404 1729 1440 1827
rect -40 1717 36 1729
rect 1364 1717 1440 1729
rect -171 1561 1571 1567
rect -171 1527 377 1561
rect 1023 1527 1571 1561
rect -171 1521 1571 1527
rect 397 1459 407 1477
rect -171 1425 407 1459
rect 459 1459 469 1477
rect 671 1459 729 1465
rect 459 1425 683 1459
rect 717 1425 763 1459
rect 671 1419 729 1425
rect 527 1391 585 1397
rect 815 1391 873 1397
rect 931 1391 941 1409
rect 523 1357 539 1391
rect 573 1357 827 1391
rect 861 1357 941 1391
rect 993 1391 1003 1409
rect 993 1357 1571 1391
rect 527 1351 585 1357
rect 815 1351 873 1357
rect 479 1315 537 1321
rect 863 1315 921 1321
rect 479 1281 491 1315
rect 525 1281 875 1315
rect 909 1281 1103 1315
rect 479 1275 537 1281
rect 863 1275 921 1281
rect 235 1213 245 1265
rect 297 1247 307 1265
rect 671 1247 729 1253
rect 297 1213 683 1247
rect 717 1213 729 1247
rect 395 1035 429 1213
rect 671 1207 729 1213
rect 567 1133 577 1185
rect 629 1175 639 1185
rect 761 1175 771 1185
rect 629 1141 771 1175
rect 629 1133 639 1141
rect 761 1133 771 1141
rect 823 1133 833 1185
rect 671 1103 729 1109
rect 971 1103 1005 1281
rect 1093 1263 1103 1281
rect 1155 1263 1165 1315
rect 671 1069 683 1103
rect 717 1069 1005 1103
rect 671 1063 729 1069
rect 479 1035 537 1041
rect 863 1035 921 1041
rect 395 1001 491 1035
rect 525 1001 875 1035
rect 909 1001 971 1035
rect 479 995 537 1001
rect 863 995 921 1001
rect 527 959 585 965
rect 815 959 873 965
rect 397 907 407 959
rect 459 925 539 959
rect 573 925 827 959
rect 861 925 877 959
rect 459 907 469 925
rect 527 919 585 925
rect 815 919 873 925
rect 671 891 729 897
rect 637 857 683 891
rect 717 857 941 891
rect 671 851 729 857
rect 931 839 941 857
rect 993 839 1003 891
rect -171 789 1571 795
rect -171 755 377 789
rect 1023 755 1571 789
rect -171 749 1571 755
rect 286 476 344 482
rect 478 476 536 482
rect 664 476 674 485
rect 726 476 736 485
rect 862 476 920 482
rect 1054 476 1112 482
rect 286 442 298 476
rect 332 442 490 476
rect 524 442 674 476
rect 726 442 874 476
rect 908 442 1066 476
rect 1100 442 1112 476
rect 286 436 344 442
rect 478 436 536 442
rect 664 433 674 442
rect 726 433 736 442
rect 862 436 920 442
rect 1054 436 1112 442
rect 382 371 440 376
rect 574 371 632 376
rect 766 371 824 376
rect 940 371 998 376
rect -171 370 1050 371
rect -171 337 394 370
rect 348 336 394 337
rect 428 336 586 370
rect 620 336 778 370
rect 812 336 952 370
rect 986 336 1050 370
rect 382 330 440 336
rect 574 330 632 336
rect 766 330 824 336
rect 940 330 998 336
rect -147 269 1571 275
rect -147 235 184 269
rect 1214 235 1571 269
rect -147 229 1571 235
<< via1 >>
rect 369 3991 421 3999
rect 369 3957 378 3991
rect 378 3957 412 3991
rect 412 3957 421 3991
rect 369 3947 421 3957
rect 863 3947 915 3999
rect 977 3992 1029 4001
rect 977 3958 987 3992
rect 987 3958 1021 3992
rect 1021 3958 1029 3992
rect 977 3949 1029 3958
rect 527 3832 579 3884
rect 360 3148 412 3157
rect 360 3114 371 3148
rect 371 3114 405 3148
rect 405 3114 412 3148
rect 360 3105 412 3114
rect 984 3148 1036 3158
rect 984 3114 995 3148
rect 995 3114 1029 3148
rect 1029 3114 1036 3148
rect 984 3106 1036 3114
rect 673 2977 727 2985
rect 673 2943 727 2977
rect 673 2933 727 2943
rect 407 2841 459 2893
rect 941 2773 993 2825
rect -21 2578 -4 2630
rect -4 2578 30 2630
rect 30 2578 31 2630
rect 245 2602 297 2654
rect 577 2582 629 2592
rect 771 2582 823 2592
rect 577 2548 587 2582
rect 587 2548 621 2582
rect 621 2548 629 2582
rect 771 2548 779 2582
rect 779 2548 813 2582
rect 813 2548 823 2582
rect 577 2540 629 2548
rect 771 2540 823 2548
rect 1159 2670 1211 2722
rect 407 2305 459 2357
rect 1159 2314 1211 2366
rect 245 2212 297 2264
rect 941 2237 993 2289
rect 1419 2303 1452 2355
rect 1452 2303 1471 2355
rect 1158 1945 1210 1997
rect 302 1871 320 1905
rect 320 1871 354 1905
rect 302 1853 354 1871
rect 416 1871 450 1905
rect 450 1871 468 1905
rect 416 1853 468 1871
rect 674 1797 726 1849
rect 836 1807 888 1859
rect 932 1871 950 1905
rect 950 1871 984 1905
rect 932 1853 984 1871
rect 1046 1871 1080 1905
rect 1080 1871 1098 1905
rect 1046 1853 1098 1871
rect 407 1425 459 1477
rect 941 1357 993 1409
rect 245 1213 297 1265
rect 577 1175 629 1185
rect 771 1175 823 1185
rect 577 1141 587 1175
rect 587 1141 621 1175
rect 621 1141 629 1175
rect 771 1141 779 1175
rect 779 1141 813 1175
rect 813 1141 823 1175
rect 577 1133 629 1141
rect 771 1133 823 1141
rect 1103 1263 1155 1315
rect 407 907 459 959
rect 941 839 993 891
rect 674 476 726 485
rect 674 442 682 476
rect 682 442 716 476
rect 716 442 726 476
rect 674 433 726 442
<< metal2 >>
rect 369 3999 421 4009
rect 863 3999 915 4009
rect 421 3947 863 3999
rect 369 3937 421 3947
rect 863 3937 915 3947
rect 977 4001 1029 4011
rect 527 3884 579 3894
rect 977 3884 1029 3949
rect 579 3832 1029 3884
rect 527 3822 579 3832
rect 360 3157 412 3167
rect 245 3105 360 3151
rect 984 3158 1036 3168
rect 412 3105 428 3151
rect 245 3099 428 3105
rect 973 3106 984 3154
rect 1036 3106 1211 3154
rect 973 3102 1211 3106
rect 245 2654 297 3099
rect 360 3095 412 3099
rect 984 3096 1036 3102
rect 673 2985 727 2995
rect -21 2630 31 2640
rect -21 1769 31 2578
rect 245 2264 297 2602
rect 407 2893 459 2903
rect 407 2357 459 2841
rect 673 2592 727 2933
rect 941 2825 993 2835
rect 571 2540 577 2592
rect 629 2540 771 2592
rect 823 2540 829 2592
rect 407 2295 459 2305
rect 941 2289 993 2773
rect 941 2227 993 2237
rect 1159 2722 1211 3102
rect 1159 2366 1211 2670
rect 245 2007 297 2212
rect 1159 2007 1211 2314
rect 245 1973 1098 2007
rect 302 1905 354 1973
rect 240 1853 302 1881
rect 240 1847 354 1853
rect 416 1905 984 1929
rect 468 1895 932 1905
rect 836 1859 888 1867
rect 416 1769 468 1853
rect -21 1735 468 1769
rect 674 1849 726 1859
rect -21 1726 31 1735
rect 245 1265 297 1735
rect 674 1711 726 1797
rect 932 1847 984 1853
rect 1046 1905 1098 1973
rect 1046 1847 1098 1853
rect 1158 1997 1211 2007
rect 1210 1945 1211 1997
rect 1419 2355 1471 2365
rect 1158 1935 1210 1945
rect 836 1791 888 1807
rect 1158 1791 1194 1935
rect 836 1755 1194 1791
rect 1419 1711 1471 2303
rect 674 1677 1471 1711
rect 245 1203 297 1213
rect 407 1477 459 1487
rect 407 959 459 1425
rect 941 1409 993 1419
rect 571 1133 577 1185
rect 629 1133 771 1185
rect 823 1133 829 1185
rect 407 897 459 907
rect 673 755 727 1133
rect 941 891 993 1357
rect 1103 1315 1155 1677
rect 1419 1667 1471 1677
rect 1103 1253 1155 1263
rect 941 829 993 839
rect 674 485 726 755
rect 674 423 726 433
<< labels >>
flabel metal1 283 4868 283 4868 5 FreeSans 400 0 0 0 outp
port 4 s
flabel metal1 1117 4868 1117 4868 5 FreeSans 400 0 0 0 outn
port 5 s
flabel metal1 -166 2489 -166 2489 3 FreeSans 400 0 0 0 clk
port 1 e
flabel metal1 1564 2214 1564 2214 1 FreeSans 400 0 0 0 clk
port 1 n
flabel metal1 -123 1858 -123 1858 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 1582 1855 1582 1855 7 FreeSans 400 0 0 0 VSS
port 7 w power bidirectional
flabel metal1 -166 1544 -166 1544 3 FreeSans 400 0 0 0 VSS
port 7 e power bidirectional
flabel metal1 -164 771 -164 771 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 -134 250 -134 250 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 -165 1442 -165 1442 1 FreeSans 400 0 0 0 ip
port 2 n
flabel metal1 1563 1373 1563 1373 1 FreeSans 400 0 0 0 in
port 3 n
flabel metal1 -160 353 -160 353 1 FreeSans 400 0 0 0 clk
port 1 n
flabel metal1 156 4865 156 4865 5 FreeSans 400 0 0 0 VSS
port 7 s power bidirectional
flabel metal1 1243 4868 1243 4868 5 FreeSans 400 0 0 0 VSS
port 7 s power bidirectional
flabel metal1 700 4864 700 4864 1 FreeSans 800 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 683 3106 717 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VPWR
flabel metal1 1227 3106 1261 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VGND
flabel locali 683 3106 717 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VPWR
flabel locali 1227 3106 1261 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VGND
flabel locali 1125 3289 1159 3323 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/X
flabel locali 853 3289 887 3323 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/X
flabel locali 785 3289 819 3323 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/X
flabel locali 989 3106 1023 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/A
flabel nwell 683 3106 717 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VPB
flabel pwell 1227 3106 1261 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VNB
rlabel comment 1244 3077 1244 3077 2 sky130_fd_sc_hd__buf_2_0/buf_2
rlabel metal1 1196 3077 1292 3445 7 sky130_fd_sc_hd__buf_2_0/VGND
rlabel metal1 652 3077 748 3445 7 sky130_fd_sc_hd__buf_2_0/VPWR
flabel metal1 683 3106 717 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VPWR
flabel metal1 139 3106 173 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VGND
flabel locali 683 3106 717 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VPWR
flabel locali 139 3106 173 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VGND
flabel locali 241 3289 275 3323 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/X
flabel locali 513 3289 547 3323 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/X
flabel locali 581 3289 615 3323 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/X
flabel locali 377 3106 411 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/A
flabel nwell 683 3106 717 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VPB
flabel pwell 139 3106 173 3140 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VNB
rlabel comment 156 3077 156 3077 8 sky130_fd_sc_hd__buf_2_1/buf_2
rlabel metal1 108 3077 204 3445 3 sky130_fd_sc_hd__buf_2_1/VGND
rlabel metal1 652 3077 748 3445 3 sky130_fd_sc_hd__buf_2_1/VPWR
flabel locali 377 3841 411 3875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/Y
flabel locali 445 3841 479 3875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/Y
flabel locali 377 3565 411 3599 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/A
flabel locali 377 3657 411 3691 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/A
flabel locali 377 3933 411 3967 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 377 4025 411 4059 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 377 4209 411 4243 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 377 4117 411 4151 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel nwell 683 4209 717 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VPB
flabel pwell 139 4209 173 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VNB
flabel metal1 139 4209 173 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VGND
flabel metal1 683 4209 717 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VPWR
rlabel comment 156 4273 156 4273 6 sky130_fd_sc_hd__nand2_4_0/nand2_4
rlabel metal1 108 3445 204 4273 3 sky130_fd_sc_hd__nand2_4_0/VGND
rlabel metal1 652 3445 748 4273 3 sky130_fd_sc_hd__nand2_4_0/VPWR
flabel locali 989 3841 1023 3875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/Y
flabel locali 921 3841 955 3875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/Y
flabel locali 989 3565 1023 3599 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/A
flabel locali 989 3657 1023 3691 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/A
flabel locali 989 3933 1023 3967 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 989 4025 1023 4059 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 989 4209 1023 4243 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 989 4117 1023 4151 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel nwell 683 4209 717 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VPB
flabel pwell 1227 4209 1261 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VNB
flabel metal1 1227 4209 1261 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VGND
flabel metal1 683 4209 717 4243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VPWR
rlabel comment 1244 4273 1244 4273 4 sky130_fd_sc_hd__nand2_4_1/nand2_4
rlabel metal1 1196 3445 1292 4273 7 sky130_fd_sc_hd__nand2_4_1/VGND
rlabel metal1 652 3445 748 4273 7 sky130_fd_sc_hd__nand2_4_1/VPWR
flabel metal1 139 4670 173 4704 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VGND
flabel metal1 683 4670 717 4704 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VPWR
flabel nwell 683 4670 717 4704 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VPB
flabel pwell 139 4670 173 4704 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VNB
rlabel comment 156 4733 156 4733 6 sky130_fd_sc_hd__decap_4_0/decap_4
rlabel metal1 108 4365 204 4733 3 sky130_fd_sc_hd__decap_4_0/VGND
rlabel metal1 652 4365 748 4733 3 sky130_fd_sc_hd__decap_4_0/VPWR
flabel metal1 1227 4394 1261 4428 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VGND
flabel metal1 683 4394 717 4428 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VPWR
flabel nwell 683 4394 717 4428 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VPB
flabel pwell 1227 4394 1261 4428 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VNB
rlabel comment 1244 4365 1244 4365 2 sky130_fd_sc_hd__decap_4_1/decap_4
rlabel metal1 1196 4365 1292 4733 7 sky130_fd_sc_hd__decap_4_1/VGND
rlabel metal1 652 4365 748 4733 7 sky130_fd_sc_hd__decap_4_1/VPWR
flabel metal1 680 4290 709 4343 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 138 4293 176 4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment 156 4365 156 4365 6 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
rlabel metal1 108 4273 204 4365 3 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel metal1 652 4273 748 4365 3 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 691 4295 720 4348 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 1224 4294 1262 4345 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment 1244 4273 1244 4273 2 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
rlabel metal1 1196 4273 1292 4365 7 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel metal1 652 4273 748 4365 7 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
<< end >>
