magic
tech sky130A
magscale 1 2
timestamp 1654124673
<< error_p >>
rect -1901 172 -1843 178
rect -1709 172 -1651 178
rect -1517 172 -1459 178
rect -1325 172 -1267 178
rect -1133 172 -1075 178
rect -941 172 -883 178
rect -749 172 -691 178
rect -557 172 -499 178
rect -365 172 -307 178
rect -173 172 -115 178
rect 19 172 77 178
rect 211 172 269 178
rect 403 172 461 178
rect 595 172 653 178
rect 787 172 845 178
rect 979 172 1037 178
rect 1171 172 1229 178
rect 1363 172 1421 178
rect 1555 172 1613 178
rect 1747 172 1805 178
rect 1939 172 1997 178
rect -1901 138 -1889 172
rect -1709 138 -1697 172
rect -1517 138 -1505 172
rect -1325 138 -1313 172
rect -1133 138 -1121 172
rect -941 138 -929 172
rect -749 138 -737 172
rect -557 138 -545 172
rect -365 138 -353 172
rect -173 138 -161 172
rect 19 138 31 172
rect 211 138 223 172
rect 403 138 415 172
rect 595 138 607 172
rect 787 138 799 172
rect 979 138 991 172
rect 1171 138 1183 172
rect 1363 138 1375 172
rect 1555 138 1567 172
rect 1747 138 1759 172
rect 1939 138 1951 172
rect -1901 132 -1843 138
rect -1709 132 -1651 138
rect -1517 132 -1459 138
rect -1325 132 -1267 138
rect -1133 132 -1075 138
rect -941 132 -883 138
rect -749 132 -691 138
rect -557 132 -499 138
rect -365 132 -307 138
rect -173 132 -115 138
rect 19 132 77 138
rect 211 132 269 138
rect 403 132 461 138
rect 595 132 653 138
rect 787 132 845 138
rect 979 132 1037 138
rect 1171 132 1229 138
rect 1363 132 1421 138
rect 1555 132 1613 138
rect 1747 132 1805 138
rect 1939 132 1997 138
rect -1997 -138 -1939 -132
rect -1805 -138 -1747 -132
rect -1613 -138 -1555 -132
rect -1421 -138 -1363 -132
rect -1229 -138 -1171 -132
rect -1037 -138 -979 -132
rect -845 -138 -787 -132
rect -653 -138 -595 -132
rect -461 -138 -403 -132
rect -269 -138 -211 -132
rect -77 -138 -19 -132
rect 115 -138 173 -132
rect 307 -138 365 -132
rect 499 -138 557 -132
rect 691 -138 749 -132
rect 883 -138 941 -132
rect 1075 -138 1133 -132
rect 1267 -138 1325 -132
rect 1459 -138 1517 -132
rect 1651 -138 1709 -132
rect 1843 -138 1901 -132
rect -1997 -172 -1985 -138
rect -1805 -172 -1793 -138
rect -1613 -172 -1601 -138
rect -1421 -172 -1409 -138
rect -1229 -172 -1217 -138
rect -1037 -172 -1025 -138
rect -845 -172 -833 -138
rect -653 -172 -641 -138
rect -461 -172 -449 -138
rect -269 -172 -257 -138
rect -77 -172 -65 -138
rect 115 -172 127 -138
rect 307 -172 319 -138
rect 499 -172 511 -138
rect 691 -172 703 -138
rect 883 -172 895 -138
rect 1075 -172 1087 -138
rect 1267 -172 1279 -138
rect 1459 -172 1471 -138
rect 1651 -172 1663 -138
rect 1843 -172 1855 -138
rect -1997 -178 -1939 -172
rect -1805 -178 -1747 -172
rect -1613 -178 -1555 -172
rect -1421 -178 -1363 -172
rect -1229 -178 -1171 -172
rect -1037 -178 -979 -172
rect -845 -178 -787 -172
rect -653 -178 -595 -172
rect -461 -178 -403 -172
rect -269 -178 -211 -172
rect -77 -178 -19 -172
rect 115 -178 173 -172
rect 307 -178 365 -172
rect 499 -178 557 -172
rect 691 -178 749 -172
rect 883 -178 941 -172
rect 1075 -178 1133 -172
rect 1267 -178 1325 -172
rect 1459 -178 1517 -172
rect 1651 -178 1709 -172
rect 1843 -178 1901 -172
<< nmos >>
rect -1983 -100 -1953 100
rect -1887 -100 -1857 100
rect -1791 -100 -1761 100
rect -1695 -100 -1665 100
rect -1599 -100 -1569 100
rect -1503 -100 -1473 100
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
rect 1473 -100 1503 100
rect 1569 -100 1599 100
rect 1665 -100 1695 100
rect 1761 -100 1791 100
rect 1857 -100 1887 100
rect 1953 -100 1983 100
<< ndiff >>
rect -2045 88 -1983 100
rect -2045 -88 -2033 88
rect -1999 -88 -1983 88
rect -2045 -100 -1983 -88
rect -1953 88 -1887 100
rect -1953 -88 -1937 88
rect -1903 -88 -1887 88
rect -1953 -100 -1887 -88
rect -1857 88 -1791 100
rect -1857 -88 -1841 88
rect -1807 -88 -1791 88
rect -1857 -100 -1791 -88
rect -1761 88 -1695 100
rect -1761 -88 -1745 88
rect -1711 -88 -1695 88
rect -1761 -100 -1695 -88
rect -1665 88 -1599 100
rect -1665 -88 -1649 88
rect -1615 -88 -1599 88
rect -1665 -100 -1599 -88
rect -1569 88 -1503 100
rect -1569 -88 -1553 88
rect -1519 -88 -1503 88
rect -1569 -100 -1503 -88
rect -1473 88 -1407 100
rect -1473 -88 -1457 88
rect -1423 -88 -1407 88
rect -1473 -100 -1407 -88
rect -1377 88 -1311 100
rect -1377 -88 -1361 88
rect -1327 -88 -1311 88
rect -1377 -100 -1311 -88
rect -1281 88 -1215 100
rect -1281 -88 -1265 88
rect -1231 -88 -1215 88
rect -1281 -100 -1215 -88
rect -1185 88 -1119 100
rect -1185 -88 -1169 88
rect -1135 -88 -1119 88
rect -1185 -100 -1119 -88
rect -1089 88 -1023 100
rect -1089 -88 -1073 88
rect -1039 -88 -1023 88
rect -1089 -100 -1023 -88
rect -993 88 -927 100
rect -993 -88 -977 88
rect -943 -88 -927 88
rect -993 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 993 100
rect 927 -88 943 88
rect 977 -88 993 88
rect 927 -100 993 -88
rect 1023 88 1089 100
rect 1023 -88 1039 88
rect 1073 -88 1089 88
rect 1023 -100 1089 -88
rect 1119 88 1185 100
rect 1119 -88 1135 88
rect 1169 -88 1185 88
rect 1119 -100 1185 -88
rect 1215 88 1281 100
rect 1215 -88 1231 88
rect 1265 -88 1281 88
rect 1215 -100 1281 -88
rect 1311 88 1377 100
rect 1311 -88 1327 88
rect 1361 -88 1377 88
rect 1311 -100 1377 -88
rect 1407 88 1473 100
rect 1407 -88 1423 88
rect 1457 -88 1473 88
rect 1407 -100 1473 -88
rect 1503 88 1569 100
rect 1503 -88 1519 88
rect 1553 -88 1569 88
rect 1503 -100 1569 -88
rect 1599 88 1665 100
rect 1599 -88 1615 88
rect 1649 -88 1665 88
rect 1599 -100 1665 -88
rect 1695 88 1761 100
rect 1695 -88 1711 88
rect 1745 -88 1761 88
rect 1695 -100 1761 -88
rect 1791 88 1857 100
rect 1791 -88 1807 88
rect 1841 -88 1857 88
rect 1791 -100 1857 -88
rect 1887 88 1953 100
rect 1887 -88 1903 88
rect 1937 -88 1953 88
rect 1887 -100 1953 -88
rect 1983 88 2045 100
rect 1983 -88 1999 88
rect 2033 -88 2045 88
rect 1983 -100 2045 -88
<< ndiffc >>
rect -2033 -88 -1999 88
rect -1937 -88 -1903 88
rect -1841 -88 -1807 88
rect -1745 -88 -1711 88
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
rect 1711 -88 1745 88
rect 1807 -88 1841 88
rect 1903 -88 1937 88
rect 1999 -88 2033 88
<< poly >>
rect -1905 172 -1839 188
rect -1905 138 -1889 172
rect -1855 138 -1839 172
rect -1983 100 -1953 126
rect -1905 122 -1839 138
rect -1713 172 -1647 188
rect -1713 138 -1697 172
rect -1663 138 -1647 172
rect -1887 100 -1857 122
rect -1791 100 -1761 126
rect -1713 122 -1647 138
rect -1521 172 -1455 188
rect -1521 138 -1505 172
rect -1471 138 -1455 172
rect -1695 100 -1665 122
rect -1599 100 -1569 126
rect -1521 122 -1455 138
rect -1329 172 -1263 188
rect -1329 138 -1313 172
rect -1279 138 -1263 172
rect -1503 100 -1473 122
rect -1407 100 -1377 126
rect -1329 122 -1263 138
rect -1137 172 -1071 188
rect -1137 138 -1121 172
rect -1087 138 -1071 172
rect -1311 100 -1281 122
rect -1215 100 -1185 126
rect -1137 122 -1071 138
rect -945 172 -879 188
rect -945 138 -929 172
rect -895 138 -879 172
rect -1119 100 -1089 122
rect -1023 100 -993 126
rect -945 122 -879 138
rect -753 172 -687 188
rect -753 138 -737 172
rect -703 138 -687 172
rect -927 100 -897 122
rect -831 100 -801 126
rect -753 122 -687 138
rect -561 172 -495 188
rect -561 138 -545 172
rect -511 138 -495 172
rect -735 100 -705 122
rect -639 100 -609 126
rect -561 122 -495 138
rect -369 172 -303 188
rect -369 138 -353 172
rect -319 138 -303 172
rect -543 100 -513 122
rect -447 100 -417 126
rect -369 122 -303 138
rect -177 172 -111 188
rect -177 138 -161 172
rect -127 138 -111 172
rect -351 100 -321 122
rect -255 100 -225 126
rect -177 122 -111 138
rect 15 172 81 188
rect 15 138 31 172
rect 65 138 81 172
rect -159 100 -129 122
rect -63 100 -33 126
rect 15 122 81 138
rect 207 172 273 188
rect 207 138 223 172
rect 257 138 273 172
rect 33 100 63 122
rect 129 100 159 126
rect 207 122 273 138
rect 399 172 465 188
rect 399 138 415 172
rect 449 138 465 172
rect 225 100 255 122
rect 321 100 351 126
rect 399 122 465 138
rect 591 172 657 188
rect 591 138 607 172
rect 641 138 657 172
rect 417 100 447 122
rect 513 100 543 126
rect 591 122 657 138
rect 783 172 849 188
rect 783 138 799 172
rect 833 138 849 172
rect 609 100 639 122
rect 705 100 735 126
rect 783 122 849 138
rect 975 172 1041 188
rect 975 138 991 172
rect 1025 138 1041 172
rect 801 100 831 122
rect 897 100 927 126
rect 975 122 1041 138
rect 1167 172 1233 188
rect 1167 138 1183 172
rect 1217 138 1233 172
rect 993 100 1023 122
rect 1089 100 1119 126
rect 1167 122 1233 138
rect 1359 172 1425 188
rect 1359 138 1375 172
rect 1409 138 1425 172
rect 1185 100 1215 122
rect 1281 100 1311 126
rect 1359 122 1425 138
rect 1551 172 1617 188
rect 1551 138 1567 172
rect 1601 138 1617 172
rect 1377 100 1407 122
rect 1473 100 1503 126
rect 1551 122 1617 138
rect 1743 172 1809 188
rect 1743 138 1759 172
rect 1793 138 1809 172
rect 1569 100 1599 122
rect 1665 100 1695 126
rect 1743 122 1809 138
rect 1935 172 2001 188
rect 1935 138 1951 172
rect 1985 138 2001 172
rect 1761 100 1791 122
rect 1857 100 1887 126
rect 1935 122 2001 138
rect 1953 100 1983 122
rect -1983 -122 -1953 -100
rect -2001 -138 -1935 -122
rect -1887 -126 -1857 -100
rect -1791 -122 -1761 -100
rect -2001 -172 -1985 -138
rect -1951 -172 -1935 -138
rect -2001 -188 -1935 -172
rect -1809 -138 -1743 -122
rect -1695 -126 -1665 -100
rect -1599 -122 -1569 -100
rect -1809 -172 -1793 -138
rect -1759 -172 -1743 -138
rect -1809 -188 -1743 -172
rect -1617 -138 -1551 -122
rect -1503 -126 -1473 -100
rect -1407 -122 -1377 -100
rect -1617 -172 -1601 -138
rect -1567 -172 -1551 -138
rect -1617 -188 -1551 -172
rect -1425 -138 -1359 -122
rect -1311 -126 -1281 -100
rect -1215 -122 -1185 -100
rect -1425 -172 -1409 -138
rect -1375 -172 -1359 -138
rect -1425 -188 -1359 -172
rect -1233 -138 -1167 -122
rect -1119 -126 -1089 -100
rect -1023 -122 -993 -100
rect -1233 -172 -1217 -138
rect -1183 -172 -1167 -138
rect -1233 -188 -1167 -172
rect -1041 -138 -975 -122
rect -927 -126 -897 -100
rect -831 -122 -801 -100
rect -1041 -172 -1025 -138
rect -991 -172 -975 -138
rect -1041 -188 -975 -172
rect -849 -138 -783 -122
rect -735 -126 -705 -100
rect -639 -122 -609 -100
rect -849 -172 -833 -138
rect -799 -172 -783 -138
rect -849 -188 -783 -172
rect -657 -138 -591 -122
rect -543 -126 -513 -100
rect -447 -122 -417 -100
rect -657 -172 -641 -138
rect -607 -172 -591 -138
rect -657 -188 -591 -172
rect -465 -138 -399 -122
rect -351 -126 -321 -100
rect -255 -122 -225 -100
rect -465 -172 -449 -138
rect -415 -172 -399 -138
rect -465 -188 -399 -172
rect -273 -138 -207 -122
rect -159 -126 -129 -100
rect -63 -122 -33 -100
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -273 -188 -207 -172
rect -81 -138 -15 -122
rect 33 -126 63 -100
rect 129 -122 159 -100
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect -81 -188 -15 -172
rect 111 -138 177 -122
rect 225 -126 255 -100
rect 321 -122 351 -100
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 111 -188 177 -172
rect 303 -138 369 -122
rect 417 -126 447 -100
rect 513 -122 543 -100
rect 303 -172 319 -138
rect 353 -172 369 -138
rect 303 -188 369 -172
rect 495 -138 561 -122
rect 609 -126 639 -100
rect 705 -122 735 -100
rect 495 -172 511 -138
rect 545 -172 561 -138
rect 495 -188 561 -172
rect 687 -138 753 -122
rect 801 -126 831 -100
rect 897 -122 927 -100
rect 687 -172 703 -138
rect 737 -172 753 -138
rect 687 -188 753 -172
rect 879 -138 945 -122
rect 993 -126 1023 -100
rect 1089 -122 1119 -100
rect 879 -172 895 -138
rect 929 -172 945 -138
rect 879 -188 945 -172
rect 1071 -138 1137 -122
rect 1185 -126 1215 -100
rect 1281 -122 1311 -100
rect 1071 -172 1087 -138
rect 1121 -172 1137 -138
rect 1071 -188 1137 -172
rect 1263 -138 1329 -122
rect 1377 -126 1407 -100
rect 1473 -122 1503 -100
rect 1263 -172 1279 -138
rect 1313 -172 1329 -138
rect 1263 -188 1329 -172
rect 1455 -138 1521 -122
rect 1569 -126 1599 -100
rect 1665 -122 1695 -100
rect 1455 -172 1471 -138
rect 1505 -172 1521 -138
rect 1455 -188 1521 -172
rect 1647 -138 1713 -122
rect 1761 -126 1791 -100
rect 1857 -122 1887 -100
rect 1647 -172 1663 -138
rect 1697 -172 1713 -138
rect 1647 -188 1713 -172
rect 1839 -138 1905 -122
rect 1953 -126 1983 -100
rect 1839 -172 1855 -138
rect 1889 -172 1905 -138
rect 1839 -188 1905 -172
<< polycont >>
rect -1889 138 -1855 172
rect -1697 138 -1663 172
rect -1505 138 -1471 172
rect -1313 138 -1279 172
rect -1121 138 -1087 172
rect -929 138 -895 172
rect -737 138 -703 172
rect -545 138 -511 172
rect -353 138 -319 172
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect 415 138 449 172
rect 607 138 641 172
rect 799 138 833 172
rect 991 138 1025 172
rect 1183 138 1217 172
rect 1375 138 1409 172
rect 1567 138 1601 172
rect 1759 138 1793 172
rect 1951 138 1985 172
rect -1985 -172 -1951 -138
rect -1793 -172 -1759 -138
rect -1601 -172 -1567 -138
rect -1409 -172 -1375 -138
rect -1217 -172 -1183 -138
rect -1025 -172 -991 -138
rect -833 -172 -799 -138
rect -641 -172 -607 -138
rect -449 -172 -415 -138
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
rect 319 -172 353 -138
rect 511 -172 545 -138
rect 703 -172 737 -138
rect 895 -172 929 -138
rect 1087 -172 1121 -138
rect 1279 -172 1313 -138
rect 1471 -172 1505 -138
rect 1663 -172 1697 -138
rect 1855 -172 1889 -138
<< locali >>
rect -1905 138 -1889 172
rect -1855 138 -1839 172
rect -1713 138 -1697 172
rect -1663 138 -1647 172
rect -1521 138 -1505 172
rect -1471 138 -1455 172
rect -1329 138 -1313 172
rect -1279 138 -1263 172
rect -1137 138 -1121 172
rect -1087 138 -1071 172
rect -945 138 -929 172
rect -895 138 -879 172
rect -753 138 -737 172
rect -703 138 -687 172
rect -561 138 -545 172
rect -511 138 -495 172
rect -369 138 -353 172
rect -319 138 -303 172
rect -177 138 -161 172
rect -127 138 -111 172
rect 15 138 31 172
rect 65 138 81 172
rect 207 138 223 172
rect 257 138 273 172
rect 399 138 415 172
rect 449 138 465 172
rect 591 138 607 172
rect 641 138 657 172
rect 783 138 799 172
rect 833 138 849 172
rect 975 138 991 172
rect 1025 138 1041 172
rect 1167 138 1183 172
rect 1217 138 1233 172
rect 1359 138 1375 172
rect 1409 138 1425 172
rect 1551 138 1567 172
rect 1601 138 1617 172
rect 1743 138 1759 172
rect 1793 138 1809 172
rect 1935 138 1951 172
rect 1985 138 2001 172
rect -2033 88 -1999 104
rect -2033 -104 -1999 -88
rect -1937 88 -1903 104
rect -1937 -104 -1903 -88
rect -1841 88 -1807 104
rect -1841 -104 -1807 -88
rect -1745 88 -1711 104
rect -1745 -104 -1711 -88
rect -1649 88 -1615 104
rect -1649 -104 -1615 -88
rect -1553 88 -1519 104
rect -1553 -104 -1519 -88
rect -1457 88 -1423 104
rect -1457 -104 -1423 -88
rect -1361 88 -1327 104
rect -1361 -104 -1327 -88
rect -1265 88 -1231 104
rect -1265 -104 -1231 -88
rect -1169 88 -1135 104
rect -1169 -104 -1135 -88
rect -1073 88 -1039 104
rect -1073 -104 -1039 -88
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect 1039 88 1073 104
rect 1039 -104 1073 -88
rect 1135 88 1169 104
rect 1135 -104 1169 -88
rect 1231 88 1265 104
rect 1231 -104 1265 -88
rect 1327 88 1361 104
rect 1327 -104 1361 -88
rect 1423 88 1457 104
rect 1423 -104 1457 -88
rect 1519 88 1553 104
rect 1519 -104 1553 -88
rect 1615 88 1649 104
rect 1615 -104 1649 -88
rect 1711 88 1745 104
rect 1711 -104 1745 -88
rect 1807 88 1841 104
rect 1807 -104 1841 -88
rect 1903 88 1937 104
rect 1903 -104 1937 -88
rect 1999 88 2033 104
rect 1999 -104 2033 -88
rect -2001 -172 -1985 -138
rect -1951 -172 -1935 -138
rect -1809 -172 -1793 -138
rect -1759 -172 -1743 -138
rect -1617 -172 -1601 -138
rect -1567 -172 -1551 -138
rect -1425 -172 -1409 -138
rect -1375 -172 -1359 -138
rect -1233 -172 -1217 -138
rect -1183 -172 -1167 -138
rect -1041 -172 -1025 -138
rect -991 -172 -975 -138
rect -849 -172 -833 -138
rect -799 -172 -783 -138
rect -657 -172 -641 -138
rect -607 -172 -591 -138
rect -465 -172 -449 -138
rect -415 -172 -399 -138
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 303 -172 319 -138
rect 353 -172 369 -138
rect 495 -172 511 -138
rect 545 -172 561 -138
rect 687 -172 703 -138
rect 737 -172 753 -138
rect 879 -172 895 -138
rect 929 -172 945 -138
rect 1071 -172 1087 -138
rect 1121 -172 1137 -138
rect 1263 -172 1279 -138
rect 1313 -172 1329 -138
rect 1455 -172 1471 -138
rect 1505 -172 1521 -138
rect 1647 -172 1663 -138
rect 1697 -172 1713 -138
rect 1839 -172 1855 -138
rect 1889 -172 1905 -138
<< viali >>
rect -1889 138 -1855 172
rect -1697 138 -1663 172
rect -1505 138 -1471 172
rect -1313 138 -1279 172
rect -1121 138 -1087 172
rect -929 138 -895 172
rect -737 138 -703 172
rect -545 138 -511 172
rect -353 138 -319 172
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect 415 138 449 172
rect 607 138 641 172
rect 799 138 833 172
rect 991 138 1025 172
rect 1183 138 1217 172
rect 1375 138 1409 172
rect 1567 138 1601 172
rect 1759 138 1793 172
rect 1951 138 1985 172
rect -2033 -88 -1999 88
rect -1937 -88 -1903 88
rect -1841 -88 -1807 88
rect -1745 -88 -1711 88
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
rect 1711 -88 1745 88
rect 1807 -88 1841 88
rect 1903 -88 1937 88
rect 1999 -88 2033 88
rect -1985 -172 -1951 -138
rect -1793 -172 -1759 -138
rect -1601 -172 -1567 -138
rect -1409 -172 -1375 -138
rect -1217 -172 -1183 -138
rect -1025 -172 -991 -138
rect -833 -172 -799 -138
rect -641 -172 -607 -138
rect -449 -172 -415 -138
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
rect 319 -172 353 -138
rect 511 -172 545 -138
rect 703 -172 737 -138
rect 895 -172 929 -138
rect 1087 -172 1121 -138
rect 1279 -172 1313 -138
rect 1471 -172 1505 -138
rect 1663 -172 1697 -138
rect 1855 -172 1889 -138
<< metal1 >>
rect -1901 172 -1843 178
rect -1901 138 -1889 172
rect -1855 138 -1843 172
rect -1901 132 -1843 138
rect -1709 172 -1651 178
rect -1709 138 -1697 172
rect -1663 138 -1651 172
rect -1709 132 -1651 138
rect -1517 172 -1459 178
rect -1517 138 -1505 172
rect -1471 138 -1459 172
rect -1517 132 -1459 138
rect -1325 172 -1267 178
rect -1325 138 -1313 172
rect -1279 138 -1267 172
rect -1325 132 -1267 138
rect -1133 172 -1075 178
rect -1133 138 -1121 172
rect -1087 138 -1075 172
rect -1133 132 -1075 138
rect -941 172 -883 178
rect -941 138 -929 172
rect -895 138 -883 172
rect -941 132 -883 138
rect -749 172 -691 178
rect -749 138 -737 172
rect -703 138 -691 172
rect -749 132 -691 138
rect -557 172 -499 178
rect -557 138 -545 172
rect -511 138 -499 172
rect -557 132 -499 138
rect -365 172 -307 178
rect -365 138 -353 172
rect -319 138 -307 172
rect -365 132 -307 138
rect -173 172 -115 178
rect -173 138 -161 172
rect -127 138 -115 172
rect -173 132 -115 138
rect 19 172 77 178
rect 19 138 31 172
rect 65 138 77 172
rect 19 132 77 138
rect 211 172 269 178
rect 211 138 223 172
rect 257 138 269 172
rect 211 132 269 138
rect 403 172 461 178
rect 403 138 415 172
rect 449 138 461 172
rect 403 132 461 138
rect 595 172 653 178
rect 595 138 607 172
rect 641 138 653 172
rect 595 132 653 138
rect 787 172 845 178
rect 787 138 799 172
rect 833 138 845 172
rect 787 132 845 138
rect 979 172 1037 178
rect 979 138 991 172
rect 1025 138 1037 172
rect 979 132 1037 138
rect 1171 172 1229 178
rect 1171 138 1183 172
rect 1217 138 1229 172
rect 1171 132 1229 138
rect 1363 172 1421 178
rect 1363 138 1375 172
rect 1409 138 1421 172
rect 1363 132 1421 138
rect 1555 172 1613 178
rect 1555 138 1567 172
rect 1601 138 1613 172
rect 1555 132 1613 138
rect 1747 172 1805 178
rect 1747 138 1759 172
rect 1793 138 1805 172
rect 1747 132 1805 138
rect 1939 172 1997 178
rect 1939 138 1951 172
rect 1985 138 1997 172
rect 1939 132 1997 138
rect -2039 88 -1993 100
rect -2039 -88 -2033 88
rect -1999 -88 -1993 88
rect -2039 -100 -1993 -88
rect -1943 88 -1897 100
rect -1943 -88 -1937 88
rect -1903 -88 -1897 88
rect -1943 -100 -1897 -88
rect -1847 88 -1801 100
rect -1847 -88 -1841 88
rect -1807 -88 -1801 88
rect -1847 -100 -1801 -88
rect -1751 88 -1705 100
rect -1751 -88 -1745 88
rect -1711 -88 -1705 88
rect -1751 -100 -1705 -88
rect -1655 88 -1609 100
rect -1655 -88 -1649 88
rect -1615 -88 -1609 88
rect -1655 -100 -1609 -88
rect -1559 88 -1513 100
rect -1559 -88 -1553 88
rect -1519 -88 -1513 88
rect -1559 -100 -1513 -88
rect -1463 88 -1417 100
rect -1463 -88 -1457 88
rect -1423 -88 -1417 88
rect -1463 -100 -1417 -88
rect -1367 88 -1321 100
rect -1367 -88 -1361 88
rect -1327 -88 -1321 88
rect -1367 -100 -1321 -88
rect -1271 88 -1225 100
rect -1271 -88 -1265 88
rect -1231 -88 -1225 88
rect -1271 -100 -1225 -88
rect -1175 88 -1129 100
rect -1175 -88 -1169 88
rect -1135 -88 -1129 88
rect -1175 -100 -1129 -88
rect -1079 88 -1033 100
rect -1079 -88 -1073 88
rect -1039 -88 -1033 88
rect -1079 -100 -1033 -88
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -887 88 -841 100
rect -887 -88 -881 88
rect -847 -88 -841 88
rect -887 -100 -841 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 841 88 887 100
rect 841 -88 847 88
rect 881 -88 887 88
rect 841 -100 887 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect 1033 88 1079 100
rect 1033 -88 1039 88
rect 1073 -88 1079 88
rect 1033 -100 1079 -88
rect 1129 88 1175 100
rect 1129 -88 1135 88
rect 1169 -88 1175 88
rect 1129 -100 1175 -88
rect 1225 88 1271 100
rect 1225 -88 1231 88
rect 1265 -88 1271 88
rect 1225 -100 1271 -88
rect 1321 88 1367 100
rect 1321 -88 1327 88
rect 1361 -88 1367 88
rect 1321 -100 1367 -88
rect 1417 88 1463 100
rect 1417 -88 1423 88
rect 1457 -88 1463 88
rect 1417 -100 1463 -88
rect 1513 88 1559 100
rect 1513 -88 1519 88
rect 1553 -88 1559 88
rect 1513 -100 1559 -88
rect 1609 88 1655 100
rect 1609 -88 1615 88
rect 1649 -88 1655 88
rect 1609 -100 1655 -88
rect 1705 88 1751 100
rect 1705 -88 1711 88
rect 1745 -88 1751 88
rect 1705 -100 1751 -88
rect 1801 88 1847 100
rect 1801 -88 1807 88
rect 1841 -88 1847 88
rect 1801 -100 1847 -88
rect 1897 88 1943 100
rect 1897 -88 1903 88
rect 1937 -88 1943 88
rect 1897 -100 1943 -88
rect 1993 88 2039 100
rect 1993 -88 1999 88
rect 2033 -88 2039 88
rect 1993 -100 2039 -88
rect -1997 -138 -1939 -132
rect -1997 -172 -1985 -138
rect -1951 -172 -1939 -138
rect -1997 -178 -1939 -172
rect -1805 -138 -1747 -132
rect -1805 -172 -1793 -138
rect -1759 -172 -1747 -138
rect -1805 -178 -1747 -172
rect -1613 -138 -1555 -132
rect -1613 -172 -1601 -138
rect -1567 -172 -1555 -138
rect -1613 -178 -1555 -172
rect -1421 -138 -1363 -132
rect -1421 -172 -1409 -138
rect -1375 -172 -1363 -138
rect -1421 -178 -1363 -172
rect -1229 -138 -1171 -132
rect -1229 -172 -1217 -138
rect -1183 -172 -1171 -138
rect -1229 -178 -1171 -172
rect -1037 -138 -979 -132
rect -1037 -172 -1025 -138
rect -991 -172 -979 -138
rect -1037 -178 -979 -172
rect -845 -138 -787 -132
rect -845 -172 -833 -138
rect -799 -172 -787 -138
rect -845 -178 -787 -172
rect -653 -138 -595 -132
rect -653 -172 -641 -138
rect -607 -172 -595 -138
rect -653 -178 -595 -172
rect -461 -138 -403 -132
rect -461 -172 -449 -138
rect -415 -172 -403 -138
rect -461 -178 -403 -172
rect -269 -138 -211 -132
rect -269 -172 -257 -138
rect -223 -172 -211 -138
rect -269 -178 -211 -172
rect -77 -138 -19 -132
rect -77 -172 -65 -138
rect -31 -172 -19 -138
rect -77 -178 -19 -172
rect 115 -138 173 -132
rect 115 -172 127 -138
rect 161 -172 173 -138
rect 115 -178 173 -172
rect 307 -138 365 -132
rect 307 -172 319 -138
rect 353 -172 365 -138
rect 307 -178 365 -172
rect 499 -138 557 -132
rect 499 -172 511 -138
rect 545 -172 557 -138
rect 499 -178 557 -172
rect 691 -138 749 -132
rect 691 -172 703 -138
rect 737 -172 749 -138
rect 691 -178 749 -172
rect 883 -138 941 -132
rect 883 -172 895 -138
rect 929 -172 941 -138
rect 883 -178 941 -172
rect 1075 -138 1133 -132
rect 1075 -172 1087 -138
rect 1121 -172 1133 -138
rect 1075 -178 1133 -172
rect 1267 -138 1325 -132
rect 1267 -172 1279 -138
rect 1313 -172 1325 -138
rect 1267 -178 1325 -172
rect 1459 -138 1517 -132
rect 1459 -172 1471 -138
rect 1505 -172 1517 -138
rect 1459 -178 1517 -172
rect 1651 -138 1709 -132
rect 1651 -172 1663 -138
rect 1697 -172 1709 -138
rect 1651 -178 1709 -172
rect 1843 -138 1901 -132
rect 1843 -172 1855 -138
rect 1889 -172 1901 -138
rect 1843 -178 1901 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 42 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
