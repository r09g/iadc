magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -77 138 -19 144
rect 19 138 77 144
rect -77 104 -65 138
rect 19 104 31 138
rect -77 98 -19 104
rect 19 98 77 104
rect -77 -102 -19 -96
rect 19 -102 77 -96
rect -77 -136 -65 -102
rect 19 -136 31 -102
rect -77 -142 -19 -136
rect 19 -142 77 -136
<< pwell >>
rect -301 -264 301 266
<< nmos >>
rect -111 -64 -81 66
rect -15 -64 15 66
rect 81 -64 111 66
<< ndiff >>
rect -173 52 -111 66
rect -173 18 -161 52
rect -127 18 -111 52
rect -173 -16 -111 18
rect -173 -50 -161 -16
rect -127 -50 -111 -16
rect -173 -64 -111 -50
rect -81 52 -15 66
rect -81 18 -65 52
rect -31 18 -15 52
rect -81 -16 -15 18
rect -81 -50 -65 -16
rect -31 -50 -15 -16
rect -81 -64 -15 -50
rect 15 52 81 66
rect 15 18 31 52
rect 65 18 81 52
rect 15 -16 81 18
rect 15 -50 31 -16
rect 65 -50 81 -16
rect 15 -64 81 -50
rect 111 52 173 66
rect 111 18 127 52
rect 161 18 173 52
rect 111 -16 173 18
rect 111 -50 127 -16
rect 161 -50 173 -16
rect 111 -64 173 -50
<< ndiffc >>
rect -161 18 -127 52
rect -161 -50 -127 -16
rect -65 18 -31 52
rect -65 -50 -31 -16
rect 31 18 65 52
rect 31 -50 65 -16
rect 127 18 161 52
rect 127 -50 161 -16
<< psubdiff >>
rect -275 206 -153 240
rect -119 206 -85 240
rect -51 206 -17 240
rect 17 206 51 240
rect 85 206 119 240
rect 153 206 275 240
rect -275 120 -241 206
rect 241 120 275 206
rect -275 52 -241 86
rect -275 -16 -241 18
rect -275 -84 -241 -50
rect 241 52 275 86
rect 241 -16 275 18
rect 241 -84 275 -50
rect -275 -204 -241 -118
rect 241 -204 275 -118
rect -275 -238 -153 -204
rect -119 -238 -85 -204
rect -51 -238 -17 -204
rect 17 -238 51 -204
rect 85 -238 119 -204
rect 153 -238 275 -204
<< psubdiffcont >>
rect -153 206 -119 240
rect -85 206 -51 240
rect -17 206 17 240
rect 51 206 85 240
rect 119 206 153 240
rect -275 86 -241 120
rect 241 86 275 120
rect -275 18 -241 52
rect -275 -50 -241 -16
rect 241 18 275 52
rect 241 -50 275 -16
rect -275 -118 -241 -84
rect 241 -118 275 -84
rect -153 -238 -119 -204
rect -85 -238 -51 -204
rect -17 -238 17 -204
rect 51 -238 85 -204
rect 119 -238 153 -204
<< poly >>
rect -129 138 129 154
rect -129 104 -65 138
rect -31 104 31 138
rect 65 104 129 138
rect -129 88 129 104
rect -111 66 -81 88
rect -15 66 15 88
rect 81 66 111 88
rect -111 -86 -81 -64
rect -15 -86 15 -64
rect 81 -86 111 -64
rect -129 -102 129 -86
rect -129 -136 -65 -102
rect -31 -136 31 -102
rect 65 -136 129 -102
rect -129 -152 129 -136
<< polycont >>
rect -65 104 -31 138
rect 31 104 65 138
rect -65 -136 -31 -102
rect 31 -136 65 -102
<< locali >>
rect -275 206 -153 240
rect -119 206 -85 240
rect -51 206 -17 240
rect 17 206 51 240
rect 85 206 119 240
rect 153 206 275 240
rect -275 120 -241 206
rect -81 104 -65 138
rect -31 104 31 138
rect 65 104 81 138
rect 241 120 275 206
rect -275 52 -241 86
rect -275 -16 -241 18
rect -275 -84 -241 -50
rect -161 54 -127 70
rect -161 -16 -127 18
rect -161 -68 -127 -52
rect -65 54 -31 70
rect -65 -16 -31 18
rect -65 -68 -31 -52
rect 31 54 65 70
rect 31 -16 65 18
rect 31 -68 65 -52
rect 127 54 161 70
rect 127 -16 161 18
rect 127 -68 161 -52
rect 241 52 275 86
rect 241 -16 275 18
rect 241 -84 275 -50
rect -275 -204 -241 -118
rect -81 -136 -65 -102
rect -31 -136 31 -102
rect 65 -136 81 -102
rect 241 -204 275 -118
rect -275 -238 -153 -204
rect -119 -238 -85 -204
rect -51 -238 -17 -204
rect 17 -238 51 -204
rect 85 -238 119 -204
rect 153 -238 275 -204
<< viali >>
rect -65 104 -31 138
rect 31 104 65 138
rect -161 52 -127 54
rect -161 20 -127 52
rect -161 -50 -127 -18
rect -161 -52 -127 -50
rect -65 52 -31 54
rect -65 20 -31 52
rect -65 -50 -31 -18
rect -65 -52 -31 -50
rect 31 52 65 54
rect 31 20 65 52
rect 31 -50 65 -18
rect 31 -52 65 -50
rect 127 52 161 54
rect 127 20 161 52
rect 127 -50 161 -18
rect 127 -52 161 -50
rect -65 -136 -31 -102
rect 31 -136 65 -102
<< metal1 >>
rect -77 138 -19 144
rect -77 104 -65 138
rect -31 104 -19 138
rect -77 98 -19 104
rect 19 138 77 144
rect 19 104 31 138
rect 65 104 77 138
rect 19 98 77 104
rect -167 54 -121 66
rect -167 20 -161 54
rect -127 20 -121 54
rect -167 18 -121 20
rect -71 54 -25 66
rect -71 20 -65 54
rect -31 20 -25 54
rect -71 18 -25 20
rect 25 54 71 66
rect 25 20 31 54
rect 65 20 71 54
rect 25 18 71 20
rect 121 54 167 66
rect 121 20 127 54
rect 161 20 167 54
rect 121 18 167 20
rect -277 -18 277 18
rect -167 -52 -161 -18
rect -127 -52 -121 -18
rect -167 -64 -121 -52
rect -71 -52 -65 -18
rect -31 -52 -25 -18
rect -71 -64 -25 -52
rect 25 -52 31 -18
rect 65 -52 71 -18
rect 25 -64 71 -52
rect 121 -52 127 -18
rect 161 -52 167 -18
rect 121 -64 167 -52
rect -77 -102 -19 -96
rect -77 -136 -65 -102
rect -31 -136 -19 -102
rect -77 -142 -19 -136
rect 19 -102 77 -96
rect 19 -136 31 -102
rect 65 -136 77 -102
rect 19 -142 77 -136
<< properties >>
string FIXED_BBOX -258 -222 258 222
<< end >>
