magic
tech sky130A
magscale 1 2
timestamp 1653453365
<< pwell >>
rect -647 -263 647 201
<< nmos >>
rect -447 -53 -417 53
rect -351 -53 -321 53
rect -255 -53 -225 53
rect -159 -53 -129 53
rect -63 -53 -33 53
rect 33 -53 63 53
rect 129 -53 159 53
rect 225 -53 255 53
rect 321 -53 351 53
rect 417 -53 447 53
<< ndiff >>
rect -509 41 -447 53
rect -509 -41 -497 41
rect -463 -41 -447 41
rect -509 -53 -447 -41
rect -417 41 -351 53
rect -417 -41 -401 41
rect -367 -41 -351 41
rect -417 -53 -351 -41
rect -321 41 -255 53
rect -321 -41 -305 41
rect -271 -41 -255 41
rect -321 -53 -255 -41
rect -225 41 -159 53
rect -225 -41 -209 41
rect -175 -41 -159 41
rect -225 -53 -159 -41
rect -129 41 -63 53
rect -129 -41 -113 41
rect -79 -41 -63 41
rect -129 -53 -63 -41
rect -33 41 33 53
rect -33 -41 -17 41
rect 17 -41 33 41
rect -33 -53 33 -41
rect 63 41 129 53
rect 63 -41 79 41
rect 113 -41 129 41
rect 63 -53 129 -41
rect 159 41 225 53
rect 159 -41 175 41
rect 209 -41 225 41
rect 159 -53 225 -41
rect 255 41 321 53
rect 255 -41 271 41
rect 305 -41 321 41
rect 255 -53 321 -41
rect 351 41 417 53
rect 351 -41 367 41
rect 401 -41 417 41
rect 351 -53 417 -41
rect 447 41 509 53
rect 447 -41 463 41
rect 497 -41 509 41
rect 447 -53 509 -41
<< ndiffc >>
rect -497 -41 -463 41
rect -401 -41 -367 41
rect -305 -41 -271 41
rect -209 -41 -175 41
rect -113 -41 -79 41
rect -17 -41 17 41
rect 79 -41 113 41
rect 175 -41 209 41
rect 271 -41 305 41
rect 367 -41 401 41
rect 463 -41 497 41
<< psubdiff >>
rect -611 131 -515 165
rect 515 131 611 165
rect -611 69 -577 131
rect 577 69 611 131
rect -611 -193 -577 -131
rect 577 -193 611 -131
rect -611 -227 -515 -193
rect 515 -227 611 -193
<< psubdiffcont >>
rect -515 131 515 165
rect -611 -131 -577 69
rect 577 -131 611 69
rect -515 -227 515 -193
<< poly >>
rect -447 53 -417 79
rect -351 53 -321 79
rect -255 53 -225 79
rect -159 53 -129 79
rect -63 53 -33 79
rect 33 53 63 79
rect 129 53 159 79
rect 225 53 255 79
rect 321 53 351 79
rect 417 53 447 79
rect -447 -75 -417 -53
rect -351 -75 -321 -53
rect -255 -75 -225 -53
rect -159 -75 -129 -53
rect -63 -75 -33 -53
rect 33 -75 63 -53
rect 129 -75 159 -53
rect 225 -75 255 -53
rect 321 -75 351 -53
rect 417 -75 447 -53
rect -513 -94 513 -75
rect -513 -128 -497 -94
rect -463 -128 -305 -94
rect -271 -128 -113 -94
rect -79 -128 79 -94
rect 113 -128 271 -94
rect 305 -128 463 -94
rect 497 -128 513 -94
rect -513 -141 513 -128
<< polycont >>
rect -497 -128 -463 -94
rect -305 -128 -271 -94
rect -113 -128 -79 -94
rect 79 -128 113 -94
rect 271 -128 305 -94
rect 463 -128 497 -94
<< locali >>
rect -611 131 -515 165
rect 515 131 611 165
rect -611 69 -577 131
rect 577 69 611 131
rect -497 41 -463 57
rect -497 -57 -463 -41
rect -401 41 -367 57
rect -401 -57 -367 -41
rect -305 41 -271 57
rect -305 -57 -271 -41
rect -209 41 -175 57
rect -209 -57 -175 -41
rect -113 41 -79 57
rect -113 -57 -79 -41
rect -17 41 17 57
rect -17 -57 17 -41
rect 79 41 113 57
rect 79 -57 113 -41
rect 175 41 209 57
rect 175 -57 209 -41
rect 271 41 305 57
rect 271 -57 305 -41
rect 367 41 401 57
rect 367 -57 401 -41
rect 463 41 497 57
rect 463 -57 497 -41
rect -513 -128 -497 -94
rect -463 -128 -447 -94
rect -321 -128 -305 -94
rect -271 -128 -255 -94
rect -129 -128 -113 -94
rect -79 -128 -63 -94
rect 63 -128 79 -94
rect 113 -128 129 -94
rect 255 -128 271 -94
rect 305 -128 321 -94
rect 447 -128 463 -94
rect 497 -128 513 -94
rect -611 -193 -577 -131
rect 577 -193 611 -131
rect -611 -227 -515 -193
rect 515 -227 611 -193
<< viali >>
rect -497 -41 -463 41
rect -401 -41 -367 41
rect -305 -41 -271 41
rect -209 -41 -175 41
rect -113 -41 -79 41
rect -17 -41 17 41
rect 79 -41 113 41
rect 175 -41 209 41
rect 271 -41 305 41
rect 367 -41 401 41
rect 463 -41 497 41
rect -497 -128 -463 -94
rect -305 -128 -271 -94
rect -113 -128 -79 -94
rect 79 -128 113 -94
rect 271 -128 305 -94
rect 463 -128 497 -94
<< metal1 >>
rect -503 41 -457 53
rect -503 -41 -497 41
rect -463 -41 -457 41
rect -503 -53 -457 -41
rect -407 41 -361 53
rect -407 -41 -401 41
rect -367 -41 -361 41
rect -407 -53 -361 -41
rect -311 41 -265 53
rect -311 -41 -305 41
rect -271 -41 -265 41
rect -311 -53 -265 -41
rect -215 41 -169 53
rect -215 -41 -209 41
rect -175 -41 -169 41
rect -215 -53 -169 -41
rect -119 41 -73 53
rect -119 -41 -113 41
rect -79 -41 -73 41
rect -119 -53 -73 -41
rect -23 41 23 53
rect -23 -41 -17 41
rect 17 -41 23 41
rect -23 -53 23 -41
rect 73 41 119 53
rect 73 -41 79 41
rect 113 -41 119 41
rect 73 -53 119 -41
rect 169 41 215 53
rect 169 -41 175 41
rect 209 -41 215 41
rect 169 -53 215 -41
rect 265 41 311 53
rect 265 -41 271 41
rect 305 -41 311 41
rect 265 -53 311 -41
rect 361 41 407 53
rect 361 -41 367 41
rect 401 -41 407 41
rect 361 -53 407 -41
rect 457 41 503 53
rect 457 -41 463 41
rect 497 -41 503 41
rect 457 -53 503 -41
rect -513 -94 -447 -81
rect -513 -128 -497 -94
rect -463 -128 -447 -94
rect -513 -141 -447 -128
rect -321 -94 -255 -81
rect -321 -128 -305 -94
rect -271 -128 -255 -94
rect -321 -141 -255 -128
rect -129 -94 -63 -81
rect -129 -128 -113 -94
rect -79 -128 -63 -94
rect -129 -141 -63 -128
rect 63 -94 129 -81
rect 63 -128 79 -94
rect 113 -128 129 -94
rect 63 -141 129 -128
rect 255 -94 321 -81
rect 255 -128 271 -94
rect 305 -128 321 -94
rect 255 -141 321 -128
rect 447 -94 513 -81
rect 447 -128 463 -94
rect 497 -128 513 -94
rect 447 -141 513 -128
<< properties >>
string FIXED_BBOX -594 -210 594 210
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.53 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
