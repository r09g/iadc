* NGSPICE file created from comparator_flat.ext - technology: sky130A

.subckt comparator_flat clk ip in outp outn VDD VSS
X0 VSS outp a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=4.2359e+12p pd=4.436e+07u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1 VDD sky130_fd_sc_hd__nand2_4_1/A outn VDD sky130_fd_pr__pfet_01v8_hvt ad=6.2558e+12p pd=6.098e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X2 VDD a_177_3251# sky130_fd_sc_hd__nand2_4_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 outn sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=6.375e+11p pd=6.55e+06u as=0p ps=0u w=500000u l=150000u
X5 VDD clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.4e+11p ps=6.56e+06u w=500000u l=150000u
X6 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=3.24e+06u as=8.05e+11p ps=8.22e+06u w=500000u l=150000u
X7 a_282_408# in a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=1.5015e+12p pd=1.504e+07u as=8.05e+11p ps=8.22e+06u w=500000u l=150000u
X8 VSS outp a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VDD sky130_fd_sc_hd__buf_2_0/A a_721_3251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X12 a_1067_3524# sky130_fd_sc_hd__nand2_4_1/A outn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X13 outp sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X14 VSS a_177_3251# sky130_fd_sc_hd__nand2_4_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X16 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=3.24e+06u as=0p ps=0u w=500000u l=150000u
X17 VDD outp outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 outn outp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 outp sky130_fd_sc_hd__nand2_4_0/A a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X20 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X21 outn outp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VDD sky130_fd_sc_hd__buf_2_1/A a_177_3251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X24 a_475_1219# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X25 VDD outn outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VDD sky130_fd_sc_hd__nand2_4_1/A outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VSS a_721_3251# sky130_fd_sc_hd__nand2_4_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X28 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X30 a_282_408# ip a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X31 a_282_408# ip a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X32 a_n16_2554# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X33 a_475_1219# in a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X34 a_282_408# in a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X35 VSS VSS a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X36 a_203_3524# outn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X38 a_n16_2554# ip a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X39 outn sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 VDD sky130_fd_sc_hd__nand2_4_0/A outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X42 VSS sky130_fd_sc_hd__buf_2_1/A a_177_3251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X43 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X44 outp sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 sky130_fd_sc_hd__buf_2_1/A clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X46 sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X47 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X48 VDD a_721_3251# sky130_fd_sc_hd__nand2_4_1/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X49 VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X50 a_203_3524# sky130_fd_sc_hd__nand2_4_0/A outp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X51 VDD clk a_n16_2554# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
X52 a_475_1219# clk VDD VDD sky130_fd_pr__pfet_01v8 ad=1.425e+11p pd=1.57e+06u as=0p ps=0u w=500000u l=150000u
X53 a_n16_2554# ip a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X54 outp sky130_fd_sc_hd__nand2_4_0/A a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X55 a_1067_3524# outp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X56 outp outn VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 VDD outn outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 outn sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X60 VSS VSS a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X61 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X62 a_n16_2554# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X63 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X64 outp outn VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 VSS outn a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X66 a_203_3524# outn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X67 VDD sky130_fd_sc_hd__nand2_4_0/A outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_1067_3524# sky130_fd_sc_hd__nand2_4_1/A outn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X69 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X70 VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X71 outn sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X72 a_282_408# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X73 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X74 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X75 VDD outp outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 VSS outn a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X77 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 VDD VDD sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X79 a_475_1219# in a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X80 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X81 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X82 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X83 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X84 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X85 a_203_3524# sky130_fd_sc_hd__nand2_4_0/A outp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X86 a_475_1219# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X87 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X88 a_1067_3524# outp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X89 VSS sky130_fd_sc_hd__buf_2_0/A a_721_3251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X90 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X91 VSS VSS a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
C0 outp a_203_3524# 0.60fF
C1 sky130_fd_sc_hd__buf_2_1/A a_177_3251# 0.26fF
C2 a_177_3251# a_721_3251# 0.06fF
C3 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_1/A 0.10fF
C4 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__buf_2_0/A 0.07fF
C5 a_475_1219# a_177_3251# 0.00fF
C6 outp sky130_fd_sc_hd__nand2_4_1/A 0.19fF
C7 outn a_177_3251# 0.02fF
C8 sky130_fd_sc_hd__nand2_4_0/A a_1067_3524# 0.01fF
C9 outp a_1067_3524# 0.39fF
C10 a_177_3251# a_n16_2554# 0.00fF
C11 VDD sky130_fd_sc_hd__buf_2_1/A 3.64fF
C12 VDD a_721_3251# 0.48fF
C13 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# 0.32fF
C14 a_177_3251# sky130_fd_sc_hd__buf_2_0/A 0.02fF
C15 VDD a_475_1219# 0.30fF
C16 VDD ip 0.04fF
C17 sky130_fd_sc_hd__buf_2_1/A a_721_3251# 0.02fF
C18 outp a_177_3251# 0.04fF
C19 VDD outn 2.38fF
C20 sky130_fd_sc_hd__buf_2_1/A a_475_1219# 0.65fF
C21 a_475_1219# a_721_3251# 0.00fF
C22 sky130_fd_sc_hd__buf_2_1/A ip 0.22fF
C23 sky130_fd_sc_hd__buf_2_1/A outn 0.05fF
C24 outn a_721_3251# 0.04fF
C25 ip a_475_1219# 0.29fF
C26 VDD a_n16_2554# 0.44fF
C27 VDD sky130_fd_sc_hd__nand2_4_0/A 0.81fF
C28 sky130_fd_sc_hd__buf_2_1/A a_n16_2554# 1.44fF
C29 VDD sky130_fd_sc_hd__buf_2_0/A 3.75fF
C30 a_721_3251# a_n16_2554# 0.00fF
C31 VDD clk 0.56fF
C32 VDD outp 2.35fF
C33 in VDD 0.04fF
C34 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__nand2_4_0/A 0.07fF
C35 a_475_1219# a_n16_2554# 1.23fF
C36 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A 5.69fF
C37 ip a_n16_2554# 0.97fF
C38 a_721_3251# sky130_fd_sc_hd__buf_2_0/A 0.26fF
C39 sky130_fd_sc_hd__nand2_4_0/A a_475_1219# 0.00fF
C40 clk sky130_fd_sc_hd__buf_2_1/A 0.05fF
C41 outp sky130_fd_sc_hd__buf_2_1/A 0.05fF
C42 outp a_721_3251# 0.02fF
C43 in sky130_fd_sc_hd__buf_2_1/A 0.15fF
C44 a_475_1219# sky130_fd_sc_hd__buf_2_0/A 1.33fF
C45 ip sky130_fd_sc_hd__buf_2_0/A 0.17fF
C46 sky130_fd_sc_hd__nand2_4_0/A outn 0.19fF
C47 clk a_475_1219# 0.13fF
C48 in a_475_1219# 1.03fF
C49 outn sky130_fd_sc_hd__buf_2_0/A 0.04fF
C50 clk ip 0.09fF
C51 in ip 0.93fF
C52 outp outn 1.74fF
C53 a_203_3524# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C54 sky130_fd_sc_hd__nand2_4_0/A a_n16_2554# 0.00fF
C55 sky130_fd_sc_hd__buf_2_0/A a_n16_2554# 0.91fF
C56 clk a_n16_2554# 0.15fF
C57 in a_n16_2554# 0.32fF
C58 a_203_3524# a_1067_3524# 0.03fF
C59 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__buf_2_0/A 0.02fF
C60 outp sky130_fd_sc_hd__nand2_4_0/A 0.56fF
C61 clk sky130_fd_sc_hd__buf_2_0/A 0.04fF
C62 outp sky130_fd_sc_hd__buf_2_0/A 0.05fF
C63 in sky130_fd_sc_hd__buf_2_0/A 0.21fF
C64 sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# 0.14fF
C65 in clk 0.07fF
C66 a_203_3524# a_177_3251# 0.02fF
C67 VDD a_282_408# 0.02fF
C68 sky130_fd_sc_hd__buf_2_1/A a_282_408# 0.09fF
C69 a_282_408# a_475_1219# 0.73fF
C70 ip a_282_408# 0.24fF
C71 VDD a_203_3524# 0.08fF
C72 a_282_408# a_n16_2554# 0.71fF
C73 VDD sky130_fd_sc_hd__nand2_4_1/A 0.76fF
C74 a_282_408# sky130_fd_sc_hd__buf_2_0/A 0.09fF
C75 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C76 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# 0.32fF
C77 outn a_203_3524# 0.41fF
C78 clk a_282_408# 0.48fF
C79 VDD a_1067_3524# 0.08fF
C80 in a_282_408# 0.28fF
C81 a_475_1219# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C82 outn sky130_fd_sc_hd__nand2_4_1/A 0.54fF
C83 a_721_3251# a_1067_3524# 0.02fF
C84 outn a_1067_3524# 0.52fF
C85 sky130_fd_sc_hd__nand2_4_0/A a_203_3524# 0.16fF
C86 VDD a_177_3251# 0.50fF
C87 sky130_fd_sc_hd__nand2_4_1/A a_n16_2554# 0.00fF
C88 clk VSS 2.24fF
C89 in VSS 1.70fF
C90 ip VSS 1.89fF
C91 a_282_408# VSS 1.97fF
C92 a_475_1219# VSS 1.53fF
C93 a_n16_2554# VSS 1.70fF
C94 sky130_fd_sc_hd__buf_2_0/A VSS 2.01fF
C95 sky130_fd_sc_hd__buf_2_1/A VSS 1.88fF
C96 a_721_3251# VSS 0.41fF
C97 a_177_3251# VSS 0.44fF
C98 sky130_fd_sc_hd__nand2_4_1/A VSS 0.69fF
C99 sky130_fd_sc_hd__nand2_4_0/A VSS 0.71fF
C100 a_1067_3524# VSS 1.03fF
C101 outp VSS 1.55fF
C102 outn VSS 1.51fF
C103 a_203_3524# VSS 1.11fF
C104 VDD VSS 11.21fF
.ends

