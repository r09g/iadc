* NGSPICE file created from ota_w_test_v2.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_YVTR7C a_n207_n140# a_n1039_n205# a_29_n205# a_327_n140#
+ a_n683_n205# a_n1275_n140# a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_1097_n205#
+ a_n505_n205# a_n741_n140# a_563_n205# a_861_n140# w_n1311_n241# a_919_n205# a_n327_n205#
+ a_n563_n140# a_385_n205# a_683_n140# a_n919_n140# a_n149_n205# a_1039_n140# a_n385_n140#
+ a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_327_n140# a_207_n205# a_149_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_149_n140# a_29_n205# a_n29_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_861_n140# a_741_n205# a_683_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_n140# a_n327_n205# a_n385_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1097_n205# a_1097_n205# a_1039_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n741_n140# a_n861_n205# a_n919_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n1097_n140# a_n1275_n140# a_n1275_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_683_n140# a_563_n205# a_505_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1039_n140# a_919_n205# a_861_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n29_n140# a_n149_n205# a_n207_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n563_n140# a_n683_n205# a_n741_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1275_n140# a_n1039_n205# 0.07fF
C1 a_207_n205# a_n861_n205# 0.01fF
C2 w_n1311_n241# a_n1039_n205# 0.20fF
C3 a_n149_n205# a_29_n205# 0.10fF
C4 a_n1039_n205# a_n861_n205# 0.10fF
C5 a_n327_n205# a_n149_n205# 0.10fF
C6 a_861_n140# a_505_n140# 0.03fF
C7 w_n1311_n241# a_741_n205# 0.15fF
C8 a_n683_n205# a_n149_n205# 0.02fF
C9 a_n861_n205# a_741_n205# 0.01fF
C10 a_861_n140# a_149_n140# 0.01fF
C11 a_n505_n205# a_1097_n205# 0.00fF
C12 a_861_n140# a_1039_n140# 0.06fF
C13 a_563_n205# a_n149_n205# 0.01fF
C14 a_505_n140# a_n919_n140# 0.01fF
C15 a_149_n140# a_n919_n140# 0.01fF
C16 a_n505_n205# a_385_n205# 0.01fF
C17 a_861_n140# a_n563_n140# 0.01fF
C18 a_n149_n205# a_207_n205# 0.03fF
C19 a_149_n140# a_505_n140# 0.03fF
C20 a_1039_n140# a_505_n140# 0.02fF
C21 a_861_n140# a_683_n140# 0.06fF
C22 w_n1311_n241# a_919_n205# 0.14fF
C23 a_861_n140# a_n29_n140# 0.01fF
C24 a_861_n140# a_1097_n205# 0.03fF
C25 a_n149_n205# a_n1039_n205# 0.01fF
C26 a_n505_n205# a_29_n205# 0.02fF
C27 a_1039_n140# a_149_n140# 0.01fF
C28 a_861_n140# a_327_n140# 0.02fF
C29 a_n563_n140# a_n919_n140# 0.03fF
C30 a_n505_n205# a_n327_n205# 0.10fF
C31 a_n683_n205# a_n505_n205# 0.10fF
C32 a_683_n140# a_n919_n140# 0.01fF
C33 a_n149_n205# a_741_n205# 0.01fF
C34 a_n563_n140# a_505_n140# 0.01fF
C35 a_n29_n140# a_n919_n140# 0.01fF
C36 a_n207_n140# a_n741_n140# 0.02fF
C37 a_505_n140# a_683_n140# 0.06fF
C38 a_327_n140# a_n919_n140# 0.01fF
C39 a_n505_n205# a_563_n205# 0.01fF
C40 a_505_n140# a_n29_n140# 0.02fF
C41 a_n563_n140# a_149_n140# 0.01fF
C42 a_1039_n140# a_n563_n140# 0.01fF
C43 a_1097_n205# a_505_n140# 0.01fF
C44 a_n1275_n140# a_n741_n140# 0.02fF
C45 a_149_n140# a_683_n140# 0.02fF
C46 a_327_n140# a_505_n140# 0.06fF
C47 a_149_n140# a_n29_n140# 0.06fF
C48 a_1039_n140# a_683_n140# 0.03fF
C49 w_n1311_n241# a_n741_n140# 0.02fF
C50 a_n385_n140# a_n741_n140# 0.03fF
C51 a_1097_n205# a_149_n140# 0.01fF
C52 a_1039_n140# a_n29_n140# 0.01fF
C53 a_1039_n140# a_1097_n205# 0.06fF
C54 a_149_n140# a_327_n140# 0.06fF
C55 a_n505_n205# a_207_n205# 0.01fF
C56 a_1039_n140# a_327_n140# 0.01fF
C57 a_n1097_n140# a_n741_n140# 0.03fF
C58 a_n1275_n140# a_n207_n140# 0.01fF
C59 a_n149_n205# a_919_n205# 0.01fF
C60 a_n505_n205# a_n1039_n205# 0.02fF
C61 a_n563_n140# a_683_n140# 0.01fF
C62 w_n1311_n241# a_n207_n140# 0.02fF
C63 a_n563_n140# a_n29_n140# 0.02fF
C64 a_n385_n140# a_n207_n140# 0.06fF
C65 a_683_n140# a_n29_n140# 0.01fF
C66 a_n563_n140# a_327_n140# 0.01fF
C67 a_n505_n205# a_741_n205# 0.01fF
C68 a_1097_n205# a_683_n140# 0.02fF
C69 w_n1311_n241# a_n1275_n140# 0.33fF
C70 a_n1097_n140# a_n207_n140# 0.01fF
C71 a_1097_n205# a_n29_n140# 0.01fF
C72 a_n385_n140# a_n1275_n140# 0.01fF
C73 a_327_n140# a_683_n140# 0.03fF
C74 a_327_n140# a_n29_n140# 0.03fF
C75 a_n1275_n140# a_n861_n205# 0.02fF
C76 a_n385_n140# w_n1311_n241# 0.02fF
C77 a_1097_n205# a_327_n140# 0.01fF
C78 w_n1311_n241# a_n861_n205# 0.20fF
C79 a_n1097_n140# a_n1275_n140# 0.06fF
C80 a_n1097_n140# w_n1311_n241# 0.02fF
C81 a_1097_n205# a_385_n205# 0.01fF
C82 a_n1097_n140# a_n385_n140# 0.01fF
C83 a_n505_n205# a_919_n205# 0.01fF
C84 a_1097_n205# a_29_n205# 0.01fF
C85 a_1097_n205# a_n327_n205# 0.00fF
C86 a_n149_n205# a_n1275_n140# 0.01fF
C87 a_385_n205# a_29_n205# 0.03fF
C88 a_1097_n205# a_563_n205# 0.01fF
C89 a_385_n205# a_n327_n205# 0.01fF
C90 a_n149_n205# w_n1311_n241# 0.19fF
C91 a_n683_n205# a_385_n205# 0.01fF
C92 a_n149_n205# a_n861_n205# 0.01fF
C93 a_385_n205# a_563_n205# 0.10fF
C94 a_1097_n205# a_207_n205# 0.01fF
C95 a_n327_n205# a_29_n205# 0.03fF
C96 a_n683_n205# a_29_n205# 0.01fF
C97 a_n683_n205# a_n327_n205# 0.03fF
C98 a_385_n205# a_207_n205# 0.10fF
C99 a_563_n205# a_29_n205# 0.02fF
C100 a_563_n205# a_n327_n205# 0.01fF
C101 a_1097_n205# a_741_n205# 0.02fF
C102 a_n683_n205# a_563_n205# 0.01fF
C103 a_385_n205# a_n1039_n205# 0.01fF
C104 a_n505_n205# a_n1275_n140# 0.01fF
C105 a_861_n140# a_n741_n140# 0.01fF
C106 a_n505_n205# w_n1311_n241# 0.20fF
C107 a_29_n205# a_207_n205# 0.10fF
C108 a_385_n205# a_741_n205# 0.03fF
C109 a_n505_n205# a_n861_n205# 0.03fF
C110 a_n327_n205# a_207_n205# 0.02fF
C111 a_n683_n205# a_207_n205# 0.01fF
C112 a_n919_n140# a_n741_n140# 0.06fF
C113 a_29_n205# a_n1039_n205# 0.01fF
C114 a_861_n140# a_n207_n140# 0.01fF
C115 a_n327_n205# a_n1039_n205# 0.01fF
C116 a_505_n140# a_n741_n140# 0.01fF
C117 a_n683_n205# a_n1039_n205# 0.03fF
C118 a_563_n205# a_207_n205# 0.03fF
C119 a_29_n205# a_741_n205# 0.01fF
C120 a_1097_n205# a_919_n205# 0.07fF
C121 a_n327_n205# a_741_n205# 0.01fF
C122 a_149_n140# a_n741_n140# 0.01fF
C123 a_n207_n140# a_n919_n140# 0.01fF
C124 a_563_n205# a_n1039_n205# 0.01fF
C125 a_n683_n205# a_741_n205# 0.01fF
C126 a_861_n140# w_n1311_n241# 0.01fF
C127 a_861_n140# a_n385_n140# 0.01fF
C128 a_505_n140# a_n207_n140# 0.01fF
C129 a_563_n205# a_741_n205# 0.10fF
C130 a_385_n205# a_919_n205# 0.02fF
C131 a_n1275_n140# a_n919_n140# 0.03fF
C132 a_149_n140# a_n207_n140# 0.03fF
C133 w_n1311_n241# a_n919_n140# 0.02fF
C134 a_207_n205# a_n1039_n205# 0.01fF
C135 a_n563_n140# a_n741_n140# 0.06fF
C136 a_n385_n140# a_n919_n140# 0.02fF
C137 a_1039_n140# a_n207_n140# 0.01fF
C138 a_n505_n205# a_n149_n205# 0.03fF
C139 a_683_n140# a_n741_n140# 0.01fF
C140 w_n1311_n241# a_505_n140# 0.02fF
C141 a_n385_n140# a_505_n140# 0.01fF
C142 a_n29_n140# a_n741_n140# 0.01fF
C143 a_n1275_n140# a_149_n140# 0.01fF
C144 a_207_n205# a_741_n205# 0.02fF
C145 a_29_n205# a_919_n205# 0.01fF
C146 a_n1097_n140# a_n919_n140# 0.06fF
C147 a_n327_n205# a_919_n205# 0.01fF
C148 a_327_n140# a_n741_n140# 0.01fF
C149 w_n1311_n241# a_149_n140# 0.02fF
C150 a_n385_n140# a_149_n140# 0.02fF
C151 a_n683_n205# a_919_n205# 0.01fF
C152 a_n563_n140# a_n207_n140# 0.03fF
C153 a_1039_n140# w_n1311_n241# 0.01fF
C154 a_n1097_n140# a_505_n140# 0.01fF
C155 a_1039_n140# a_n385_n140# 0.01fF
C156 a_683_n140# a_n207_n140# 0.01fF
C157 a_563_n205# a_919_n205# 0.03fF
C158 a_n207_n140# a_n29_n140# 0.06fF
C159 a_n1097_n140# a_149_n140# 0.01fF
C160 a_1097_n205# a_n207_n140# 0.01fF
C161 a_n563_n140# a_n1275_n140# 0.01fF
C162 a_327_n140# a_n207_n140# 0.02fF
C163 a_n563_n140# w_n1311_n241# 0.02fF
C164 a_n563_n140# a_n385_n140# 0.06fF
C165 a_n1275_n140# a_n29_n140# 0.01fF
C166 w_n1311_n241# a_683_n140# 0.02fF
C167 a_n385_n140# a_683_n140# 0.01fF
C168 w_n1311_n241# a_n29_n140# 0.02fF
C169 a_207_n205# a_919_n205# 0.01fF
C170 a_n1275_n140# a_327_n140# 0.01fF
C171 a_n385_n140# a_n29_n140# 0.03fF
C172 a_1097_n205# w_n1311_n241# 0.28fF
C173 a_n1097_n140# a_n563_n140# 0.02fF
C174 a_1097_n205# a_n385_n140# 0.01fF
C175 w_n1311_n241# a_327_n140# 0.02fF
C176 a_n385_n140# a_327_n140# 0.01fF
C177 a_385_n205# a_n1275_n140# 0.00fF
C178 a_n1097_n140# a_n29_n140# 0.01fF
C179 a_385_n205# w_n1311_n241# 0.17fF
C180 a_n1097_n140# a_327_n140# 0.01fF
C181 a_741_n205# a_919_n205# 0.10fF
C182 a_385_n205# a_n861_n205# 0.01fF
C183 a_n1275_n140# a_29_n205# 0.00fF
C184 a_n327_n205# a_n1275_n140# 0.01fF
C185 w_n1311_n241# a_29_n205# 0.19fF
C186 a_n683_n205# a_n1275_n140# 0.01fF
C187 a_n327_n205# w_n1311_n241# 0.20fF
C188 a_29_n205# a_n861_n205# 0.01fF
C189 a_n683_n205# w_n1311_n241# 0.20fF
C190 a_n327_n205# a_n861_n205# 0.02fF
C191 a_n683_n205# a_n861_n205# 0.10fF
C192 a_563_n205# w_n1311_n241# 0.16fF
C193 a_1097_n205# a_n149_n205# 0.00fF
C194 a_563_n205# a_n861_n205# 0.01fF
C195 a_n1275_n140# a_207_n205# 0.00fF
C196 a_385_n205# a_n149_n205# 0.02fF
C197 w_n1311_n241# a_207_n205# 0.18fF
C198 w_n1311_n241# VSUBS 3.79fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AKSJZW a_n149_n195# a_n207_n140# a_207_n195# a_327_n140#
+ a_n1275_n140# a_n861_n195# a_n29_n140# a_149_n140# a_n1097_n140# a_n1039_n195# a_29_n195#
+ a_n683_n195# a_n741_n140# a_741_n195# a_861_n140# a_1097_n195# a_n563_n140# a_n505_n195#
+ a_563_n195# a_683_n140# a_n919_n140# a_919_n195# a_1039_n140# a_n385_n140# a_n327_n195#
+ a_385_n195# a_505_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n195# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n195# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n195# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n195# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_327_n140# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_861_n140# a_741_n195# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n207_n140# a_n327_n195# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_1097_n195# a_1097_n195# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n195# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1275_n140# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n195# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n195# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n207_n140# a_683_n140# 0.01fF
C1 a_n149_n195# a_n861_n195# 0.01fF
C2 a_n207_n140# a_861_n140# 0.01fF
C3 a_505_n140# a_n563_n140# 0.01fF
C4 a_149_n140# a_327_n140# 0.06fF
C5 a_149_n140# a_683_n140# 0.02fF
C6 a_n385_n140# a_n29_n140# 0.03fF
C7 a_861_n140# a_149_n140# 0.01fF
C8 a_n1275_n140# a_n919_n140# 0.03fF
C9 a_919_n195# a_n505_n195# 0.01fF
C10 a_505_n140# a_n1097_n140# 0.01fF
C11 a_n1275_n140# a_n505_n195# 0.01fF
C12 a_n207_n140# a_n919_n140# 0.01fF
C13 a_n563_n140# a_327_n140# 0.01fF
C14 a_1097_n195# a_505_n140# 0.01fF
C15 a_n563_n140# a_683_n140# 0.01fF
C16 a_741_n195# a_n861_n195# 0.01fF
C17 a_n1039_n195# a_n505_n195# 0.02fF
C18 a_n563_n140# a_861_n140# 0.01fF
C19 a_n207_n140# a_n1275_n140# 0.01fF
C20 a_505_n140# a_1039_n140# 0.02fF
C21 a_n1039_n195# a_n1275_n140# 0.06fF
C22 a_149_n140# a_n919_n140# 0.01fF
C23 a_n1097_n140# a_327_n140# 0.01fF
C24 a_1097_n195# a_327_n140# 0.01fF
C25 a_1097_n195# a_683_n140# 0.02fF
C26 a_n683_n195# a_n505_n195# 0.10fF
C27 a_n683_n195# a_919_n195# 0.01fF
C28 a_149_n140# a_n1275_n140# 0.01fF
C29 a_1097_n195# a_861_n140# 0.03fF
C30 a_n563_n140# a_n919_n140# 0.03fF
C31 a_n683_n195# a_n1275_n140# 0.01fF
C32 a_327_n140# a_1039_n140# 0.01fF
C33 a_n207_n140# a_149_n140# 0.03fF
C34 a_n327_n195# a_n505_n195# 0.10fF
C35 a_1039_n140# a_683_n140# 0.03fF
C36 a_n327_n195# a_919_n195# 0.01fF
C37 a_n683_n195# a_n1039_n195# 0.03fF
C38 a_861_n140# a_1039_n140# 0.06fF
C39 a_n327_n195# a_n1275_n140# 0.01fF
C40 a_n563_n140# a_n1275_n140# 0.01fF
C41 a_505_n140# a_n741_n140# 0.01fF
C42 a_n1097_n140# a_n919_n140# 0.06fF
C43 a_29_n195# a_n505_n195# 0.02fF
C44 a_n207_n140# a_n563_n140# 0.03fF
C45 a_n327_n195# a_n1039_n195# 0.01fF
C46 a_29_n195# a_919_n195# 0.01fF
C47 a_29_n195# a_n1275_n140# 0.00fF
C48 a_1097_n195# a_n505_n195# 0.00fF
C49 a_n1097_n140# a_n1275_n140# 0.06fF
C50 a_1097_n195# a_919_n195# 0.06fF
C51 a_29_n195# a_n1039_n195# 0.01fF
C52 a_207_n195# a_n505_n195# 0.01fF
C53 a_327_n140# a_n741_n140# 0.01fF
C54 a_n563_n140# a_149_n140# 0.01fF
C55 a_n207_n140# a_n1097_n140# 0.01fF
C56 a_919_n195# a_207_n195# 0.01fF
C57 a_n741_n140# a_683_n140# 0.01fF
C58 a_385_n195# a_n505_n195# 0.01fF
C59 a_n327_n195# a_n683_n195# 0.03fF
C60 a_385_n195# a_919_n195# 0.02fF
C61 a_563_n195# a_n505_n195# 0.01fF
C62 a_207_n195# a_n1275_n140# 0.00fF
C63 a_1097_n195# a_n207_n140# 0.01fF
C64 a_861_n140# a_n741_n140# 0.01fF
C65 a_563_n195# a_919_n195# 0.03fF
C66 a_385_n195# a_n1275_n140# 0.00fF
C67 a_n1039_n195# a_207_n195# 0.01fF
C68 a_n683_n195# a_29_n195# 0.01fF
C69 a_149_n140# a_n1097_n140# 0.01fF
C70 a_n207_n140# a_1039_n140# 0.01fF
C71 a_385_n195# a_n1039_n195# 0.01fF
C72 a_563_n195# a_n1039_n195# 0.01fF
C73 a_505_n140# a_n29_n140# 0.02fF
C74 a_1097_n195# a_149_n140# 0.01fF
C75 a_n327_n195# a_29_n195# 0.03fF
C76 a_n919_n140# a_n741_n140# 0.06fF
C77 a_n563_n140# a_n1097_n140# 0.02fF
C78 a_n683_n195# a_207_n195# 0.01fF
C79 a_149_n140# a_1039_n140# 0.01fF
C80 a_n683_n195# a_385_n195# 0.01fF
C81 a_1097_n195# a_n327_n195# 0.00fF
C82 a_563_n195# a_n683_n195# 0.01fF
C83 a_n29_n140# a_327_n140# 0.03fF
C84 a_n327_n195# a_207_n195# 0.02fF
C85 a_n1275_n140# a_n741_n140# 0.02fF
C86 a_n29_n140# a_683_n140# 0.01fF
C87 a_n327_n195# a_385_n195# 0.01fF
C88 a_n149_n195# a_n505_n195# 0.03fF
C89 a_n207_n140# a_n741_n140# 0.02fF
C90 a_n563_n140# a_1039_n140# 0.01fF
C91 a_563_n195# a_n327_n195# 0.01fF
C92 a_1097_n195# a_29_n195# 0.01fF
C93 a_n29_n140# a_861_n140# 0.01fF
C94 a_919_n195# a_n149_n195# 0.01fF
C95 a_n1275_n140# a_n149_n195# 0.01fF
C96 a_29_n195# a_207_n195# 0.10fF
C97 a_n385_n140# a_505_n140# 0.01fF
C98 a_29_n195# a_385_n195# 0.03fF
C99 a_563_n195# a_29_n195# 0.02fF
C100 a_n1039_n195# a_n149_n195# 0.01fF
C101 a_149_n140# a_n741_n140# 0.01fF
C102 a_1097_n195# a_207_n195# 0.01fF
C103 a_1097_n195# a_385_n195# 0.01fF
C104 a_1097_n195# a_1039_n140# 0.06fF
C105 a_563_n195# a_1097_n195# 0.01fF
C106 a_n29_n140# a_n919_n140# 0.01fF
C107 a_385_n195# a_207_n195# 0.10fF
C108 a_n385_n140# a_327_n140# 0.01fF
C109 a_563_n195# a_207_n195# 0.03fF
C110 a_n385_n140# a_683_n140# 0.01fF
C111 a_n563_n140# a_n741_n140# 0.06fF
C112 a_741_n195# a_n505_n195# 0.01fF
C113 a_n683_n195# a_n149_n195# 0.02fF
C114 a_563_n195# a_385_n195# 0.10fF
C115 a_741_n195# a_919_n195# 0.10fF
C116 a_n385_n140# a_861_n140# 0.01fF
C117 a_n29_n140# a_n1275_n140# 0.01fF
C118 a_n29_n140# a_n207_n140# 0.06fF
C119 a_n327_n195# a_n149_n195# 0.10fF
C120 a_n1097_n140# a_n741_n140# 0.03fF
C121 a_29_n195# a_n149_n195# 0.10fF
C122 a_n29_n140# a_149_n140# 0.06fF
C123 a_n385_n140# a_n919_n140# 0.02fF
C124 a_n683_n195# a_741_n195# 0.01fF
C125 a_1097_n195# a_n149_n195# 0.00fF
C126 a_207_n195# a_n149_n195# 0.03fF
C127 a_n385_n140# a_n1275_n140# 0.01fF
C128 a_n29_n140# a_n563_n140# 0.02fF
C129 a_385_n195# a_n149_n195# 0.02fF
C130 a_n327_n195# a_741_n195# 0.01fF
C131 a_n861_n195# a_n505_n195# 0.03fF
C132 a_563_n195# a_n149_n195# 0.01fF
C133 a_n385_n140# a_n207_n140# 0.06fF
C134 a_n1275_n140# a_n861_n195# 0.02fF
C135 a_29_n195# a_741_n195# 0.01fF
C136 a_n29_n140# a_n1097_n140# 0.01fF
C137 a_n1039_n195# a_n861_n195# 0.10fF
C138 a_n385_n140# a_149_n140# 0.02fF
C139 a_1097_n195# a_n29_n140# 0.01fF
C140 a_1097_n195# a_741_n195# 0.02fF
C141 a_741_n195# a_207_n195# 0.02fF
C142 a_n29_n140# a_1039_n140# 0.01fF
C143 a_385_n195# a_741_n195# 0.03fF
C144 a_n385_n140# a_n563_n140# 0.06fF
C145 a_n683_n195# a_n861_n195# 0.10fF
C146 a_563_n195# a_741_n195# 0.10fF
C147 a_n327_n195# a_n861_n195# 0.02fF
C148 a_n385_n140# a_n1097_n140# 0.01fF
C149 a_505_n140# a_327_n140# 0.06fF
C150 a_505_n140# a_683_n140# 0.06fF
C151 a_n385_n140# a_1097_n195# 0.01fF
C152 a_29_n195# a_n861_n195# 0.01fF
C153 a_505_n140# a_861_n140# 0.03fF
C154 a_n29_n140# a_n741_n140# 0.01fF
C155 a_n385_n140# a_1039_n140# 0.01fF
C156 a_327_n140# a_683_n140# 0.03fF
C157 a_207_n195# a_n861_n195# 0.01fF
C158 a_385_n195# a_n861_n195# 0.01fF
C159 a_741_n195# a_n149_n195# 0.01fF
C160 a_861_n140# a_327_n140# 0.02fF
C161 a_563_n195# a_n861_n195# 0.01fF
C162 a_861_n140# a_683_n140# 0.06fF
C163 a_505_n140# a_n919_n140# 0.01fF
C164 a_n385_n140# a_n741_n140# 0.03fF
C165 a_505_n140# a_n207_n140# 0.01fF
C166 a_327_n140# a_n919_n140# 0.01fF
C167 a_n919_n140# a_683_n140# 0.01fF
C168 a_n1275_n140# a_327_n140# 0.01fF
C169 a_505_n140# a_149_n140# 0.03fF
C170 a_n207_n140# a_327_n140# 0.02fF
C171 a_1039_n140# VSUBS 0.01fF
C172 a_861_n140# VSUBS 0.01fF
C173 a_683_n140# VSUBS 0.02fF
C174 a_505_n140# VSUBS 0.02fF
C175 a_327_n140# VSUBS 0.02fF
C176 a_149_n140# VSUBS 0.02fF
C177 a_n29_n140# VSUBS 0.02fF
C178 a_n207_n140# VSUBS 0.02fF
C179 a_n385_n140# VSUBS 0.02fF
C180 a_n563_n140# VSUBS 0.02fF
C181 a_n741_n140# VSUBS 0.02fF
C182 a_n919_n140# VSUBS 0.02fF
C183 a_n1097_n140# VSUBS 0.02fF
C184 a_1097_n195# VSUBS 0.31fF
C185 a_919_n195# VSUBS 0.19fF
C186 a_741_n195# VSUBS 0.20fF
C187 a_563_n195# VSUBS 0.21fF
C188 a_385_n195# VSUBS 0.22fF
C189 a_207_n195# VSUBS 0.23fF
C190 a_29_n195# VSUBS 0.23fF
C191 a_n149_n195# VSUBS 0.24fF
C192 a_n327_n195# VSUBS 0.24fF
C193 a_n505_n195# VSUBS 0.24fF
C194 a_n683_n195# VSUBS 0.24fF
C195 a_n861_n195# VSUBS 0.24fF
C196 a_n1039_n195# VSUBS 0.24fF
C197 a_n1275_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_K7HVMB a_664_n120# a_n608_n120# a_n86_n120# a_72_n208#
+ a_240_n120# a_n184_n120# a_n562_142# a_n510_n120# a_28_n120# a_n298_n120# a_126_n120#
+ a_452_n120# a_n396_n120# a_284_142# a_n138_142# a_550_n120# a_496_n208# a_338_n120#
+ a_n350_n208# a_n820_n120# VSUBS
X0 a_n820_n120# a_n820_n120# a_n820_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X1 a_n510_n120# a_n562_142# a_n608_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X2 a_664_n120# a_664_n120# a_664_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X3 a_n298_n120# a_n350_n208# a_n396_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X4 a_550_n120# a_496_n208# a_452_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X5 a_126_n120# a_72_n208# a_28_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X6 a_n86_n120# a_n138_142# a_n184_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X7 a_338_n120# a_284_142# a_240_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
C0 a_n820_n120# a_452_n120# 0.01fF
C1 a_n820_n120# a_664_n120# 0.02fF
C2 a_n350_n208# a_n138_142# 0.01fF
C3 a_n608_n120# a_550_n120# 0.01fF
C4 a_n350_n208# a_n562_142# 0.01fF
C5 a_72_n208# a_284_142# 0.01fF
C6 a_n298_n120# a_n608_n120# 0.03fF
C7 a_n820_n120# a_240_n120# 0.01fF
C8 a_n298_n120# a_550_n120# 0.01fF
C9 a_n820_n120# a_n510_n120# 0.06fF
C10 a_664_n120# a_n138_142# 0.00fF
C11 a_n396_n120# a_n820_n120# 0.04fF
C12 a_664_n120# a_n562_142# 0.00fF
C13 a_n820_n120# a_126_n120# 0.02fF
C14 a_n820_n120# a_28_n120# 0.02fF
C15 a_n86_n120# a_n820_n120# 0.02fF
C16 a_n510_n120# a_n562_142# 0.00fF
C17 a_n298_n120# a_n350_n208# 0.00fF
C18 a_452_n120# a_n608_n120# 0.01fF
C19 a_664_n120# a_n608_n120# 0.01fF
C20 a_n86_n120# a_n138_142# 0.00fF
C21 a_452_n120# a_550_n120# 0.11fF
C22 a_664_n120# a_550_n120# 0.13fF
C23 a_452_n120# a_n298_n120# 0.01fF
C24 a_664_n120# a_n298_n120# 0.01fF
C25 a_240_n120# a_n608_n120# 0.01fF
C26 a_n820_n120# a_496_n208# 0.00fF
C27 a_n510_n120# a_n608_n120# 0.11fF
C28 a_240_n120# a_550_n120# 0.03fF
C29 a_240_n120# a_n298_n120# 0.01fF
C30 a_n510_n120# a_550_n120# 0.01fF
C31 a_n396_n120# a_n608_n120# 0.04fF
C32 a_n298_n120# a_n510_n120# 0.04fF
C33 a_n820_n120# a_338_n120# 0.01fF
C34 a_n396_n120# a_550_n120# 0.01fF
C35 a_126_n120# a_n608_n120# 0.01fF
C36 a_n396_n120# a_n298_n120# 0.11fF
C37 a_28_n120# a_n608_n120# 0.01fF
C38 a_126_n120# a_550_n120# 0.02fF
C39 a_n138_142# a_496_n208# 0.00fF
C40 a_664_n120# a_n350_n208# 0.00fF
C41 a_n86_n120# a_n608_n120# 0.01fF
C42 a_496_n208# a_n562_142# 0.00fF
C43 a_n298_n120# a_126_n120# 0.02fF
C44 a_28_n120# a_550_n120# 0.01fF
C45 a_n86_n120# a_550_n120# 0.01fF
C46 a_28_n120# a_n298_n120# 0.02fF
C47 a_n86_n120# a_n298_n120# 0.04fF
C48 a_452_n120# a_664_n120# 0.06fF
C49 a_n820_n120# a_284_142# 0.00fF
C50 a_n820_n120# a_n184_n120# 0.03fF
C51 a_452_n120# a_240_n120# 0.04fF
C52 a_240_n120# a_664_n120# 0.03fF
C53 a_452_n120# a_n510_n120# 0.01fF
C54 a_664_n120# a_n510_n120# 0.01fF
C55 a_n396_n120# a_452_n120# 0.01fF
C56 a_n396_n120# a_664_n120# 0.01fF
C57 a_284_142# a_n138_142# 0.01fF
C58 a_452_n120# a_126_n120# 0.02fF
C59 a_n608_n120# a_338_n120# 0.01fF
C60 a_664_n120# a_126_n120# 0.03fF
C61 a_240_n120# a_n510_n120# 0.01fF
C62 a_284_142# a_n562_142# 0.01fF
C63 a_452_n120# a_28_n120# 0.02fF
C64 a_664_n120# a_28_n120# 0.02fF
C65 a_338_n120# a_550_n120# 0.04fF
C66 a_n86_n120# a_452_n120# 0.01fF
C67 a_n396_n120# a_240_n120# 0.01fF
C68 a_n86_n120# a_664_n120# 0.02fF
C69 a_n298_n120# a_338_n120# 0.01fF
C70 a_n396_n120# a_n510_n120# 0.09fF
C71 a_240_n120# a_126_n120# 0.09fF
C72 a_72_n208# a_n820_n120# 0.00fF
C73 a_240_n120# a_28_n120# 0.04fF
C74 a_126_n120# a_n510_n120# 0.01fF
C75 a_n86_n120# a_240_n120# 0.02fF
C76 a_28_n120# a_n510_n120# 0.01fF
C77 a_n350_n208# a_496_n208# 0.01fF
C78 a_n86_n120# a_n510_n120# 0.02fF
C79 a_n396_n120# a_126_n120# 0.01fF
C80 a_n396_n120# a_28_n120# 0.02fF
C81 a_n86_n120# a_n396_n120# 0.03fF
C82 a_28_n120# a_126_n120# 0.11fF
C83 a_n184_n120# a_n608_n120# 0.02fF
C84 a_72_n208# a_n138_142# 0.01fF
C85 a_n86_n120# a_126_n120# 0.04fF
C86 a_452_n120# a_496_n208# 0.00fF
C87 a_72_n208# a_n562_142# 0.00fF
C88 a_664_n120# a_496_n208# 0.01fF
C89 a_n184_n120# a_550_n120# 0.01fF
C90 a_n86_n120# a_28_n120# 0.09fF
C91 a_n184_n120# a_n298_n120# 0.09fF
C92 a_452_n120# a_338_n120# 0.09fF
C93 a_664_n120# a_338_n120# 0.04fF
C94 a_240_n120# a_338_n120# 0.11fF
C95 a_284_142# a_n350_n208# 0.00fF
C96 a_n510_n120# a_338_n120# 0.01fF
C97 a_n396_n120# a_338_n120# 0.01fF
C98 a_126_n120# a_338_n120# 0.04fF
C99 a_284_142# a_664_n120# 0.01fF
C100 a_28_n120# a_338_n120# 0.03fF
C101 a_452_n120# a_n184_n120# 0.01fF
C102 a_664_n120# a_n184_n120# 0.02fF
C103 a_n86_n120# a_338_n120# 0.02fF
C104 a_284_142# a_240_n120# 0.00fF
C105 a_240_n120# a_n184_n120# 0.02fF
C106 a_n184_n120# a_n510_n120# 0.02fF
C107 a_72_n208# a_n350_n208# 0.01fF
C108 a_n396_n120# a_n184_n120# 0.04fF
C109 a_n184_n120# a_126_n120# 0.03fF
C110 a_28_n120# a_n184_n120# 0.04fF
C111 a_72_n208# a_664_n120# 0.00fF
C112 a_n86_n120# a_n184_n120# 0.11fF
C113 a_n820_n120# a_n138_142# 0.00fF
C114 a_n820_n120# a_n562_142# 0.01fF
C115 a_284_142# a_496_n208# 0.01fF
C116 a_72_n208# a_28_n120# 0.00fF
C117 a_n138_142# a_n562_142# 0.01fF
C118 a_n184_n120# a_338_n120# 0.01fF
C119 a_n820_n120# a_n608_n120# 0.13fF
C120 a_n820_n120# a_550_n120# 0.01fF
C121 a_n820_n120# a_n298_n120# 0.03fF
C122 a_72_n208# a_496_n208# 0.01fF
C123 a_n820_n120# a_n350_n208# 0.01fF
C124 a_550_n120# VSUBS 0.01fF
C125 a_452_n120# VSUBS 0.01fF
C126 a_338_n120# VSUBS 0.01fF
C127 a_240_n120# VSUBS 0.01fF
C128 a_126_n120# VSUBS 0.02fF
C129 a_28_n120# VSUBS 0.01fF
C130 a_n86_n120# VSUBS 0.01fF
C131 a_n184_n120# VSUBS 0.02fF
C132 a_n298_n120# VSUBS 0.02fF
C133 a_n396_n120# VSUBS 0.02fF
C134 a_n510_n120# VSUBS 0.02fF
C135 a_n608_n120# VSUBS 0.02fF
C136 a_496_n208# VSUBS 0.11fF
C137 a_664_n120# VSUBS 0.17fF
C138 a_72_n208# VSUBS 0.10fF
C139 a_284_142# VSUBS 0.10fF
C140 a_n350_n208# VSUBS 0.12fF
C141 a_n138_142# VSUBS 0.11fF
C142 a_n820_n120# VSUBS 0.20fF
C143 a_n562_142# VSUBS 0.14fF
.ends

.subckt sky130_fd_pr__nfet_01v8_S6RQQZ a_n149_n194# a_n207_n140# a_207_n194# a_1453_n194#
+ a_n1217_n194# a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140#
+ a_n1097_n140# a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194#
+ a_861_n140# a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140#
+ a_n919_n140# a_919_n194# a_n1631_n140# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194#
+ a_n1395_n194# a_505_n140# a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n1453_n140# a_n1631_n140# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1453_n194# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n505_n194# a_n1631_n140# 0.01fF
C1 a_n207_n140# a_n563_n140# 0.03fF
C2 a_861_n140# a_1217_n140# 0.03fF
C3 a_683_n140# a_149_n140# 0.02fF
C4 a_327_n140# a_n29_n140# 0.03fF
C5 a_n207_n140# a_n385_n140# 0.06fF
C6 a_683_n140# a_861_n140# 0.06fF
C7 a_n1039_n194# a_n861_n194# 0.10fF
C8 a_n1039_n194# a_563_n194# 0.01fF
C9 a_n563_n140# a_1039_n140# 0.01fF
C10 a_n1097_n140# a_n919_n140# 0.06fF
C11 a_n1039_n194# a_n1217_n194# 0.10fF
C12 a_n1275_n140# a_n29_n140# 0.01fF
C13 a_n1097_n140# a_n563_n140# 0.02fF
C14 a_n1453_n140# a_n1275_n140# 0.06fF
C15 a_n385_n140# a_1039_n140# 0.01fF
C16 a_563_n194# a_1097_n194# 0.02fF
C17 a_n385_n140# a_n1097_n140# 0.01fF
C18 a_n1039_n194# a_n1395_n194# 0.03fF
C19 a_563_n194# a_n861_n194# 0.01fF
C20 a_n207_n140# a_1395_n140# 0.01fF
C21 a_n1217_n194# a_n861_n194# 0.03fF
C22 a_327_n140# a_1217_n140# 0.01fF
C23 a_n1275_n140# a_n1631_n140# 0.03fF
C24 a_327_n140# a_683_n140# 0.03fF
C25 a_n1395_n194# a_n861_n194# 0.02fF
C26 a_1395_n140# a_1039_n140# 0.03fF
C27 a_n741_n140# a_505_n140# 0.01fF
C28 a_n1395_n194# a_n1217_n194# 0.10fF
C29 a_n1039_n194# a_n683_n194# 0.03fF
C30 a_n1453_n140# a_n29_n140# 0.01fF
C31 a_1453_n194# a_1395_n140# 0.06fF
C32 a_n207_n140# a_1039_n140# 0.01fF
C33 a_1453_n194# a_1097_n194# 0.02fF
C34 a_n919_n140# a_505_n140# 0.01fF
C35 a_n207_n140# a_n1097_n140# 0.01fF
C36 a_n29_n140# a_n1631_n140# 0.01fF
C37 a_n1039_n194# a_n327_n194# 0.01fF
C38 a_n683_n194# a_n861_n194# 0.10fF
C39 a_505_n140# a_n563_n140# 0.01fF
C40 a_n1453_n140# a_n1631_n140# 0.06fF
C41 a_n683_n194# a_563_n194# 0.01fF
C42 a_1453_n194# a_563_n194# 0.01fF
C43 a_n385_n140# a_505_n140# 0.01fF
C44 a_n683_n194# a_n1217_n194# 0.02fF
C45 a_n29_n140# a_1217_n140# 0.01fF
C46 a_n327_n194# a_1097_n194# 0.01fF
C47 a_n741_n140# a_149_n140# 0.01fF
C48 a_n741_n140# a_861_n140# 0.01fF
C49 a_919_n194# a_1097_n194# 0.10fF
C50 a_n327_n194# a_n861_n194# 0.02fF
C51 a_n29_n140# a_683_n140# 0.01fF
C52 a_n683_n194# a_n1395_n194# 0.01fF
C53 a_n1039_n194# a_n149_n194# 0.01fF
C54 a_n327_n194# a_563_n194# 0.01fF
C55 a_741_n194# a_1097_n194# 0.03fF
C56 a_n1039_n194# a_29_n194# 0.01fF
C57 a_n327_n194# a_n1217_n194# 0.01fF
C58 a_563_n194# a_919_n194# 0.03fF
C59 a_207_n194# a_n1039_n194# 0.01fF
C60 a_741_n194# a_n861_n194# 0.01fF
C61 a_n149_n194# a_1097_n194# 0.01fF
C62 a_1395_n140# a_505_n140# 0.01fF
C63 a_741_n194# a_563_n194# 0.10fF
C64 a_1453_n194# a_1039_n140# 0.02fF
C65 a_n327_n194# a_n1395_n194# 0.01fF
C66 a_29_n194# a_1097_n194# 0.01fF
C67 a_n919_n140# a_149_n140# 0.01fF
C68 a_n149_n194# a_n861_n194# 0.01fF
C69 a_207_n194# a_1097_n194# 0.01fF
C70 a_n563_n140# a_149_n140# 0.01fF
C71 a_563_n194# a_n149_n194# 0.01fF
C72 a_29_n194# a_n861_n194# 0.01fF
C73 a_861_n140# a_n563_n140# 0.01fF
C74 a_29_n194# a_563_n194# 0.02fF
C75 a_207_n194# a_n861_n194# 0.01fF
C76 a_n149_n194# a_n1217_n194# 0.01fF
C77 a_n385_n140# a_149_n140# 0.02fF
C78 a_207_n194# a_563_n194# 0.03fF
C79 a_683_n140# a_1217_n140# 0.02fF
C80 a_29_n194# a_n1217_n194# 0.01fF
C81 a_n385_n140# a_861_n140# 0.01fF
C82 a_n741_n140# a_327_n140# 0.01fF
C83 a_207_n194# a_n1217_n194# 0.01fF
C84 a_n1395_n194# a_n149_n194# 0.01fF
C85 a_n207_n140# a_505_n140# 0.01fF
C86 a_29_n194# a_n1395_n194# 0.01fF
C87 a_207_n194# a_n1395_n194# 0.01fF
C88 a_n741_n140# a_n1275_n140# 0.02fF
C89 a_1395_n140# a_149_n140# 0.01fF
C90 a_n683_n194# a_n327_n194# 0.03fF
C91 a_861_n140# a_1395_n140# 0.02fF
C92 a_505_n140# a_1039_n140# 0.02fF
C93 a_n683_n194# a_919_n194# 0.01fF
C94 a_1097_n194# a_1275_n194# 0.10fF
C95 a_1453_n194# a_919_n194# 0.01fF
C96 a_327_n140# a_n919_n140# 0.01fF
C97 a_n1097_n140# a_505_n140# 0.01fF
C98 a_327_n140# a_n563_n140# 0.01fF
C99 a_n1039_n194# a_n505_n194# 0.02fF
C100 a_741_n194# a_n683_n194# 0.01fF
C101 a_741_n194# a_1453_n194# 0.01fF
C102 a_563_n194# a_1275_n194# 0.01fF
C103 a_327_n140# a_n385_n140# 0.01fF
C104 a_n1275_n140# a_n919_n140# 0.03fF
C105 a_n683_n194# a_n149_n194# 0.02fF
C106 a_1097_n194# a_n505_n194# 0.01fF
C107 a_n327_n194# a_919_n194# 0.01fF
C108 a_1453_n194# a_n149_n194# 0.00fF
C109 a_n1275_n140# a_n563_n140# 0.01fF
C110 a_n683_n194# a_29_n194# 0.01fF
C111 a_1453_n194# a_29_n194# 0.00fF
C112 a_n207_n140# a_149_n140# 0.03fF
C113 a_n505_n194# a_n861_n194# 0.03fF
C114 a_1453_n194# a_505_n140# 0.01fF
C115 a_207_n194# a_n683_n194# 0.01fF
C116 a_207_n194# a_1453_n194# 0.00fF
C117 a_741_n194# a_n327_n194# 0.01fF
C118 a_n1275_n140# a_n385_n140# 0.01fF
C119 a_563_n194# a_n505_n194# 0.01fF
C120 a_n207_n140# a_861_n140# 0.01fF
C121 a_741_n194# a_919_n194# 0.10fF
C122 a_n741_n140# a_n29_n140# 0.01fF
C123 a_n1217_n194# a_n505_n194# 0.01fF
C124 a_n327_n194# a_n149_n194# 0.10fF
C125 a_n1453_n140# a_n741_n140# 0.01fF
C126 a_327_n140# a_1395_n140# 0.01fF
C127 a_n327_n194# a_29_n194# 0.03fF
C128 a_n149_n194# a_919_n194# 0.01fF
C129 a_1039_n140# a_149_n140# 0.01fF
C130 a_207_n194# a_n327_n194# 0.02fF
C131 a_n1395_n194# a_n505_n194# 0.01fF
C132 a_29_n194# a_919_n194# 0.01fF
C133 a_n1097_n140# a_149_n140# 0.01fF
C134 a_861_n140# a_1039_n140# 0.06fF
C135 a_741_n194# a_n149_n194# 0.01fF
C136 a_207_n194# a_919_n194# 0.01fF
C137 a_n1039_n194# a_385_n194# 0.01fF
C138 a_n741_n140# a_n1631_n140# 0.01fF
C139 a_741_n194# a_29_n194# 0.01fF
C140 a_207_n194# a_741_n194# 0.02fF
C141 a_n29_n140# a_n919_n140# 0.01fF
C142 a_29_n194# a_n149_n194# 0.10fF
C143 a_385_n194# a_1097_n194# 0.01fF
C144 a_n29_n140# a_n563_n140# 0.02fF
C145 a_n1453_n140# a_n919_n140# 0.02fF
C146 a_207_n194# a_n149_n194# 0.03fF
C147 a_1453_n194# a_149_n140# 0.01fF
C148 a_n1453_n140# a_n563_n140# 0.01fF
C149 a_1453_n194# a_1275_n194# 0.06fF
C150 a_385_n194# a_n861_n194# 0.01fF
C151 a_327_n140# a_n207_n140# 0.02fF
C152 a_207_n194# a_29_n194# 0.10fF
C153 a_n29_n140# a_n385_n140# 0.03fF
C154 a_1453_n194# a_861_n140# 0.01fF
C155 a_385_n194# a_563_n194# 0.10fF
C156 a_n741_n140# a_683_n140# 0.01fF
C157 a_n1453_n140# a_n385_n140# 0.01fF
C158 a_385_n194# a_n1217_n194# 0.01fF
C159 a_n919_n140# a_n1631_n140# 0.01fF
C160 a_n1275_n140# a_n207_n140# 0.01fF
C161 a_n683_n194# a_n505_n194# 0.10fF
C162 a_n1631_n140# a_n563_n140# 0.01fF
C163 a_n327_n194# a_1275_n194# 0.01fF
C164 a_327_n140# a_1039_n140# 0.01fF
C165 a_919_n194# a_1275_n194# 0.03fF
C166 a_327_n140# a_n1097_n140# 0.01fF
C167 a_n385_n140# a_n1631_n140# 0.01fF
C168 a_n29_n140# a_1395_n140# 0.01fF
C169 a_741_n194# a_1275_n194# 0.02fF
C170 a_n327_n194# a_n505_n194# 0.10fF
C171 a_683_n140# a_n919_n140# 0.01fF
C172 a_n385_n140# a_1217_n140# 0.01fF
C173 a_n1275_n140# a_n1097_n140# 0.06fF
C174 a_683_n140# a_n563_n140# 0.01fF
C175 a_919_n194# a_n505_n194# 0.01fF
C176 a_n149_n194# a_1275_n194# 0.01fF
C177 a_29_n194# a_1275_n194# 0.01fF
C178 a_327_n140# a_1453_n194# 0.01fF
C179 a_n1039_n194# a_n1631_n140# 0.01fF
C180 a_505_n140# a_149_n140# 0.03fF
C181 a_683_n140# a_n385_n140# 0.01fF
C182 a_207_n194# a_1275_n194# 0.01fF
C183 a_741_n194# a_n505_n194# 0.01fF
C184 a_861_n140# a_505_n140# 0.03fF
C185 a_n149_n194# a_n505_n194# 0.03fF
C186 a_n683_n194# a_385_n194# 0.01fF
C187 a_29_n194# a_n505_n194# 0.02fF
C188 a_n207_n140# a_n29_n140# 0.06fF
C189 a_1453_n194# a_385_n194# 0.01fF
C190 a_1395_n140# a_1217_n140# 0.06fF
C191 a_n1631_n140# a_n861_n194# 0.01fF
C192 a_n1453_n140# a_n207_n140# 0.01fF
C193 a_207_n194# a_n505_n194# 0.01fF
C194 a_683_n140# a_1395_n140# 0.01fF
C195 a_n1217_n194# a_n1631_n140# 0.02fF
C196 a_n29_n140# a_1039_n140# 0.01fF
C197 a_n327_n194# a_385_n194# 0.01fF
C198 a_n207_n140# a_n1631_n140# 0.01fF
C199 a_n29_n140# a_n1097_n140# 0.01fF
C200 a_n1395_n194# a_n1631_n140# 0.06fF
C201 a_385_n194# a_919_n194# 0.02fF
C202 a_n1453_n140# a_n1097_n140# 0.03fF
C203 a_327_n140# a_505_n140# 0.06fF
C204 a_861_n140# a_149_n140# 0.01fF
C205 a_741_n194# a_385_n194# 0.03fF
C206 a_n207_n140# a_1217_n140# 0.01fF
C207 a_385_n194# a_n149_n194# 0.02fF
C208 a_n207_n140# a_683_n140# 0.01fF
C209 a_n1097_n140# a_n1631_n140# 0.02fF
C210 a_1453_n194# a_n29_n140# 0.01fF
C211 a_29_n194# a_385_n194# 0.03fF
C212 a_207_n194# a_385_n194# 0.10fF
C213 a_1039_n140# a_1217_n140# 0.06fF
C214 a_683_n140# a_1039_n140# 0.03fF
C215 a_n683_n194# a_n1631_n140# 0.01fF
C216 a_n741_n140# a_n919_n140# 0.06fF
C217 a_327_n140# a_149_n140# 0.06fF
C218 a_n741_n140# a_n563_n140# 0.06fF
C219 a_1453_n194# a_1217_n140# 0.03fF
C220 a_327_n140# a_861_n140# 0.02fF
C221 a_n327_n194# a_n1631_n140# 0.00fF
C222 a_n741_n140# a_n385_n140# 0.03fF
C223 a_1453_n194# a_683_n140# 0.01fF
C224 a_n1275_n140# a_149_n140# 0.01fF
C225 a_n29_n140# a_505_n140# 0.02fF
C226 a_385_n194# a_1275_n194# 0.01fF
C227 a_n919_n140# a_n563_n140# 0.03fF
C228 a_n149_n194# a_n1631_n140# 0.00fF
C229 a_385_n194# a_n505_n194# 0.01fF
C230 a_29_n194# a_n1631_n140# 0.00fF
C231 a_n385_n140# a_n919_n140# 0.02fF
C232 a_n385_n140# a_n563_n140# 0.06fF
C233 a_505_n140# a_1217_n140# 0.01fF
C234 a_683_n140# a_505_n140# 0.06fF
C235 a_n1275_n140# a_327_n140# 0.01fF
C236 a_n29_n140# a_149_n140# 0.06fF
C237 a_n1453_n140# a_149_n140# 0.01fF
C238 a_n29_n140# a_861_n140# 0.01fF
C239 a_n741_n140# a_n207_n140# 0.02fF
C240 a_n741_n140# a_n1097_n140# 0.03fF
C241 a_1217_n140# a_149_n140# 0.01fF
C242 a_n207_n140# a_n919_n140# 0.01fF
C243 a_1395_n140# VSUBS 0.01fF
C244 a_1217_n140# VSUBS 0.01fF
C245 a_1039_n140# VSUBS 0.02fF
C246 a_861_n140# VSUBS 0.02fF
C247 a_683_n140# VSUBS 0.02fF
C248 a_505_n140# VSUBS 0.02fF
C249 a_327_n140# VSUBS 0.02fF
C250 a_149_n140# VSUBS 0.02fF
C251 a_n29_n140# VSUBS 0.02fF
C252 a_n207_n140# VSUBS 0.02fF
C253 a_n385_n140# VSUBS 0.02fF
C254 a_n563_n140# VSUBS 0.02fF
C255 a_n741_n140# VSUBS 0.02fF
C256 a_n919_n140# VSUBS 0.02fF
C257 a_n1097_n140# VSUBS 0.02fF
C258 a_n1275_n140# VSUBS 0.02fF
C259 a_n1453_n140# VSUBS 0.02fF
C260 a_1453_n194# VSUBS 0.31fF
C261 a_1275_n194# VSUBS 0.19fF
C262 a_1097_n194# VSUBS 0.20fF
C263 a_919_n194# VSUBS 0.21fF
C264 a_741_n194# VSUBS 0.22fF
C265 a_563_n194# VSUBS 0.23fF
C266 a_385_n194# VSUBS 0.23fF
C267 a_207_n194# VSUBS 0.24fF
C268 a_29_n194# VSUBS 0.24fF
C269 a_n149_n194# VSUBS 0.24fF
C270 a_n327_n194# VSUBS 0.24fF
C271 a_n505_n194# VSUBS 0.24fF
C272 a_n683_n194# VSUBS 0.24fF
C273 a_n861_n194# VSUBS 0.24fF
C274 a_n1039_n194# VSUBS 0.24fF
C275 a_n1217_n194# VSUBS 0.24fF
C276 a_n1395_n194# VSUBS 0.24fF
C277 a_n1631_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6RUDQZ a_n594_n195# a_n1008_n140# a_n652_n140# a_652_n195#
+ a_772_n140# a_n60_n195# a_n474_n140# a_n416_n195# a_474_n195# a_594_n140# a_n296_n140#
+ a_n238_n195# a_60_n140# a_296_n195# a_416_n140# a_n118_n140# a_118_n195# a_238_n140#
+ a_n772_n195# a_n830_n140# a_830_n195# VSUBS
X0 a_772_n140# a_652_n195# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n195# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n195# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n195# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n195# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_830_n195# a_830_n195# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n1008_n140# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n195# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n195# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n195# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n195# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_474_n195# a_830_n195# 0.02fF
C1 a_n594_n195# a_n1008_n140# 0.02fF
C2 a_n416_n195# a_118_n195# 0.02fF
C3 a_n60_n195# a_296_n195# 0.03fF
C4 a_474_n195# a_652_n195# 0.10fF
C5 a_n416_n195# a_n594_n195# 0.10fF
C6 a_n830_n140# a_60_n140# 0.01fF
C7 a_830_n195# a_n772_n195# 0.00fF
C8 a_n474_n140# a_n652_n140# 0.06fF
C9 a_n474_n140# a_830_n195# 0.01fF
C10 a_652_n195# a_n772_n195# 0.01fF
C11 a_n118_n140# a_n296_n140# 0.06fF
C12 a_n830_n140# a_594_n140# 0.01fF
C13 a_60_n140# a_n652_n140# 0.01fF
C14 a_n60_n195# a_n1008_n140# 0.01fF
C15 a_772_n140# a_n830_n140# 0.01fF
C16 a_60_n140# a_830_n195# 0.01fF
C17 a_n60_n195# a_n416_n195# 0.03fF
C18 a_n296_n140# a_n1008_n140# 0.01fF
C19 a_594_n140# a_n652_n140# 0.01fF
C20 a_n474_n140# a_416_n140# 0.01fF
C21 a_594_n140# a_830_n195# 0.03fF
C22 a_772_n140# a_n652_n140# 0.01fF
C23 a_772_n140# a_830_n195# 0.06fF
C24 a_474_n195# a_n772_n195# 0.01fF
C25 a_60_n140# a_416_n140# 0.03fF
C26 a_n238_n195# a_830_n195# 0.01fF
C27 a_652_n195# a_n238_n195# 0.01fF
C28 a_296_n195# a_n1008_n140# 0.00fF
C29 a_n830_n140# a_238_n140# 0.01fF
C30 a_n118_n140# a_n1008_n140# 0.01fF
C31 a_594_n140# a_416_n140# 0.06fF
C32 a_296_n195# a_n416_n195# 0.01fF
C33 a_772_n140# a_416_n140# 0.03fF
C34 a_n652_n140# a_238_n140# 0.01fF
C35 a_60_n140# a_n474_n140# 0.02fF
C36 a_830_n195# a_118_n195# 0.01fF
C37 a_238_n140# a_830_n195# 0.01fF
C38 a_n594_n195# a_830_n195# 0.00fF
C39 a_652_n195# a_118_n195# 0.02fF
C40 a_n416_n195# a_n1008_n140# 0.01fF
C41 a_652_n195# a_n594_n195# 0.01fF
C42 a_n474_n140# a_594_n140# 0.01fF
C43 a_474_n195# a_n238_n195# 0.01fF
C44 a_n830_n140# a_n296_n140# 0.02fF
C45 a_772_n140# a_n474_n140# 0.01fF
C46 a_n238_n195# a_n772_n195# 0.02fF
C47 a_416_n140# a_238_n140# 0.06fF
C48 a_60_n140# a_594_n140# 0.02fF
C49 a_n60_n195# a_830_n195# 0.01fF
C50 a_772_n140# a_60_n140# 0.01fF
C51 a_n60_n195# a_652_n195# 0.01fF
C52 a_n296_n140# a_n652_n140# 0.03fF
C53 a_n296_n140# a_830_n195# 0.01fF
C54 a_474_n195# a_118_n195# 0.03fF
C55 a_474_n195# a_n594_n195# 0.01fF
C56 a_772_n140# a_594_n140# 0.06fF
C57 a_n118_n140# a_n830_n140# 0.01fF
C58 a_n772_n195# a_118_n195# 0.01fF
C59 a_n594_n195# a_n772_n195# 0.10fF
C60 a_n474_n140# a_238_n140# 0.01fF
C61 a_n296_n140# a_416_n140# 0.01fF
C62 a_296_n195# a_830_n195# 0.01fF
C63 a_n118_n140# a_n652_n140# 0.02fF
C64 a_n830_n140# a_n1008_n140# 0.06fF
C65 a_n118_n140# a_830_n195# 0.01fF
C66 a_60_n140# a_238_n140# 0.06fF
C67 a_n60_n195# a_474_n195# 0.02fF
C68 a_296_n195# a_652_n195# 0.03fF
C69 a_n60_n195# a_n772_n195# 0.01fF
C70 a_594_n140# a_238_n140# 0.03fF
C71 a_n652_n140# a_n1008_n140# 0.03fF
C72 a_772_n140# a_238_n140# 0.02fF
C73 a_652_n195# a_n1008_n140# 0.00fF
C74 a_n296_n140# a_n474_n140# 0.06fF
C75 a_n416_n195# a_830_n195# 0.00fF
C76 a_n118_n140# a_416_n140# 0.02fF
C77 a_n238_n195# a_118_n195# 0.03fF
C78 a_n416_n195# a_652_n195# 0.01fF
C79 a_n594_n195# a_n238_n195# 0.03fF
C80 a_n296_n140# a_60_n140# 0.03fF
C81 a_474_n195# a_296_n195# 0.10fF
C82 a_416_n140# a_n1008_n140# 0.01fF
C83 a_296_n195# a_n772_n195# 0.01fF
C84 a_n296_n140# a_594_n140# 0.01fF
C85 a_n118_n140# a_n474_n140# 0.03fF
C86 a_772_n140# a_n296_n140# 0.01fF
C87 a_n60_n195# a_n238_n195# 0.10fF
C88 a_n594_n195# a_118_n195# 0.01fF
C89 a_474_n195# a_n1008_n140# 0.00fF
C90 a_474_n195# a_n416_n195# 0.01fF
C91 a_n118_n140# a_60_n140# 0.06fF
C92 a_n772_n195# a_n1008_n140# 0.06fF
C93 a_n474_n140# a_n1008_n140# 0.02fF
C94 a_n416_n195# a_n772_n195# 0.03fF
C95 a_n118_n140# a_594_n140# 0.01fF
C96 a_n830_n140# a_n652_n140# 0.06fF
C97 a_n60_n195# a_118_n195# 0.10fF
C98 a_60_n140# a_n1008_n140# 0.01fF
C99 a_n60_n195# a_n594_n195# 0.02fF
C100 a_n118_n140# a_772_n140# 0.01fF
C101 a_n296_n140# a_238_n140# 0.02fF
C102 a_296_n195# a_n238_n195# 0.02fF
C103 a_594_n140# a_n1008_n140# 0.01fF
C104 a_n652_n140# a_830_n195# 0.01fF
C105 a_652_n195# a_830_n195# 0.06fF
C106 a_n830_n140# a_416_n140# 0.01fF
C107 a_n238_n195# a_n1008_n140# 0.01fF
C108 a_296_n195# a_118_n195# 0.10fF
C109 a_n416_n195# a_n238_n195# 0.10fF
C110 a_n118_n140# a_238_n140# 0.03fF
C111 a_296_n195# a_n594_n195# 0.01fF
C112 a_n652_n140# a_416_n140# 0.01fF
C113 a_416_n140# a_830_n195# 0.02fF
C114 a_n830_n140# a_n474_n140# 0.03fF
C115 a_n1008_n140# a_118_n195# 0.01fF
C116 a_238_n140# a_n1008_n140# 0.01fF
C117 a_772_n140# VSUBS 0.01fF
C118 a_594_n140# VSUBS 0.01fF
C119 a_416_n140# VSUBS 0.02fF
C120 a_238_n140# VSUBS 0.02fF
C121 a_60_n140# VSUBS 0.02fF
C122 a_n118_n140# VSUBS 0.02fF
C123 a_n296_n140# VSUBS 0.02fF
C124 a_n474_n140# VSUBS 0.02fF
C125 a_n652_n140# VSUBS 0.02fF
C126 a_n830_n140# VSUBS 0.02fF
C127 a_830_n195# VSUBS 0.31fF
C128 a_652_n195# VSUBS 0.19fF
C129 a_474_n195# VSUBS 0.20fF
C130 a_296_n195# VSUBS 0.21fF
C131 a_118_n195# VSUBS 0.22fF
C132 a_n60_n195# VSUBS 0.23fF
C133 a_n238_n195# VSUBS 0.23fF
C134 a_n416_n195# VSUBS 0.24fF
C135 a_n594_n195# VSUBS 0.24fF
C136 a_n772_n195# VSUBS 0.24fF
C137 a_n1008_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_SD55Q9 a_352_607# a_232_552# a_644_607# a_174_607#
+ a_60_607# a_n232_n389# a_466_607# a_524_552# a_n524_n389# a_n410_n887# a_n702_n887#
+ a_n994_n887# a_644_n389# a_352_n389# a_524_54# a_60_n389# a_n60_54# a_n352_54# a_n232_n887#
+ a_n352_n444# a_n524_n887# a_174_n389# a_n60_n444# a_n644_n444# a_466_n389# a_644_n887#
+ a_352_n887# a_n118_n389# a_60_n887# a_n352_n942# a_174_n887# a_n60_n942# a_n644_n942#
+ a_232_n444# a_466_n887# a_n118_n887# a_524_n444# a_n118_109# a_n410_109# a_n644_54#
+ a_758_n887# a_n232_109# a_n702_109# a_n524_109# a_n352_552# a_352_109# a_232_54#
+ a_n644_552# a_644_109# a_174_109# a_60_109# a_n60_552# a_232_n942# a_466_109# a_n410_607#
+ a_524_n942# a_n410_n389# a_n118_607# a_n702_n389# a_n232_607# a_n702_607# a_n524_607#
+ VSUBS
X0 a_60_n389# a_n60_n444# a_n118_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_644_n887# a_524_n942# a_466_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_644_607# a_524_552# a_466_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n524_607# a_n644_552# a_n702_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_352_n389# a_232_n444# a_174_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_644_n389# a_524_n444# a_466_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n232_n887# a_n352_n942# a_n410_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_644_109# a_524_54# a_466_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n524_n887# a_n644_n942# a_n702_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_352_607# a_232_552# a_174_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n524_109# a_n644_54# a_n702_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n232_607# a_n352_552# a_n410_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n232_n389# a_n352_n444# a_n410_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n524_n389# a_n644_n444# a_n702_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_60_607# a_n60_552# a_n118_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_352_109# a_232_54# a_174_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n232_109# a_n352_54# a_n410_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_60_n887# a_n60_n942# a_n118_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_60_109# a_n60_54# a_n118_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_352_n887# a_232_n942# a_174_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n410_109# a_n410_607# 0.01fF
C1 a_n232_109# a_n524_109# 0.07fF
C2 a_n702_n887# a_352_n887# 0.02fF
C3 a_466_109# a_60_109# 0.05fF
C4 a_352_n389# a_n118_n389# 0.04fF
C5 a_n524_607# a_466_607# 0.02fF
C6 a_n118_n389# a_n118_607# 0.00fF
C7 a_n410_n389# a_60_n389# 0.04fF
C8 a_644_n887# a_n118_n887# 0.03fF
C9 a_174_109# a_n118_109# 0.07fF
C10 a_n232_109# a_n410_109# 0.13fF
C11 a_758_n887# a_n232_n389# 0.04fF
C12 a_758_n887# a_60_n887# 0.05fF
C13 a_n994_n887# a_232_n444# 0.01fF
C14 a_466_109# a_644_109# 0.13fF
C15 a_n702_109# a_758_n887# 0.02fF
C16 a_n524_607# a_n702_607# 0.13fF
C17 a_n524_n389# a_n410_n389# 0.25fF
C18 a_n524_n887# a_644_n887# 0.02fF
C19 a_n410_n887# a_352_n887# 0.03fF
C20 a_524_n444# a_n644_n444# 0.01fF
C21 a_644_n887# a_644_607# 0.00fF
C22 a_n352_n942# a_524_n942# 0.01fF
C23 a_232_54# a_524_54# 0.04fF
C24 a_n524_607# a_n410_607# 0.25fF
C25 a_644_n887# a_644_109# 0.00fF
C26 a_466_607# a_n702_607# 0.02fF
C27 a_n644_n942# a_758_n887# 0.01fF
C28 a_644_n887# a_n232_n887# 0.02fF
C29 a_174_607# a_174_n389# 0.00fF
C30 a_n644_n942# a_n644_54# 0.03fF
C31 a_n702_n389# a_n702_607# 0.00fF
C32 a_n118_109# a_n994_n887# 0.05fF
C33 a_n352_54# a_n60_54# 0.04fF
C34 a_n352_54# a_n994_n887# 0.02fF
C35 a_n524_607# a_n232_607# 0.07fF
C36 a_352_n887# a_60_n887# 0.07fF
C37 a_n410_607# a_466_607# 0.02fF
C38 a_n994_n887# a_466_n887# 0.03fF
C39 a_644_n389# a_n410_n389# 0.02fF
C40 a_60_n389# a_60_109# 0.01fF
C41 a_n524_n887# a_n524_n389# 0.01fF
C42 a_758_n887# a_524_54# 0.05fF
C43 a_n410_607# a_n702_607# 0.07fF
C44 a_n644_54# a_524_54# 0.01fF
C45 a_758_n887# a_524_n444# 0.06fF
C46 a_n644_n942# a_n60_n942# 0.02fF
C47 a_758_n887# a_n524_109# 0.03fF
C48 a_n232_607# a_466_607# 0.03fF
C49 a_352_n389# a_n994_n887# 0.03fF
C50 a_n994_n887# a_n118_607# 0.05fF
C51 a_466_n389# a_n118_n389# 0.03fF
C52 a_n410_n389# a_174_n389# 0.03fF
C53 a_174_109# a_466_109# 0.07fF
C54 a_n232_607# a_n702_607# 0.04fF
C55 a_758_n887# a_n410_109# 0.03fF
C56 a_n410_n389# a_n410_n887# 0.01fF
C57 a_n60_n444# a_n644_n444# 0.02fF
C58 a_n524_607# a_60_607# 0.03fF
C59 a_n702_109# a_352_109# 0.02fF
C60 a_n994_n887# a_n352_n444# 0.02fF
C61 a_n232_607# a_n410_607# 0.13fF
C62 a_n118_n389# a_60_n389# 0.13fF
C63 a_n702_n887# a_n118_n887# 0.03fF
C64 a_n702_n887# a_n524_n887# 0.13fF
C65 a_n524_n389# a_n118_n389# 0.05fF
C66 a_n410_n389# a_n232_n389# 0.13fF
C67 a_466_109# a_n994_n887# 0.03fF
C68 a_n994_n887# a_n352_n942# 0.02fF
C69 a_n232_109# a_n232_607# 0.01fF
C70 a_60_607# a_466_607# 0.05fF
C71 a_n524_607# a_758_n887# 0.03fF
C72 a_644_n389# a_644_607# 0.00fF
C73 a_n644_552# a_n644_n942# 0.01fF
C74 a_n410_n887# a_n118_n887# 0.07fF
C75 a_60_607# a_n702_607# 0.03fF
C76 a_644_n389# a_644_109# 0.01fF
C77 a_758_n887# a_n60_n444# 0.01fF
C78 a_n524_n887# a_n410_n887# 0.25fF
C79 a_n702_n887# a_n232_n887# 0.04fF
C80 a_n994_n887# a_644_n887# 0.02fF
C81 a_758_n887# a_466_607# 0.12fF
C82 a_758_n887# a_n702_n389# 0.02fF
C83 a_232_n444# a_n352_n444# 0.02fF
C84 a_n644_n942# a_232_n942# 0.01fF
C85 a_60_607# a_n410_607# 0.04fF
C86 a_466_n389# a_n994_n887# 0.03fF
C87 a_n118_109# a_n118_607# 0.01fF
C88 a_758_n887# a_n702_607# 0.02fF
C89 a_n118_n887# a_60_n887# 0.13fF
C90 a_n410_n887# a_n232_n887# 0.13fF
C91 a_352_109# a_n524_109# 0.02fF
C92 a_644_n389# a_n118_n389# 0.03fF
C93 a_n524_n887# a_60_n887# 0.03fF
C94 a_n60_n942# a_n60_n444# 0.15fF
C95 a_n524_607# a_352_607# 0.02fF
C96 a_60_607# a_n232_607# 0.07fF
C97 a_n410_109# a_352_109# 0.03fF
C98 a_60_n887# a_60_109# 0.00fF
C99 a_758_n887# a_n410_607# 0.03fF
C100 a_n702_109# a_60_109# 0.03fF
C101 a_n994_n887# a_60_n389# 0.04fF
C102 a_174_607# a_n524_607# 0.03fF
C103 a_n118_n389# a_174_n389# 0.07fF
C104 a_n352_54# a_n352_n444# 0.15fF
C105 a_n232_n389# a_n232_n887# 0.01fF
C106 a_352_607# a_466_607# 0.25fF
C107 a_n702_109# a_644_109# 0.01fF
C108 a_n232_n887# a_60_n887# 0.07fF
C109 a_n994_n887# a_n524_n389# 0.12fF
C110 a_n410_n389# a_n410_109# 0.01fF
C111 a_758_n887# a_n232_109# 0.04fF
C112 a_n118_109# a_466_109# 0.03fF
C113 a_758_n887# a_n232_607# 0.04fF
C114 a_352_607# a_n702_607# 0.02fF
C115 a_n352_54# a_n352_n942# 0.03fF
C116 a_174_607# a_466_607# 0.07fF
C117 a_n60_552# a_n60_n444# 0.03fF
C118 a_466_109# a_466_n887# 0.00fF
C119 a_n232_n389# a_n118_n389# 0.25fF
C120 a_174_607# a_n702_607# 0.02fF
C121 a_352_607# a_n410_607# 0.03fF
C122 a_758_n887# a_n644_n444# 0.01fF
C123 a_n644_54# a_n644_n444# 0.15fF
C124 a_n524_n887# a_n524_109# 0.00fF
C125 a_174_109# a_174_n389# 0.01fF
C126 a_n644_n942# a_524_n942# 0.01fF
C127 a_758_n887# a_174_n887# 0.06fF
C128 a_758_n887# a_232_54# 0.02fF
C129 a_n644_54# a_232_54# 0.01fF
C130 a_174_607# a_n410_607# 0.03fF
C131 a_n524_109# a_60_109# 0.03fF
C132 a_644_n389# a_n994_n887# 0.02fF
C133 a_n232_607# a_352_607# 0.03fF
C134 a_466_n887# a_644_n887# 0.13fF
C135 a_n702_n887# a_n994_n887# 0.33fF
C136 a_758_n887# a_60_607# 0.05fF
C137 a_644_109# a_n524_109# 0.02fF
C138 a_n410_109# a_60_109# 0.04fF
C139 a_466_n389# a_466_n887# 0.01fF
C140 a_n410_n389# a_n702_n389# 0.07fF
C141 a_n352_n942# a_n352_n444# 0.15fF
C142 a_174_607# a_n232_607# 0.05fF
C143 a_524_n942# a_524_54# 0.03fF
C144 a_n994_n887# a_174_n389# 0.04fF
C145 a_n410_109# a_644_109# 0.02fF
C146 a_524_n444# a_524_n942# 0.15fF
C147 a_n702_109# a_174_109# 0.02fF
C148 a_n994_n887# a_n410_n887# 0.08fF
C149 a_524_54# a_524_552# 0.15fF
C150 a_232_552# a_232_54# 0.15fF
C151 a_524_n444# a_524_552# 0.03fF
C152 a_352_n389# a_466_n389# 0.25fF
C153 a_758_n887# a_n644_54# 0.01fF
C154 a_174_n887# a_352_n887# 0.13fF
C155 a_n524_607# a_n524_n887# 0.00fF
C156 a_n232_109# a_352_109# 0.03fF
C157 a_n410_n389# a_n410_607# 0.00fF
C158 a_60_607# a_352_607# 0.07fF
C159 a_174_607# a_174_n887# 0.00fF
C160 a_n524_607# a_644_607# 0.02fF
C161 a_n994_n887# a_n232_n389# 0.06fF
C162 a_n994_n887# a_60_n887# 0.04fF
C163 a_352_n389# a_60_n389# 0.07fF
C164 a_n702_109# a_n994_n887# 0.33fF
C165 a_758_n887# a_232_552# 0.02fF
C166 a_758_n887# a_n60_n942# 0.01fF
C167 a_174_607# a_60_607# 0.25fF
C168 a_352_n389# a_n524_n389# 0.02fF
C169 a_466_n389# a_466_109# 0.01fF
C170 a_758_n887# a_352_n887# 0.08fF
C171 a_758_n887# a_352_607# 0.08fF
C172 a_466_607# a_644_607# 0.13fF
C173 a_n644_552# a_n644_n444# 0.03fF
C174 a_n644_n942# a_n994_n887# 0.05fF
C175 a_174_109# a_n524_109# 0.03fF
C176 a_644_607# a_n702_607# 0.01fF
C177 a_174_607# a_758_n887# 0.06fF
C178 a_174_109# a_n410_109# 0.03fF
C179 a_n702_n887# a_466_n887# 0.02fF
C180 a_n60_54# a_524_54# 0.02fF
C181 a_758_n887# a_n60_552# 0.01fF
C182 a_n410_607# a_644_607# 0.02fF
C183 a_232_54# a_232_n942# 0.03fF
C184 a_n994_n887# a_524_54# 0.01fF
C185 a_n994_n887# a_524_n444# 0.01fF
C186 a_644_n389# a_352_n389# 0.07fF
C187 a_758_n887# a_n352_552# 0.01fF
C188 a_n994_n887# a_n524_109# 0.12fF
C189 a_352_607# a_352_n887# 0.00fF
C190 a_n702_n389# a_n118_n389# 0.03fF
C191 a_758_n887# a_352_109# 0.08fF
C192 a_n232_109# a_60_109# 0.07fF
C193 a_n644_552# a_758_n887# 0.01fF
C194 a_n644_552# a_n644_54# 0.15fF
C195 a_466_n887# a_n410_n887# 0.02fF
C196 a_n232_607# a_644_607# 0.02fF
C197 a_n232_109# a_644_109# 0.02fF
C198 a_n994_n887# a_n410_109# 0.08fF
C199 a_n232_109# a_n232_n887# 0.00fF
C200 a_174_607# a_352_607# 0.13fF
C201 a_n702_109# a_n118_109# 0.03fF
C202 a_352_n389# a_174_n389# 0.13fF
C203 a_466_n389# a_60_n389# 0.05fF
C204 a_758_n887# a_n410_n389# 0.03fF
C205 a_n232_607# a_n232_n887# 0.00fF
C206 a_232_552# a_n60_552# 0.04fF
C207 a_n60_n942# a_n60_552# 0.01fF
C208 a_174_n887# a_n118_n887# 0.07fF
C209 a_758_n887# a_232_n942# 0.02fF
C210 a_466_n389# a_n524_n389# 0.02fF
C211 a_232_552# a_n352_552# 0.02fF
C212 a_n524_n887# a_174_n887# 0.03fF
C213 a_466_n887# a_60_n887# 0.05fF
C214 a_n644_552# a_232_552# 0.01fF
C215 a_352_n887# a_352_109# 0.00fF
C216 a_524_n444# a_232_n444# 0.04fF
C217 a_352_607# a_352_109# 0.01fF
C218 a_352_n389# a_n232_n389# 0.03fF
C219 a_n524_607# a_n994_n887# 0.12fF
C220 a_n524_n389# a_60_n389# 0.03fF
C221 a_60_607# a_60_109# 0.01fF
C222 a_n232_n887# a_174_n887# 0.05fF
C223 a_n60_54# a_n60_n444# 0.15fF
C224 a_60_607# a_644_607# 0.03fF
C225 a_232_552# a_232_n942# 0.01fF
C226 a_n60_n942# a_232_n942# 0.04fF
C227 a_n994_n887# a_n60_n444# 0.01fF
C228 a_758_n887# a_n118_n887# 0.04fF
C229 a_644_n389# a_644_n887# 0.01fF
C230 a_n702_n887# a_644_n887# 0.01fF
C231 a_758_n887# a_n524_n887# 0.03fF
C232 a_n352_552# a_n60_552# 0.04fF
C233 a_n994_n887# a_466_607# 0.03fF
C234 a_n118_109# a_n524_109# 0.05fF
C235 a_n994_n887# a_n702_n389# 0.33fF
C236 a_644_n389# a_466_n389# 0.13fF
C237 a_n352_54# a_524_54# 0.01fF
C238 a_n644_552# a_n60_552# 0.02fF
C239 a_758_n887# a_60_109# 0.05fF
C240 a_758_n887# a_644_607# 0.33fF
C241 a_n994_n887# a_n702_607# 0.33fF
C242 a_174_109# a_n232_109# 0.05fF
C243 a_644_n887# a_n410_n887# 0.02fF
C244 a_n644_552# a_n352_552# 0.04fF
C245 a_758_n887# a_644_109# 0.33fF
C246 a_n118_109# a_n410_109# 0.07fF
C247 a_758_n887# a_n232_n887# 0.04fF
C248 a_n702_109# a_466_109# 0.02fF
C249 a_466_n389# a_174_n389# 0.07fF
C250 a_352_n887# a_n118_n887# 0.04fF
C251 a_644_n389# a_60_n389# 0.03fF
C252 a_n994_n887# a_n410_607# 0.08fF
C253 a_758_n887# a_524_n942# 0.05fF
C254 a_n60_n444# a_232_n444# 0.04fF
C255 a_n524_n887# a_352_n887# 0.02fF
C256 a_644_n389# a_n524_n389# 0.02fF
C257 a_758_n887# a_524_552# 0.05fF
C258 a_644_n887# a_60_n887# 0.03fF
C259 a_n232_109# a_n994_n887# 0.06fF
C260 a_n644_n942# a_n352_n942# 0.04fF
C261 a_758_n887# a_n118_n389# 0.04fF
C262 a_60_n389# a_174_n389# 0.25fF
C263 a_n994_n887# a_n232_607# 0.06fF
C264 a_352_607# a_644_607# 0.07fF
C265 a_174_109# a_174_n887# 0.00fF
C266 a_466_n389# a_n232_n389# 0.03fF
C267 a_n524_n389# a_174_n389# 0.03fF
C268 a_n232_n887# a_352_n887# 0.03fF
C269 a_524_n444# a_n352_n444# 0.01fF
C270 a_n60_n942# a_524_n942# 0.02fF
C271 a_174_607# a_644_607# 0.04fF
C272 a_232_552# a_524_552# 0.04fF
C273 a_n994_n887# a_n644_n444# 0.05fF
C274 a_n60_54# a_232_54# 0.04fF
C275 a_466_109# a_n524_109# 0.02fF
C276 a_n232_n389# a_60_n389# 0.07fF
C277 a_60_n389# a_60_n887# 0.01fF
C278 a_n994_n887# a_174_n887# 0.04fF
C279 a_n994_n887# a_232_54# 0.01fF
C280 a_758_n887# a_174_109# 0.06fF
C281 a_n524_n389# a_n232_n389# 0.07fF
C282 a_n524_607# a_n118_607# 0.05fF
C283 a_352_109# a_60_109# 0.07fF
C284 a_466_109# a_n410_109# 0.02fF
C285 a_60_607# a_n994_n887# 0.04fF
C286 a_466_n887# a_466_607# 0.00fF
C287 a_644_109# a_352_109# 0.07fF
C288 a_644_n389# a_174_n389# 0.04fF
C289 a_n60_552# a_524_552# 0.02fF
C290 a_n702_n887# a_n410_n887# 0.07fF
C291 a_466_607# a_n118_607# 0.03fF
C292 a_352_n389# a_n702_n389# 0.02fF
C293 a_758_n887# a_n60_54# 0.01fF
C294 a_n60_54# a_n644_54# 0.02fF
C295 a_758_n887# a_n994_n887# 0.07fF
C296 a_n232_109# a_n118_109# 0.25fF
C297 a_n352_552# a_524_552# 0.01fF
C298 a_n644_54# a_n994_n887# 0.05fF
C299 a_n60_n444# a_n352_n444# 0.04fF
C300 a_232_n444# a_n644_n444# 0.01fF
C301 a_n118_607# a_n702_607# 0.03fF
C302 a_n644_552# a_524_552# 0.01fF
C303 a_232_54# a_232_n444# 0.15fF
C304 a_644_n389# a_n232_n389# 0.02fF
C305 a_n702_n887# a_60_n887# 0.03fF
C306 a_n524_n887# a_n118_n887# 0.05fF
C307 a_n702_109# a_n702_n887# 0.00fF
C308 a_n410_607# a_n118_607# 0.07fF
C309 a_232_n942# a_524_n942# 0.04fF
C310 a_n60_54# a_n60_n942# 0.03fF
C311 a_174_607# a_174_109# 0.01fF
C312 a_n410_n389# a_n118_n389# 0.07fF
C313 a_n524_n389# a_n524_109# 0.01fF
C314 a_466_109# a_466_607# 0.01fF
C315 a_232_552# a_n994_n887# 0.01fF
C316 a_n994_n887# a_n60_n942# 0.01fF
C317 a_n232_n389# a_174_n389# 0.05fF
C318 a_n994_n887# a_352_n887# 0.03fF
C319 a_n232_n887# a_n118_n887# 0.25fF
C320 a_n232_607# a_n118_607# 0.25fF
C321 a_n994_n887# a_352_607# 0.03fF
C322 a_n410_n887# a_60_n887# 0.04fF
C323 a_n352_54# a_232_54# 0.02fF
C324 a_758_n887# a_232_n444# 0.02fF
C325 a_n524_n887# a_n232_n887# 0.07fF
C326 a_174_109# a_352_109# 0.13fF
C327 a_644_109# a_60_109# 0.03fF
C328 a_174_607# a_n994_n887# 0.04fF
C329 a_466_n887# a_174_n887# 0.07fF
C330 a_644_109# a_644_607# 0.01fF
C331 a_n60_54# a_n60_552# 0.15fF
C332 a_466_n389# a_466_607# 0.00fF
C333 a_466_n389# a_n702_n389# 0.02fF
C334 a_n118_n389# a_n118_n887# 0.01fF
C335 a_n994_n887# a_n60_552# 0.01fF
C336 a_758_n887# a_n118_109# 0.04fF
C337 a_n232_109# a_466_109# 0.03fF
C338 a_232_552# a_232_n444# 0.03fF
C339 a_n524_607# a_n524_n389# 0.00fF
C340 a_n352_552# a_n994_n887# 0.02fF
C341 a_n352_54# a_758_n887# 0.01fF
C342 a_n352_54# a_n644_54# 0.04fF
C343 a_n994_n887# a_352_109# 0.03fF
C344 a_60_607# a_n118_607# 0.13fF
C345 a_n644_552# a_n994_n887# 0.05fF
C346 a_n644_n444# a_n352_n444# 0.04fF
C347 a_n702_n389# a_60_n389# 0.03fF
C348 a_758_n887# a_466_n887# 0.12fF
C349 a_n994_n887# a_n410_n389# 0.08fF
C350 a_n524_n389# a_n702_n389# 0.13fF
C351 a_524_n942# a_524_552# 0.01fF
C352 a_n994_n887# a_232_n942# 0.01fF
C353 a_758_n887# a_352_n389# 0.08fF
C354 a_758_n887# a_n118_607# 0.04fF
C355 a_n410_109# a_n410_n887# 0.00fF
C356 a_174_109# a_60_109# 0.25fF
C357 a_n702_109# a_n524_109# 0.13fF
C358 a_758_n887# a_n352_n444# 0.01fF
C359 a_644_n887# a_174_n887# 0.04fF
C360 a_466_n887# a_352_n887# 0.25fF
C361 a_174_109# a_644_109# 0.04fF
C362 a_n994_n887# a_n118_n887# 0.05fF
C363 a_n702_109# a_n410_109# 0.07fF
C364 a_758_n887# a_466_109# 0.12fF
C365 a_352_n389# a_352_n887# 0.01fF
C366 a_758_n887# a_n352_n942# 0.01fF
C367 a_n524_n887# a_n994_n887# 0.12fF
C368 a_644_n389# a_n702_n389# 0.01fF
C369 a_352_n389# a_352_607# 0.00fF
C370 a_n702_n887# a_n702_n389# 0.01fF
C371 a_352_607# a_n118_607# 0.04fF
C372 a_232_n942# a_232_n444# 0.15fF
C373 a_n118_109# a_352_109# 0.04fF
C374 a_n994_n887# a_60_109# 0.04fF
C375 a_n702_n887# a_n702_607# 0.00fF
C376 a_n352_54# a_n352_552# 0.15fF
C377 a_n994_n887# a_644_607# 0.02fF
C378 a_174_607# a_n118_607# 0.07fF
C379 a_n994_n887# a_644_109# 0.02fF
C380 a_n702_n389# a_174_n389# 0.02fF
C381 a_758_n887# a_644_n887# 0.33fF
C382 a_n994_n887# a_n232_n887# 0.06fF
C383 a_524_n444# a_524_54# 0.15fF
C384 a_n352_n942# a_n60_n942# 0.04fF
C385 a_60_607# a_60_n389# 0.00fF
C386 a_758_n887# a_466_n389# 0.12fF
C387 a_n994_n887# a_524_n942# 0.01fF
C388 a_n994_n887# a_524_552# 0.01fF
C389 a_352_n389# a_352_109# 0.01fF
C390 a_n994_n887# a_n118_n389# 0.05fF
C391 a_n410_109# a_n524_109# 0.25fF
C392 a_n410_n887# a_n410_607# 0.00fF
C393 a_n702_n389# a_n232_n389# 0.04fF
C394 a_n702_109# a_n702_n389# 0.01fF
C395 a_758_n887# a_60_n389# 0.05fF
C396 a_352_n389# a_n410_n389# 0.03fF
C397 a_644_n887# a_352_n887# 0.07fF
C398 a_n352_552# a_n352_n444# 0.03fF
C399 a_n702_109# a_n702_607# 0.01fF
C400 a_n118_109# a_n118_n887# 0.00fF
C401 a_758_n887# a_n524_n389# 0.03fF
C402 a_n352_552# a_n352_n942# 0.01fF
C403 a_n702_n887# a_174_n887# 0.02fF
C404 a_466_109# a_352_109# 0.25fF
C405 a_n118_109# a_60_109# 0.13fF
C406 a_466_n887# a_n118_n887# 0.03fF
C407 a_n524_607# a_n524_109# 0.01fF
C408 a_174_109# a_n994_n887# 0.04fF
C409 a_n118_109# a_644_109# 0.03fF
C410 a_n232_109# a_n232_n389# 0.01fF
C411 a_524_n444# a_n60_n444# 0.02fF
C412 a_n524_n887# a_466_n887# 0.02fF
C413 a_n702_109# a_n232_109# 0.04fF
C414 a_n232_607# a_n232_n389# 0.00fF
C415 a_174_n887# a_174_n389# 0.01fF
C416 a_n410_n887# a_174_n887# 0.03fF
C417 a_n118_n887# a_n118_607# 0.00fF
C418 a_n352_n942# a_232_n942# 0.02fF
C419 a_644_n389# a_758_n887# 0.33fF
C420 a_n60_54# a_n994_n887# 0.01fF
C421 a_466_n887# a_n232_n887# 0.03fF
C422 a_758_n887# a_n702_n887# 0.02fF
C423 a_644_607# a_n118_607# 0.03fF
C424 a_n118_109# a_n118_n389# 0.01fF
C425 a_174_n887# a_60_n887# 0.25fF
C426 a_758_n887# a_174_n389# 0.06fF
C427 a_466_n389# a_n410_n389# 0.02fF
C428 a_758_n887# a_n410_n887# 0.03fF
C429 a_60_607# a_60_n887# 0.00fF
C430 a_n644_n942# a_n644_n444# 0.15fF
C431 a_644_n887# VSUBS 0.01fF
C432 a_466_n887# VSUBS 0.01fF
C433 a_352_n887# VSUBS 0.01fF
C434 a_174_n887# VSUBS 0.01fF
C435 a_60_n887# VSUBS 0.01fF
C436 a_n118_n887# VSUBS 0.01fF
C437 a_n232_n887# VSUBS 0.01fF
C438 a_n410_n887# VSUBS 0.01fF
C439 a_n524_n887# VSUBS 0.01fF
C440 a_n702_n887# VSUBS 0.01fF
C441 a_524_n942# VSUBS 0.17fF
C442 a_232_n942# VSUBS 0.19fF
C443 a_n60_n942# VSUBS 0.20fF
C444 a_n352_n942# VSUBS 0.21fF
C445 a_n644_n942# VSUBS 0.22fF
C446 a_644_n389# VSUBS 0.01fF
C447 a_466_n389# VSUBS 0.01fF
C448 a_352_n389# VSUBS 0.01fF
C449 a_174_n389# VSUBS 0.01fF
C450 a_60_n389# VSUBS 0.01fF
C451 a_n118_n389# VSUBS 0.01fF
C452 a_n232_n389# VSUBS 0.01fF
C453 a_n410_n389# VSUBS 0.01fF
C454 a_n524_n389# VSUBS 0.01fF
C455 a_n702_n389# VSUBS 0.01fF
C456 a_524_n444# VSUBS 0.16fF
C457 a_232_n444# VSUBS 0.17fF
C458 a_n60_n444# VSUBS 0.18fF
C459 a_n352_n444# VSUBS 0.19fF
C460 a_n644_n444# VSUBS 0.20fF
C461 a_644_109# VSUBS 0.01fF
C462 a_466_109# VSUBS 0.01fF
C463 a_352_109# VSUBS 0.01fF
C464 a_174_109# VSUBS 0.01fF
C465 a_60_109# VSUBS 0.01fF
C466 a_n118_109# VSUBS 0.01fF
C467 a_n232_109# VSUBS 0.01fF
C468 a_n410_109# VSUBS 0.01fF
C469 a_n524_109# VSUBS 0.01fF
C470 a_n702_109# VSUBS 0.01fF
C471 a_524_54# VSUBS 0.17fF
C472 a_232_54# VSUBS 0.18fF
C473 a_n60_54# VSUBS 0.19fF
C474 a_n352_54# VSUBS 0.20fF
C475 a_n644_54# VSUBS 0.21fF
C476 a_644_607# VSUBS 0.02fF
C477 a_466_607# VSUBS 0.02fF
C478 a_352_607# VSUBS 0.02fF
C479 a_174_607# VSUBS 0.02fF
C480 a_60_607# VSUBS 0.02fF
C481 a_n118_607# VSUBS 0.02fF
C482 a_n232_607# VSUBS 0.02fF
C483 a_n410_607# VSUBS 0.02fF
C484 a_n524_607# VSUBS 0.02fF
C485 a_n702_607# VSUBS 0.02fF
C486 a_758_n887# VSUBS 1.42fF
C487 a_524_552# VSUBS 0.20fF
C488 a_232_552# VSUBS 0.22fF
C489 a_n60_552# VSUBS 0.23fF
C490 a_n352_552# VSUBS 0.24fF
C491 a_n644_552# VSUBS 0.25fF
C492 a_n994_n887# VSUBS 1.65fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EZNTQN a_n830_109# a_n772_54# a_118_552# a_n652_n887#
+ a_n772_n444# a_n652_109# a_594_n389# a_60_607# a_772_n887# a_n474_109# a_n772_552#
+ a_772_109# a_n296_109# a_n594_552# a_118_n942# a_n296_n389# a_594_109# a_n594_54#
+ a_n474_n887# a_60_n389# a_n594_n444# a_n60_54# a_n830_607# a_n772_n942# a_416_n389#
+ a_652_n444# a_n416_54# a_n652_607# a_594_n887# a_n474_607# a_n60_n444# a_772_607#
+ a_n296_607# a_594_607# a_652_552# a_n296_n887# a_n118_n389# a_n238_54# a_474_552#
+ a_60_n887# a_n594_n942# a_n416_n444# a_238_n389# a_474_n444# a_296_552# a_416_n887#
+ a_652_n942# a_652_54# a_n830_n389# a_n60_n942# a_n118_n887# a_n238_n444# a_n118_109#
+ a_n416_552# a_296_n444# a_416_109# a_474_54# a_n416_n942# a_238_109# a_n238_552#
+ a_238_n887# a_474_n942# a_n1110_n1061# a_n652_n389# a_n830_n887# a_60_109# a_772_n389#
+ a_296_54# a_n60_552# a_n238_n942# a_n118_607# a_296_n942# a_118_n444# a_416_607#
+ a_n474_n389# a_118_54# a_238_607#
X0 a_n652_109# a_n772_54# a_n830_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_60_n389# a_n60_n444# a_n118_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_594_n389# a_474_n444# a_416_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1110_n1061# a_n1110_n1061# a_772_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n830_n887# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n474_n887# a_n594_n942# a_n652_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_594_607# a_474_552# a_416_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_109# a_n416_54# a_n474_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_416_n887# a_296_n942# a_238_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n474_607# a_n594_552# a_n652_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n296_n887# a_n416_n942# a_n474_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1110_n1061# a_n1110_n1061# a_772_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1110_n1061# a_n1110_n1061# a_772_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_238_607# a_118_552# a_60_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_238_n887# a_118_n942# a_60_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n830_n389# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n474_n389# a_n594_n444# a_n652_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n830_607# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n118_607# a_n238_552# a_n296_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_594_109# a_474_54# a_416_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_416_n389# a_296_n444# a_238_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_772_n887# a_652_n942# a_594_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n474_109# a_n594_54# a_n652_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n296_n389# a_n416_n444# a_n474_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1110_n1061# a_n1110_n1061# a_772_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_238_109# a_118_54# a_60_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_238_n389# a_118_n444# a_60_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_607# a_296_552# a_238_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n830_109# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n118_109# a_n238_54# a_n296_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n118_n887# a_n238_n942# a_n296_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_60_607# a_n60_552# a_n118_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_772_n389# a_652_n444# a_594_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_772_607# a_652_552# a_594_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_n652_n887# a_n772_n942# a_n830_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_594_n887# a_474_n942# a_416_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_n652_607# a_n772_552# a_n830_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_60_n887# a_n60_n942# a_n118_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_416_109# a_296_54# a_238_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n118_n389# a_n238_n444# a_n296_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_60_109# a_n60_54# a_n118_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X41 a_n296_607# a_n416_552# a_n474_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X42 a_772_109# a_652_54# a_594_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_n652_n389# a_n772_n444# a_n830_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n238_54# a_118_54# 0.03fF
C1 a_416_607# a_60_607# 0.03fF
C2 a_n652_607# a_772_607# 0.01fF
C3 a_296_54# a_296_n942# 0.03fF
C4 a_n60_n942# a_n60_54# 0.03fF
C5 a_594_607# a_594_n887# 0.00fF
C6 a_n772_54# a_n416_54# 0.03fF
C7 a_n238_54# a_n60_54# 0.10fF
C8 a_n118_109# a_n118_607# 0.00fF
C9 a_n60_552# a_652_552# 0.01fF
C10 a_594_607# a_416_607# 0.06fF
C11 a_n594_n444# a_n416_n444# 0.10fF
C12 a_n474_607# a_238_607# 0.01fF
C13 a_n60_n942# a_n594_n942# 0.02fF
C14 a_652_54# a_474_54# 0.10fF
C15 a_n296_n887# a_238_n887# 0.02fF
C16 a_n830_n389# a_n296_n389# 0.02fF
C17 a_296_552# a_296_n444# 0.03fF
C18 a_n594_n444# a_n772_n444# 0.10fF
C19 a_652_54# a_118_54# 0.02fF
C20 a_n772_54# a_n772_n942# 0.03fF
C21 a_n118_n887# a_n830_n887# 0.01fF
C22 a_n652_109# a_n830_109# 0.06fF
C23 a_416_n389# a_n474_n389# 0.01fF
C24 a_652_552# a_n594_552# 0.01fF
C25 a_238_n389# a_n830_n389# 0.01fF
C26 a_n60_54# a_652_54# 0.01fF
C27 a_416_n389# a_416_n887# 0.00fF
C28 a_n118_n887# a_n118_607# 0.00fF
C29 a_772_n887# a_594_n887# 0.06fF
C30 a_118_n942# a_n772_n942# 0.01fF
C31 a_n118_n887# a_n118_109# 0.00fF
C32 a_n772_n444# a_n416_n444# 0.03fF
C33 a_n652_n887# a_60_n887# 0.01fF
C34 a_296_552# a_n60_552# 0.03fF
C35 a_n830_109# a_594_109# 0.01fF
C36 a_n238_552# a_n60_552# 0.10fF
C37 a_n474_109# a_n474_607# 0.00fF
C38 a_474_n942# a_n772_n942# 0.01fF
C39 a_772_109# a_n118_109# 0.01fF
C40 a_n416_n942# a_n594_n942# 0.10fF
C41 a_474_552# a_474_n942# 0.01fF
C42 a_n296_n389# a_n296_607# 0.00fF
C43 a_n652_607# a_416_607# 0.01fF
C44 a_296_54# a_296_n444# 0.15fF
C45 a_n118_607# a_238_607# 0.03fF
C46 a_n60_552# a_n416_552# 0.03fF
C47 a_n652_n389# a_60_n389# 0.01fF
C48 a_n830_607# a_772_607# 0.01fF
C49 a_n594_n942# a_296_n942# 0.01fF
C50 a_n830_n389# a_594_n389# 0.01fF
C51 a_n474_n887# a_n474_607# 0.00fF
C52 a_296_552# a_n594_552# 0.01fF
C53 a_118_n444# a_118_54# 0.15fF
C54 a_n238_552# a_n594_552# 0.03fF
C55 a_n652_109# a_n652_n887# 0.00fF
C56 a_118_552# a_118_n942# 0.01fF
C57 a_n296_n887# a_772_n887# 0.01fF
C58 a_238_n389# a_n296_n389# 0.02fF
C59 a_n238_n942# a_118_n942# 0.03fF
C60 a_416_109# a_n118_109# 0.02fF
C61 a_n594_n444# a_n238_n444# 0.03fF
C62 a_n416_n942# a_n416_n444# 0.15fF
C63 a_n416_552# a_n594_552# 0.10fF
C64 a_n594_n942# a_652_n942# 0.01fF
C65 a_60_n887# a_238_n887# 0.06fF
C66 a_n238_n942# a_474_n942# 0.01fF
C67 a_416_n389# a_416_607# 0.00fF
C68 a_n772_n444# a_n772_552# 0.03fF
C69 a_n652_n887# a_238_n887# 0.01fF
C70 a_60_n887# a_60_607# 0.00fF
C71 a_n474_109# a_n118_109# 0.03fF
C72 a_n830_n389# a_n118_n389# 0.01fF
C73 a_n416_n942# a_n60_n942# 0.03fF
C74 a_474_n444# a_474_54# 0.15fF
C75 a_n296_607# a_60_607# 0.03fF
C76 a_n474_607# a_n474_n389# 0.00fF
C77 a_n238_54# a_652_54# 0.01fF
C78 a_n474_n887# a_n830_n887# 0.03fF
C79 a_n594_n444# a_118_n444# 0.01fF
C80 a_n474_607# a_772_607# 0.01fF
C81 a_n238_n444# a_n416_n444# 0.10fF
C82 a_n652_109# a_594_109# 0.01fF
C83 a_594_607# a_n296_607# 0.01fF
C84 a_n652_n389# a_772_n389# 0.01fF
C85 a_238_n389# a_238_n887# 0.00fF
C86 a_416_109# a_772_109# 0.03fF
C87 a_n296_n389# a_594_n389# 0.01fF
C88 a_n60_n942# a_296_n942# 0.03fF
C89 a_n238_n444# a_n772_n444# 0.02fF
C90 a_296_54# a_n594_54# 0.01fF
C91 a_416_607# a_n830_607# 0.01fF
C92 a_238_n389# a_594_n389# 0.03fF
C93 a_60_109# a_n118_109# 0.06fF
C94 a_118_n444# a_n416_n444# 0.02fF
C95 a_n238_n444# a_n238_54# 0.15fF
C96 a_n594_n444# a_296_n444# 0.01fF
C97 a_772_109# a_772_n389# 0.00fF
C98 a_n474_109# a_772_109# 0.01fF
C99 a_n60_54# a_n60_552# 0.15fF
C100 a_n60_n942# a_652_n942# 0.01fF
C101 a_772_n389# a_60_n389# 0.01fF
C102 a_238_109# a_n118_109# 0.03fF
C103 a_n594_n444# a_474_n444# 0.01fF
C104 a_118_n444# a_n772_n444# 0.01fF
C105 a_60_n887# a_772_n887# 0.01fF
C106 a_n830_n887# a_416_n887# 0.01fF
C107 a_652_n444# a_n594_n444# 0.01fF
C108 a_n296_n389# a_n118_n389# 0.06fF
C109 a_594_n389# a_594_109# 0.00fF
C110 a_n118_607# a_772_607# 0.01fF
C111 a_n118_n887# a_n474_n887# 0.03fF
C112 a_n416_n942# a_296_n942# 0.01fF
C113 a_n652_n887# a_772_n887# 0.01fF
C114 a_474_54# a_n594_54# 0.01fF
C115 a_474_552# a_118_552# 0.03fF
C116 a_238_n389# a_n118_n389# 0.03fF
C117 a_594_607# a_594_109# 0.00fF
C118 a_296_n444# a_n416_n444# 0.01fF
C119 a_n238_n942# a_n772_n942# 0.02fF
C120 a_118_54# a_n594_54# 0.01fF
C121 a_n652_607# a_n296_607# 0.03fF
C122 a_772_109# a_60_109# 0.01fF
C123 a_n830_n389# a_416_n389# 0.01fF
C124 a_474_n444# a_n416_n444# 0.01fF
C125 a_60_109# a_60_n389# 0.00fF
C126 a_n474_607# a_416_607# 0.01fF
C127 a_416_109# a_n474_109# 0.01fF
C128 a_n652_n389# a_n474_n389# 0.06fF
C129 a_652_n444# a_n416_n444# 0.01fF
C130 a_n652_607# a_n652_n887# 0.00fF
C131 a_652_54# a_652_n942# 0.03fF
C132 a_296_n444# a_n772_n444# 0.01fF
C133 a_n416_n942# a_652_n942# 0.01fF
C134 a_n60_54# a_n594_54# 0.02fF
C135 a_238_109# a_772_109# 0.02fF
C136 a_594_607# a_60_607# 0.02fF
C137 a_594_607# a_594_n389# 0.00fF
C138 a_n594_n942# a_n594_552# 0.01fF
C139 a_474_n444# a_n772_n444# 0.01fF
C140 a_296_54# a_n772_54# 0.01fF
C141 a_652_n444# a_n772_n444# 0.01fF
C142 a_n594_n444# a_n594_552# 0.03fF
C143 a_652_n942# a_296_n942# 0.03fF
C144 a_n652_109# a_n652_607# 0.00fF
C145 a_n594_n942# a_n594_54# 0.03fF
C146 a_n118_n887# a_416_n887# 0.02fF
C147 a_n474_n389# a_60_n389# 0.02fF
C148 a_238_109# a_238_607# 0.00fF
C149 a_772_109# a_772_607# 0.00fF
C150 a_n60_54# a_n60_n444# 0.15fF
C151 a_n830_109# a_n830_607# 0.00fF
C152 a_416_109# a_60_109# 0.03fF
C153 a_n594_n444# a_n594_54# 0.15fF
C154 a_n118_n389# a_594_n389# 0.01fF
C155 a_n830_n887# a_594_n887# 0.01fF
C156 a_238_n887# a_772_n887# 0.02fF
C157 a_n830_n389# a_n830_607# 0.00fF
C158 a_474_552# a_652_552# 0.10fF
C159 a_n60_n942# a_n60_552# 0.01fF
C160 a_n238_n444# a_118_n444# 0.03fF
C161 a_238_109# a_416_109# 0.06fF
C162 a_n474_109# a_n474_n887# 0.00fF
C163 a_416_n389# a_n296_n389# 0.01fF
C164 a_416_607# a_n118_607# 0.02fF
C165 a_772_607# a_238_607# 0.02fF
C166 a_n118_109# a_n296_109# 0.06fF
C167 a_n474_109# a_60_109# 0.02fF
C168 a_n772_54# a_474_54# 0.01fF
C169 a_n772_54# a_118_54# 0.01fF
C170 a_n594_n444# a_n60_n444# 0.02fF
C171 a_238_n389# a_416_n389# 0.06fF
C172 a_652_n444# a_652_54# 0.15fF
C173 a_n652_607# a_60_607# 0.01fF
C174 a_238_109# a_n474_109# 0.01fF
C175 a_296_n444# a_296_n942# 0.15fF
C176 a_416_109# a_416_n887# 0.00fF
C177 a_n772_54# a_n60_54# 0.01fF
C178 a_118_552# a_652_552# 0.02fF
C179 a_n830_607# a_n296_607# 0.02fF
C180 a_n416_54# a_n416_552# 0.15fF
C181 a_118_n942# a_118_54# 0.03fF
C182 a_n238_n444# a_296_n444# 0.02fF
C183 a_n60_552# a_n772_552# 0.01fF
C184 a_594_607# a_n652_607# 0.01fF
C185 a_n296_n887# a_n830_n887# 0.02fF
C186 a_474_n942# a_474_54# 0.03fF
C187 a_296_552# a_474_552# 0.10fF
C188 a_n238_n444# a_474_n444# 0.01fF
C189 a_n474_109# a_n474_n389# 0.00fF
C190 a_772_n389# a_n474_n389# 0.01fF
C191 a_n238_552# a_474_552# 0.01fF
C192 a_n238_54# a_n594_54# 0.03fF
C193 a_n60_n444# a_n416_n444# 0.03fF
C194 a_772_n389# a_772_607# 0.00fF
C195 a_652_n444# a_n238_n444# 0.01fF
C196 a_n118_n887# a_594_n887# 0.01fF
C197 a_772_109# a_n296_109# 0.01fF
C198 a_296_54# a_n416_54# 0.01fF
C199 a_238_109# a_60_109# 0.06fF
C200 a_n772_n444# a_n60_n444# 0.01fF
C201 a_118_n444# a_296_n444# 0.10fF
C202 a_652_n444# a_652_n942# 0.15fF
C203 a_474_552# a_n416_552# 0.01fF
C204 a_n772_552# a_n594_552# 0.10fF
C205 a_416_n389# a_594_n389# 0.06fF
C206 a_n594_n942# a_118_n942# 0.01fF
C207 a_n60_n942# a_n60_n444# 0.15fF
C208 a_118_n444# a_474_n444# 0.03fF
C209 a_n474_n887# a_n474_n389# 0.00fF
C210 a_652_n444# a_118_n444# 0.02fF
C211 a_296_552# a_118_552# 0.10fF
C212 a_n474_n887# a_416_n887# 0.01fF
C213 a_n830_109# a_n830_n887# 0.00fF
C214 a_n238_552# a_118_552# 0.03fF
C215 a_474_n942# a_n594_n942# 0.01fF
C216 a_652_54# a_n594_54# 0.01fF
C217 a_n474_607# a_n296_607# 0.06fF
C218 a_416_607# a_238_607# 0.06fF
C219 a_n830_n389# a_n830_n887# 0.00fF
C220 a_n238_n942# a_n238_552# 0.01fF
C221 a_416_109# a_n296_109# 0.01fF
C222 a_n296_n887# a_n118_n887# 0.06fF
C223 a_416_109# a_416_607# 0.00fF
C224 a_118_552# a_n416_552# 0.02fF
C225 a_n830_109# a_n118_109# 0.01fF
C226 a_n416_54# a_474_54# 0.01fF
C227 a_474_n444# a_296_n444# 0.10fF
C228 a_n772_54# a_n772_n444# 0.15fF
C229 a_416_n389# a_n118_n389# 0.02fF
C230 a_n830_607# a_60_607# 0.01fF
C231 a_n416_54# a_118_54# 0.02fF
C232 a_652_n444# a_296_n444# 0.03fF
C233 a_n474_109# a_n296_109# 0.06fF
C234 a_n772_54# a_n238_54# 0.02fF
C235 a_652_n444# a_474_n444# 0.10fF
C236 a_n416_54# a_n60_54# 0.03fF
C237 a_594_607# a_n830_607# 0.01fF
C238 a_n830_n887# a_60_n887# 0.01fF
C239 a_n830_n389# a_n652_n389# 0.06fF
C240 a_n60_n942# a_118_n942# 0.10fF
C241 a_296_552# a_652_552# 0.03fF
C242 a_n238_552# a_652_552# 0.01fF
C243 a_474_552# a_474_54# 0.15fF
C244 a_n652_n887# a_n830_n887# 0.06fF
C245 a_n118_607# a_n296_607# 0.06fF
C246 a_n238_n444# a_n60_n444# 0.10fF
C247 a_474_n942# a_n60_n942# 0.02fF
C248 a_n830_109# a_772_109# 0.01fF
C249 a_n474_n887# a_594_n887# 0.01fF
C250 a_60_109# a_n296_109# 0.03fF
C251 a_n772_54# a_n772_552# 0.15fF
C252 a_n416_552# a_652_552# 0.01fF
C253 a_n772_54# a_652_54# 0.01fF
C254 a_n830_n389# a_60_n389# 0.01fF
C255 a_n474_607# a_60_607# 0.02fF
C256 a_238_109# a_n296_109# 0.02fF
C257 a_118_n444# a_n60_n444# 0.10fF
C258 a_n594_n942# a_n772_n942# 0.10fF
C259 a_n416_n942# a_118_n942# 0.02fF
C260 a_594_607# a_n474_607# 0.01fF
C261 a_n652_n887# a_n652_n389# 0.00fF
C262 a_118_552# a_118_54# 0.15fF
C263 a_n652_109# a_n118_109# 0.02fF
C264 a_n118_n887# a_60_n887# 0.06fF
C265 a_n652_n389# a_n296_n389# 0.03fF
C266 a_296_552# a_n238_552# 0.02fF
C267 a_n416_54# a_n416_n444# 0.15fF
C268 a_n830_109# a_416_109# 0.01fF
C269 a_n416_n942# a_474_n942# 0.01fF
C270 a_n652_607# a_n830_607# 0.06fF
C271 a_n830_n887# a_238_n887# 0.01fF
C272 a_60_n389# a_60_n887# 0.00fF
C273 a_118_n942# a_296_n942# 0.10fF
C274 a_n60_552# a_n594_552# 0.02fF
C275 a_n296_n887# a_n474_n887# 0.06fF
C276 a_n118_n887# a_n652_n887# 0.02fF
C277 a_238_n389# a_n652_n389# 0.01fF
C278 a_416_607# a_772_607# 0.03fF
C279 a_416_n887# a_594_n887# 0.06fF
C280 a_n652_109# a_n652_n389# 0.00fF
C281 a_416_607# a_416_n887# 0.00fF
C282 a_296_552# a_n416_552# 0.01fF
C283 a_296_n444# a_n60_n444# 0.03fF
C284 a_n238_552# a_n416_552# 0.10fF
C285 a_474_n942# a_296_n942# 0.10fF
C286 a_n118_109# a_594_109# 0.01fF
C287 a_n830_109# a_n474_109# 0.03fF
C288 a_n296_n389# a_60_n389# 0.03fF
C289 a_n238_54# a_n416_54# 0.10fF
C290 a_474_n444# a_n60_n444# 0.02fF
C291 a_n830_n389# a_772_n389# 0.01fF
C292 a_n118_607# a_60_607# 0.06fF
C293 a_n296_607# a_238_607# 0.02fF
C294 a_118_n942# a_652_n942# 0.02fF
C295 a_652_n444# a_n60_n444# 0.01fF
C296 a_n238_n942# a_n594_n942# 0.03fF
C297 a_n652_109# a_772_109# 0.01fF
C298 a_238_n389# a_60_n389# 0.06fF
C299 a_n772_n444# a_n772_n942# 0.15fF
C300 a_594_607# a_n118_607# 0.01fF
C301 a_474_n942# a_652_n942# 0.10fF
C302 a_296_54# a_296_552# 0.15fF
C303 a_118_n444# a_118_n942# 0.15fF
C304 a_n60_n942# a_n772_n942# 0.01fF
C305 a_n652_607# a_n474_607# 0.06fF
C306 a_n594_552# a_n594_54# 0.15fF
C307 a_n60_552# a_n60_n444# 0.03fF
C308 a_n296_n887# a_416_n887# 0.01fF
C309 a_n652_n389# a_594_n389# 0.01fF
C310 a_238_n389# a_238_607# 0.00fF
C311 a_n830_109# a_60_109# 0.01fF
C312 a_n416_54# a_652_54# 0.01fF
C313 a_n416_54# a_n416_n942# 0.03fF
C314 a_772_109# a_594_109# 0.06fF
C315 a_n118_n887# a_238_n887# 0.03fF
C316 a_n118_607# a_n118_n389# 0.00fF
C317 a_238_109# a_n830_109# 0.01fF
C318 a_n830_n887# a_772_n887# 0.01fF
C319 a_n652_109# a_416_109# 0.01fF
C320 a_n118_109# a_n118_n389# 0.00fF
C321 a_n772_552# a_n772_n942# 0.01fF
C322 a_60_n389# a_60_607# 0.00fF
C323 a_n296_n389# a_772_n389# 0.01fF
C324 a_60_n389# a_594_n389# 0.02fF
C325 a_n416_n942# a_n772_n942# 0.03fF
C326 a_474_552# a_n772_552# 0.01fF
C327 a_238_n887# a_238_607# 0.00fF
C328 a_n474_n887# a_60_n887# 0.02fF
C329 a_n238_n942# a_n60_n942# 0.10fF
C330 a_n830_n389# a_n474_n389# 0.03fF
C331 a_n652_n389# a_n118_n389# 0.02fF
C332 a_238_n389# a_772_n389# 0.02fF
C333 a_474_n444# a_474_n942# 0.15fF
C334 a_n652_109# a_n474_109# 0.06fF
C335 a_60_109# a_60_n887# 0.00fF
C336 a_n238_n942# a_n238_54# 0.03fF
C337 a_416_109# a_594_109# 0.06fF
C338 a_n652_607# a_n118_607# 0.02fF
C339 a_n652_n887# a_n474_n887# 0.06fF
C340 a_238_607# a_60_607# 0.06fF
C341 a_296_n942# a_n772_n942# 0.01fF
C342 a_n118_n887# a_n118_n389# 0.00fF
C343 a_594_607# a_238_607# 0.03fF
C344 a_n296_n887# a_n296_109# 0.00fF
C345 a_n296_n887# a_594_n887# 0.01fF
C346 a_n474_109# a_594_109# 0.01fF
C347 a_118_552# a_n772_552# 0.01fF
C348 a_60_n389# a_n118_n389# 0.06fF
C349 a_n118_n887# a_772_n887# 0.01fF
C350 a_n652_607# a_n652_n389# 0.00fF
C351 a_652_n942# a_n772_n942# 0.01fF
C352 a_n652_109# a_60_109# 0.01fF
C353 a_296_54# a_474_54# 0.10fF
C354 a_n474_607# a_n830_607# 0.03fF
C355 a_772_109# a_772_n887# 0.00fF
C356 a_n238_n942# a_n416_n942# 0.10fF
C357 a_n772_54# a_n594_54# 0.10fF
C358 a_296_54# a_118_54# 0.10fF
C359 a_n296_607# a_772_607# 0.01fF
C360 a_60_n887# a_416_n887# 0.03fF
C361 a_238_109# a_238_n389# 0.00fF
C362 a_772_n389# a_594_n389# 0.06fF
C363 a_n652_109# a_238_109# 0.01fF
C364 a_n296_n389# a_n474_n389# 0.06fF
C365 a_296_54# a_n60_54# 0.03fF
C366 a_n652_n887# a_416_n887# 0.01fF
C367 a_n238_n942# a_296_n942# 0.02fF
C368 a_60_109# a_594_109# 0.02fF
C369 a_n474_n887# a_238_n887# 0.01fF
C370 a_n830_109# a_n296_109# 0.02fF
C371 a_238_n389# a_n474_n389# 0.01fF
C372 a_n238_n942# a_n238_n444# 0.15fF
C373 a_238_109# a_594_109# 0.03fF
C374 a_416_n389# a_n652_n389# 0.01fF
C375 a_n772_552# a_652_552# 0.01fF
C376 a_n830_607# a_n830_n887# 0.00fF
C377 a_60_109# a_60_607# 0.00fF
C378 a_652_54# a_652_552# 0.15fF
C379 a_n238_n942# a_652_n942# 0.01fF
C380 a_n652_607# a_238_607# 0.01fF
C381 a_238_109# a_238_n887# 0.00fF
C382 a_118_n444# a_118_552# 0.03fF
C383 a_474_54# a_118_54# 0.03fF
C384 a_772_n389# a_n118_n389# 0.01fF
C385 a_n416_552# a_n416_n444# 0.03fF
C386 a_n830_607# a_n118_607# 0.01fF
C387 a_474_n444# a_474_552# 0.03fF
C388 a_n238_54# a_n238_552# 0.15fF
C389 a_n60_54# a_474_54# 0.02fF
C390 a_772_n389# a_772_n887# 0.00fF
C391 a_n60_54# a_118_54# 0.10fF
C392 a_416_n389# a_60_n389# 0.03fF
C393 a_n296_607# a_n296_109# 0.00fF
C394 a_238_n887# a_416_n887# 0.06fF
C395 a_60_n887# a_594_n887# 0.02fF
C396 a_n474_n389# a_594_n389# 0.01fF
C397 a_416_607# a_n296_607# 0.01fF
C398 a_474_552# a_n60_552# 0.02fF
C399 a_772_607# a_60_607# 0.01fF
C400 a_n652_n887# a_594_n887# 0.01fF
C401 a_652_n942# a_652_552# 0.01fF
C402 a_n296_n389# a_n296_109# 0.00fF
C403 a_n474_n887# a_772_n887# 0.01fF
C404 a_296_552# a_n772_552# 0.01fF
C405 a_n238_552# a_n772_552# 0.02fF
C406 a_n416_54# a_n594_54# 0.10fF
C407 a_594_607# a_772_607# 0.06fF
C408 a_416_109# a_416_n389# 0.00fF
C409 a_n652_109# a_n296_109# 0.03fF
C410 a_n474_607# a_n118_607# 0.03fF
C411 a_296_54# a_n238_54# 0.02fF
C412 a_474_552# a_n594_552# 0.01fF
C413 a_n416_552# a_n772_552# 0.03fF
C414 a_296_552# a_296_n942# 0.01fF
C415 a_n416_n942# a_n416_552# 0.01fF
C416 a_118_552# a_n60_552# 0.10fF
C417 a_n474_n389# a_n118_n389# 0.03fF
C418 a_n296_n887# a_60_n887# 0.03fF
C419 a_474_n942# a_118_n942# 0.03fF
C420 a_n296_n887# a_n296_607# 0.00fF
C421 a_n830_109# a_n830_n389# 0.00fF
C422 a_n238_n444# a_n238_552# 0.03fF
C423 a_416_n389# a_772_n389# 0.03fF
C424 a_n296_109# a_594_109# 0.01fF
C425 a_n830_607# a_238_607# 0.01fF
C426 a_n296_n887# a_n652_n887# 0.03fF
C427 a_n594_n444# a_n594_n942# 0.15fF
C428 a_594_n887# a_594_109# 0.00fF
C429 a_772_n887# a_772_607# 0.00fF
C430 a_n296_n887# a_n296_n389# 0.00fF
C431 a_238_n887# a_594_n887# 0.03fF
C432 a_296_54# a_652_54# 0.03fF
C433 a_772_n887# a_416_n887# 0.03fF
C434 a_118_552# a_n594_552# 0.01fF
C435 a_n238_54# a_474_54# 0.01fF
C436 a_652_n444# a_652_552# 0.03fF
C437 a_594_n887# a_594_n389# 0.00fF
C438 a_772_n887# a_n1110_n1061# 0.10fF
C439 a_594_n887# a_n1110_n1061# 0.06fF
C440 a_416_n887# a_n1110_n1061# 0.05fF
C441 a_238_n887# a_n1110_n1061# 0.05fF
C442 a_60_n887# a_n1110_n1061# 0.04fF
C443 a_n118_n887# a_n1110_n1061# 0.04fF
C444 a_n296_n887# a_n1110_n1061# 0.05fF
C445 a_n474_n887# a_n1110_n1061# 0.05fF
C446 a_n652_n887# a_n1110_n1061# 0.06fF
C447 a_n830_n887# a_n1110_n1061# 0.10fF
C448 a_652_n942# a_n1110_n1061# 0.27fF
C449 a_474_n942# a_n1110_n1061# 0.24fF
C450 a_296_n942# a_n1110_n1061# 0.24fF
C451 a_118_n942# a_n1110_n1061# 0.24fF
C452 a_n60_n942# a_n1110_n1061# 0.25fF
C453 a_n238_n942# a_n1110_n1061# 0.26fF
C454 a_n416_n942# a_n1110_n1061# 0.26fF
C455 a_n594_n942# a_n1110_n1061# 0.27fF
C456 a_n772_n942# a_n1110_n1061# 0.32fF
C457 a_772_n389# a_n1110_n1061# 0.10fF
C458 a_594_n389# a_n1110_n1061# 0.06fF
C459 a_416_n389# a_n1110_n1061# 0.05fF
C460 a_238_n389# a_n1110_n1061# 0.04fF
C461 a_60_n389# a_n1110_n1061# 0.04fF
C462 a_n118_n389# a_n1110_n1061# 0.04fF
C463 a_n296_n389# a_n1110_n1061# 0.04fF
C464 a_n474_n389# a_n1110_n1061# 0.05fF
C465 a_n652_n389# a_n1110_n1061# 0.06fF
C466 a_n830_n389# a_n1110_n1061# 0.10fF
C467 a_652_n444# a_n1110_n1061# 0.22fF
C468 a_474_n444# a_n1110_n1061# 0.19fF
C469 a_296_n444# a_n1110_n1061# 0.19fF
C470 a_118_n444# a_n1110_n1061# 0.19fF
C471 a_n60_n444# a_n1110_n1061# 0.20fF
C472 a_n238_n444# a_n1110_n1061# 0.21fF
C473 a_n416_n444# a_n1110_n1061# 0.21fF
C474 a_n594_n444# a_n1110_n1061# 0.22fF
C475 a_n772_n444# a_n1110_n1061# 0.27fF
C476 a_772_109# a_n1110_n1061# 0.10fF
C477 a_594_109# a_n1110_n1061# 0.06fF
C478 a_416_109# a_n1110_n1061# 0.05fF
C479 a_238_109# a_n1110_n1061# 0.05fF
C480 a_60_109# a_n1110_n1061# 0.04fF
C481 a_n118_109# a_n1110_n1061# 0.04fF
C482 a_n296_109# a_n1110_n1061# 0.05fF
C483 a_n474_109# a_n1110_n1061# 0.05fF
C484 a_n652_109# a_n1110_n1061# 0.06fF
C485 a_n830_109# a_n1110_n1061# 0.10fF
C486 a_652_54# a_n1110_n1061# 0.23fF
C487 a_474_54# a_n1110_n1061# 0.20fF
C488 a_296_54# a_n1110_n1061# 0.20fF
C489 a_118_54# a_n1110_n1061# 0.21fF
C490 a_n60_54# a_n1110_n1061# 0.21fF
C491 a_n238_54# a_n1110_n1061# 0.22fF
C492 a_n416_54# a_n1110_n1061# 0.23fF
C493 a_n594_54# a_n1110_n1061# 0.24fF
C494 a_n772_54# a_n1110_n1061# 0.28fF
C495 a_772_607# a_n1110_n1061# 0.10fF
C496 a_594_607# a_n1110_n1061# 0.06fF
C497 a_416_607# a_n1110_n1061# 0.06fF
C498 a_238_607# a_n1110_n1061# 0.05fF
C499 a_60_607# a_n1110_n1061# 0.05fF
C500 a_n118_607# a_n1110_n1061# 0.05fF
C501 a_n296_607# a_n1110_n1061# 0.05fF
C502 a_n474_607# a_n1110_n1061# 0.06fF
C503 a_n652_607# a_n1110_n1061# 0.07fF
C504 a_n830_607# a_n1110_n1061# 0.10fF
C505 a_652_552# a_n1110_n1061# 0.30fF
C506 a_474_552# a_n1110_n1061# 0.27fF
C507 a_296_552# a_n1110_n1061# 0.27fF
C508 a_118_552# a_n1110_n1061# 0.27fF
C509 a_n60_552# a_n1110_n1061# 0.28fF
C510 a_n238_552# a_n1110_n1061# 0.29fF
C511 a_n416_552# a_n1110_n1061# 0.29fF
C512 a_n594_552# a_n1110_n1061# 0.30fF
C513 a_n772_552# a_n1110_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_JJWXCM a_n207_n140# a_29_n204# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n204# a_563_n204# a_n741_n140# a_n327_n204# a_385_n204# a_n563_n140#
+ a_n149_n204# w_n777_n240# a_n385_n140# a_207_n204# a_505_n140# VSUBS
X0 a_n385_n140# a_n505_n204# a_n563_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n204# a_149_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n204# a_n29_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n327_n204# a_n385_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_563_n204# a_563_n204# a_505_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n29_n140# a_n149_n204# a_n207_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_505_n140# a_385_n204# a_327_n140# w_n777_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n385_n140# a_n741_n140# 0.03fF
C1 a_n327_n204# a_n741_n140# 0.02fF
C2 a_385_n204# a_n741_n140# 0.01fF
C3 a_n149_n204# a_n741_n140# 0.01fF
C4 a_n327_n204# a_385_n204# 0.01fF
C5 a_n505_n204# a_207_n204# 0.01fF
C6 a_n149_n204# a_n327_n204# 0.10fF
C7 a_n149_n204# a_385_n204# 0.02fF
C8 a_n741_n140# a_207_n204# 0.01fF
C9 a_327_n140# a_n563_n140# 0.02fF
C10 a_n327_n204# a_207_n204# 0.02fF
C11 a_385_n204# a_207_n204# 0.10fF
C12 a_n149_n204# a_207_n204# 0.03fF
C13 a_n563_n140# a_149_n140# 0.03fF
C14 a_n563_n140# a_563_n204# 0.01fF
C15 a_n29_n140# a_n563_n140# 0.04fF
C16 a_n207_n140# a_n563_n140# 0.06fF
C17 a_n563_n140# w_n777_n240# 0.02fF
C18 a_563_n204# a_29_n204# 0.01fF
C19 a_29_n204# w_n777_n240# 0.16fF
C20 a_n563_n140# a_505_n140# 0.02fF
C21 a_327_n140# a_149_n140# 0.13fF
C22 a_327_n140# a_563_n204# 0.03fF
C23 a_327_n140# a_n29_n140# 0.06fF
C24 a_n207_n140# a_327_n140# 0.04fF
C25 a_327_n140# w_n777_n240# 0.02fF
C26 a_149_n140# a_563_n204# 0.02fF
C27 a_n505_n204# a_29_n204# 0.02fF
C28 a_n29_n140# a_149_n140# 0.13fF
C29 a_n207_n140# a_149_n140# 0.06fF
C30 a_n29_n140# a_563_n204# 0.01fF
C31 a_149_n140# w_n777_n240# 0.02fF
C32 a_n207_n140# a_563_n204# 0.01fF
C33 a_563_n204# w_n777_n240# 0.28fF
C34 a_n207_n140# a_n29_n140# 0.13fF
C35 a_n29_n140# w_n777_n240# 0.02fF
C36 a_n385_n140# a_n563_n140# 0.13fF
C37 a_n207_n140# w_n777_n240# 0.02fF
C38 a_n563_n140# a_n741_n140# 0.06fF
C39 a_327_n140# a_505_n140# 0.13fF
C40 a_29_n204# a_n741_n140# 0.01fF
C41 a_n327_n204# a_29_n204# 0.03fF
C42 a_149_n140# a_505_n140# 0.06fF
C43 a_563_n204# a_505_n140# 0.06fF
C44 a_385_n204# a_29_n204# 0.03fF
C45 a_n29_n140# a_505_n140# 0.04fF
C46 a_n207_n140# a_505_n140# 0.03fF
C47 w_n777_n240# a_505_n140# 0.02fF
C48 a_n149_n204# a_29_n204# 0.10fF
C49 a_n505_n204# a_563_n204# 0.01fF
C50 a_327_n140# a_n385_n140# 0.03fF
C51 a_n505_n204# w_n777_n240# 0.19fF
C52 a_n385_n140# a_149_n140# 0.04fF
C53 a_327_n140# a_n741_n140# 0.01fF
C54 a_n385_n140# a_563_n204# 0.01fF
C55 a_n29_n140# a_n385_n140# 0.06fF
C56 a_n207_n140# a_n385_n140# 0.13fF
C57 a_n385_n140# w_n777_n240# 0.02fF
C58 a_29_n204# a_207_n204# 0.10fF
C59 a_149_n140# a_n741_n140# 0.01fF
C60 a_563_n204# a_n741_n140# 0.01fF
C61 a_n29_n140# a_n741_n140# 0.01fF
C62 a_n207_n140# a_n741_n140# 0.02fF
C63 a_n741_n140# w_n777_n240# 0.33fF
C64 a_n327_n204# a_563_n204# 0.01fF
C65 a_385_n204# a_563_n204# 0.07fF
C66 a_n327_n204# w_n777_n240# 0.18fF
C67 a_385_n204# w_n777_n240# 0.14fF
C68 a_n149_n204# a_563_n204# 0.01fF
C69 a_n149_n204# w_n777_n240# 0.17fF
C70 a_n385_n140# a_505_n140# 0.02fF
C71 a_n741_n140# a_505_n140# 0.01fF
C72 a_563_n204# a_207_n204# 0.02fF
C73 a_n505_n204# a_n741_n140# 0.07fF
C74 w_n777_n240# a_207_n204# 0.15fF
C75 a_n505_n204# a_n327_n204# 0.10fF
C76 a_n505_n204# a_385_n204# 0.01fF
C77 a_n149_n204# a_n505_n204# 0.03fF
C78 w_n777_n240# VSUBS 2.24fF
.ends

.subckt sky130_fd_pr__nfet_01v8_LJREPQ a_n149_n195# a_n207_n140# a_207_n195# a_n29_n140#
+ a_149_n140# a_29_n195# a_n385_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_207_n195# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n385_n140# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n149_n195# a_n385_n140# 0.06fF
C1 a_n149_n195# a_29_n195# 0.10fF
C2 a_n149_n195# a_207_n195# 0.02fF
C3 a_29_n195# a_n385_n140# 0.02fF
C4 a_207_n195# a_n385_n140# 0.03fF
C5 a_207_n195# a_29_n195# 0.06fF
C6 a_n29_n140# a_n385_n140# 0.03fF
C7 a_n29_n140# a_207_n195# 0.03fF
C8 a_149_n140# a_n385_n140# 0.02fF
C9 a_149_n140# a_207_n195# 0.06fF
C10 a_149_n140# a_n29_n140# 0.06fF
C11 a_n207_n140# a_n385_n140# 0.06fF
C12 a_207_n195# a_n207_n140# 0.02fF
C13 a_n29_n140# a_n207_n140# 0.06fF
C14 a_149_n140# a_n207_n140# 0.03fF
C15 a_149_n140# VSUBS 0.01fF
C16 a_n29_n140# VSUBS 0.01fF
C17 a_n207_n140# VSUBS 0.02fF
C18 a_207_n195# VSUBS 0.31fF
C19 a_29_n195# VSUBS 0.19fF
C20 a_n149_n195# VSUBS 0.20fF
C21 a_n385_n140# VSUBS 0.33fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SAWXCM a_n207_n140# a_29_n204# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n204# a_563_n204# a_n741_n140# a_n327_n204# a_385_n204# a_n563_n140#
+ a_n149_n204# w_n777_n240# a_n385_n140# a_207_n204# a_505_n140# VSUBS
X0 a_505_n140# a_385_n204# a_327_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n385_n140# a_n505_n204# a_n563_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_327_n140# a_207_n204# a_149_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_149_n140# a_29_n204# a_n29_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n204# a_n385_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_563_n204# a_563_n204# a_505_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n29_n140# a_n149_n204# a_n207_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n385_n140# a_563_n204# 0.01fF
C1 a_505_n140# a_n29_n140# 0.04fF
C2 a_505_n140# a_n741_n140# 0.01fF
C3 a_149_n140# a_n207_n140# 0.06fF
C4 a_n385_n140# a_n563_n140# 0.13fF
C5 a_385_n204# a_n505_n204# 0.01fF
C6 a_29_n204# a_207_n204# 0.10fF
C7 a_29_n204# a_563_n204# 0.01fF
C8 a_n327_n204# a_n149_n204# 0.10fF
C9 a_n505_n204# a_207_n204# 0.01fF
C10 a_n385_n140# w_n777_n240# 0.02fF
C11 a_n505_n204# a_563_n204# 0.01fF
C12 a_149_n140# a_505_n140# 0.06fF
C13 a_29_n204# w_n777_n240# 0.16fF
C14 a_n505_n204# w_n777_n240# 0.19fF
C15 a_327_n140# a_563_n204# 0.03fF
C16 a_n563_n140# a_327_n140# 0.02fF
C17 a_385_n204# a_n741_n140# 0.01fF
C18 a_n207_n140# a_505_n140# 0.03fF
C19 w_n777_n240# a_327_n140# 0.02fF
C20 a_207_n204# a_n741_n140# 0.01fF
C21 a_n505_n204# a_29_n204# 0.02fF
C22 a_563_n204# a_n29_n140# 0.01fF
C23 a_n741_n140# a_563_n204# 0.01fF
C24 a_n563_n140# a_n29_n140# 0.04fF
C25 a_n563_n140# a_n741_n140# 0.06fF
C26 a_n385_n140# a_327_n140# 0.03fF
C27 a_385_n204# a_n149_n204# 0.02fF
C28 w_n777_n240# a_n29_n140# 0.02fF
C29 w_n777_n240# a_n741_n140# 0.33fF
C30 a_149_n140# a_563_n204# 0.02fF
C31 a_149_n140# a_n563_n140# 0.03fF
C32 a_n149_n204# a_207_n204# 0.03fF
C33 a_n149_n204# a_563_n204# 0.01fF
C34 a_n385_n140# a_n29_n140# 0.06fF
C35 a_n385_n140# a_n741_n140# 0.03fF
C36 a_n327_n204# a_385_n204# 0.01fF
C37 a_149_n140# w_n777_n240# 0.02fF
C38 a_29_n204# a_n741_n140# 0.01fF
C39 a_n149_n204# w_n777_n240# 0.17fF
C40 a_n207_n140# a_563_n204# 0.01fF
C41 a_n327_n204# a_207_n204# 0.02fF
C42 a_n327_n204# a_563_n204# 0.01fF
C43 a_n505_n204# a_n741_n140# 0.07fF
C44 a_149_n140# a_n385_n140# 0.04fF
C45 a_n207_n140# a_n563_n140# 0.06fF
C46 a_n207_n140# w_n777_n240# 0.02fF
C47 a_n149_n204# a_29_n204# 0.10fF
C48 a_505_n140# a_563_n204# 0.06fF
C49 a_n327_n204# w_n777_n240# 0.18fF
C50 a_327_n140# a_n29_n140# 0.06fF
C51 a_505_n140# a_n563_n140# 0.02fF
C52 a_327_n140# a_n741_n140# 0.01fF
C53 a_n149_n204# a_n505_n204# 0.03fF
C54 a_n385_n140# a_n207_n140# 0.13fF
C55 a_505_n140# w_n777_n240# 0.02fF
C56 a_n327_n204# a_29_n204# 0.03fF
C57 a_n741_n140# a_n29_n140# 0.01fF
C58 a_149_n140# a_327_n140# 0.13fF
C59 a_n385_n140# a_505_n140# 0.02fF
C60 a_n327_n204# a_n505_n204# 0.10fF
C61 a_385_n204# a_207_n204# 0.10fF
C62 a_149_n140# a_n29_n140# 0.13fF
C63 a_149_n140# a_n741_n140# 0.01fF
C64 a_385_n204# a_563_n204# 0.07fF
C65 a_n149_n204# a_n741_n140# 0.01fF
C66 a_n207_n140# a_327_n140# 0.04fF
C67 a_207_n204# a_563_n204# 0.02fF
C68 a_n563_n140# a_563_n204# 0.01fF
C69 a_385_n204# w_n777_n240# 0.14fF
C70 a_505_n140# a_327_n140# 0.13fF
C71 a_n207_n140# a_n29_n140# 0.13fF
C72 a_n207_n140# a_n741_n140# 0.02fF
C73 a_n327_n204# a_n741_n140# 0.02fF
C74 a_207_n204# w_n777_n240# 0.15fF
C75 w_n777_n240# a_563_n204# 0.28fF
C76 a_n563_n140# w_n777_n240# 0.02fF
C77 a_385_n204# a_29_n204# 0.03fF
C78 w_n777_n240# VSUBS 2.24fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_28TRYY a_n149_54# a_n1097_109# a_919_n444# a_29_54#
+ a_1097_n942# a_n29_n389# a_n327_n444# a_n207_n887# a_n1555_n1061# a_n1097_n389#
+ a_385_n444# a_149_n389# a_563_54# a_n505_n942# a_n207_109# a_n1275_n887# a_n505_552#
+ a_563_n942# a_327_n887# a_505_109# a_n741_n389# a_n327_552# a_n1217_54# a_327_109#
+ a_n1275_607# a_n149_552# a_861_n389# a_149_109# a_n1097_607# a_385_54# a_n149_n444#
+ a_919_n942# a_n29_109# a_n29_n887# a_n327_n942# a_207_n444# a_n1097_n887# a_385_n942#
+ a_149_n887# a_1097_552# a_n207_607# a_n1039_54# a_207_54# a_n1217_n444# a_n563_n389#
+ a_1217_n389# a_505_607# a_n861_n444# a_n741_n887# a_n861_54# a_327_607# a_683_n389#
+ a_207_552# a_149_607# a_861_n887# a_n919_n389# a_n741_109# a_n149_n942# a_n919_109#
+ a_n29_607# a_919_54# a_n1217_552# a_1217_109# a_n563_109# a_n1039_n444# a_n385_n389#
+ a_n861_552# a_n683_54# a_207_n942# a_n1039_552# a_1039_109# a_29_n444# a_1039_n389#
+ a_861_109# a_n385_109# a_n683_n444# a_n1217_n942# a_n563_n887# a_29_552# a_n683_552#
+ a_1217_n887# a_683_109# a_n861_n942# a_741_n444# a_505_n389# a_683_n887# a_n505_54#
+ a_n919_n887# a_n741_607# a_n919_607# a_1217_607# a_1097_54# a_1097_n444# a_n563_607#
+ a_n207_n389# a_n1039_n942# a_n385_n887# a_1039_607# a_1039_n887# a_861_607# a_29_n942#
+ a_n385_607# a_n327_54# a_n505_n444# a_n683_n942# a_741_552# a_n1275_n389# a_919_552#
+ a_683_607# a_563_n444# a_327_n389# a_563_552# a_741_n942# a_505_n887# a_741_54#
+ a_n1275_109# a_385_552#
X0 a_n919_607# a_n1039_552# a_n1097_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1039_607# a_919_552# a_861_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_109# a_29_54# a_n29_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1097_n887# a_n1217_n942# a_n1275_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_683_n887# a_563_n942# a_505_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n207_n389# a_n327_n444# a_n385_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_607# a_n327_552# a_n385_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n1275_109# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=3.248e+12p ps=2.704e+07u w=1.4e+06u l=600000u
X8 a_683_109# a_563_54# a_505_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_1217_n389# a_1097_n444# a_1039_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1275_n389# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n563_109# a_n683_54# a_n741_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1555_n1061# a_n1555_n1061# a_1217_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_n741_n389# a_n861_n444# a_n919_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n29_n887# a_n149_n942# a_n207_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n919_109# a_n1039_54# a_n1097_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_327_109# a_207_54# a_149_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1039_109# a_919_54# a_861_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1097_n389# a_n1217_n444# a_n1275_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_683_n389# a_563_n444# a_505_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_1039_n389# a_919_n444# a_861_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_505_607# a_385_552# a_327_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n207_109# a_n327_54# a_n385_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_n563_n887# a_n683_n942# a_n741_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_1217_607# a_1097_552# a_1039_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n919_n887# a_n1039_n942# a_n1097_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_505_n887# a_385_n942# a_327_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_861_607# a_741_552# a_683_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_n29_n389# a_n149_n444# a_n207_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n385_n887# a_n505_n942# a_n563_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n741_607# a_n861_552# a_n919_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_n1555_n1061# a_n1555_n1061# a_1217_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X32 a_n29_607# a_n149_552# a_n207_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_505_109# a_385_54# a_327_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_327_n887# a_207_n942# a_149_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X35 a_n563_n389# a_n683_n444# a_n741_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_149_n887# a_29_n942# a_n29_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_n1097_607# a_n1217_552# a_n1275_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X38 a_1217_109# a_1097_54# a_1039_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n919_n389# a_n1039_n444# a_n1097_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_505_n389# a_385_n444# a_327_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X41 a_n385_607# a_n505_552# a_n563_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X42 a_861_109# a_741_54# a_683_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_861_n887# a_741_n942# a_683_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X44 a_n385_n389# a_n505_n444# a_n563_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X45 a_n741_109# a_n861_54# a_n919_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X46 a_n1555_n1061# a_n1555_n1061# a_1217_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X47 a_n29_109# a_n149_54# a_n207_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X48 a_327_n389# a_207_n444# a_149_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X49 a_149_n389# a_29_n444# a_n29_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X50 a_149_607# a_29_552# a_n29_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X51 a_n1097_109# a_n1217_54# a_n1275_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X52 a_n207_n887# a_n327_n942# a_n385_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X53 a_n1275_607# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X54 a_683_607# a_563_552# a_505_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X55 a_n385_109# a_n505_54# a_n563_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X56 a_861_n389# a_741_n444# a_683_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X57 a_1217_n887# a_1097_n942# a_1039_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X58 a_n1275_n887# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X59 a_n563_607# a_n683_552# a_n741_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X60 a_n1555_n1061# a_n1555_n1061# a_1217_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X61 a_n741_n887# a_n861_n942# a_n919_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X62 a_327_607# a_207_552# a_149_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X63 a_1039_n887# a_919_n942# a_861_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n207_109# a_149_109# 0.03fF
C1 a_n505_n444# a_n505_54# 0.15fF
C2 a_n919_607# a_n919_n389# 0.00fF
C3 a_n1039_n444# a_n149_n444# 0.01fF
C4 a_n207_n389# a_n563_n389# 0.03fF
C5 a_n327_552# a_n327_54# 0.15fF
C6 a_n683_n444# a_n683_n942# 0.15fF
C7 a_n1097_109# a_n563_109# 0.02fF
C8 a_n327_n444# a_n861_n444# 0.02fF
C9 a_n29_n887# a_n1097_n887# 0.01fF
C10 a_n207_n887# a_1217_n887# 0.01fF
C11 a_n861_n942# a_n683_n942# 0.10fF
C12 a_n919_n389# a_n1275_n389# 0.03fF
C13 a_n741_109# a_n385_109# 0.03fF
C14 a_n207_109# a_n29_109# 0.06fF
C15 a_1217_109# a_1217_n389# 0.00fF
C16 a_741_552# a_29_552# 0.01fF
C17 a_505_n389# a_n919_n389# 0.01fF
C18 a_327_109# a_n1275_109# 0.01fF
C19 a_919_54# a_1097_54# 0.10fF
C20 a_385_n444# a_n1217_n444# 0.01fF
C21 a_327_109# a_1217_109# 0.01fF
C22 a_n505_552# a_n505_n942# 0.01fF
C23 a_n327_552# a_741_552# 0.01fF
C24 a_919_n942# a_n505_n942# 0.01fF
C25 a_n683_54# a_385_54# 0.01fF
C26 a_n505_552# a_n1217_552# 0.01fF
C27 a_741_n942# a_n505_n942# 0.01fF
C28 a_n563_n887# a_n563_607# 0.00fF
C29 a_683_109# a_505_109# 0.06fF
C30 a_505_607# a_1039_607# 0.02fF
C31 a_149_n389# a_n563_n389# 0.01fF
C32 a_919_54# a_741_54# 0.10fF
C33 a_n207_n389# a_n741_n389# 0.02fF
C34 a_861_109# a_n385_109# 0.01fF
C35 a_683_109# a_149_109# 0.02fF
C36 a_207_n444# a_n149_n444# 0.03fF
C37 a_1039_109# a_861_109# 0.06fF
C38 a_741_n444# a_741_n942# 0.15fF
C39 a_1097_n942# a_1097_54# 0.03fF
C40 a_1039_607# a_n563_607# 0.01fF
C41 a_385_n942# a_n1217_n942# 0.01fF
C42 a_149_n887# a_n1097_n887# 0.01fF
C43 a_n207_607# a_n207_n389# 0.00fF
C44 a_385_n942# a_29_n942# 0.03fF
C45 a_n327_n444# a_n327_54# 0.15fF
C46 a_n29_109# a_683_109# 0.01fF
C47 a_n919_109# a_n919_n887# 0.00fF
C48 a_919_54# a_563_54# 0.03fF
C49 a_n385_n887# a_505_n887# 0.01fF
C50 a_207_n444# a_n1039_n444# 0.01fF
C51 a_505_607# a_n919_607# 0.01fF
C52 a_n29_n887# a_n29_109# 0.00fF
C53 a_327_n887# a_n919_n887# 0.01fF
C54 a_n385_607# a_1217_607# 0.01fF
C55 a_741_54# a_1097_54# 0.03fF
C56 a_n861_54# a_n505_54# 0.03fF
C57 a_n741_n389# a_149_n389# 0.01fF
C58 a_n683_n444# a_n1217_n444# 0.02fF
C59 a_1217_109# a_505_109# 0.01fF
C60 a_385_552# a_741_552# 0.03fF
C61 a_919_552# a_741_552# 0.10fF
C62 a_149_n887# a_149_n389# 0.00fF
C63 a_n1275_109# a_149_109# 0.01fF
C64 a_505_n887# a_683_n887# 0.06fF
C65 a_n1097_n389# a_n1097_607# 0.00fF
C66 a_1217_109# a_149_109# 0.01fF
C67 a_n919_607# a_n563_607# 0.03fF
C68 a_29_n942# a_29_552# 0.01fF
C69 a_505_n389# a_505_607# 0.00fF
C70 a_n1217_n942# a_n861_n942# 0.03fF
C71 a_n149_n942# a_n683_n942# 0.02fF
C72 a_29_n942# a_n861_n942# 0.01fF
C73 a_n741_109# a_n1097_109# 0.03fF
C74 a_563_54# a_1097_54# 0.02fF
C75 a_n1275_109# a_n29_109# 0.01fF
C76 a_741_n444# a_n149_n444# 0.01fF
C77 a_n385_109# a_n385_n389# 0.00fF
C78 a_n861_552# a_n1217_552# 0.03fF
C79 a_1217_109# a_n29_109# 0.01fF
C80 a_n1039_54# a_n505_54# 0.02fF
C81 a_1217_n887# a_1217_607# 0.00fF
C82 a_n505_n444# a_563_n444# 0.01fF
C83 a_149_n887# a_149_109# 0.00fF
C84 a_n1097_n389# a_n563_n389# 0.02fF
C85 a_741_552# a_1097_552# 0.03fF
C86 a_563_n942# a_n683_n942# 0.01fF
C87 a_919_54# a_207_54# 0.01fF
C88 a_683_n389# a_1217_n389# 0.02fF
C89 a_327_109# a_n919_109# 0.01fF
C90 a_1097_n942# a_n505_n942# 0.01fF
C91 a_327_607# a_327_109# 0.00fF
C92 a_n385_n389# a_n29_n389# 0.03fF
C93 a_563_54# a_741_54# 0.10fF
C94 a_n1039_54# a_n861_54# 0.10fF
C95 a_919_n444# a_563_n444# 0.03fF
C96 a_683_n887# a_683_607# 0.00fF
C97 a_n29_n887# a_505_n887# 0.02fF
C98 a_n207_n389# a_683_n389# 0.01fF
C99 a_29_n444# a_n149_n444# 0.10fF
C100 a_n683_54# a_n149_54# 0.02fF
C101 a_n563_n887# a_n207_n887# 0.03fF
C102 a_327_n887# a_327_109# 0.00fF
C103 a_1039_109# a_1039_607# 0.00fF
C104 a_n385_n389# a_n1275_n389# 0.01fF
C105 a_385_n444# a_n505_n444# 0.01fF
C106 a_n919_n887# a_n741_n887# 0.06fF
C107 a_n505_54# a_385_54# 0.01fF
C108 a_n1275_n887# a_n919_n887# 0.03fF
C109 a_741_552# a_n149_552# 0.01fF
C110 a_1097_n444# a_n149_n444# 0.01fF
C111 a_1039_109# a_n385_109# 0.01fF
C112 a_207_552# a_n683_552# 0.01fF
C113 a_505_n389# a_n385_n389# 0.01fF
C114 a_n683_54# a_n683_n444# 0.15fF
C115 a_n327_n444# a_n1217_n444# 0.01fF
C116 a_327_n887# a_n1097_n887# 0.01fF
C117 a_327_n389# a_1217_n389# 0.01fF
C118 a_n1097_n389# a_n741_n389# 0.03fF
C119 a_683_607# a_683_109# 0.00fF
C120 a_385_n444# a_919_n444# 0.02fF
C121 a_207_54# a_1097_54# 0.01fF
C122 a_29_n444# a_n1039_n444# 0.01fF
C123 a_327_109# a_327_n389# 0.00fF
C124 a_149_607# a_149_n389# 0.00fF
C125 a_327_n389# a_n207_n389# 0.02fF
C126 a_n861_54# a_385_54# 0.01fF
C127 a_n1039_n942# a_n683_n942# 0.03fF
C128 a_n385_n887# a_683_n887# 0.01fF
C129 a_741_n444# a_741_54# 0.15fF
C130 a_683_n389# a_149_n389# 0.02fF
C131 a_n683_552# a_n1039_552# 0.03fF
C132 a_505_607# a_1217_607# 0.01fF
C133 a_741_n444# a_207_n444# 0.02fF
C134 a_207_54# a_741_54# 0.02fF
C135 a_1039_n389# a_1217_n389# 0.06fF
C136 a_149_n887# a_505_n887# 0.03fF
C137 a_505_109# a_n919_109# 0.01fF
C138 a_n207_109# a_683_109# 0.01fF
C139 a_149_607# a_149_109# 0.00fF
C140 a_n1217_54# a_n1217_552# 0.15fF
C141 a_n149_n942# a_n1217_n942# 0.01fF
C142 a_1097_n942# a_1097_n444# 0.15fF
C143 a_207_54# a_207_n444# 0.15fF
C144 a_n207_n389# a_1039_n389# 0.01fF
C145 a_n149_n942# a_29_n942# 0.10fF
C146 a_n29_109# a_n29_607# 0.00fF
C147 a_n919_109# a_149_109# 0.01fF
C148 a_1097_n444# a_1097_54# 0.15fF
C149 a_n1039_54# a_385_54# 0.01fF
C150 a_n29_n389# a_n1275_n389# 0.01fF
C151 a_n861_n444# a_n149_n444# 0.01fF
C152 a_563_552# a_n683_552# 0.01fF
C153 a_327_n389# a_149_n389# 0.06fF
C154 a_207_54# a_563_54# 0.03fF
C155 a_n683_n444# a_n505_n444# 0.10fF
C156 a_505_n389# a_n29_n389# 0.02fF
C157 a_207_n444# a_29_n444# 0.10fF
C158 a_n385_n887# a_n29_n887# 0.03fF
C159 a_n29_109# a_n919_109# 0.01fF
C160 a_207_54# a_n1217_54# 0.01fF
C161 a_919_n942# a_n683_n942# 0.01fF
C162 a_683_n887# a_683_109# 0.00fF
C163 a_563_n942# a_29_n942# 0.02fF
C164 a_741_n942# a_n683_n942# 0.01fF
C165 a_n861_n444# a_n861_552# 0.03fF
C166 a_n919_n389# a_n919_n887# 0.00fF
C167 a_327_109# a_n563_109# 0.01fF
C168 a_861_n389# a_1217_n389# 0.03fF
C169 a_n505_552# a_741_552# 0.01fF
C170 a_29_54# a_919_54# 0.01fF
C171 a_n1039_54# a_n1039_552# 0.15fF
C172 a_n1097_n887# a_n741_n887# 0.03fF
C173 a_919_n444# a_n683_n444# 0.01fF
C174 a_207_552# a_207_n942# 0.01fF
C175 a_n1275_n887# a_n1097_n887# 0.06fF
C176 a_207_n444# a_1097_n444# 0.01fF
C177 a_n29_n887# a_683_n887# 0.01fF
C178 a_n861_n444# a_n1039_n444# 0.10fF
C179 a_n207_n389# a_861_n389# 0.01fF
C180 a_741_n942# a_741_552# 0.01fF
C181 a_n1275_109# a_n207_109# 0.01fF
C182 a_1039_n389# a_149_n389# 0.01fF
C183 a_n207_109# a_1217_109# 0.01fF
C184 a_n385_109# a_n1097_109# 0.01fF
C185 a_n207_607# a_683_607# 0.01fF
C186 a_207_n942# a_n327_n942# 0.02fF
C187 a_n505_54# a_n149_54# 0.03fF
C188 a_207_552# a_n1039_552# 0.01fF
C189 a_n1217_n942# a_n1039_n942# 0.10fF
C190 a_919_54# a_n327_54# 0.01fF
C191 a_29_n942# a_n1039_n942# 0.01fF
C192 a_1039_607# a_1217_607# 0.06fF
C193 a_149_n887# a_n385_n887# 0.02fF
C194 a_29_54# a_1097_54# 0.01fF
C195 a_741_n444# a_29_n444# 0.01fF
C196 a_861_n389# a_149_n389# 0.01fF
C197 a_n207_607# a_n207_109# 0.00fF
C198 a_n861_54# a_n149_54# 0.01fF
C199 a_683_607# a_n741_607# 0.01fF
C200 a_207_n444# a_n861_n444# 0.01fF
C201 a_n683_552# a_29_552# 0.01fF
C202 a_n327_n444# a_n505_n444# 0.10fF
C203 a_n683_n444# a_n683_552# 0.03fF
C204 a_1217_n389# a_1217_n887# 0.00fF
C205 a_207_552# a_563_552# 0.03fF
C206 a_505_109# a_n563_109# 0.01fF
C207 a_n207_n389# a_n919_n389# 0.01fF
C208 a_149_n887# a_683_n887# 0.02fF
C209 a_327_n887# a_505_n887# 0.06fF
C210 a_327_n389# a_n1097_n389# 0.01fF
C211 a_1217_109# a_683_109# 0.02fF
C212 a_29_54# a_741_54# 0.01fF
C213 a_149_109# a_n563_109# 0.01fF
C214 a_741_n444# a_1097_n444# 0.03fF
C215 a_n327_552# a_n683_552# 0.03fF
C216 a_683_607# a_n29_607# 0.01fF
C217 a_919_n444# a_n327_n444# 0.01fF
C218 a_919_552# a_919_n444# 0.03fF
C219 a_385_n444# a_385_54# 0.15fF
C220 a_n861_54# a_n861_n942# 0.03fF
C221 a_741_552# a_n861_552# 0.01fF
C222 a_683_607# a_861_607# 0.06fF
C223 a_n1039_54# a_n149_54# 0.01fF
C224 a_149_607# a_683_607# 0.02fF
C225 a_n327_54# a_1097_54# 0.01fF
C226 a_n29_109# a_n563_109# 0.02fF
C227 a_29_n942# a_919_n942# 0.01fF
C228 a_741_n942# a_29_n942# 0.01fF
C229 a_563_552# a_n1039_552# 0.01fF
C230 a_327_607# a_683_607# 0.03fF
C231 a_861_n887# a_505_n887# 0.03fF
C232 a_29_54# a_563_54# 0.02fF
C233 a_563_552# a_563_n444# 0.03fF
C234 a_1097_n444# a_29_n444# 0.01fF
C235 a_683_n389# a_683_607# 0.00fF
C236 a_29_54# a_n1217_54# 0.01fF
C237 a_327_109# a_n741_109# 0.01fF
C238 a_n207_607# a_n1097_607# 0.01fF
C239 a_207_n942# a_385_n942# 0.10fF
C240 a_n919_n389# a_149_n389# 0.01fF
C241 a_n741_n389# a_n563_n389# 0.06fF
C242 a_149_n887# a_n29_n887# 0.06fF
C243 a_741_54# a_n327_54# 0.01fF
C244 a_385_n942# a_385_54# 0.03fF
C245 a_385_n444# a_563_n444# 0.10fF
C246 a_741_n444# a_n861_n444# 0.01fF
C247 a_n207_109# a_n919_109# 0.01fF
C248 a_n149_54# a_385_54# 0.02fF
C249 a_385_n942# a_n327_n942# 0.01fF
C250 a_385_552# a_n683_552# 0.01fF
C251 a_563_54# a_n327_54# 0.01fF
C252 a_n149_n444# a_n1217_n444# 0.01fF
C253 a_741_552# a_741_54# 0.15fF
C254 a_327_109# a_861_109# 0.02fF
C255 a_919_552# a_n683_552# 0.01fF
C256 a_505_n887# a_n741_n887# 0.01fF
C257 a_n1097_607# a_n741_607# 0.03fF
C258 a_n1217_54# a_n327_54# 0.01fF
C259 a_207_552# a_29_552# 0.10fF
C260 a_n563_n887# a_n919_n887# 0.03fF
C261 a_207_n942# a_n861_n942# 0.01fF
C262 a_327_n887# a_n385_n887# 0.01fF
C263 a_n861_n444# a_29_n444# 0.01fF
C264 a_29_54# a_207_54# 0.10fF
C265 a_207_552# a_n327_552# 0.02fF
C266 a_683_n887# a_683_n389# 0.00fF
C267 a_n29_607# a_n1097_607# 0.01fF
C268 a_327_n887# a_683_n887# 0.03fF
C269 a_n1039_n444# a_n1217_n444# 0.10fF
C270 a_149_607# a_n1097_607# 0.01fF
C271 a_n741_109# a_505_109# 0.01fF
C272 a_n327_n942# a_n861_n942# 0.02fF
C273 a_29_54# a_29_n444# 0.15fF
C274 a_n505_n942# a_n683_n942# 0.10fF
C275 a_29_552# a_n1039_552# 0.01fF
C276 a_385_n444# a_385_n942# 0.15fF
C277 a_683_109# a_n919_109# 0.01fF
C278 a_n29_n887# a_n29_607# 0.00fF
C279 a_n741_109# a_149_109# 0.01fF
C280 a_327_607# a_n1097_607# 0.01fF
C281 a_861_n887# a_n385_n887# 0.01fF
C282 a_n327_552# a_n327_n942# 0.01fF
C283 a_n683_n444# a_563_n444# 0.01fF
C284 a_683_n389# a_683_109# 0.00fF
C285 a_n1097_n389# a_n919_n389# 0.06fF
C286 a_n327_552# a_n1039_552# 0.01fF
C287 a_29_n942# a_1097_n942# 0.01fF
C288 a_207_54# a_n327_54# 0.02fF
C289 a_n741_109# a_n29_109# 0.01fF
C290 a_563_552# a_29_552# 0.02fF
C291 a_n385_n389# a_1217_n389# 0.01fF
C292 a_861_n887# a_683_n887# 0.06fF
C293 a_1039_n887# a_505_n887# 0.02fF
C294 a_n149_552# a_n683_552# 0.02fF
C295 a_n505_552# a_n505_n444# 0.03fF
C296 a_861_109# a_505_109# 0.03fF
C297 a_n919_607# a_n919_n887# 0.00fF
C298 a_n207_n887# a_n919_n887# 0.01fF
C299 a_683_n389# a_n563_n389# 0.01fF
C300 a_n207_n389# a_n385_n389# 0.06fF
C301 a_n327_552# a_563_552# 0.01fF
C302 a_n741_n389# a_n741_607# 0.00fF
C303 a_327_n887# a_n29_n887# 0.03fF
C304 a_861_109# a_149_109# 0.01fF
C305 a_741_n444# a_741_552# 0.03fF
C306 a_505_607# a_505_109# 0.00fF
C307 a_385_n444# a_n683_n444# 0.01fF
C308 a_919_54# a_n683_54# 0.01fF
C309 a_385_552# a_207_552# 0.10fF
C310 a_207_n444# a_n1217_n444# 0.01fF
C311 a_919_552# a_207_552# 0.01fF
C312 a_385_552# a_385_54# 0.15fF
C313 a_505_n887# a_1217_n887# 0.01fF
C314 a_n385_n887# a_n741_n887# 0.03fF
C315 a_n207_109# a_n563_109# 0.03fF
C316 a_n1275_109# a_n919_109# 0.03fF
C317 a_n563_n887# a_n1097_n887# 0.02fF
C318 a_919_n444# a_919_n942# 0.15fF
C319 a_n385_n887# a_n1275_n887# 0.01fF
C320 a_861_109# a_n29_109# 0.01fF
C321 a_n207_607# a_n741_607# 0.02fF
C322 a_683_607# a_n385_607# 0.01fF
C323 a_n1217_54# a_n1217_n444# 0.15fF
C324 a_683_n887# a_n741_n887# 0.01fF
C325 a_861_n887# a_n29_n887# 0.01fF
C326 a_327_n389# a_n563_n389# 0.01fF
C327 a_327_109# a_n385_109# 0.01fF
C328 a_n327_n444# a_n327_n942# 0.15fF
C329 a_149_n887# a_149_607# 0.00fF
C330 a_n1217_n942# a_n1217_54# 0.03fF
C331 a_207_n942# a_n149_n942# 0.03fF
C332 a_n207_607# a_n29_607# 0.06fF
C333 a_385_n942# a_n861_n942# 0.01fF
C334 a_207_552# a_1097_552# 0.01fF
C335 a_n1097_607# a_n1275_607# 0.06fF
C336 a_385_552# a_n1039_552# 0.01fF
C337 a_n385_n389# a_149_n389# 0.02fF
C338 a_683_n389# a_n741_n389# 0.01fF
C339 a_1039_109# a_327_109# 0.01fF
C340 a_n327_n444# a_563_n444# 0.01fF
C341 a_1217_n389# a_n29_n389# 0.01fF
C342 a_n207_607# a_861_607# 0.01fF
C343 a_n207_607# a_149_607# 0.03fF
C344 a_563_n942# a_207_n942# 0.03fF
C345 a_n505_n444# a_n149_n444# 0.03fF
C346 a_149_n887# a_327_n887# 0.06fF
C347 a_n1217_n444# a_n1217_552# 0.03fF
C348 a_n207_n389# a_n29_n389# 0.06fF
C349 a_n1217_n942# a_n505_n942# 0.01fF
C350 a_327_607# a_n207_607# 0.02fF
C351 a_1039_n389# a_n563_n389# 0.01fF
C352 a_385_552# a_563_552# 0.10fF
C353 a_29_n942# a_n505_n942# 0.02fF
C354 a_n149_n942# a_n327_n942# 0.10fF
C355 a_n505_552# a_n505_54# 0.15fF
C356 a_919_552# a_563_552# 0.03fF
C357 a_n385_n887# a_n385_607# 0.00fF
C358 a_683_109# a_n563_109# 0.01fF
C359 a_n207_n887# a_n207_n389# 0.00fF
C360 a_n1217_n942# a_n1217_552# 0.01fF
C361 a_n505_552# a_n683_552# 0.10fF
C362 a_1039_n887# a_n385_n887# 0.01fF
C363 a_n683_54# a_741_54# 0.01fF
C364 a_n29_607# a_n741_607# 0.01fF
C365 a_n1039_54# a_n1039_n942# 0.03fF
C366 a_505_n389# a_1217_n389# 0.01fF
C367 a_385_552# a_385_n444# 0.03fF
C368 a_n29_n887# a_n741_n887# 0.01fF
C369 a_207_552# a_n149_552# 0.03fF
C370 a_n207_n389# a_n1275_n389# 0.01fF
C371 a_919_n444# a_n149_n444# 0.01fF
C372 a_327_n389# a_n741_n389# 0.01fF
C373 a_385_n444# a_n327_n444# 0.01fF
C374 a_n207_n887# a_n1097_n887# 0.01fF
C375 a_n29_n887# a_n1275_n887# 0.01fF
C376 a_n327_552# a_29_552# 0.03fF
C377 a_919_54# a_919_n444# 0.15fF
C378 a_563_n942# a_n327_n942# 0.01fF
C379 a_861_607# a_n741_607# 0.01fF
C380 a_505_n389# a_n207_n389# 0.01fF
C381 a_149_607# a_n741_607# 0.01fF
C382 a_505_607# a_505_n887# 0.00fF
C383 a_n563_n389# a_n563_109# 0.00fF
C384 a_n1275_109# a_n1275_607# 0.00fF
C385 a_861_n887# a_149_n887# 0.01fF
C386 a_n505_n444# a_n1039_n444# 0.02fF
C387 a_1039_n887# a_683_n887# 0.03fF
C388 a_563_n942# a_563_n444# 0.15fF
C389 a_563_552# a_1097_552# 0.02fF
C390 a_327_607# a_n741_607# 0.01fF
C391 a_n385_n887# a_1217_n887# 0.01fF
C392 a_29_54# a_n327_54# 0.03fF
C393 a_n683_54# a_563_54# 0.01fF
C394 a_861_n389# a_n563_n389# 0.01fF
C395 a_29_n444# a_n1217_n444# 0.01fF
C396 a_n29_607# a_861_607# 0.01fF
C397 a_n385_109# a_505_109# 0.01fF
C398 a_n683_54# a_n1217_54# 0.02fF
C399 a_n29_n389# a_149_n389# 0.06fF
C400 a_149_607# a_n29_607# 0.06fF
C401 a_n1097_607# a_n385_607# 0.01fF
C402 a_n1275_109# a_n1275_n887# 0.00fF
C403 a_385_552# a_385_n942# 0.01fF
C404 a_n149_552# a_n1039_552# 0.01fF
C405 a_n385_109# a_149_109# 0.02fF
C406 a_207_n942# a_n1039_n942# 0.01fF
C407 a_1039_109# a_505_109# 0.02fF
C408 a_327_607# a_n29_607# 0.03fF
C409 a_n1275_109# a_n563_109# 0.01fF
C410 a_563_n942# a_563_552# 0.01fF
C411 a_149_607# a_861_607# 0.01fF
C412 a_29_n942# a_29_n444# 0.15fF
C413 a_683_n887# a_1217_n887# 0.02fF
C414 a_1039_109# a_149_109# 0.01fF
C415 a_149_n389# a_n1275_n389# 0.01fF
C416 a_n741_109# a_n207_109# 0.02fF
C417 a_n385_n389# a_n1097_n389# 0.01fF
C418 a_327_607# a_861_607# 0.02fF
C419 a_327_607# a_149_607# 0.06fF
C420 a_n741_n389# a_n741_n887# 0.00fF
C421 a_n385_109# a_n29_109# 0.03fF
C422 a_505_n389# a_149_n389# 0.03fF
C423 a_505_607# a_683_607# 0.06fF
C424 a_563_552# a_n149_552# 0.01fF
C425 a_149_n887# a_n741_n887# 0.01fF
C426 a_n207_607# a_n1275_607# 0.01fF
C427 a_1039_n887# a_n29_n887# 0.01fF
C428 a_327_109# a_n1097_109# 0.01fF
C429 a_919_54# a_n505_54# 0.01fF
C430 a_149_n887# a_n1275_n887# 0.01fF
C431 a_1039_109# a_n29_109# 0.01fF
C432 a_n1039_n942# a_n327_n942# 0.01fF
C433 a_385_n942# a_n149_n942# 0.02fF
C434 a_207_n444# a_n505_n444# 0.01fF
C435 a_385_552# a_29_552# 0.03fF
C436 a_919_552# a_29_552# 0.01fF
C437 a_861_n389# a_n741_n389# 0.01fF
C438 a_n1039_n942# a_n1039_552# 0.01fF
C439 a_n683_n444# a_n327_n444# 0.03fF
C440 a_327_607# a_327_n887# 0.00fF
C441 a_683_607# a_n563_607# 0.01fF
C442 a_n1097_109# a_n1097_n887# 0.00fF
C443 a_505_n389# a_505_109# 0.00fF
C444 a_n29_109# a_n29_n389# 0.00fF
C445 a_n861_552# a_n683_552# 0.10fF
C446 a_207_552# a_n505_552# 0.01fF
C447 a_n563_n887# a_505_n887# 0.01fF
C448 a_n919_n389# a_n563_n389# 0.03fF
C449 a_385_552# a_n327_552# 0.01fF
C450 a_861_109# a_n207_109# 0.01fF
C451 a_207_n942# a_919_n942# 0.01fF
C452 a_n149_n942# a_n149_54# 0.03fF
C453 a_919_552# a_n327_552# 0.01fF
C454 a_n327_552# a_n327_n444# 0.03fF
C455 a_207_54# a_n683_54# 0.01fF
C456 a_919_n444# a_207_n444# 0.01fF
C457 a_n29_n887# a_1217_n887# 0.01fF
C458 a_563_n942# a_385_n942# 0.10fF
C459 a_741_n942# a_207_n942# 0.02fF
C460 a_n861_54# a_n861_552# 0.15fF
C461 a_1217_n389# a_1217_607# 0.00fF
C462 a_861_n887# a_861_607# 0.00fF
C463 a_n741_607# a_n1275_607# 0.02fF
C464 a_327_607# a_327_n389# 0.00fF
C465 a_n861_n444# a_n1217_n444# 0.03fF
C466 a_1097_552# a_29_552# 0.01fF
C467 a_n741_109# a_683_109# 0.01fF
C468 a_327_n389# a_683_n389# 0.03fF
C469 a_n505_54# a_1097_54# 0.01fF
C470 a_n149_n942# a_n861_n942# 0.01fF
C471 a_n505_n942# a_n505_n444# 0.15fF
C472 a_919_n942# a_n327_n942# 0.01fF
C473 a_n1097_n389# a_n29_n389# 0.01fF
C474 a_n741_607# a_n741_n887# 0.00fF
C475 a_n29_607# a_n1275_607# 0.01fF
C476 a_n505_552# a_n1039_552# 0.02fF
C477 a_741_n942# a_n327_n942# 0.01fF
C478 a_327_n887# a_327_n389# 0.00fF
C479 a_n327_552# a_1097_552# 0.01fF
C480 a_1039_n887# a_149_n887# 0.01fF
C481 a_861_n887# a_327_n887# 0.02fF
C482 a_1217_109# a_1217_n887# 0.00fF
C483 a_n149_552# a_n149_54# 0.15fF
C484 a_149_607# a_n1275_607# 0.01fF
C485 a_n207_607# a_n385_607# 0.06fF
C486 a_n1097_n389# a_n1275_n389# 0.06fF
C487 a_563_n942# a_n861_n942# 0.01fF
C488 a_n741_n389# a_n919_n389# 0.06fF
C489 a_n1097_109# a_505_109# 0.01fF
C490 a_741_54# a_n505_54# 0.01fF
C491 a_741_n444# a_n505_n444# 0.01fF
C492 a_683_n389# a_1039_n389# 0.03fF
C493 a_29_54# a_29_n942# 0.03fF
C494 a_327_607# a_n1275_607# 0.01fF
C495 a_563_552# a_n505_552# 0.01fF
C496 a_505_n389# a_n1097_n389# 0.01fF
C497 a_861_109# a_683_109# 0.06fF
C498 a_n1097_109# a_149_109# 0.01fF
C499 a_n149_552# a_29_552# 0.10fF
C500 a_n1039_54# a_n1039_n444# 0.15fF
C501 a_385_n942# a_n1039_n942# 0.01fF
C502 a_n207_n887# a_505_n887# 0.01fF
C503 a_505_607# a_n1097_607# 0.01fF
C504 a_149_n887# a_1217_n887# 0.01fF
C505 a_683_607# a_1039_607# 0.03fF
C506 a_385_552# a_919_552# 0.02fF
C507 a_n861_54# a_741_54# 0.01fF
C508 a_n1275_109# a_n741_109# 0.02fF
C509 a_741_n444# a_919_n444# 0.10fF
C510 a_n327_552# a_n149_552# 0.10fF
C511 a_919_54# a_385_54# 0.02fF
C512 a_n919_109# a_n563_109# 0.03fF
C513 a_n1097_109# a_n29_109# 0.01fF
C514 a_563_54# a_n505_54# 0.01fF
C515 a_861_n389# a_861_607# 0.00fF
C516 a_n385_n887# a_n385_n389# 0.00fF
C517 a_n1097_607# a_n563_607# 0.02fF
C518 a_n1217_54# a_n505_54# 0.01fF
C519 a_n505_n444# a_29_n444# 0.02fF
C520 a_505_n389# a_505_n887# 0.00fF
C521 a_327_n887# a_n741_n887# 0.01fF
C522 a_n741_607# a_n385_607# 0.03fF
C523 a_207_552# a_n861_552# 0.01fF
C524 a_n563_n887# a_n385_n887# 0.06fF
C525 a_327_n887# a_n1275_n887# 0.01fF
C526 a_327_n389# a_1039_n389# 0.01fF
C527 a_n741_109# a_n741_n389# 0.00fF
C528 a_683_n389# a_861_n389# 0.06fF
C529 a_n861_54# a_563_54# 0.01fF
C530 a_385_552# a_1097_552# 0.01fF
C531 a_919_552# a_1097_552# 0.10fF
C532 a_n29_607# a_n385_607# 0.03fF
C533 a_919_n444# a_29_n444# 0.01fF
C534 a_n861_54# a_n1217_54# 0.03fF
C535 a_n505_n444# a_1097_n444# 0.01fF
C536 a_n149_n444# a_563_n444# 0.01fF
C537 a_n1039_n942# a_n861_n942# 0.10fF
C538 a_n505_n942# a_n505_54# 0.03fF
C539 a_n563_n887# a_683_n887# 0.01fF
C540 a_n1217_n942# a_n683_n942# 0.02fF
C541 a_861_109# a_1217_109# 0.03fF
C542 a_683_607# a_n919_607# 0.01fF
C543 a_n563_607# a_n563_n389# 0.00fF
C544 a_385_n942# a_919_n942# 0.02fF
C545 a_207_n942# a_1097_n942# 0.01fF
C546 a_29_n942# a_n683_n942# 0.01fF
C547 a_861_607# a_n385_607# 0.01fF
C548 a_n1097_109# a_n1097_n389# 0.00fF
C549 a_741_n942# a_385_n942# 0.03fF
C550 a_149_607# a_n385_607# 0.02fF
C551 a_n207_109# a_n385_109# 0.06fF
C552 a_861_n887# a_n741_n887# 0.01fF
C553 a_29_54# a_n683_54# 0.01fF
C554 a_n683_552# a_n1217_552# 0.02fF
C555 a_n861_552# a_n1039_552# 0.10fF
C556 a_919_n444# a_1097_n444# 0.10fF
C557 a_385_54# a_1097_54# 0.01fF
C558 a_n385_109# a_n385_n887# 0.00fF
C559 a_1039_109# a_n207_109# 0.01fF
C560 a_327_607# a_n385_607# 0.01fF
C561 a_n1039_54# a_563_54# 0.01fF
C562 a_327_n389# a_861_n389# 0.02fF
C563 a_n1039_54# a_n1217_54# 0.10fF
C564 a_n1039_n444# a_n1039_552# 0.03fF
C565 a_861_n887# a_861_n389# 0.00fF
C566 a_1097_n942# a_n327_n942# 0.01fF
C567 a_385_552# a_n149_552# 0.02fF
C568 a_n505_552# a_29_552# 0.02fF
C569 a_n1039_n444# a_563_n444# 0.01fF
C570 a_385_n444# a_n149_n444# 0.02fF
C571 a_207_54# a_n505_54# 0.01fF
C572 a_919_552# a_n149_552# 0.01fF
C573 a_563_552# a_n861_552# 0.01fF
C574 a_n207_109# a_n207_n887# 0.00fF
C575 a_n919_n389# a_n919_109# 0.00fF
C576 a_741_54# a_385_54# 0.03fF
C577 a_1039_n887# a_327_n887# 0.01fF
C578 a_207_n942# a_207_n444# 0.15fF
C579 a_n1275_n887# a_n1275_607# 0.00fF
C580 a_n563_n887# a_n29_n887# 0.02fF
C581 a_683_n389# a_n919_n389# 0.01fF
C582 a_n327_552# a_n505_552# 0.10fF
C583 a_n385_n887# a_n207_n887# 0.06fF
C584 a_563_n942# a_n149_n942# 0.01fF
C585 a_n741_109# a_n741_607# 0.00fF
C586 a_207_552# a_207_n444# 0.03fF
C587 a_n385_n389# a_n563_n389# 0.06fF
C588 a_741_n942# a_n861_n942# 0.01fF
C589 a_n563_n887# a_n563_n389# 0.00fF
C590 a_n861_n444# a_n505_n444# 0.03fF
C591 a_n207_607# a_505_607# 0.01fF
C592 a_207_54# a_n861_54# 0.01fF
C593 a_861_n389# a_1039_n389# 0.06fF
C594 a_n683_54# a_n327_54# 0.03fF
C595 a_n1275_n887# a_n741_n887# 0.02fF
C596 a_n1097_n887# a_n919_n887# 0.06fF
C597 a_n385_109# a_683_109# 0.01fF
C598 a_n149_552# a_1097_552# 0.01fF
C599 a_n149_n942# a_n149_552# 0.01fF
C600 a_n207_n887# a_683_n887# 0.01fF
C601 a_327_n887# a_1217_n887# 0.01fF
C602 a_563_54# a_385_54# 0.10fF
C603 a_385_n444# a_n1039_n444# 0.01fF
C604 a_n683_54# a_n683_n942# 0.03fF
C605 a_n207_607# a_n563_607# 0.03fF
C606 a_n1217_54# a_385_54# 0.01fF
C607 a_861_n887# a_1039_n887# 0.06fF
C608 a_1039_109# a_683_109# 0.03fF
C609 a_327_n389# a_n919_n389# 0.01fF
C610 a_207_n444# a_563_n444# 0.03fF
C611 a_n741_109# a_n919_109# 0.06fF
C612 a_n149_n444# a_n149_54# 0.15fF
C613 a_207_54# a_n1039_54# 0.01fF
C614 a_207_n942# a_n505_n942# 0.01fF
C615 a_919_54# a_n149_54# 0.01fF
C616 a_n1217_n942# a_n1217_n444# 0.15fF
C617 a_n919_607# a_n1097_607# 0.06fF
C618 a_505_607# a_n741_607# 0.01fF
C619 a_n385_607# a_n1275_607# 0.01fF
C620 a_n385_n389# a_n741_n389# 0.03fF
C621 a_1039_n887# a_1039_n389# 0.00fF
C622 a_861_n887# a_1217_n887# 0.03fF
C623 a_563_54# a_563_n444# 0.15fF
C624 a_207_552# a_n1217_552# 0.01fF
C625 a_n29_n887# a_n29_n389# 0.00fF
C626 a_n683_n444# a_n149_n444# 0.02fF
C627 a_29_n942# a_n1217_n942# 0.01fF
C628 a_n149_n942# a_n1039_n942# 0.01fF
C629 a_149_n887# a_n563_n887# 0.01fF
C630 a_n207_n389# a_1217_n389# 0.01fF
C631 a_505_607# a_n29_607# 0.02fF
C632 a_385_n942# a_1097_n942# 0.01fF
C633 a_n29_n389# a_n563_n389# 0.02fF
C634 a_n563_607# a_n741_607# 0.06fF
C635 a_861_109# a_861_607# 0.00fF
C636 a_385_552# a_n505_552# 0.01fF
C637 a_n1275_109# a_n385_109# 0.01fF
C638 a_n207_109# a_n1097_109# 0.01fF
C639 a_n207_n887# a_n29_n887# 0.06fF
C640 a_919_552# a_n505_552# 0.01fF
C641 a_n505_n942# a_n327_n942# 0.10fF
C642 a_1217_109# a_n385_109# 0.01fF
C643 a_385_n444# a_207_n444# 0.10fF
C644 a_n861_552# a_29_552# 0.01fF
C645 a_505_607# a_861_607# 0.03fF
C646 a_563_552# a_563_54# 0.15fF
C647 a_919_552# a_919_n942# 0.01fF
C648 a_683_607# a_1217_607# 0.02fF
C649 a_149_607# a_505_607# 0.03fF
C650 a_207_54# a_207_n942# 0.03fF
C651 a_1039_109# a_1217_109# 0.06fF
C652 a_563_n942# a_n1039_n942# 0.01fF
C653 a_n861_552# a_n861_n942# 0.01fF
C654 a_207_54# a_207_552# 0.15fF
C655 a_n29_607# a_n563_607# 0.02fF
C656 a_207_54# a_385_54# 0.10fF
C657 a_n563_n389# a_n1275_n389# 0.01fF
C658 a_327_607# a_505_607# 0.06fF
C659 a_n327_552# a_n861_552# 0.02fF
C660 a_n149_54# a_1097_54# 0.01fF
C661 a_n1217_552# a_n1039_552# 0.10fF
C662 a_505_n389# a_n563_n389# 0.01fF
C663 a_861_607# a_n563_607# 0.01fF
C664 a_n683_n444# a_n1039_n444# 0.03fF
C665 a_149_607# a_n563_607# 0.01fF
C666 a_n207_607# a_1039_607# 0.01fF
C667 a_n505_552# a_1097_552# 0.01fF
C668 a_n861_54# a_n861_n444# 0.15fF
C669 a_327_607# a_n563_607# 0.01fF
C670 a_29_54# a_n505_54# 0.02fF
C671 a_741_n444# a_563_n444# 0.10fF
C672 a_n149_n942# a_919_n942# 0.01fF
C673 a_n1275_109# a_n1275_n389# 0.00fF
C674 a_1217_n389# a_149_n389# 0.01fF
C675 a_741_n942# a_n149_n942# 0.01fF
C676 a_n741_n389# a_n29_n389# 0.01fF
C677 a_741_54# a_n149_54# 0.01fF
C678 a_n207_n389# a_149_n389# 0.03fF
C679 a_n1097_109# a_n1097_607# 0.00fF
C680 a_861_n887# a_861_109# 0.00fF
C681 a_29_54# a_n861_54# 0.01fF
C682 a_149_n887# a_n207_n887# 0.03fF
C683 a_563_n942# a_919_n942# 0.03fF
C684 a_563_n942# a_741_n942# 0.10fF
C685 a_n741_n389# a_n1275_n389# 0.02fF
C686 a_n741_109# a_n741_n887# 0.00fF
C687 a_29_n444# a_563_n444# 0.02fF
C688 a_n505_552# a_n149_552# 0.03fF
C689 a_n327_n444# a_n149_n444# 0.10fF
C690 a_327_109# a_505_109# 0.06fF
C691 a_n207_607# a_n919_607# 0.01fF
C692 a_385_n444# a_741_n444# 0.03fF
C693 a_563_54# a_n149_54# 0.01fF
C694 a_505_n389# a_n741_n389# 0.01fF
C695 a_n207_607# a_n207_n887# 0.00fF
C696 a_n741_109# a_n563_109# 0.06fF
C697 a_919_54# a_919_552# 0.15fF
C698 a_n683_n444# a_207_n444# 0.01fF
C699 a_327_109# a_149_109# 0.06fF
C700 a_n1217_54# a_n149_54# 0.01fF
C701 a_n505_54# a_n327_54# 0.10fF
C702 a_385_n942# a_n505_n942# 0.01fF
C703 a_683_n389# a_n385_n389# 0.01fF
C704 a_385_552# a_n861_552# 0.01fF
C705 a_29_54# a_n1039_54# 0.01fF
C706 a_n29_607# a_1039_607# 0.01fF
C707 a_1097_n444# a_563_n444# 0.02fF
C708 a_505_n887# a_n919_n887# 0.01fF
C709 a_1039_n887# a_1217_n887# 0.06fF
C710 a_n683_552# a_n683_n942# 0.01fF
C711 a_327_109# a_n29_109# 0.03fF
C712 a_1039_607# a_861_607# 0.06fF
C713 a_n861_54# a_n327_54# 0.02fF
C714 a_149_607# a_1039_607# 0.01fF
C715 a_327_n887# a_n563_n887# 0.01fF
C716 a_n149_n942# a_n149_n444# 0.15fF
C717 a_385_n444# a_29_n444# 0.03fF
C718 a_n327_n444# a_n1039_n444# 0.01fF
C719 a_n1275_109# a_n1097_109# 0.06fF
C720 a_n505_n444# a_n1217_n444# 0.01fF
C721 a_327_607# a_1039_607# 0.01fF
C722 a_861_109# a_n563_109# 0.01fF
C723 a_n563_607# a_n1275_607# 0.01fF
C724 a_n919_607# a_n741_607# 0.06fF
C725 a_741_552# a_n683_552# 0.01fF
C726 a_n385_109# a_n919_109# 0.02fF
C727 a_861_109# a_861_n389# 0.00fF
C728 a_327_n389# a_n385_n389# 0.01fF
C729 a_385_n444# a_1097_n444# 0.01fF
C730 a_n29_607# a_n29_n389# 0.00fF
C731 a_n505_n942# a_n861_n942# 0.03fF
C732 a_149_n389# a_149_109# 0.00fF
C733 a_29_552# a_n1217_552# 0.01fF
C734 a_n29_607# a_n919_607# 0.01fF
C735 a_n1039_54# a_n327_54# 0.01fF
C736 a_29_54# a_385_54# 0.03fF
C737 a_861_n887# a_n563_n887# 0.01fF
C738 a_n207_n389# a_n1097_n389# 0.01fF
C739 a_207_54# a_n149_54# 0.03fF
C740 a_n563_607# a_n563_109# 0.00fF
C741 a_n149_552# a_n149_n444# 0.03fF
C742 a_n327_552# a_n1217_552# 0.01fF
C743 a_149_607# a_n919_607# 0.01fF
C744 a_n861_n444# a_563_n444# 0.01fF
C745 a_741_n444# a_n683_n444# 0.01fF
C746 a_1097_n942# a_1097_552# 0.01fF
C747 a_n149_n942# a_1097_n942# 0.01fF
C748 a_n919_607# a_n919_109# 0.00fF
C749 a_n1097_n887# a_n1097_n389# 0.00fF
C750 a_683_n389# a_n29_n389# 0.01fF
C751 a_505_109# a_149_109# 0.03fF
C752 a_327_607# a_n919_607# 0.01fF
C753 a_1217_109# a_1217_607# 0.00fF
C754 a_n385_n389# a_1039_n389# 0.01fF
C755 a_1097_552# a_1097_54# 0.15fF
C756 a_207_n444# a_n327_n444# 0.02fF
C757 a_n149_552# a_n861_552# 0.01fF
C758 a_505_607# a_n385_607# 0.01fF
C759 a_327_n887# a_n207_n887# 0.02fF
C760 a_563_n942# a_1097_n942# 0.02fF
C761 a_741_n942# a_919_n942# 0.10fF
C762 a_n29_109# a_505_109# 0.02fF
C763 a_29_n444# a_29_552# 0.03fF
C764 a_n327_54# a_385_54# 0.01fF
C765 a_n683_n444# a_29_n444# 0.01fF
C766 a_n29_109# a_149_109# 0.06fF
C767 a_505_n887# a_n1097_n887# 0.01fF
C768 a_505_n389# a_683_n389# 0.06fF
C769 a_385_n444# a_n861_n444# 0.01fF
C770 a_n385_n887# a_n919_n887# 0.02fF
C771 a_n563_n887# a_n741_n887# 0.06fF
C772 a_207_n942# a_n683_n942# 0.01fF
C773 a_1039_n389# a_1039_607# 0.00fF
C774 a_n563_607# a_n385_607# 0.06fF
C775 a_n1097_n389# a_149_n389# 0.01fF
C776 a_n563_n887# a_n1275_n887# 0.01fF
C777 a_327_n389# a_n29_n389# 0.03fF
C778 a_n563_n887# a_n563_109# 0.00fF
C779 a_861_n389# a_n385_n389# 0.01fF
C780 a_n207_607# a_1217_607# 0.01fF
C781 a_683_n887# a_n919_n887# 0.01fF
C782 a_n327_n942# a_n327_54# 0.03fF
C783 a_861_n887# a_n207_n887# 0.01fF
C784 a_207_552# a_741_552# 0.02fF
C785 a_1039_109# a_1039_n389# 0.00fF
C786 a_327_n389# a_n1275_n389# 0.01fF
C787 a_385_552# a_n1217_552# 0.01fF
C788 a_n327_n942# a_n683_n942# 0.03fF
C789 a_n1039_n942# a_n1039_n444# 0.15fF
C790 a_327_n389# a_505_n389# 0.06fF
C791 a_1039_n389# a_n29_n389# 0.01fF
C792 a_861_109# a_n741_109# 0.01fF
C793 a_n1097_109# a_n919_109# 0.06fF
C794 a_n385_109# a_n563_109# 0.06fF
C795 a_563_n942# a_563_54# 0.03fF
C796 a_741_n444# a_n327_n444# 0.01fF
C797 a_n919_607# a_n1275_607# 0.03fF
C798 a_n385_n389# a_n385_607# 0.00fF
C799 a_919_54# a_919_n942# 0.03fF
C800 a_505_n887# a_505_109# 0.00fF
C801 a_n149_n942# a_n505_n942# 0.03fF
C802 a_1039_109# a_n563_109# 0.01fF
C803 a_n505_552# a_n861_552# 0.03fF
C804 a_n1275_n389# a_n1275_607# 0.00fF
C805 a_327_109# a_n207_109# 0.02fF
C806 a_1039_n887# a_n563_n887# 0.01fF
C807 a_n207_109# a_n207_n389# 0.00fF
C808 a_505_n389# a_1039_n389# 0.02fF
C809 a_n207_n887# a_n741_n887# 0.02fF
C810 a_n29_n887# a_n919_n887# 0.01fF
C811 a_n29_607# a_1217_607# 0.01fF
C812 a_n207_n887# a_n1275_n887# 0.01fF
C813 a_n683_n444# a_n861_n444# 0.10fF
C814 a_n385_n389# a_n919_n389# 0.02fF
C815 a_29_54# a_n149_54# 0.10fF
C816 a_563_n942# a_n505_n942# 0.01fF
C817 a_n861_n444# a_n861_n942# 0.15fF
C818 a_n327_n444# a_29_n444# 0.03fF
C819 a_861_n389# a_n29_n389# 0.01fF
C820 a_1039_607# a_n385_607# 0.01fF
C821 a_n1275_n887# a_n1275_n389# 0.00fF
C822 a_563_552# a_741_552# 0.10fF
C823 a_861_607# a_1217_607# 0.03fF
C824 a_n683_54# a_n505_54# 0.10fF
C825 a_149_607# a_1217_607# 0.01fF
C826 a_1039_n887# a_1039_607# 0.00fF
C827 a_n683_54# a_n683_552# 0.15fF
C828 a_n385_n887# a_n1097_n887# 0.01fF
C829 a_919_n444# a_n505_n444# 0.01fF
C830 a_n385_109# a_n385_607# 0.00fF
C831 a_29_54# a_29_552# 0.15fF
C832 a_327_607# a_1217_607# 0.01fF
C833 a_919_n942# a_1097_n942# 0.10fF
C834 a_741_n942# a_1097_n942# 0.03fF
C835 a_n327_n444# a_1097_n444# 0.01fF
C836 a_n149_552# a_n1217_552# 0.01fF
C837 a_n683_54# a_n861_54# 0.10fF
C838 a_207_n942# a_n1217_n942# 0.01fF
C839 a_505_n389# a_861_n389# 0.03fF
C840 a_1039_n887# a_1039_109# 0.00fF
C841 a_207_n942# a_29_n942# 0.10fF
C842 a_385_n942# a_n683_n942# 0.01fF
C843 a_327_109# a_683_109# 0.03fF
C844 a_n149_54# a_n327_54# 0.10fF
C845 a_505_607# a_n563_607# 0.01fF
C846 a_n919_607# a_n385_607# 0.02fF
C847 a_149_n887# a_n919_n887# 0.01fF
C848 a_741_n942# a_741_54# 0.03fF
C849 a_1097_n444# a_1097_552# 0.03fF
C850 a_1039_n887# a_n207_n887# 0.01fF
C851 a_n1097_n887# a_n1097_607# 0.00fF
C852 a_n1039_n942# a_n505_n942# 0.02fF
C853 a_n1217_n942# a_n327_n942# 0.01fF
C854 a_n207_109# a_505_109# 0.01fF
C855 a_n1039_54# a_n683_54# 0.03fF
C856 a_29_n942# a_n327_n942# 0.03fF
C857 a_n919_n389# a_n29_n389# 0.01fF
C858 a_1217_n887# a_n1555_n1061# 0.10fF
C859 a_1039_n887# a_n1555_n1061# 0.05fF
C860 a_861_n887# a_n1555_n1061# 0.04fF
C861 a_683_n887# a_n1555_n1061# 0.03fF
C862 a_505_n887# a_n1555_n1061# 0.03fF
C863 a_327_n887# a_n1555_n1061# 0.03fF
C864 a_149_n887# a_n1555_n1061# 0.03fF
C865 a_n29_n887# a_n1555_n1061# 0.03fF
C866 a_n207_n887# a_n1555_n1061# 0.03fF
C867 a_n385_n887# a_n1555_n1061# 0.03fF
C868 a_n563_n887# a_n1555_n1061# 0.03fF
C869 a_n741_n887# a_n1555_n1061# 0.03fF
C870 a_n919_n887# a_n1555_n1061# 0.04fF
C871 a_n1097_n887# a_n1555_n1061# 0.05fF
C872 a_n1275_n887# a_n1555_n1061# 0.10fF
C873 a_1097_n942# a_n1555_n1061# 0.27fF
C874 a_919_n942# a_n1555_n1061# 0.23fF
C875 a_741_n942# a_n1555_n1061# 0.23fF
C876 a_563_n942# a_n1555_n1061# 0.24fF
C877 a_385_n942# a_n1555_n1061# 0.24fF
C878 a_207_n942# a_n1555_n1061# 0.25fF
C879 a_29_n942# a_n1555_n1061# 0.26fF
C880 a_n149_n942# a_n1555_n1061# 0.26fF
C881 a_n327_n942# a_n1555_n1061# 0.26fF
C882 a_n505_n942# a_n1555_n1061# 0.26fF
C883 a_n683_n942# a_n1555_n1061# 0.26fF
C884 a_n861_n942# a_n1555_n1061# 0.26fF
C885 a_n1039_n942# a_n1555_n1061# 0.27fF
C886 a_n1217_n942# a_n1555_n1061# 0.32fF
C887 a_1217_n389# a_n1555_n1061# 0.10fF
C888 a_1039_n389# a_n1555_n1061# 0.05fF
C889 a_861_n389# a_n1555_n1061# 0.04fF
C890 a_683_n389# a_n1555_n1061# 0.03fF
C891 a_505_n389# a_n1555_n1061# 0.03fF
C892 a_327_n389# a_n1555_n1061# 0.02fF
C893 a_149_n389# a_n1555_n1061# 0.03fF
C894 a_n29_n389# a_n1555_n1061# 0.03fF
C895 a_n207_n389# a_n1555_n1061# 0.03fF
C896 a_n385_n389# a_n1555_n1061# 0.02fF
C897 a_n563_n389# a_n1555_n1061# 0.03fF
C898 a_n741_n389# a_n1555_n1061# 0.03fF
C899 a_n919_n389# a_n1555_n1061# 0.04fF
C900 a_n1097_n389# a_n1555_n1061# 0.05fF
C901 a_n1275_n389# a_n1555_n1061# 0.10fF
C902 a_1097_n444# a_n1555_n1061# 0.22fF
C903 a_919_n444# a_n1555_n1061# 0.18fF
C904 a_741_n444# a_n1555_n1061# 0.18fF
C905 a_563_n444# a_n1555_n1061# 0.19fF
C906 a_385_n444# a_n1555_n1061# 0.19fF
C907 a_207_n444# a_n1555_n1061# 0.20fF
C908 a_29_n444# a_n1555_n1061# 0.21fF
C909 a_n149_n444# a_n1555_n1061# 0.21fF
C910 a_n327_n444# a_n1555_n1061# 0.21fF
C911 a_n505_n444# a_n1555_n1061# 0.21fF
C912 a_n683_n444# a_n1555_n1061# 0.21fF
C913 a_n861_n444# a_n1555_n1061# 0.21fF
C914 a_n1039_n444# a_n1555_n1061# 0.22fF
C915 a_n1217_n444# a_n1555_n1061# 0.27fF
C916 a_1217_109# a_n1555_n1061# 0.10fF
C917 a_1039_109# a_n1555_n1061# 0.05fF
C918 a_861_109# a_n1555_n1061# 0.04fF
C919 a_683_109# a_n1555_n1061# 0.03fF
C920 a_505_109# a_n1555_n1061# 0.03fF
C921 a_327_109# a_n1555_n1061# 0.03fF
C922 a_149_109# a_n1555_n1061# 0.03fF
C923 a_n29_109# a_n1555_n1061# 0.03fF
C924 a_n207_109# a_n1555_n1061# 0.03fF
C925 a_n385_109# a_n1555_n1061# 0.03fF
C926 a_n563_109# a_n1555_n1061# 0.03fF
C927 a_n741_109# a_n1555_n1061# 0.03fF
C928 a_n919_109# a_n1555_n1061# 0.04fF
C929 a_n1097_109# a_n1555_n1061# 0.06fF
C930 a_n1275_109# a_n1555_n1061# 0.10fF
C931 a_1097_54# a_n1555_n1061# 0.23fF
C932 a_919_54# a_n1555_n1061# 0.20fF
C933 a_741_54# a_n1555_n1061# 0.20fF
C934 a_563_54# a_n1555_n1061# 0.20fF
C935 a_385_54# a_n1555_n1061# 0.21fF
C936 a_207_54# a_n1555_n1061# 0.21fF
C937 a_29_54# a_n1555_n1061# 0.22fF
C938 a_n149_54# a_n1555_n1061# 0.22fF
C939 a_n327_54# a_n1555_n1061# 0.22fF
C940 a_n505_54# a_n1555_n1061# 0.22fF
C941 a_n683_54# a_n1555_n1061# 0.22fF
C942 a_n861_54# a_n1555_n1061# 0.23fF
C943 a_n1039_54# a_n1555_n1061# 0.23fF
C944 a_n1217_54# a_n1555_n1061# 0.28fF
C945 a_1217_607# a_n1555_n1061# 0.10fF
C946 a_1039_607# a_n1555_n1061# 0.06fF
C947 a_861_607# a_n1555_n1061# 0.05fF
C948 a_683_607# a_n1555_n1061# 0.04fF
C949 a_505_607# a_n1555_n1061# 0.03fF
C950 a_327_607# a_n1555_n1061# 0.03fF
C951 a_149_607# a_n1555_n1061# 0.03fF
C952 a_n29_607# a_n1555_n1061# 0.04fF
C953 a_n207_607# a_n1555_n1061# 0.03fF
C954 a_n385_607# a_n1555_n1061# 0.03fF
C955 a_n563_607# a_n1555_n1061# 0.03fF
C956 a_n741_607# a_n1555_n1061# 0.04fF
C957 a_n919_607# a_n1555_n1061# 0.05fF
C958 a_n1097_607# a_n1555_n1061# 0.06fF
C959 a_n1275_607# a_n1555_n1061# 0.10fF
C960 a_1097_552# a_n1555_n1061# 0.30fF
C961 a_919_552# a_n1555_n1061# 0.26fF
C962 a_741_552# a_n1555_n1061# 0.26fF
C963 a_563_552# a_n1555_n1061# 0.27fF
C964 a_385_552# a_n1555_n1061# 0.27fF
C965 a_207_552# a_n1555_n1061# 0.28fF
C966 a_29_552# a_n1555_n1061# 0.29fF
C967 a_n149_552# a_n1555_n1061# 0.29fF
C968 a_n327_552# a_n1555_n1061# 0.29fF
C969 a_n505_552# a_n1555_n1061# 0.29fF
C970 a_n683_552# a_n1555_n1061# 0.29fF
C971 a_n861_552# a_n1555_n1061# 0.29fF
C972 a_n1039_552# a_n1555_n1061# 0.30fF
C973 a_n1217_552# a_n1555_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EL6FQZ a_n1008_n140# a_n594_n195# a_1306_n140# a_n652_n140#
+ a_652_n195# a_772_n140# a_n1662_n195# a_n1720_n140# a_n60_n195# a_2076_n195# a_2196_n140#
+ a_n474_n140# a_1008_n195# a_n416_n195# a_1128_n140# a_474_n195# a_594_n140# a_n1484_n195#
+ a_n1542_n140# a_1720_n195# a_1840_n140# a_n296_n140# a_n1898_n140# a_n238_n195#
+ a_2018_n140# a_60_n140# a_296_n195# a_n1364_n140# a_n1306_n195# a_416_n140# a_1542_n195#
+ a_n2432_n140# a_1662_n140# a_n950_n195# a_1898_n195# a_n118_n140# a_118_n195# a_n2196_n195#
+ a_238_n140# a_n1186_n140# a_n2254_n140# a_1364_n195# a_n1128_n195# a_n772_n195#
+ a_1484_n140# a_n830_n140# a_830_n195# a_950_n140# a_n1840_n195# a_n2076_n140# a_2254_n195#
+ a_1186_n195# a_n2018_n195# VSUBS
X0 a_2254_n195# a_2254_n195# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1128_n140# a_1008_n195# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n1186_n140# a_n1306_n195# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_772_n140# a_652_n195# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_1662_n140# a_1542_n195# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n118_n140# a_n238_n195# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_2196_n140# a_2076_n195# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2254_n140# a_n2432_n140# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n652_n140# a_n772_n195# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_2018_n140# a_1898_n195# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1008_n140# a_n1128_n195# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_594_n140# a_474_n195# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_60_n140# a_n60_n195# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1484_n140# a_1364_n195# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1542_n140# a_n1662_n195# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_950_n140# a_830_n195# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n2076_n140# a_n2196_n195# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_n830_n140# a_n950_n195# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n474_n140# a_n594_n195# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_1840_n140# a_1720_n195# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_416_n140# a_296_n195# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n1898_n140# a_n2018_n195# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n296_n140# a_n416_n195# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_1306_n140# a_1186_n195# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1720_n140# a_n1840_n195# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n1364_n140# a_n1484_n195# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_238_n140# a_118_n195# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n296_n140# a_n652_n140# 0.03fF
C1 a_1898_n195# a_1186_n195# 0.01fF
C2 a_2254_n195# a_1008_n195# 0.00fF
C3 a_594_n140# a_60_n140# 0.02fF
C4 a_1186_n195# a_1008_n195# 0.10fF
C5 a_238_n140# a_n118_n140# 0.03fF
C6 a_n296_n140# a_n474_n140# 0.06fF
C7 a_1128_n140# a_950_n140# 0.06fF
C8 a_n830_n140# a_772_n140# 0.01fF
C9 a_n830_n140# a_n1720_n140# 0.01fF
C10 a_n2018_n195# a_n772_n195# 0.01fF
C11 a_n2196_n195# a_n594_n195# 0.01fF
C12 a_n1840_n195# a_n238_n195# 0.01fF
C13 a_n594_n195# a_830_n195# 0.01fF
C14 a_n416_n195# a_830_n195# 0.01fF
C15 a_n1186_n140# a_n1008_n140# 0.06fF
C16 a_1128_n140# a_1306_n140# 0.06fF
C17 a_n60_n195# a_n950_n195# 0.01fF
C18 a_n1364_n140# a_n118_n140# 0.01fF
C19 a_n1186_n140# a_n652_n140# 0.02fF
C20 a_n1542_n140# a_n1364_n140# 0.06fF
C21 a_2254_n195# a_1720_n195# 0.01fF
C22 a_238_n140# a_1662_n140# 0.01fF
C23 a_1128_n140# a_n296_n140# 0.01fF
C24 a_1720_n195# a_1186_n195# 0.02fF
C25 a_n1840_n195# a_n1128_n195# 0.01fF
C26 a_n60_n195# a_1542_n195# 0.01fF
C27 a_n60_n195# a_296_n195# 0.03fF
C28 a_n474_n140# a_n1186_n140# 0.01fF
C29 a_1128_n140# a_1484_n140# 0.03fF
C30 a_n830_n140# a_n2254_n140# 0.01fF
C31 a_1306_n140# a_950_n140# 0.03fF
C32 a_n1720_n140# a_n1008_n140# 0.01fF
C33 a_772_n140# a_n652_n140# 0.01fF
C34 a_n2018_n195# a_n2196_n195# 0.10fF
C35 a_n1720_n140# a_n652_n140# 0.01fF
C36 a_474_n195# a_1898_n195# 0.01fF
C37 a_2254_n195# a_1542_n195# 0.01fF
C38 a_1542_n195# a_1186_n195# 0.03fF
C39 a_n296_n140# a_950_n140# 0.01fF
C40 a_296_n195# a_1186_n195# 0.01fF
C41 a_474_n195# a_1008_n195# 0.02fF
C42 a_238_n140# a_594_n140# 0.03fF
C43 a_1484_n140# a_950_n140# 0.02fF
C44 a_772_n140# a_n474_n140# 0.01fF
C45 a_n2432_n140# a_n1306_n195# 0.01fF
C46 a_n1720_n140# a_n474_n140# 0.01fF
C47 a_n1840_n195# a_n594_n195# 0.01fF
C48 a_n2196_n195# a_n772_n195# 0.01fF
C49 a_n238_n195# a_1008_n195# 0.01fF
C50 a_n1840_n195# a_n416_n195# 0.01fF
C51 a_1128_n140# a_1840_n140# 0.01fF
C52 a_n296_n140# a_1306_n140# 0.01fF
C53 a_n830_n140# a_416_n140# 0.01fF
C54 a_n772_n195# a_830_n195# 0.01fF
C55 a_1484_n140# a_1306_n140# 0.06fF
C56 a_2076_n195# a_1898_n195# 0.10fF
C57 a_n1186_n140# a_n2076_n140# 0.01fF
C58 a_n2254_n140# a_n1008_n140# 0.01fF
C59 a_n1484_n195# a_n1662_n195# 0.10fF
C60 a_n2254_n140# a_n652_n140# 0.01fF
C61 a_2076_n195# a_1008_n195# 0.01fF
C62 a_n950_n195# a_n1306_n195# 0.03fF
C63 a_1128_n140# a_772_n140# 0.03fF
C64 a_474_n195# a_1720_n195# 0.01fF
C65 a_n1542_n140# a_n118_n140# 0.01fF
C66 a_n1484_n195# a_118_n195# 0.01fF
C67 a_1898_n195# a_1364_n195# 0.02fF
C68 a_1840_n140# a_950_n140# 0.01fF
C69 a_n2432_n140# a_n830_n140# 0.01fF
C70 a_1364_n195# a_1008_n195# 0.03fF
C71 a_296_n195# a_n1306_n195# 0.01fF
C72 a_474_n195# a_n950_n195# 0.01fF
C73 a_n1720_n140# a_n2076_n140# 0.03fF
C74 a_1840_n140# a_1306_n140# 0.02fF
C75 a_n2432_n140# a_n1128_n195# 0.00fF
C76 a_n1840_n195# a_n2018_n195# 0.10fF
C77 a_n1008_n140# a_416_n140# 0.01fF
C78 a_n296_n140# a_n1186_n140# 0.01fF
C79 a_474_n195# a_1542_n195# 0.01fF
C80 a_2076_n195# a_1720_n195# 0.03fF
C81 a_n238_n195# a_n950_n195# 0.01fF
C82 a_772_n140# a_950_n140# 0.06fF
C83 a_474_n195# a_296_n195# 0.10fF
C84 a_416_n140# a_n652_n140# 0.01fF
C85 a_1840_n140# a_1484_n140# 0.03fF
C86 a_n594_n195# a_1008_n195# 0.01fF
C87 a_n474_n140# a_416_n140# 0.01fF
C88 a_n1840_n195# a_n772_n195# 0.01fF
C89 a_n238_n195# a_296_n195# 0.02fF
C90 a_772_n140# a_1306_n140# 0.02fF
C91 a_n416_n195# a_1008_n195# 0.01fF
C92 a_n830_n140# a_60_n140# 0.01fF
C93 a_n830_n140# a_n1898_n140# 0.01fF
C94 a_1364_n195# a_1720_n195# 0.03fF
C95 a_2018_n140# a_1128_n140# 0.01fF
C96 a_n950_n195# a_n1128_n195# 0.10fF
C97 a_n2254_n140# a_n2076_n140# 0.06fF
C98 a_2076_n195# a_1542_n195# 0.02fF
C99 a_772_n140# a_n296_n140# 0.01fF
C100 a_n2432_n140# a_n1008_n140# 0.01fF
C101 a_n296_n140# a_n1720_n140# 0.01fF
C102 a_n118_n140# a_594_n140# 0.01fF
C103 a_772_n140# a_1484_n140# 0.01fF
C104 a_296_n195# a_n1128_n195# 0.01fF
C105 a_n1484_n195# a_n60_n195# 0.01fF
C106 a_118_n195# a_652_n195# 0.02fF
C107 a_1128_n140# a_416_n140# 0.01fF
C108 a_1542_n195# a_1364_n195# 0.10fF
C109 a_296_n195# a_1364_n195# 0.01fF
C110 a_2018_n140# a_950_n140# 0.01fF
C111 a_n1008_n140# a_60_n140# 0.01fF
C112 a_n1840_n195# a_n2196_n195# 0.03fF
C113 a_594_n140# a_1662_n140# 0.01fF
C114 a_n1008_n140# a_n1898_n140# 0.01fF
C115 a_n1720_n140# a_n1186_n140# 0.02fF
C116 a_n594_n195# a_n950_n195# 0.03fF
C117 a_2018_n140# a_1306_n140# 0.01fF
C118 a_n652_n140# a_60_n140# 0.01fF
C119 a_n416_n195# a_n950_n195# 0.02fF
C120 a_n1898_n140# a_n652_n140# 0.01fF
C121 a_772_n140# a_1840_n140# 0.01fF
C122 a_416_n140# a_950_n140# 0.02fF
C123 a_n474_n140# a_60_n140# 0.02fF
C124 a_296_n195# a_n594_n195# 0.01fF
C125 a_n60_n195# a_n1662_n195# 0.01fF
C126 a_n474_n140# a_n1898_n140# 0.01fF
C127 a_n416_n195# a_296_n195# 0.01fF
C128 a_n2432_n140# a_n2018_n195# 0.02fF
C129 a_2018_n140# a_1484_n140# 0.02fF
C130 a_n830_n140# a_238_n140# 0.01fF
C131 a_1306_n140# a_416_n140# 0.01fF
C132 a_118_n195# a_n60_n195# 0.10fF
C133 a_n2432_n140# a_n2076_n140# 0.03fF
C134 a_n1186_n140# a_n2254_n140# 0.01fF
C135 a_n2432_n140# a_n772_n195# 0.00fF
C136 a_n296_n140# a_416_n140# 0.01fF
C137 a_2196_n140# a_1662_n140# 0.02fF
C138 a_1484_n140# a_416_n140# 0.01fF
C139 a_n60_n195# a_652_n195# 0.01fF
C140 a_1128_n140# a_60_n140# 0.01fF
C141 a_n830_n140# a_n1364_n140# 0.02fF
C142 a_n2018_n195# a_n950_n195# 0.01fF
C143 a_n1484_n195# a_n1306_n195# 0.10fF
C144 a_118_n195# a_1186_n195# 0.01fF
C145 a_2254_n195# a_1662_n140# 0.01fF
C146 a_2018_n140# a_1840_n140# 0.06fF
C147 a_1898_n195# a_830_n195# 0.01fF
C148 a_n2076_n140# a_n1898_n140# 0.06fF
C149 a_2254_n195# a_652_n195# 0.00fF
C150 a_n1720_n140# a_n2254_n140# 0.02fF
C151 a_n772_n195# a_n950_n195# 0.10fF
C152 a_238_n140# a_n1008_n140# 0.01fF
C153 a_652_n195# a_1186_n195# 0.02fF
C154 a_830_n195# a_1008_n195# 0.10fF
C155 a_n1186_n140# a_416_n140# 0.01fF
C156 a_238_n140# a_n652_n140# 0.01fF
C157 a_594_n140# a_2196_n140# 0.01fF
C158 a_950_n140# a_60_n140# 0.01fF
C159 a_2018_n140# a_772_n140# 0.01fF
C160 a_n238_n195# a_n1484_n195# 0.01fF
C161 a_1840_n140# a_416_n140# 0.01fF
C162 a_296_n195# a_n772_n195# 0.01fF
C163 a_238_n140# a_n474_n140# 0.01fF
C164 a_n2432_n140# a_n2196_n195# 0.06fF
C165 a_1306_n140# a_60_n140# 0.01fF
C166 a_n1364_n140# a_n1008_n140# 0.03fF
C167 a_n1662_n195# a_n1306_n195# 0.03fF
C168 a_n1364_n140# a_n652_n140# 0.01fF
C169 a_118_n195# a_n1306_n195# 0.01fF
C170 a_n296_n140# a_60_n140# 0.03fF
C171 a_772_n140# a_416_n140# 0.03fF
C172 a_n2432_n140# a_n1186_n140# 0.01fF
C173 a_n1484_n195# a_n1128_n195# 0.03fF
C174 a_n296_n140# a_n1898_n140# 0.01fF
C175 a_830_n195# a_1720_n195# 0.01fF
C176 a_n1364_n140# a_n474_n140# 0.01fF
C177 a_1484_n140# a_60_n140# 0.01fF
C178 a_n830_n140# a_n118_n140# 0.01fF
C179 a_n2196_n195# a_n950_n195# 0.01fF
C180 a_1128_n140# a_238_n140# 0.01fF
C181 a_118_n195# a_474_n195# 0.03fF
C182 a_n60_n195# a_1186_n195# 0.01fF
C183 a_n238_n195# a_n1662_n195# 0.01fF
C184 a_n1542_n140# a_n830_n140# 0.01fF
C185 a_2254_n195# a_2196_n140# 0.06fF
C186 a_n238_n195# a_118_n195# 0.03fF
C187 a_1542_n195# a_830_n195# 0.01fF
C188 a_474_n195# a_652_n195# 0.10fF
C189 a_296_n195# a_830_n195# 0.02fF
C190 a_n2432_n140# a_n1720_n140# 0.01fF
C191 a_n1186_n140# a_60_n140# 0.01fF
C192 a_n1186_n140# a_n1898_n140# 0.01fF
C193 a_2254_n195# a_1186_n195# 0.01fF
C194 a_n1662_n195# a_n1128_n195# 0.02fF
C195 a_n1484_n195# a_n594_n195# 0.01fF
C196 a_238_n140# a_950_n140# 0.01fF
C197 a_n416_n195# a_n1484_n195# 0.01fF
C198 a_n238_n195# a_652_n195# 0.01fF
C199 a_n2432_n140# a_n1840_n195# 0.01fF
C200 a_2018_n140# a_416_n140# 0.01fF
C201 a_118_n195# a_n1128_n195# 0.01fF
C202 a_n1364_n140# a_n2076_n140# 0.01fF
C203 a_n118_n140# a_n1008_n140# 0.01fF
C204 a_238_n140# a_1306_n140# 0.01fF
C205 a_2076_n195# a_652_n195# 0.01fF
C206 a_n118_n140# a_n652_n140# 0.02fF
C207 a_118_n195# a_1364_n195# 0.01fF
C208 a_n1542_n140# a_n1008_n140# 0.02fF
C209 a_n60_n195# a_n1306_n195# 0.01fF
C210 a_772_n140# a_60_n140# 0.01fF
C211 a_n2432_n140# a_n2254_n140# 0.06fF
C212 a_n1542_n140# a_n652_n140# 0.01fF
C213 a_n1720_n140# a_n1898_n140# 0.06fF
C214 a_238_n140# a_n296_n140# 0.02fF
C215 a_n118_n140# a_n474_n140# 0.03fF
C216 a_238_n140# a_1484_n140# 0.01fF
C217 a_n830_n140# a_594_n140# 0.01fF
C218 a_n1840_n195# a_n950_n195# 0.01fF
C219 a_n1542_n140# a_n474_n140# 0.01fF
C220 a_1364_n195# a_652_n195# 0.01fF
C221 a_n60_n195# a_474_n195# 0.02fF
C222 a_n1662_n195# a_n594_n195# 0.01fF
C223 a_n416_n195# a_n1662_n195# 0.01fF
C224 a_1898_n195# a_1008_n195# 0.01fF
C225 a_n1484_n195# a_n2018_n195# 0.02fF
C226 a_n1364_n140# a_n296_n140# 0.01fF
C227 a_118_n195# a_n594_n195# 0.01fF
C228 a_n416_n195# a_118_n195# 0.02fF
C229 a_n238_n195# a_n60_n195# 0.10fF
C230 a_n2254_n140# a_n1898_n140# 0.03fF
C231 a_238_n140# a_n1186_n140# 0.01fF
C232 a_1128_n140# a_n118_n140# 0.01fF
C233 a_474_n195# a_1186_n195# 0.01fF
C234 a_n1484_n195# a_n772_n195# 0.01fF
C235 a_n594_n195# a_652_n195# 0.01fF
C236 a_n416_n195# a_652_n195# 0.01fF
C237 a_1840_n140# a_238_n140# 0.01fF
C238 a_n60_n195# a_n1128_n195# 0.01fF
C239 a_n238_n195# a_1186_n195# 0.01fF
C240 a_594_n140# a_n1008_n140# 0.01fF
C241 a_1898_n195# a_1720_n195# 0.10fF
C242 a_n1364_n140# a_n1186_n140# 0.06fF
C243 a_594_n140# a_n652_n140# 0.01fF
C244 a_1720_n195# a_1008_n195# 0.01fF
C245 a_n1542_n140# a_n2076_n140# 0.02fF
C246 a_n60_n195# a_1364_n195# 0.01fF
C247 a_n1662_n195# a_n2018_n195# 0.03fF
C248 a_2254_n195# a_2076_n195# 0.06fF
C249 a_n118_n140# a_950_n140# 0.01fF
C250 a_772_n140# a_238_n140# 0.02fF
C251 a_2076_n195# a_1186_n195# 0.01fF
C252 a_1128_n140# a_1662_n140# 0.02fF
C253 a_416_n140# a_60_n140# 0.03fF
C254 a_594_n140# a_n474_n140# 0.01fF
C255 a_n1662_n195# a_n772_n195# 0.01fF
C256 a_n118_n140# a_1306_n140# 0.01fF
C257 a_1898_n195# a_1542_n195# 0.03fF
C258 a_2254_n195# a_1364_n195# 0.01fF
C259 a_296_n195# a_1898_n195# 0.01fF
C260 a_n1484_n195# a_n2196_n195# 0.01fF
C261 a_1542_n195# a_1008_n195# 0.02fF
C262 a_1364_n195# a_1186_n195# 0.10fF
C263 a_n1364_n140# a_n1720_n140# 0.03fF
C264 a_118_n195# a_n772_n195# 0.01fF
C265 a_n60_n195# a_n594_n195# 0.02fF
C266 a_296_n195# a_1008_n195# 0.01fF
C267 a_n416_n195# a_n60_n195# 0.03fF
C268 a_n296_n140# a_n118_n140# 0.06fF
C269 a_n2432_n140# a_n950_n195# 0.00fF
C270 a_n118_n140# a_1484_n140# 0.01fF
C271 a_1662_n140# a_950_n140# 0.01fF
C272 a_n1542_n140# a_n296_n140# 0.01fF
C273 a_n238_n195# a_n1306_n195# 0.01fF
C274 a_1128_n140# a_594_n140# 0.02fF
C275 a_n2432_n140# a_n1898_n140# 0.02fF
C276 a_n772_n195# a_652_n195# 0.01fF
C277 a_1306_n140# a_1662_n140# 0.03fF
C278 a_n238_n195# a_474_n195# 0.01fF
C279 a_n416_n195# a_1186_n195# 0.01fF
C280 a_1542_n195# a_1720_n195# 0.10fF
C281 a_n1364_n140# a_n2254_n140# 0.01fF
C282 a_n1128_n195# a_n1306_n195# 0.10fF
C283 a_296_n195# a_1720_n195# 0.01fF
C284 a_n118_n140# a_n1186_n140# 0.01fF
C285 a_n1662_n195# a_n2196_n195# 0.02fF
C286 a_1484_n140# a_1662_n140# 0.06fF
C287 a_594_n140# a_950_n140# 0.03fF
C288 a_474_n195# a_2076_n195# 0.01fF
C289 a_n1542_n140# a_n1186_n140# 0.03fF
C290 a_238_n140# a_416_n140# 0.06fF
C291 a_296_n195# a_n950_n195# 0.01fF
C292 a_474_n195# a_n1128_n195# 0.01fF
C293 a_118_n195# a_830_n195# 0.01fF
C294 a_1128_n140# a_2196_n140# 0.01fF
C295 a_594_n140# a_1306_n140# 0.01fF
C296 a_296_n195# a_1542_n195# 0.01fF
C297 a_474_n195# a_1364_n195# 0.01fF
C298 a_n1840_n195# a_n1484_n195# 0.03fF
C299 a_n238_n195# a_n1128_n195# 0.01fF
C300 a_1128_n140# a_2254_n195# 0.01fF
C301 a_n60_n195# a_n772_n195# 0.01fF
C302 a_772_n140# a_n118_n140# 0.01fF
C303 a_n296_n140# a_594_n140# 0.01fF
C304 a_n1720_n140# a_n118_n140# 0.01fF
C305 a_830_n195# a_652_n195# 0.10fF
C306 a_594_n140# a_1484_n140# 0.01fF
C307 a_n594_n195# a_n1306_n195# 0.01fF
C308 a_n1542_n140# a_n1720_n140# 0.06fF
C309 a_n238_n195# a_1364_n195# 0.01fF
C310 a_n416_n195# a_n1306_n195# 0.01fF
C311 a_1840_n140# a_1662_n140# 0.06fF
C312 a_2196_n140# a_950_n140# 0.01fF
C313 a_2076_n195# a_1364_n195# 0.01fF
C314 a_474_n195# a_n594_n195# 0.01fF
C315 a_n416_n195# a_474_n195# 0.01fF
C316 a_2254_n195# a_950_n140# 0.01fF
C317 a_1306_n140# a_2196_n140# 0.01fF
C318 a_772_n140# a_1662_n140# 0.01fF
C319 a_n2432_n140# a_n1364_n140# 0.01fF
C320 a_n238_n195# a_n594_n195# 0.03fF
C321 a_n1840_n195# a_n1662_n195# 0.10fF
C322 a_n238_n195# a_n416_n195# 0.10fF
C323 a_2254_n195# a_1306_n140# 0.01fF
C324 a_n1542_n140# a_n2254_n140# 0.01fF
C325 a_1840_n140# a_594_n140# 0.01fF
C326 a_n830_n140# a_n1008_n140# 0.06fF
C327 a_1484_n140# a_2196_n140# 0.01fF
C328 a_238_n140# a_60_n140# 0.06fF
C329 a_n830_n140# a_n652_n140# 0.06fF
C330 a_n60_n195# a_830_n195# 0.01fF
C331 a_n2018_n195# a_n1306_n195# 0.01fF
C332 a_2254_n195# a_1484_n140# 0.01fF
C333 a_n830_n140# a_n474_n140# 0.03fF
C334 a_n594_n195# a_n1128_n195# 0.02fF
C335 a_n416_n195# a_n1128_n195# 0.01fF
C336 a_772_n140# a_594_n140# 0.06fF
C337 a_n1364_n140# a_60_n140# 0.01fF
C338 a_n1364_n140# a_n1898_n140# 0.02fF
C339 a_n118_n140# a_416_n140# 0.02fF
C340 a_n772_n195# a_n1306_n195# 0.02fF
C341 a_2254_n195# a_830_n195# 0.00fF
C342 a_830_n195# a_1186_n195# 0.03fF
C343 a_2018_n140# a_1662_n140# 0.03fF
C344 a_n2432_n140# a_n1484_n195# 0.01fF
C345 a_1840_n140# a_2196_n140# 0.03fF
C346 a_474_n195# a_n772_n195# 0.01fF
C347 a_n1008_n140# a_n652_n140# 0.03fF
C348 a_1840_n140# a_2254_n195# 0.02fF
C349 a_n416_n195# a_n594_n195# 0.10fF
C350 a_n238_n195# a_n772_n195# 0.02fF
C351 a_n474_n140# a_n1008_n140# 0.02fF
C352 a_772_n140# a_2196_n140# 0.01fF
C353 a_416_n140# a_1662_n140# 0.01fF
C354 a_n474_n140# a_n652_n140# 0.06fF
C355 a_n2018_n195# a_n1128_n195# 0.01fF
C356 a_n830_n140# a_n2076_n140# 0.01fF
C357 a_n2432_n140# a_n1542_n140# 0.01fF
C358 a_118_n195# a_1008_n195# 0.01fF
C359 a_n1484_n195# a_n950_n195# 0.02fF
C360 a_2018_n140# a_594_n140# 0.01fF
C361 a_772_n140# a_2254_n195# 0.01fF
C362 a_n2196_n195# a_n1306_n195# 0.01fF
C363 a_n2432_n140# a_n1662_n195# 0.01fF
C364 a_1898_n195# a_652_n195# 0.01fF
C365 a_n772_n195# a_n1128_n195# 0.03fF
C366 a_652_n195# a_1008_n195# 0.03fF
C367 a_594_n140# a_416_n140# 0.06fF
C368 a_n118_n140# a_60_n140# 0.06fF
C369 a_n1364_n140# a_238_n140# 0.01fF
C370 a_474_n195# a_830_n195# 0.03fF
C371 a_n1542_n140# a_60_n140# 0.01fF
C372 a_n1542_n140# a_n1898_n140# 0.03fF
C373 a_118_n195# a_1720_n195# 0.01fF
C374 a_n830_n140# a_n296_n140# 0.02fF
C375 a_n2018_n195# a_n594_n195# 0.01fF
C376 a_n416_n195# a_n2018_n195# 0.01fF
C377 a_1128_n140# a_n474_n140# 0.01fF
C378 a_n1662_n195# a_n950_n195# 0.01fF
C379 a_n1008_n140# a_n2076_n140# 0.01fF
C380 a_2018_n140# a_2196_n140# 0.06fF
C381 a_n238_n195# a_830_n195# 0.01fF
C382 a_n2076_n140# a_n652_n140# 0.01fF
C383 a_118_n195# a_n950_n195# 0.01fF
C384 a_652_n195# a_1720_n195# 0.01fF
C385 a_n594_n195# a_n772_n195# 0.10fF
C386 a_2018_n140# a_2254_n195# 0.03fF
C387 a_1662_n140# a_60_n140# 0.01fF
C388 a_n652_n140# a_950_n140# 0.01fF
C389 a_n416_n195# a_n772_n195# 0.03fF
C390 a_n474_n140# a_n2076_n140# 0.01fF
C391 a_2076_n195# a_830_n195# 0.01fF
C392 a_118_n195# a_1542_n195# 0.01fF
C393 a_n2196_n195# a_n1128_n195# 0.01fF
C394 a_118_n195# a_296_n195# 0.10fF
C395 a_n60_n195# a_1008_n195# 0.01fF
C396 a_n950_n195# a_652_n195# 0.01fF
C397 a_n474_n140# a_950_n140# 0.01fF
C398 a_n830_n140# a_n1186_n140# 0.03fF
C399 a_n1840_n195# a_n1306_n195# 0.02fF
C400 a_1364_n195# a_830_n195# 0.02fF
C401 a_1542_n195# a_652_n195# 0.01fF
C402 a_n296_n140# a_n1008_n140# 0.01fF
C403 a_296_n195# a_652_n195# 0.03fF
C404 a_2254_n195# a_1898_n195# 0.02fF
C405 a_2196_n140# VSUBS 0.01fF
C406 a_2018_n140# VSUBS 0.01fF
C407 a_1840_n140# VSUBS 0.02fF
C408 a_1662_n140# VSUBS 0.02fF
C409 a_1484_n140# VSUBS 0.02fF
C410 a_1306_n140# VSUBS 0.02fF
C411 a_1128_n140# VSUBS 0.02fF
C412 a_950_n140# VSUBS 0.02fF
C413 a_772_n140# VSUBS 0.02fF
C414 a_594_n140# VSUBS 0.02fF
C415 a_416_n140# VSUBS 0.02fF
C416 a_238_n140# VSUBS 0.02fF
C417 a_60_n140# VSUBS 0.02fF
C418 a_n118_n140# VSUBS 0.02fF
C419 a_n296_n140# VSUBS 0.02fF
C420 a_n474_n140# VSUBS 0.02fF
C421 a_n652_n140# VSUBS 0.02fF
C422 a_n830_n140# VSUBS 0.02fF
C423 a_n1008_n140# VSUBS 0.02fF
C424 a_n1186_n140# VSUBS 0.02fF
C425 a_n1364_n140# VSUBS 0.02fF
C426 a_n1542_n140# VSUBS 0.02fF
C427 a_n1720_n140# VSUBS 0.02fF
C428 a_n1898_n140# VSUBS 0.02fF
C429 a_n2076_n140# VSUBS 0.02fF
C430 a_n2254_n140# VSUBS 0.02fF
C431 a_2254_n195# VSUBS 0.31fF
C432 a_2076_n195# VSUBS 0.19fF
C433 a_1898_n195# VSUBS 0.20fF
C434 a_1720_n195# VSUBS 0.21fF
C435 a_1542_n195# VSUBS 0.22fF
C436 a_1364_n195# VSUBS 0.23fF
C437 a_1186_n195# VSUBS 0.23fF
C438 a_1008_n195# VSUBS 0.24fF
C439 a_830_n195# VSUBS 0.24fF
C440 a_652_n195# VSUBS 0.24fF
C441 a_474_n195# VSUBS 0.24fF
C442 a_296_n195# VSUBS 0.24fF
C443 a_118_n195# VSUBS 0.24fF
C444 a_n60_n195# VSUBS 0.24fF
C445 a_n238_n195# VSUBS 0.24fF
C446 a_n416_n195# VSUBS 0.24fF
C447 a_n594_n195# VSUBS 0.24fF
C448 a_n772_n195# VSUBS 0.24fF
C449 a_n950_n195# VSUBS 0.24fF
C450 a_n1128_n195# VSUBS 0.24fF
C451 a_n1306_n195# VSUBS 0.24fF
C452 a_n1484_n195# VSUBS 0.24fF
C453 a_n1662_n195# VSUBS 0.24fF
C454 a_n1840_n195# VSUBS 0.24fF
C455 a_n2018_n195# VSUBS 0.24fF
C456 a_n2196_n195# VSUBS 0.24fF
C457 a_n2432_n140# VSUBS 0.36fF
.ends

.subckt bias_circuit bias_c bias_e i_bias VDD m1_1243_5997# m1_3443_5997# m1_5643_5997#
+ bias_a m1_7347_1428# m1_7639_1420# m1_7169_923# m1_3551_3596# m1_7461_921# m1_7347_423#
+ m1_7639_427# bias_b VSS bias_d
Xsky130_fd_pr__nfet_01v8_6RUDQZ_0 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_1 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_2 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_3 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_SD55Q9_0 m1_7347_1428# bias_e m1_7639_1420# bias_e m1_7055_1417#
+ m1_6763_422# bias_e bias_e m1_6471_422# VSS VSS VSS m1_7639_427# m1_7347_423# bias_e
+ m1_7055_433# bias_e bias_e m1_6763_422# bias_e m1_6471_422# m1_7169_923# bias_e
+ bias_e m1_7461_921# m1_7639_427# m1_7347_423# m1_6877_922# m1_7055_433# bias_e VSS
+ bias_e bias_e bias_e VSS VSS bias_e m1_6877_922# m1_6585_923# bias_e VSS m1_6763_1422#
+ m1_6293_922# m1_6471_1426# bias_e m1_7347_1428# bias_e bias_e m1_7639_1420# m1_7169_923#
+ m1_7055_1417# bias_e bias_e m1_7461_921# bias_e bias_e m1_6585_923# bias_e m1_6293_922#
+ m1_6763_1422# bias_e m1_6471_1426# VSS sky130_fd_pr__nfet_01v8_SD55Q9
Xsky130_fd_pr__nfet_01v8_EZNTQN_0 bias_c i_bias i_bias VSS i_bias VSS i_bias VSS VSS
+ bias_c i_bias VSS VSS i_bias i_bias VSS bias_c i_bias i_bias VSS i_bias i_bias bias_c
+ i_bias VSS i_bias i_bias VSS i_bias bias_c i_bias VSS VSS bias_c i_bias VSS i_bias
+ i_bias i_bias VSS i_bias i_bias i_bias i_bias i_bias VSS i_bias i_bias i_bias i_bias
+ i_bias i_bias bias_c i_bias i_bias VSS i_bias i_bias bias_c i_bias i_bias i_bias
+ VSS VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS i_bias i_bias
+ bias_c sky130_fd_pr__nfet_01v8_EZNTQN
Xsky130_fd_pr__pfet_01v8_JJWXCM_0 bias_b bias_c m1_1243_5997# m1_1243_5997# bias_b
+ bias_c VDD VDD bias_c bias_c bias_b bias_c VDD m1_1243_5997# bias_c bias_b VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_1 m1_3551_3596# bias_c m1_3443_5997# m1_3443_5997#
+ m1_3551_3596# bias_c VDD VDD bias_c bias_c m1_3551_3596# bias_c VDD m1_3443_5997#
+ bias_c m1_3551_3596# VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_2 bias_e bias_c m1_5643_5997# m1_5643_5997# bias_e
+ bias_c VDD VDD bias_c bias_c bias_e bias_c VDD m1_5643_5997# bias_c bias_e VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__nfet_01v8_LJREPQ_0 m1_3551_3596# bias_d VSS bias_a bias_d m1_3551_3596#
+ VSS VSS sky130_fd_pr__nfet_01v8_LJREPQ
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_0 m1_1243_5997# bias_b VDD VDD m1_1243_5997# bias_b
+ VDD VDD bias_b bias_b m1_1243_5997# bias_b VDD VDD bias_b m1_1243_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_1 m1_3443_5997# bias_b VDD VDD m1_3443_5997# bias_b
+ VDD VDD bias_b bias_b m1_3443_5997# bias_b VDD VDD bias_b m1_3443_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_2 m1_5643_5997# bias_b VDD VDD m1_5643_5997# bias_b
+ VDD VDD bias_b bias_b m1_5643_5997# bias_b VDD VDD bias_b m1_5643_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__nfet_01v8_lvt_28TRYY_0 bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b VSS bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c
+ bias_b bias_c bias_b bias_b bias_c bias_b bias_b bias_b bias_b bias_c bias_b bias_b
+ bias_b bias_c bias_c bias_b bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_c bias_b bias_b bias_b
+ bias_b bias_c bias_b bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b
+ bias_b bias_b bias_c bias_b bias_b bias_b bias_c bias_b bias_b bias_c bias_b bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_c bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b
+ bias_b bias_b sky130_fd_pr__nfet_01v8_lvt_28TRYY
Xsky130_fd_pr__nfet_01v8_EL6FQZ_0 bias_d m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# bias_d VSS m1_3551_3596# m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
Xsky130_fd_pr__nfet_01v8_EL6FQZ_1 bias_d m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# bias_d VSS m1_3551_3596# m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
C0 m1_6877_922# m1_6293_922# 0.01fF
C1 m1_7055_433# m1_7639_427# 0.01fF
C2 bias_e m1_5643_5997# 0.71fF
C3 m1_6763_1422# m1_6763_422# -0.00fF
C4 bias_a m1_7169_923# 0.00fF
C5 m1_6585_923# m1_7169_923# 0.01fF
C6 bias_a m1_6763_1422# 0.00fF
C7 m1_7461_921# m1_6293_922# 0.01fF
C8 m1_7461_921# m1_6877_922# 0.01fF
C9 m1_7347_1428# m1_6763_1422# 0.01fF
C10 bias_e m1_7055_1417# 0.33fF
C11 i_bias li_3433_399# 0.03fF
C12 m1_7639_427# m1_7347_423# 0.03fF
C13 m1_6471_422# m1_7639_427# 0.01fF
C14 bias_d li_3433_399# 5.36fF
C15 bias_e m1_6763_422# 0.26fF
C16 bias_a m1_7055_1417# 0.00fF
C17 bias_e bias_a 0.24fF
C18 bias_e m1_6585_923# 0.22fF
C19 bias_c VDD 4.90fF
C20 m1_7055_433# m1_7055_1417# -0.00fF
C21 m1_3551_3596# li_3433_399# 0.03fF
C22 m1_7347_1428# m1_7055_1417# 0.03fF
C23 bias_e m1_7055_433# 0.26fF
C24 bias_e m1_7347_1428# 0.32fF
C25 bias_a m1_6763_422# 0.01fF
C26 bias_c m1_3443_5997# 0.44fF
C27 bias_a m1_6585_923# 0.00fF
C28 m1_7055_433# m1_6763_422# 0.03fF
C29 VDD m1_3443_5997# 0.84fF
C30 bias_a m1_7055_433# 0.01fF
C31 m1_6293_922# bias_d 0.00fF
C32 m1_7347_1428# bias_a 0.00fF
C33 m1_6471_1426# m1_7639_1420# 0.01fF
C34 bias_e m1_6471_422# 0.25fF
C35 bias_e m1_7347_423# 0.26fF
C36 bias_c i_bias 5.62fF
C37 bias_c bias_d 0.90fF
C38 bias_e li_3433_399# 0.02fF
C39 m1_6471_422# m1_6763_422# 0.03fF
C40 m1_6763_422# m1_7347_423# 0.01fF
C41 m1_6293_922# m1_7169_923# 0.01fF
C42 m1_6877_922# m1_7169_923# 0.03fF
C43 m1_6471_1426# bias_d 0.01fF
C44 VDD bias_d 0.07fF
C45 bias_a m1_7347_423# 0.01fF
C46 bias_a m1_6471_422# 0.01fF
C47 bias_c m1_3551_3596# 2.13fF
C48 m1_7055_433# m1_7347_423# 0.03fF
C49 m1_6471_422# m1_7055_433# 0.01fF
C50 m1_3443_5997# bias_d 0.03fF
C51 m1_7347_1428# m1_7347_423# -0.00fF
C52 bias_a li_3433_399# 7.53fF
C53 m1_6585_923# li_3433_399# 0.01fF
C54 m1_3551_3596# VDD 0.64fF
C55 m1_7461_921# m1_7169_923# 0.03fF
C56 bias_c bias_b 22.43fF
C57 m1_7639_1420# bias_d 0.00fF
C58 VDD bias_b 8.29fF
C59 m1_3551_3596# m1_3443_5997# 0.98fF
C60 m1_6471_1426# m1_6763_1422# 0.03fF
C61 m1_7639_1420# m1_7639_427# -0.00fF
C62 bias_e m1_6293_922# 0.18fF
C63 bias_e m1_6877_922# 0.22fF
C64 bias_c m1_5643_5997# 0.44fF
C65 m1_3443_5997# bias_b 0.65fF
C66 i_bias bias_d 0.00fF
C67 m1_6471_422# m1_7347_423# 0.01fF
C68 VDD m1_5643_5997# 1.16fF
C69 bias_c m1_1243_5997# 0.52fF
C70 bias_a m1_6293_922# 0.01fF
C71 m1_7639_1420# m1_6763_1422# 0.01fF
C72 m1_6293_922# m1_6585_923# 0.03fF
C73 bias_a m1_6877_922# 0.00fF
C74 m1_6877_922# m1_6585_923# 0.03fF
C75 VDD m1_1243_5997# 1.50fF
C76 bias_e bias_c 0.65fF
C77 m1_7461_921# bias_e 0.21fF
C78 m1_5643_5997# m1_3443_5997# 0.11fF
C79 m1_6471_422# li_3433_399# 0.01fF
C80 m1_6471_1426# m1_7055_1417# 0.01fF
C81 bias_e m1_6471_1426# 0.34fF
C82 bias_e VDD 0.26fF
C83 m1_3551_3596# bias_d 18.83fF
C84 m1_3443_5997# m1_1243_5997# 0.07fF
C85 bias_b i_bias 0.60fF
C86 bias_a bias_c 0.02fF
C87 m1_7461_921# bias_a 0.00fF
C88 m1_7461_921# m1_6585_923# 0.01fF
C89 bias_e m1_3443_5997# 0.02fF
C90 bias_b bias_d 0.26fF
C91 m1_6763_1422# bias_d 0.00fF
C92 bias_a m1_6471_1426# 0.01fF
C93 m1_7639_1420# m1_7055_1417# 0.01fF
C94 bias_e m1_7639_1420# 0.18fF
C95 m1_5643_5997# bias_d 0.03fF
C96 m1_3551_3596# bias_b 0.71fF
C97 m1_7347_1428# m1_6471_1426# 0.01fF
C98 bias_a m1_7639_1420# 0.00fF
C99 m1_6293_922# li_3433_399# 0.02fF
C100 m1_3551_3596# m1_5643_5997# 0.08fF
C101 m1_7055_1417# bias_d 0.00fF
C102 bias_e bias_d 0.26fF
C103 m1_7347_1428# m1_7639_1420# 0.03fF
C104 m1_3551_3596# m1_1243_5997# 0.03fF
C105 m1_5643_5997# bias_b 0.63fF
C106 bias_e m1_7639_427# 0.18fF
C107 bias_a i_bias 0.02fF
C108 m1_6471_1426# m1_6471_422# -0.00fF
C109 bias_e m1_3551_3596# 0.76fF
C110 bias_b m1_1243_5997# 0.77fF
C111 bias_a bias_d 7.33fF
C112 m1_6585_923# bias_d 0.00fF
C113 m1_7639_427# m1_6763_422# 0.01fF
C114 m1_6471_1426# li_3433_399# 0.01fF
C115 bias_e m1_7169_923# 0.22fF
C116 bias_e bias_b 0.07fF
C117 m1_6763_1422# m1_7055_1417# 0.03fF
C118 bias_a m1_7639_427# 0.01fF
C119 m1_7347_1428# bias_d 0.00fF
C120 bias_e m1_6763_1422# 0.33fF
C121 bias_a m1_3551_3596# 0.26fF
C122 m1_3551_3596# VSS -340.55fF
C123 bias_b VSS -284.38fF
C124 m1_5643_5997# VSS 38.06fF
C125 m1_3443_5997# VSS 35.86fF
C126 m1_1243_5997# VSS 25.05fF
C127 VDD VSS 131.72fF
C128 i_bias VSS -60.06fF
C129 bias_c VSS -50.79fF
C130 m1_7639_427# VSS 0.32fF
C131 m1_7347_423# VSS 0.27fF
C132 m1_7461_921# VSS 0.22fF
C133 m1_7169_923# VSS 0.20fF
C134 m1_7055_433# VSS 0.28fF
C135 m1_6763_422# VSS 0.35fF
C136 m1_6471_422# VSS 0.38fF
C137 m1_7639_1420# VSS 0.31fF
C138 m1_7347_1428# VSS 0.20fF
C139 m1_6877_922# VSS 0.21fF
C140 m1_6585_923# VSS 0.29fF
C141 m1_6293_922# VSS 0.32fF
C142 m1_7055_1417# VSS 0.20fF
C143 m1_6763_1422# VSS 0.29fF
C144 m1_6471_1426# VSS 0.30fF
C145 bias_e VSS 7.90fF
C146 bias_d VSS -76.91fF
C147 li_3433_399# VSS 5.57fF
C148 bias_a VSS -48.09fF
.ends

.subckt sky130_fd_pr__pfet_01v8_YVTMSC a_n207_n140# a_29_n205# a_327_n140# a_n683_n205#
+ a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_n505_n205# a_n741_n140# a_563_n205#
+ a_861_n140# a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_683_n140# w_n1133_n241#
+ a_n919_n140# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_861_n140# a_741_n205# a_683_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n205# a_n385_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n741_n140# a_n861_n205# a_n919_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_683_n140# a_563_n205# a_505_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_919_n205# a_919_n205# a_861_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_n29_n140# a_n149_n205# a_n207_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n563_n140# a_n683_n205# a_n741_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_n919_n140# a_n1097_n140# a_n1097_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_505_n140# a_385_n205# a_327_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n505_n205# a_n861_n205# 0.03fF
C1 a_n149_n205# a_n1097_n140# 0.01fF
C2 a_n149_n205# a_919_n205# 0.01fF
C3 a_385_n205# a_207_n205# 0.10fF
C4 a_n683_n205# a_n505_n205# 0.10fF
C5 a_n29_n140# w_n1133_n241# 0.02fF
C6 a_n919_n140# a_505_n140# 0.01fF
C7 a_n563_n140# a_n207_n140# 0.03fF
C8 a_n385_n140# a_683_n140# 0.01fF
C9 a_563_n205# a_n149_n205# 0.01fF
C10 a_n563_n140# a_n1097_n140# 0.02fF
C11 a_207_n205# a_n861_n205# 0.01fF
C12 a_n563_n140# a_n741_n140# 0.06fF
C13 a_n29_n140# a_149_n140# 0.06fF
C14 a_n563_n140# a_919_n205# 0.01fF
C15 a_919_n205# a_741_n205# 0.07fF
C16 a_n327_n205# a_n505_n205# 0.10fF
C17 a_n683_n205# a_207_n205# 0.01fF
C18 a_29_n205# a_n1097_n140# 0.01fF
C19 a_563_n205# a_741_n205# 0.10fF
C20 a_29_n205# a_919_n205# 0.01fF
C21 a_n385_n140# a_n207_n140# 0.06fF
C22 a_683_n140# a_n207_n140# 0.01fF
C23 a_n505_n205# w_n1133_n241# 0.20fF
C24 a_n1097_n140# a_n385_n140# 0.01fF
C25 a_505_n140# a_n563_n140# 0.01fF
C26 a_n741_n140# a_n385_n140# 0.03fF
C27 a_919_n205# a_n385_n140# 0.01fF
C28 a_n741_n140# a_683_n140# 0.01fF
C29 a_563_n205# a_29_n205# 0.02fF
C30 a_919_n205# a_683_n140# 0.03fF
C31 a_327_n140# w_n1133_n241# 0.02fF
C32 a_385_n205# a_n149_n205# 0.02fF
C33 a_n327_n205# a_207_n205# 0.02fF
C34 a_207_n205# w_n1133_n241# 0.17fF
C35 a_n149_n205# a_n861_n205# 0.01fF
C36 a_327_n140# a_149_n140# 0.06fF
C37 a_861_n140# w_n1133_n241# 0.01fF
C38 a_385_n205# a_741_n205# 0.03fF
C39 a_n1097_n140# a_n207_n140# 0.01fF
C40 a_n149_n205# a_n683_n205# 0.02fF
C41 a_n741_n140# a_n207_n140# 0.02fF
C42 a_505_n140# a_n385_n140# 0.01fF
C43 a_919_n205# a_n207_n140# 0.01fF
C44 a_505_n140# a_683_n140# 0.06fF
C45 a_861_n140# a_149_n140# 0.01fF
C46 a_n29_n140# a_327_n140# 0.03fF
C47 a_741_n205# a_n861_n205# 0.01fF
C48 a_n1097_n140# a_n741_n140# 0.03fF
C49 a_385_n205# a_29_n205# 0.03fF
C50 a_n919_n140# w_n1133_n241# 0.02fF
C51 a_n683_n205# a_741_n205# 0.01fF
C52 a_29_n205# a_n861_n205# 0.01fF
C53 a_n149_n205# a_n327_n205# 0.10fF
C54 a_861_n140# a_n29_n140# 0.01fF
C55 a_563_n205# a_n1097_n140# 0.00fF
C56 a_n919_n140# a_149_n140# 0.01fF
C57 a_563_n205# a_919_n205# 0.02fF
C58 a_505_n140# a_n207_n140# 0.01fF
C59 a_n149_n205# w_n1133_n241# 0.19fF
C60 a_29_n205# a_n683_n205# 0.01fF
C61 a_505_n140# a_n1097_n140# 0.01fF
C62 a_505_n140# a_n741_n140# 0.01fF
C63 a_505_n140# a_919_n205# 0.02fF
C64 a_n327_n205# a_741_n205# 0.01fF
C65 a_n919_n140# a_n29_n140# 0.01fF
C66 a_n505_n205# a_207_n205# 0.01fF
C67 a_n563_n140# w_n1133_n241# 0.02fF
C68 a_741_n205# w_n1133_n241# 0.14fF
C69 a_29_n205# a_n327_n205# 0.03fF
C70 a_385_n205# a_n1097_n140# 0.00fF
C71 a_385_n205# a_919_n205# 0.01fF
C72 a_n563_n140# a_149_n140# 0.01fF
C73 a_861_n140# a_327_n140# 0.02fF
C74 a_29_n205# w_n1133_n241# 0.18fF
C75 a_n1097_n140# a_n861_n205# 0.07fF
C76 a_563_n205# a_385_n205# 0.10fF
C77 w_n1133_n241# a_n385_n140# 0.02fF
C78 w_n1133_n241# a_683_n140# 0.01fF
C79 a_n1097_n140# a_n683_n205# 0.02fF
C80 a_n563_n140# a_n29_n140# 0.02fF
C81 a_919_n205# a_n683_n205# 0.00fF
C82 a_n919_n140# a_327_n140# 0.01fF
C83 a_563_n205# a_n861_n205# 0.01fF
C84 a_149_n140# a_n385_n140# 0.02fF
C85 a_149_n140# a_683_n140# 0.02fF
C86 a_n149_n205# a_n505_n205# 0.03fF
C87 a_563_n205# a_n683_n205# 0.01fF
C88 a_n327_n205# a_n1097_n140# 0.01fF
C89 w_n1133_n241# a_n207_n140# 0.02fF
C90 a_n327_n205# a_919_n205# 0.00fF
C91 a_n29_n140# a_n385_n140# 0.03fF
C92 a_n29_n140# a_683_n140# 0.01fF
C93 a_n1097_n140# w_n1133_n241# 0.33fF
C94 a_n505_n205# a_741_n205# 0.01fF
C95 a_n741_n140# w_n1133_n241# 0.02fF
C96 a_919_n205# w_n1133_n241# 0.28fF
C97 a_n149_n205# a_207_n205# 0.03fF
C98 a_149_n140# a_n207_n140# 0.03fF
C99 a_563_n205# a_n327_n205# 0.01fF
C100 a_385_n205# a_n861_n205# 0.01fF
C101 a_n563_n140# a_327_n140# 0.01fF
C102 a_n1097_n140# a_149_n140# 0.01fF
C103 a_29_n205# a_n505_n205# 0.02fF
C104 a_n741_n140# a_149_n140# 0.01fF
C105 a_919_n205# a_149_n140# 0.01fF
C106 a_563_n205# w_n1133_n241# 0.15fF
C107 a_385_n205# a_n683_n205# 0.01fF
C108 a_n29_n140# a_n207_n140# 0.06fF
C109 a_741_n205# a_207_n205# 0.02fF
C110 a_861_n140# a_n563_n140# 0.01fF
C111 a_n683_n205# a_n861_n205# 0.10fF
C112 a_505_n140# w_n1133_n241# 0.02fF
C113 a_n1097_n140# a_n29_n140# 0.01fF
C114 a_n741_n140# a_n29_n140# 0.01fF
C115 a_919_n205# a_n29_n140# 0.01fF
C116 a_29_n205# a_207_n205# 0.10fF
C117 a_327_n140# a_n385_n140# 0.01fF
C118 a_327_n140# a_683_n140# 0.03fF
C119 a_385_n205# a_n327_n205# 0.01fF
C120 a_505_n140# a_149_n140# 0.03fF
C121 a_n919_n140# a_n563_n140# 0.03fF
C122 a_385_n205# w_n1133_n241# 0.16fF
C123 a_n327_n205# a_n861_n205# 0.02fF
C124 a_861_n140# a_n385_n140# 0.01fF
C125 a_861_n140# a_683_n140# 0.06fF
C126 a_505_n140# a_n29_n140# 0.02fF
C127 a_n1097_n140# a_n505_n205# 0.01fF
C128 a_n861_n205# w_n1133_n241# 0.20fF
C129 a_n327_n205# a_n683_n205# 0.03fF
C130 a_327_n140# a_n207_n140# 0.02fF
C131 a_919_n205# a_n505_n205# 0.00fF
C132 a_n149_n205# a_741_n205# 0.01fF
C133 a_n1097_n140# a_327_n140# 0.01fF
C134 a_n919_n140# a_n385_n140# 0.02fF
C135 a_n683_n205# w_n1133_n241# 0.20fF
C136 a_n919_n140# a_683_n140# 0.01fF
C137 a_n741_n140# a_327_n140# 0.01fF
C138 a_919_n205# a_327_n140# 0.01fF
C139 a_563_n205# a_n505_n205# 0.01fF
C140 a_861_n140# a_n207_n140# 0.01fF
C141 a_n149_n205# a_29_n205# 0.10fF
C142 a_n1097_n140# a_207_n205# 0.00fF
C143 a_919_n205# a_207_n205# 0.01fF
C144 a_861_n140# a_n741_n140# 0.01fF
C145 a_861_n140# a_919_n205# 0.06fF
C146 a_n327_n205# w_n1133_n241# 0.19fF
C147 a_n919_n140# a_n207_n140# 0.01fF
C148 a_563_n205# a_207_n205# 0.03fF
C149 a_29_n205# a_741_n205# 0.01fF
C150 a_505_n140# a_327_n140# 0.06fF
C151 a_n919_n140# a_n1097_n140# 0.06fF
C152 a_n919_n140# a_n741_n140# 0.06fF
C153 a_n563_n140# a_n385_n140# 0.06fF
C154 a_385_n205# a_n505_n205# 0.01fF
C155 a_n563_n140# a_683_n140# 0.01fF
C156 a_861_n140# a_505_n140# 0.03fF
C157 a_149_n140# w_n1133_n241# 0.02fF
C158 w_n1133_n241# VSUBS 3.28fF
.ends

.subckt ota_w_test_v2_without_cmfb on bias_circuit_0/m1_3551_3596# li_11121_570# li_11122_5650#
+ cmc li_14138_570# VSS VDD bias_circuit_0/bias_d in li_8434_570# bias_circuit_0/bias_b
+ li_8436_5651# i_bias bias_e bias_circuit_0/m1_1243_5997# bias_circuit_0/m1_3443_5997#
+ op bias_circuit_0/bias_c bias_a ip bias_circuit_0/m1_5643_5997#
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_0 VDD bias_circuit_0/bias_b bias_circuit_0/bias_b
+ li_8436_5651# bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_8436_5651# VDD
+ li_8436_5651# VDD bias_circuit_0/bias_b li_8436_5651# bias_circuit_0/bias_b VDD
+ VDD bias_circuit_0/bias_b bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_8436_5651#
+ VDD bias_circuit_0/bias_b li_8436_5651# li_8436_5651# bias_circuit_0/bias_b VDD
+ bias_circuit_0/bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_8 bias_circuit_0/bias_d li_8434_570# bias_circuit_0/bias_d
+ on VSS bias_circuit_0/bias_d on li_8434_570# on bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on bias_circuit_0/bias_d li_8434_570# VSS li_8434_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on li_8434_570# bias_circuit_0/bias_d on on bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_1 VDD bias_circuit_0/bias_b bias_circuit_0/bias_b
+ li_11122_5650# bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_11122_5650# VDD
+ li_11122_5650# VDD bias_circuit_0/bias_b li_11122_5650# bias_circuit_0/bias_b VDD
+ VDD bias_circuit_0/bias_b bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_11122_5650#
+ VDD bias_circuit_0/bias_b li_11122_5650# li_11122_5650# bias_circuit_0/bias_b VDD
+ bias_circuit_0/bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_9 bias_circuit_0/bias_d li_11121_570# bias_circuit_0/bias_d
+ op VSS bias_circuit_0/bias_d op li_11121_570# op bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op bias_circuit_0/bias_d li_11121_570# VSS li_11121_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op li_11121_570# bias_circuit_0/bias_d op op bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_2 VDD bias_circuit_0/bias_b bias_circuit_0/bias_b
+ li_8436_5651# bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_8436_5651# VDD
+ li_8436_5651# VDD bias_circuit_0/bias_b li_8436_5651# bias_circuit_0/bias_b VDD
+ VDD bias_circuit_0/bias_b bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_8436_5651#
+ VDD bias_circuit_0/bias_b li_8436_5651# li_8436_5651# bias_circuit_0/bias_b VDD
+ bias_circuit_0/bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_3 VDD bias_circuit_0/bias_b bias_circuit_0/bias_b
+ li_11122_5650# bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_11122_5650# VDD
+ li_11122_5650# VDD bias_circuit_0/bias_b li_11122_5650# bias_circuit_0/bias_b VDD
+ VDD bias_circuit_0/bias_b bias_circuit_0/bias_b VDD bias_circuit_0/bias_b li_11122_5650#
+ VDD bias_circuit_0/bias_b li_11122_5650# li_11122_5650# bias_circuit_0/bias_b VDD
+ bias_circuit_0/bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_0 VSS li_8436_5651# li_14138_570# ip li_8436_5651#
+ li_8436_5651# ip li_14138_570# li_8436_5651# li_14138_570# li_14138_570# li_8436_5651#
+ li_8436_5651# ip ip li_14138_570# ip li_14138_570# ip VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_1 VSS li_11122_5650# li_14138_570# in li_11122_5650#
+ li_11122_5650# in li_14138_570# li_11122_5650# li_14138_570# li_14138_570# li_11122_5650#
+ li_11122_5650# in in li_14138_570# in li_14138_570# in VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_AKSJZW_10 bias_circuit_0/bias_d li_11121_570# bias_circuit_0/bias_d
+ op VSS bias_circuit_0/bias_d op li_11121_570# op bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op bias_circuit_0/bias_d li_11121_570# VSS li_11121_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op li_11121_570# bias_circuit_0/bias_d op op bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_0 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_AKSJZW_11 bias_circuit_0/bias_d li_11121_570# bias_circuit_0/bias_d
+ op VSS bias_circuit_0/bias_d op li_11121_570# op bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op bias_circuit_0/bias_d li_11121_570# VSS li_11121_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op li_11121_570# bias_circuit_0/bias_d op op bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_1 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_2 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_3 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_4 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_5 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_6 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_7 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_8 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_9 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_10 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_11 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xbias_circuit_0 bias_circuit_0/bias_c bias_e i_bias VDD bias_circuit_0/m1_1243_5997#
+ bias_circuit_0/m1_3443_5997# bias_circuit_0/m1_5643_5997# bias_a bias_circuit_0/m1_7347_1428#
+ bias_circuit_0/m1_7639_1420# bias_circuit_0/m1_7169_923# bias_circuit_0/m1_3551_3596#
+ bias_circuit_0/m1_7461_921# bias_circuit_0/m1_7347_423# bias_circuit_0/m1_7639_427#
+ bias_circuit_0/bias_b VSS bias_circuit_0/bias_d bias_circuit
Xsky130_fd_pr__pfet_01v8_YVTMSC_0 on bias_circuit_0/bias_c li_8436_5651# bias_circuit_0/bias_c
+ bias_circuit_0/bias_c li_8436_5651# on VDD bias_circuit_0/bias_c li_8436_5651# bias_circuit_0/bias_c
+ on VDD bias_circuit_0/bias_c on bias_circuit_0/bias_c li_8436_5651# VDD on bias_circuit_0/bias_c
+ li_8436_5651# bias_circuit_0/bias_c on bias_circuit_0/bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_1 on bias_circuit_0/bias_c li_8436_5651# bias_circuit_0/bias_c
+ bias_circuit_0/bias_c li_8436_5651# on VDD bias_circuit_0/bias_c li_8436_5651# bias_circuit_0/bias_c
+ on VDD bias_circuit_0/bias_c on bias_circuit_0/bias_c li_8436_5651# VDD on bias_circuit_0/bias_c
+ li_8436_5651# bias_circuit_0/bias_c on bias_circuit_0/bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_0 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_YVTMSC_2 op bias_circuit_0/bias_c li_11122_5650# bias_circuit_0/bias_c
+ bias_circuit_0/bias_c li_11122_5650# op VDD bias_circuit_0/bias_c li_11122_5650#
+ bias_circuit_0/bias_c op VDD bias_circuit_0/bias_c op bias_circuit_0/bias_c li_11122_5650#
+ VDD op bias_circuit_0/bias_c li_11122_5650# bias_circuit_0/bias_c op bias_circuit_0/bias_c
+ VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_3 op bias_circuit_0/bias_c li_11122_5650# bias_circuit_0/bias_c
+ bias_circuit_0/bias_c li_11122_5650# op VDD bias_circuit_0/bias_c li_11122_5650#
+ bias_circuit_0/bias_c op VDD bias_circuit_0/bias_c op bias_circuit_0/bias_c li_11122_5650#
+ VDD op bias_circuit_0/bias_c li_11122_5650# bias_circuit_0/bias_c op bias_circuit_0/bias_c
+ VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_2 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_1 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_3 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_4 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_5 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_6 bias_circuit_0/bias_d li_8434_570# bias_circuit_0/bias_d
+ on VSS bias_circuit_0/bias_d on li_8434_570# on bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on bias_circuit_0/bias_d li_8434_570# VSS li_8434_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on li_8434_570# bias_circuit_0/bias_d on on bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_7 bias_circuit_0/bias_d li_8434_570# bias_circuit_0/bias_d
+ on VSS bias_circuit_0/bias_d on li_8434_570# on bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on bias_circuit_0/bias_d li_8434_570# VSS li_8434_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on li_8434_570# bias_circuit_0/bias_d on on bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
C0 li_14138_570# in 1.51fF
C1 op bias_circuit_0/bias_c 4.28fF
C2 VDD li_8436_5651# 4.41fF
C3 VDD bias_circuit_0/bias_d 3.18fF
C4 li_11122_5650# ip 0.01fF
C5 bias_circuit_0/m1_3551_3596# bias_circuit_0/bias_d 0.03fF
C6 bias_circuit_0/bias_d li_11121_570# 6.33fF
C7 li_11122_5650# bias_circuit_0/bias_c 3.17fF
C8 li_14138_570# li_11121_570# 0.23fF
C9 op li_11122_5650# 2.52fF
C10 ip in 0.03fF
C11 bias_a on 0.48fF
C12 cmc li_14138_570# 26.90fF
C13 bias_circuit_0/m1_7639_427# bias_a 0.01fF
C14 li_8434_570# li_8436_5651# 0.16fF
C15 li_8434_570# bias_circuit_0/bias_d 9.32fF
C16 VDD bias_circuit_0/bias_c 6.33fF
C17 bias_circuit_0/m1_7639_1420# bias_circuit_0/bias_d 0.00fF
C18 op VDD 0.65fF
C19 li_11122_5650# in 1.09fF
C20 bias_circuit_0/m1_3551_3596# bias_circuit_0/bias_c 0.00fF
C21 li_11121_570# bias_circuit_0/bias_c 0.12fF
C22 op li_11121_570# 4.14fF
C23 li_8434_570# bias_circuit_0/m1_7461_921# 0.01fF
C24 VDD li_11122_5650# 4.00fF
C25 li_11122_5650# li_11121_570# 0.16fF
C26 m1_15613_3568# bias_a 0.01fF
C27 li_8434_570# bias_circuit_0/bias_c 0.12fF
C28 cmc li_11122_5650# 0.13fF
C29 op li_8434_570# 0.19fF
C30 cmc in 0.31fF
C31 m1_17393_3568# li_14138_570# 0.01fF
C32 bias_circuit_0/bias_b on 0.27fF
C33 VDD bias_circuit_0/m1_3551_3596# 0.15fF
C34 VDD li_11121_570# 0.02fF
C35 on li_8436_5651# 2.50fF
C36 m1_17393_3568# ip 0.00fF
C37 bias_circuit_0/bias_d on 10.14fF
C38 VDD li_8434_570# 0.03fF
C39 li_8434_570# li_11121_570# 0.53fF
C40 li_14138_570# m1_18877_3928# 0.00fF
C41 bias_a li_8436_5651# 0.14fF
C42 bias_a bias_circuit_0/bias_d 2.87fF
C43 m1_17393_3568# li_11122_5650# 0.00fF
C44 li_14138_570# bias_a 27.43fF
C45 bias_e li_8434_570# 0.00fF
C46 m1_17393_3568# in 0.01fF
C47 bias_circuit_0/bias_c on 4.65fF
C48 li_8434_570# bias_circuit_0/m1_7639_1420# 0.01fF
C49 op on 0.59fF
C50 bias_a ip 0.31fF
C51 m1_15613_3568# li_14138_570# 0.01fF
C52 li_11122_5650# on 0.12fF
C53 op bias_a 0.52fF
C54 m1_18877_3928# in 0.00fF
C55 m1_17097_3928# li_14138_570# 0.00fF
C56 m1_15613_3568# ip 0.01fF
C57 VDD on 0.64fF
C58 bias_circuit_0/bias_b li_8436_5651# 4.78fF
C59 bias_circuit_0/bias_b bias_circuit_0/bias_d 0.02fF
C60 bias_circuit_0/m1_3551_3596# on 0.00fF
C61 li_11121_570# on 0.17fF
C62 cmc m1_18877_3928# 0.01fF
C63 m1_17097_3928# ip 0.01fF
C64 bias_circuit_0/bias_d li_8436_5651# 0.66fF
C65 bias_a li_11121_570# 10.56fF
C66 li_8434_570# on 4.12fF
C67 cmc bias_a 0.77fF
C68 bias_circuit_0/m1_7639_427# li_8434_570# 0.01fF
C69 li_14138_570# li_8436_5651# 0.80fF
C70 bias_e on 0.01fF
C71 li_14138_570# bias_circuit_0/bias_d 0.02fF
C72 bias_circuit_0/bias_b bias_circuit_0/bias_c 1.94fF
C73 bias_circuit_0/m1_7639_1420# on 0.00fF
C74 op bias_circuit_0/bias_b 0.27fF
C75 li_8434_570# bias_a 10.56fF
C76 bias_e bias_a 0.00fF
C77 m1_17097_3928# in 0.00fF
C78 ip li_8436_5651# 1.22fF
C79 bias_a bias_circuit_0/m1_7639_1420# 0.00fF
C80 bias_circuit_0/bias_b li_11122_5650# 4.63fF
C81 bias_circuit_0/bias_c li_8436_5651# 4.18fF
C82 bias_circuit_0/bias_d bias_circuit_0/bias_c 2.13fF
C83 op li_8436_5651# 0.13fF
C84 li_14138_570# ip 1.47fF
C85 op bias_circuit_0/bias_d 9.36fF
C86 op li_14138_570# 0.08fF
C87 li_11122_5650# li_8436_5651# 1.48fF
C88 bias_circuit_0/bias_d li_11122_5650# 0.28fF
C89 VDD bias_circuit_0/bias_b 13.69fF
C90 li_14138_570# li_11122_5650# -0.03fF
C91 in li_8436_5651# 0.01fF
C92 m1_17393_3568# VSS 0.09fF $ **FLOATING
C93 m1_15613_3568# VSS 0.05fF $ **FLOATING
C94 m1_18877_3928# VSS 0.10fF $ **FLOATING
C95 m1_17097_3928# VSS 0.09fF $ **FLOATING
C96 on VSS 6.48fF
C97 li_11121_570# VSS 10.65fF
C98 li_11122_5650# VSS 2.59fF
C99 li_8434_570# VSS 11.16fF
C100 bias_a VSS -301.12fF
C101 li_8436_5651# VSS 6.46fF
C102 bias_circuit_0/m1_3551_3596# VSS -342.22fF
C103 bias_circuit_0/bias_b VSS -356.81fF
C104 bias_circuit_0/m1_5643_5997# VSS 38.05fF
C105 bias_circuit_0/m1_3443_5997# VSS 35.85fF
C106 bias_circuit_0/m1_1243_5997# VSS 25.03fF
C107 VDD VSS 274.60fF
C108 i_bias VSS -60.83fF
C109 bias_circuit_0/bias_c VSS -127.80fF
C110 bias_circuit_0/m1_7639_427# VSS 0.13fF
C111 bias_circuit_0/m1_7347_423# VSS 0.13fF
C112 bias_circuit_0/m1_7461_921# VSS 0.14fF
C113 bias_circuit_0/m1_7169_923# VSS 0.14fF
C114 bias_circuit_0/m1_7055_433# VSS 0.14fF
C115 bias_circuit_0/m1_6763_422# VSS 0.20fF
C116 bias_circuit_0/m1_6471_422# VSS 0.20fF
C117 bias_circuit_0/m1_7639_1420# VSS 0.13fF
C118 bias_circuit_0/m1_7347_1428# VSS 0.14fF
C119 bias_circuit_0/m1_6877_922# VSS 0.14fF
C120 bias_circuit_0/m1_6585_923# VSS 0.22fF
C121 bias_circuit_0/m1_6293_922# VSS 0.16fF
C122 bias_circuit_0/m1_7055_1417# VSS 0.14fF
C123 bias_circuit_0/m1_6763_1422# VSS 0.22fF
C124 bias_circuit_0/m1_6471_1426# VSS 0.22fF
C125 bias_e VSS 5.12fF
C126 bias_circuit_0/bias_d VSS -235.40fF
C127 bias_circuit_0/li_3433_399# VSS 4.65fF
C128 li_14138_570# VSS 41.84fF
C129 cmc VSS -93.04fF
C130 op VSS 5.27fF
C131 in VSS -27.59fF
C132 ip VSS -27.52fF
.ends

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 w_n646_n356# a_448_n136# 0.13fF
C1 w_n646_n356# a_352_n136# 0.08fF
C2 w_n646_n356# a_n416_n136# 0.08fF
C3 a_n128_n136# w_n646_n356# 0.05fF
C4 w_n646_n356# a_n224_n136# 0.06fF
C5 a_448_n136# a_n512_n234# 0.03fF
C6 a_352_n136# a_n512_n234# 0.03fF
C7 a_160_n136# a_64_n136# 0.33fF
C8 a_n512_n234# a_n416_n136# 0.03fF
C9 w_n646_n356# a_256_n136# 0.06fF
C10 a_n128_n136# a_n512_n234# 0.03fF
C11 a_n512_n234# a_n224_n136# 0.03fF
C12 a_n508_n136# a_448_n136# 0.02fF
C13 a_n320_n136# a_160_n136# 0.04fF
C14 a_n508_n136# a_352_n136# 0.02fF
C15 a_n508_n136# a_n416_n136# 0.33fF
C16 a_n508_n136# a_n128_n136# 0.05fF
C17 a_n508_n136# a_n224_n136# 0.07fF
C18 a_256_n136# a_n512_n234# 0.03fF
C19 a_n320_n136# a_64_n136# 0.05fF
C20 a_n508_n136# a_256_n136# 0.02fF
C21 a_448_n136# a_160_n136# 0.07fF
C22 a_352_n136# a_160_n136# 0.12fF
C23 a_160_n136# a_n416_n136# 0.03fF
C24 a_n32_n136# w_n646_n356# 0.05fF
C25 a_n128_n136# a_160_n136# 0.07fF
C26 a_160_n136# a_n224_n136# 0.05fF
C27 a_448_n136# a_64_n136# 0.05fF
C28 a_352_n136# a_64_n136# 0.07fF
C29 a_n416_n136# a_64_n136# 0.04fF
C30 a_n320_n136# a_448_n136# 0.02fF
C31 a_n32_n136# a_n512_n234# 0.03fF
C32 a_n320_n136# a_352_n136# 0.03fF
C33 a_256_n136# a_160_n136# 0.33fF
C34 a_n128_n136# a_64_n136# 0.12fF
C35 a_n224_n136# a_64_n136# 0.07fF
C36 a_n320_n136# a_n416_n136# 0.33fF
C37 a_n320_n136# a_n128_n136# 0.12fF
C38 a_n320_n136# a_n224_n136# 0.33fF
C39 a_n32_n136# a_n508_n136# 0.04fF
C40 a_256_n136# a_64_n136# 0.12fF
C41 a_n320_n136# a_256_n136# 0.03fF
C42 a_352_n136# a_448_n136# 0.33fF
C43 a_448_n136# a_n416_n136# 0.02fF
C44 a_352_n136# a_n416_n136# 0.02fF
C45 w_n646_n356# a_n512_n234# 1.47fF
C46 a_n128_n136# a_448_n136# 0.03fF
C47 a_448_n136# a_n224_n136# 0.03fF
C48 a_n32_n136# a_160_n136# 0.12fF
C49 a_n128_n136# a_352_n136# 0.04fF
C50 a_352_n136# a_n224_n136# 0.03fF
C51 a_n128_n136# a_n416_n136# 0.07fF
C52 a_n224_n136# a_n416_n136# 0.12fF
C53 a_n508_n136# w_n646_n356# 0.13fF
C54 a_n128_n136# a_n224_n136# 0.33fF
C55 a_448_n136# a_256_n136# 0.12fF
C56 a_n32_n136# a_64_n136# 0.33fF
C57 a_352_n136# a_256_n136# 0.33fF
C58 a_256_n136# a_n416_n136# 0.03fF
C59 a_n320_n136# a_n32_n136# 0.07fF
C60 a_n128_n136# a_256_n136# 0.05fF
C61 a_256_n136# a_n224_n136# 0.04fF
C62 a_n508_n136# a_n512_n234# 0.03fF
C63 w_n646_n356# a_160_n136# 0.06fF
C64 a_n32_n136# a_448_n136# 0.04fF
C65 w_n646_n356# a_64_n136# 0.05fF
C66 a_160_n136# a_n512_n234# 0.03fF
C67 a_n32_n136# a_352_n136# 0.05fF
C68 a_n32_n136# a_n416_n136# 0.05fF
C69 a_n320_n136# w_n646_n356# 0.06fF
C70 a_n32_n136# a_n128_n136# 0.33fF
C71 a_n32_n136# a_n224_n136# 0.12fF
C72 a_n508_n136# a_160_n136# 0.03fF
C73 a_n512_n234# a_64_n136# 0.03fF
C74 a_n320_n136# a_n512_n234# 0.03fF
C75 a_n32_n136# a_256_n136# 0.07fF
C76 a_n508_n136# a_64_n136# 0.03fF
C77 a_n320_n136# a_n508_n136# 0.12fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# a_448_n52# a_n416_n52# a_160_n52#
+ a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149# a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_160_n52# a_n508_n52# 0.01fF
C1 a_160_n52# a_n416_n52# 0.01fF
C2 a_n512_n149# a_352_n52# 0.03fF
C3 a_n508_n52# a_64_n52# 0.01fF
C4 a_n416_n52# a_64_n52# 0.02fF
C5 a_n508_n52# a_n128_n52# 0.02fF
C6 a_n128_n52# a_n416_n52# 0.03fF
C7 a_448_n52# a_n32_n52# 0.02fF
C8 a_256_n52# a_n224_n52# 0.02fF
C9 a_n224_n52# a_n320_n52# 0.13fF
C10 a_160_n52# a_64_n52# 0.13fF
C11 a_n512_n149# a_n32_n52# 0.03fF
C12 a_160_n52# a_n128_n52# 0.03fF
C13 a_n128_n52# a_64_n52# 0.05fF
C14 a_256_n52# a_448_n52# 0.05fF
C15 a_448_n52# a_n320_n52# 0.01fF
C16 a_n508_n52# a_n224_n52# 0.03fF
C17 a_n416_n52# a_n224_n52# 0.05fF
C18 a_352_n52# a_n32_n52# 0.02fF
C19 a_n512_n149# a_256_n52# 0.03fF
C20 a_n512_n149# a_n320_n52# 0.03fF
C21 a_160_n52# a_n224_n52# 0.02fF
C22 a_448_n52# a_n508_n52# 0.01fF
C23 a_448_n52# a_n416_n52# 0.01fF
C24 a_n224_n52# a_64_n52# 0.03fF
C25 a_256_n52# a_352_n52# 0.13fF
C26 a_352_n52# a_n320_n52# 0.01fF
C27 a_n128_n52# a_n224_n52# 0.13fF
C28 a_n512_n149# a_n508_n52# 0.03fF
C29 a_n512_n149# a_n416_n52# 0.03fF
C30 a_448_n52# a_160_n52# 0.03fF
C31 a_448_n52# a_64_n52# 0.02fF
C32 a_448_n52# a_n128_n52# 0.01fF
C33 a_256_n52# a_n32_n52# 0.03fF
C34 a_n512_n149# a_160_n52# 0.03fF
C35 a_n32_n52# a_n320_n52# 0.03fF
C36 a_n508_n52# a_352_n52# 0.01fF
C37 a_352_n52# a_n416_n52# 0.01fF
C38 a_n512_n149# a_64_n52# 0.03fF
C39 a_n512_n149# a_n128_n52# 0.03fF
C40 a_160_n52# a_352_n52# 0.05fF
C41 a_256_n52# a_n320_n52# 0.01fF
C42 a_n508_n52# a_n32_n52# 0.02fF
C43 a_n416_n52# a_n32_n52# 0.02fF
C44 a_352_n52# a_64_n52# 0.03fF
C45 a_448_n52# a_n224_n52# 0.01fF
C46 a_352_n52# a_n128_n52# 0.02fF
C47 a_160_n52# a_n32_n52# 0.05fF
C48 a_n512_n149# a_n224_n52# 0.03fF
C49 a_256_n52# a_n508_n52# 0.01fF
C50 a_256_n52# a_n416_n52# 0.01fF
C51 a_n32_n52# a_64_n52# 0.13fF
C52 a_n508_n52# a_n320_n52# 0.05fF
C53 a_n416_n52# a_n320_n52# 0.13fF
C54 a_n128_n52# a_n32_n52# 0.13fF
C55 a_n512_n149# a_448_n52# 0.03fF
C56 a_352_n52# a_n224_n52# 0.01fF
C57 a_256_n52# a_160_n52# 0.13fF
C58 a_160_n52# a_n320_n52# 0.02fF
C59 a_256_n52# a_64_n52# 0.05fF
C60 a_64_n52# a_n320_n52# 0.02fF
C61 a_256_n52# a_n128_n52# 0.02fF
C62 a_n508_n52# a_n416_n52# 0.13fF
C63 a_n128_n52# a_n320_n52# 0.05fF
C64 a_448_n52# a_352_n52# 0.13fF
C65 a_n32_n52# a_n224_n52# 0.05fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate en en_b VDD in out VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in out in in VSS out in out out en out nmos_tgate
C0 en out 0.01fF
C1 in out 0.77fF
C2 VDD en_b -0.11fF
C3 VDD en 0.12fF
C4 VDD in 0.70fF
C5 VDD out 0.29fF
C6 en en_b 0.07fF
C7 in en_b 0.15fF
C8 en_b out 0.01fF
C9 in en 0.13fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 m3_n630_n580# c1_n530_n480# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb cm op cmc p2_b p2 p1 on unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_8/in
+ transmission_gate_4/out bias_a VDD transmission_gate_3/out transmission_gate_7/in
+ VSS p1_b
Xtransmission_gate_10 p1 p1_b VDD transmission_gate_3/out on VSS transmission_gate
Xtransmission_gate_11 p1 p1_b VDD transmission_gate_4/out op VSS transmission_gate
Xtransmission_gate_0 p1 p1_b VDD cm transmission_gate_7/in VSS transmission_gate
Xtransmission_gate_1 p1 p1_b VDD cm transmission_gate_6/in VSS transmission_gate
Xtransmission_gate_2 p1 p1_b VDD bias_a transmission_gate_8/in VSS transmission_gate
Xtransmission_gate_3 p2 p2_b VDD cm transmission_gate_3/out VSS transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 p2_b VDD cm transmission_gate_4/out VSS transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 p2_b VDD bias_a transmission_gate_9/in VSS transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 p2_b VDD transmission_gate_6/in op VSS transmission_gate
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 p2_b VDD transmission_gate_7/in on VSS transmission_gate
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 p2_b VDD transmission_gate_8/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 p1_b VDD transmission_gate_9/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 cmc unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C1 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_27/c1_n530_n480# -0.37fF
C2 transmission_gate_6/in on 0.40fF
C3 transmission_gate_8/in op 0.82fF
C4 op transmission_gate_3/out 0.56fF
C5 unit_cap_mim_m3m4_32/c1_n530_n480# on 0.06fF
C6 unit_cap_mim_m3m4_28/m3_n630_n580# transmission_gate_8/in 0.10fF
C7 cmc unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C8 unit_cap_mim_m3m4_29/c1_n530_n480# op 0.03fF
C9 unit_cap_mim_m3m4_27/m3_n630_n580# transmission_gate_6/in 0.14fF
C10 transmission_gate_8/in unit_cap_mim_m3m4_20/m3_n630_n580# 0.17fF
C11 unit_cap_mim_m3m4_30/c1_n530_n480# transmission_gate_4/out -0.25fF
C12 p2_b p1_b 2.92fF
C13 p2 unit_cap_mim_m3m4_17/m3_n630_n580# 0.04fF
C14 unit_cap_mim_m3m4_26/c1_n530_n480# on 0.06fF
C15 p1 p2_b 2.16fF
C16 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C17 VDD transmission_gate_4/out -0.03fF
C18 op unit_cap_mim_m3m4_23/c1_n530_n480# 0.13fF
C19 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580# -0.29fF
C20 unit_cap_mim_m3m4_30/m3_n630_n580# p1_b 0.01fF
C21 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C22 transmission_gate_6/in unit_cap_mim_m3m4_27/c1_n530_n480# -0.12fF
C23 p1 unit_cap_mim_m3m4_30/m3_n630_n580# 0.06fF
C24 transmission_gate_8/in transmission_gate_4/out 0.26fF
C25 transmission_gate_3/out transmission_gate_4/out 0.37fF
C26 cm p1_b 1.15fF
C27 VDD transmission_gate_8/in 0.00fF
C28 transmission_gate_9/in p1_b 0.59fF
C29 VDD transmission_gate_3/out -0.01fF
C30 p1 cm 1.50fF
C31 transmission_gate_7/in op 2.63fF
C32 p1 transmission_gate_9/in 0.70fF
C33 unit_cap_mim_m3m4_25/m3_n630_n580# transmission_gate_9/in 0.38fF
C34 p2 p2_b 6.60fF
C35 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C36 op unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C37 transmission_gate_8/in transmission_gate_3/out 0.23fF
C38 unit_cap_mim_m3m4_31/c1_n530_n480# op 0.05fF
C39 unit_cap_mim_m3m4_35/m3_n630_n580# transmission_gate_8/in -0.17fF
C40 cmc p1_b 0.52fF
C41 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580# -0.20fF
C42 p1 cmc 0.49fF
C43 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580# -0.20fF
C44 on p1_b 0.45fF
C45 transmission_gate_7/in unit_cap_mim_m3m4_20/m3_n630_n580# -0.57fF
C46 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C47 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_3/out -0.11fF
C48 unit_cap_mim_m3m4_16/m3_n630_n580# transmission_gate_4/out -0.29fF
C49 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C50 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580# -0.14fF
C51 bias_a p2_b 0.48fF
C52 p1 on 0.49fF
C53 transmission_gate_6/in unit_cap_mim_m3m4_18/m3_n630_n580# 0.06fF
C54 unit_cap_mim_m3m4_23/c1_n530_n480# transmission_gate_4/out 0.06fF
C55 p2 cm 1.33fF
C56 p2 transmission_gate_9/in 0.14fF
C57 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C58 unit_cap_mim_m3m4_21/m3_n630_n580# p1_b 0.05fF
C59 p1 unit_cap_mim_m3m4_21/m3_n630_n580# 0.06fF
C60 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C61 bias_a cm 0.91fF
C62 transmission_gate_9/in bias_a 0.02fF
C63 transmission_gate_7/in transmission_gate_4/out 0.61fF
C64 transmission_gate_3/out unit_cap_mim_m3m4_23/c1_n530_n480# -0.13fF
C65 p2 cmc 0.25fF
C66 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C67 transmission_gate_7/in VDD -0.11fF
C68 unit_cap_mim_m3m4_28/c1_n530_n480# transmission_gate_6/in 0.05fF
C69 p2 on 0.24fF
C70 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_23/c1_n530_n480# -0.19fF
C71 unit_cap_mim_m3m4_31/c1_n530_n480# transmission_gate_4/out 0.06fF
C72 unit_cap_mim_m3m4_27/c1_n530_n480# p1_b 0.06fF
C73 transmission_gate_8/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C74 transmission_gate_7/in transmission_gate_8/in 0.73fF
C75 transmission_gate_7/in transmission_gate_3/out 0.29fF
C76 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_24/m3_n630_n580# 0.10fF
C77 p1 unit_cap_mim_m3m4_27/c1_n530_n480# 0.11fF
C78 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C79 transmission_gate_6/in p1_b 0.41fF
C80 p1 transmission_gate_6/in 0.37fF
C81 op p2_b 0.42fF
C82 unit_cap_mim_m3m4_16/c1_n530_n480# transmission_gate_4/out 0.06fF
C83 unit_cap_mim_m3m4_18/m3_n630_n580# p1_b 0.06fF
C84 p2 unit_cap_mim_m3m4_27/c1_n530_n480# 0.04fF
C85 p1 unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C86 unit_cap_mim_m3m4_30/m3_n630_n580# op 0.55fF
C87 unit_cap_mim_m3m4_26/c1_n530_n480# p1_b 0.06fF
C88 cmc unit_cap_mim_m3m4_26/m3_n630_n580# 0.10fF
C89 p1 unit_cap_mim_m3m4_26/c1_n530_n480# 0.11fF
C90 p2 transmission_gate_6/in 0.61fF
C91 op transmission_gate_9/in 0.67fF
C92 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.12fF
C93 transmission_gate_7/in unit_cap_mim_m3m4_19/m3_n630_n580# -0.29fF
C94 unit_cap_mim_m3m4_17/m3_n630_n580# transmission_gate_3/out -0.21fF
C95 unit_cap_mim_m3m4_28/c1_n530_n480# p1_b 0.06fF
C96 transmission_gate_6/in bias_a 0.05fF
C97 p1 unit_cap_mim_m3m4_28/c1_n530_n480# 0.11fF
C98 cmc op 4.14fF
C99 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C100 op unit_cap_mim_m3m4_22/c1_n530_n480# 0.07fF
C101 p2_b transmission_gate_4/out 0.06fF
C102 op on 1.84fF
C103 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580# -0.21fF
C104 VDD p2_b 1.69fF
C105 p2 unit_cap_mim_m3m4_26/c1_n530_n480# 0.04fF
C106 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_30/c1_n530_n480# -0.12fF
C107 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.17fF
C108 unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_4/out -0.62fF
C109 unit_cap_mim_m3m4_27/m3_n630_n580# op 0.49fF
C110 transmission_gate_8/in p2_b 0.40fF
C111 p1 p1_b 8.88fF
C112 transmission_gate_3/out p2_b 0.10fF
C113 unit_cap_mim_m3m4_20/m3_n630_n580# on 0.60fF
C114 p2 unit_cap_mim_m3m4_28/c1_n530_n480# 0.04fF
C115 cm transmission_gate_4/out 0.08fF
C116 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.12fF
C117 transmission_gate_9/in transmission_gate_4/out 3.08fF
C118 unit_cap_mim_m3m4_24/c1_n530_n480# p1_b 0.06fF
C119 VDD cm 1.33fF
C120 VDD transmission_gate_9/in -0.09fF
C121 transmission_gate_8/in unit_cap_mim_m3m4_34/m3_n630_n580# 0.57fF
C122 p1 unit_cap_mim_m3m4_24/c1_n530_n480# 0.11fF
C123 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_34/m3_n630_n580# 0.17fF
C124 op unit_cap_mim_m3m4_31/m3_n630_n580# 0.03fF
C125 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580# -0.21fF
C126 transmission_gate_7/in unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C127 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_20/m3_n630_n580# 0.17fF
C128 cmc transmission_gate_4/out 0.10fF
C129 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.12fF
C130 transmission_gate_8/in cm 0.03fF
C131 transmission_gate_8/in transmission_gate_9/in 3.35fF
C132 cm transmission_gate_3/out 0.19fF
C133 transmission_gate_9/in transmission_gate_3/out 1.28fF
C134 op unit_cap_mim_m3m4_27/c1_n530_n480# 0.02fF
C135 VDD cmc 0.82fF
C136 on transmission_gate_4/out 3.23fF
C137 p2 p1_b 5.94fF
C138 VDD on -0.02fF
C139 transmission_gate_9/in unit_cap_mim_m3m4_23/m3_n630_n580# 0.17fF
C140 p1 p2 2.82fF
C141 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_33/c1_n530_n480# -0.19fF
C142 transmission_gate_8/in unit_cap_mim_m3m4_21/c1_n530_n480# -0.31fF
C143 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C144 cmc transmission_gate_8/in 8.39fF
C145 cmc transmission_gate_3/out 1.02fF
C146 transmission_gate_6/in op 0.59fF
C147 bias_a p1_b 0.52fF
C148 transmission_gate_8/in on 0.86fF
C149 unit_cap_mim_m3m4_24/c1_n530_n480# p2 0.04fF
C150 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_20/c1_n530_n480# -0.19fF
C151 transmission_gate_3/out on 0.39fF
C152 p1 bias_a 0.81fF
C153 unit_cap_mim_m3m4_28/m3_n630_n580# transmission_gate_6/in -0.12fF
C154 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580# -0.36fF
C155 transmission_gate_9/in unit_cap_mim_m3m4_24/m3_n630_n580# 0.16fF
C156 transmission_gate_9/in unit_cap_mim_m3m4_16/m3_n630_n580# 0.17fF
C157 transmission_gate_7/in p2_b 0.41fF
C158 unit_cap_mim_m3m4_23/m3_n630_n580# on 0.48fF
C159 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C160 unit_cap_mim_m3m4_31/m3_n630_n580# transmission_gate_4/out 0.53fF
C161 unit_cap_mim_m3m4_21/m3_n630_n580# transmission_gate_8/in -0.97fF
C162 unit_cap_mim_m3m4_29/m3_n630_n580# transmission_gate_6/in -0.62fF
C163 transmission_gate_7/in cm 0.11fF
C164 transmission_gate_7/in transmission_gate_9/in 0.02fF
C165 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C166 p2 bias_a 0.60fF
C167 on unit_cap_mim_m3m4_23/c1_n530_n480# 0.21fF
C168 transmission_gate_6/in transmission_gate_4/out 0.46fF
C169 unit_cap_mim_m3m4_28/c1_n530_n480# op 0.18fF
C170 VDD transmission_gate_6/in 0.06fF
C171 transmission_gate_7/in cmc 0.07fF
C172 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580# -0.32fF
C173 transmission_gate_7/in on 3.11fF
C174 unit_cap_mim_m3m4_25/c1_n530_n480# p1_b 0.06fF
C175 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.17fF
C176 transmission_gate_6/in transmission_gate_8/in -0.36fF
C177 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C178 transmission_gate_6/in transmission_gate_3/out 0.76fF
C179 unit_cap_mim_m3m4_25/c1_n530_n480# p1 0.11fF
C180 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580# -0.32fF
C181 op p1_b 0.28fF
C182 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C183 unit_cap_mim_m3m4_18/c1_n530_n480# on 0.06fF
C184 unit_cap_mim_m3m4_29/c1_n530_n480# transmission_gate_6/in -0.25fF
C185 p1 op 0.52fF
C186 unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_9/in -0.62fF
C187 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.17fF
C188 unit_cap_mim_m3m4_20/m3_n630_n580# p1_b 0.05fF
C189 p1 unit_cap_mim_m3m4_20/m3_n630_n580# 0.06fF
C190 unit_cap_mim_m3m4_25/c1_n530_n480# p2 0.04fF
C191 unit_cap_mim_m3m4_29/m3_n630_n580# p1_b 0.05fF
C192 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C193 unit_cap_mim_m3m4_22/m3_n630_n580# cmc 0.69fF
C194 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480# -0.19fF
C195 p1 unit_cap_mim_m3m4_29/m3_n630_n580# 0.06fF
C196 transmission_gate_7/in unit_cap_mim_m3m4_20/c1_n530_n480# -0.19fF
C197 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# -0.26fF
C198 p2 op 0.16fF
C199 unit_cap_mim_m3m4_17/m3_n630_n580# cmc 0.17fF
C200 cmc unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C201 transmission_gate_7/in transmission_gate_6/in 0.45fF
C202 p1_b transmission_gate_4/out 0.55fF
C203 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C204 VDD p1_b 1.00fF
C205 p1 transmission_gate_4/out 0.80fF
C206 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C207 cm p2_b 1.01fF
C208 p1 VDD 1.10fF
C209 transmission_gate_9/in p2_b 0.02fF
C210 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C211 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C212 transmission_gate_8/in p1_b 0.17fF
C213 transmission_gate_3/out p1_b 0.59fF
C214 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C215 unit_cap_mim_m3m4_35/m3_n630_n580# p1_b 0.01fF
C216 p1 transmission_gate_8/in 0.39fF
C217 p1 transmission_gate_3/out 0.71fF
C218 cmc p2_b 0.12fF
C219 p1 unit_cap_mim_m3m4_35/m3_n630_n580# 0.07fF
C220 unit_cap_mim_m3m4_23/m3_n630_n580# p1_b 0.05fF
C221 on p2_b 0.37fF
C222 unit_cap_mim_m3m4_29/c1_n530_n480# p1_b 0.06fF
C223 p1 unit_cap_mim_m3m4_23/m3_n630_n580# 0.06fF
C224 unit_cap_mim_m3m4_17/c1_n530_n480# op 0.06fF
C225 transmission_gate_9/in cm 0.04fF
C226 unit_cap_mim_m3m4_29/c1_n530_n480# p1 0.11fF
C227 p2 transmission_gate_4/out 0.15fF
C228 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480# -0.20fF
C229 VDD p2 4.16fF
C230 unit_cap_mim_m3m4_24/m3_n630_n580# p1_b 0.06fF
C231 unit_cap_mim_m3m4_16/m3_n630_n580# p1_b 0.06fF
C232 transmission_gate_7/in unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C233 cmc transmission_gate_9/in 6.93fF
C234 p1 unit_cap_mim_m3m4_24/m3_n630_n580# 0.08fF
C235 bias_a transmission_gate_4/out 0.09fF
C236 p1 unit_cap_mim_m3m4_16/m3_n630_n580# 0.08fF
C237 transmission_gate_9/in unit_cap_mim_m3m4_22/c1_n530_n480# -0.25fF
C238 p2 transmission_gate_8/in 0.63fF
C239 p2 transmission_gate_3/out 0.15fF
C240 VDD bias_a 0.69fF
C241 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_24/m3_n630_n580# 0.17fF
C242 transmission_gate_9/in on 1.03fF
C243 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580# -0.30fF
C244 cmc unit_cap_mim_m3m4_21/c1_n530_n480# 0.12fF
C245 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C246 unit_cap_mim_m3m4_29/c1_n530_n480# p2 0.04fF
C247 transmission_gate_8/in bias_a 0.03fF
C248 unit_cap_mim_m3m4_21/c1_n530_n480# on 0.06fF
C249 bias_a transmission_gate_3/out 0.05fF
C250 cmc unit_cap_mim_m3m4_22/c1_n530_n480# 0.12fF
C251 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C252 cmc on 1.98fF
C253 unit_cap_mim_m3m4_19/m3_n630_n580# p1_b 0.06fF
C254 transmission_gate_7/in p1_b 0.40fF
C255 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C256 p1 unit_cap_mim_m3m4_19/m3_n630_n580# 0.08fF
C257 p1 transmission_gate_7/in 0.39fF
C258 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.17fF
C259 p2 unit_cap_mim_m3m4_24/m3_n630_n580# 0.05fF
C260 p2 unit_cap_mim_m3m4_16/m3_n630_n580# 0.05fF
C261 unit_cap_mim_m3m4_28/m3_n630_n580# op 0.67fF
C262 unit_cap_mim_m3m4_27/m3_n630_n580# cmc 0.10fF
C263 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_21/c1_n530_n480# -0.19fF
C264 transmission_gate_6/in p2_b 0.42fF
C265 transmission_gate_9/in unit_cap_mim_m3m4_31/m3_n630_n580# 0.12fF
C266 unit_cap_mim_m3m4_21/m3_n630_n580# cmc 0.68fF
C267 unit_cap_mim_m3m4_29/m3_n630_n580# op 0.39fF
C268 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.17fF
C269 unit_cap_mim_m3m4_25/c1_n530_n480# transmission_gate_4/out 0.06fF
C270 transmission_gate_7/in p2 0.60fF
C271 transmission_gate_7/in unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C272 unit_cap_mim_m3m4_30/c1_n530_n480# op 0.17fF
C273 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C274 transmission_gate_6/in cm 0.19fF
C275 transmission_gate_6/in transmission_gate_9/in 0.09fF
C276 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_20/m3_n630_n580# 0.10fF
C277 unit_cap_mim_m3m4_22/m3_n630_n580# p1_b 0.05fF
C278 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C279 op transmission_gate_4/out 1.08fF
C280 p1 unit_cap_mim_m3m4_22/m3_n630_n580# 0.06fF
C281 transmission_gate_7/in bias_a 0.09fF
C282 on unit_cap_mim_m3m4_20/c1_n530_n480# 0.15fF
C283 VDD op -0.48fF
C284 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_35/c1_n530_n480# -0.13fF
C285 unit_cap_mim_m3m4_17/m3_n630_n580# p1_b 0.06fF
C286 transmission_gate_6/in cmc 1.17fF
C287 p1 unit_cap_mim_m3m4_17/m3_n630_n580# 0.08fF
C288 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C289 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C290 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.39fF
C291 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C292 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.51fF
C293 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C294 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.74fF
C295 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C296 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.51fF
C297 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.52fF
C298 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.56fF
C299 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.60fF
C300 cmc VSS -29.29fF
C301 transmission_gate_9/in VSS 3.31fF
C302 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.54fF
C303 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.61fF
C304 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C305 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C306 p2 VSS 101.65fF
C307 p2_b VSS 36.06fF
C308 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.84fF
C309 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C310 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.40fF
C311 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C312 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.03fF
C313 transmission_gate_4/out VSS -4.34fF
C314 transmission_gate_3/out VSS 0.32fF
C315 p1 VSS 85.98fF
C316 transmission_gate_8/in VSS 3.12fF
C317 bias_a VSS 6.68fF
C318 transmission_gate_6/in VSS -13.34fF
C319 transmission_gate_7/in VSS 9.47fF
C320 cm VSS 5.76fF
C321 op VSS -0.11fF
C322 p1_b VSS 109.11fF
C323 VDD VSS 69.52fF
C324 on VSS -13.19fF
.ends

.subckt ota_w_test_v2 ip in p1 p1_b p2 p2_b op on i_bias cm bias_a bias_b bias_c bias_d
+ cmc VDD VSS
Xota_w_test_v2_without_cmfb_0 on ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596#
+ ota_w_test_v2_without_cmfb_0/li_11121_570# ota_w_test_v2_without_cmfb_0/li_11122_5650#
+ cmc ota_w_test_v2_without_cmfb_0/li_14138_570# VSS VDD bias_d in ota_w_test_v2_without_cmfb_0/li_8434_570#
+ bias_b ota_w_test_v2_without_cmfb_0/li_8436_5651# i_bias cm ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997#
+ ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# op bias_c bias_a ip ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997#
+ ota_w_test_v2_without_cmfb
Xsc_cmfb_0 cm op cmc p2_b p2 p1 on sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_8/in
+ sc_cmfb_0/transmission_gate_4/out bias_a VDD sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_7/in
+ VSS p1_b sc_cmfb
C0 VDD on 0.18fF
C1 p1_b p1 0.00fF
C2 sc_cmfb_0/transmission_gate_4/out p1 0.05fF
C3 bias_d on 7.34fF
C4 bias_a sc_cmfb_0/transmission_gate_7/in 0.00fF
C5 p2_b p1 0.00fF
C6 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.02fF
C7 ota_w_test_v2_without_cmfb_0/li_11122_5650# on 0.22fF
C8 VDD sc_cmfb_0/transmission_gate_3/out -0.00fF
C9 bias_b cm 3.45fF
C10 bias_a cm 3.09fF
C11 sc_cmfb_0/transmission_gate_8/in p1 0.00fF
C12 bias_b VDD 0.16fF
C13 bias_a VDD 0.02fF
C14 p1_b sc_cmfb_0/transmission_gate_4/out 0.00fF
C15 ota_w_test_v2_without_cmfb_0/li_14138_570# in -0.00fF
C16 bias_a bias_d -0.00fF
C17 ota_w_test_v2_without_cmfb_0/li_14138_570# ip 0.00fF
C18 bias_b ota_w_test_v2_without_cmfb_0/li_11122_5650# -0.00fF
C19 i_bias bias_c 0.00fF
C20 ota_w_test_v2_without_cmfb_0/li_11121_570# on 0.01fF
C21 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VDD 0.00fF
C22 cmc cm -2.78fF
C23 cmc op 0.19fF
C24 p1 on 0.01fF
C25 cmc VDD -0.01fF
C26 sc_cmfb_0/transmission_gate_7/in cm 0.00fF
C27 ota_w_test_v2_without_cmfb_0/li_8436_5651# bias_c -0.00fF
C28 VDD sc_cmfb_0/transmission_gate_7/in 0.00fF
C29 ota_w_test_v2_without_cmfb_0/li_8434_570# on 0.00fF
C30 ota_w_test_v2_without_cmfb_0/li_14138_570# ota_w_test_v2_without_cmfb_0/li_8436_5651# 0.00fF
C31 op cm 1.43fF
C32 VDD cm -0.01fF
C33 VDD op 2.85fF
C34 bias_a p1 0.00fF
C35 bias_d cm 4.24fF
C36 on ota_w_test_v2_without_cmfb_0/li_8436_5651# 0.37fF
C37 bias_d op -0.00fF
C38 p1_b on 0.01fF
C39 op ota_w_test_v2_without_cmfb_0/li_11122_5650# 0.36fF
C40 VDD ota_w_test_v2_without_cmfb_0/li_11122_5650# 0.23fF
C41 p1_b sc_cmfb_0/transmission_gate_3/out -0.00fF
C42 p1_b bias_a 0.00fF
C43 on bias_c -0.00fF
C44 op ip 0.01fF
C45 ota_w_test_v2_without_cmfb_0/li_11121_570# cm 0.39fF
C46 ota_w_test_v2_without_cmfb_0/li_11121_570# op 0.00fF
C47 ota_w_test_v2_without_cmfb_0/li_14138_570# on 0.01fF
C48 bias_a sc_cmfb_0/transmission_gate_8/in 0.00fF
C49 bias_d ota_w_test_v2_without_cmfb_0/li_11121_570# -0.00fF
C50 op p1 0.01fF
C51 bias_b bias_c 0.26fF
C52 ota_w_test_v2_without_cmfb_0/li_8434_570# cm 0.38fF
C53 bias_a bias_c 2.52fF
C54 bias_d ota_w_test_v2_without_cmfb_0/li_8434_570# -0.00fF
C55 VDD ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.00fF
C56 on sc_cmfb_0/transmission_gate_3/out 0.00fF
C57 p1_b cm 0.01fF
C58 op ota_w_test_v2_without_cmfb_0/li_8436_5651# 0.40fF
C59 VDD ota_w_test_v2_without_cmfb_0/li_8436_5651# -0.00fF
C60 p1_b op 0.00fF
C61 sc_cmfb_0/transmission_gate_4/out op 0.00fF
C62 p1_b VDD -0.00fF
C63 sc_cmfb_0/transmission_gate_4/out VDD 0.04fF
C64 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VDD 0.00fF
C65 ota_w_test_v2_without_cmfb_0/li_11122_5650# ota_w_test_v2_without_cmfb_0/li_8436_5651# -0.00fF
C66 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# cm 0.23fF
C67 VDD sc_cmfb_0/transmission_gate_8/in -0.03fF
C68 cmc ota_w_test_v2_without_cmfb_0/li_14138_570# 0.03fF
C69 bias_b bias_a 0.15fF
C70 cm bias_c 2.51fF
C71 op bias_c 1.56fF
C72 cmc on 0.13fF
C73 ip ota_w_test_v2_without_cmfb_0/li_8436_5651# -0.00fF
C74 ota_w_test_v2_without_cmfb_0/li_14138_570# cm 1.29fF
C75 ota_w_test_v2_without_cmfb_0/li_14138_570# op 0.00fF
C76 ota_w_test_v2_without_cmfb_0/li_11122_5650# bias_c 0.00fF
C77 on cm 3.11fF
C78 op on 3.35fF
C79 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C80 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C81 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C82 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C83 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C84 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C85 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C86 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C87 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C88 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.37fF
C89 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C90 sc_cmfb_0/transmission_gate_9/in VSS 1.93fF
C91 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C92 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C93 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C94 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C95 p2 VSS 101.39fF
C96 p2_b VSS 34.70fF
C97 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C98 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C99 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C100 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C101 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.86fF
C102 sc_cmfb_0/transmission_gate_4/out VSS -5.46fF
C103 sc_cmfb_0/transmission_gate_3/out VSS -0.76fF
C104 p1 VSS 85.48fF
C105 sc_cmfb_0/transmission_gate_8/in VSS 1.87fF
C106 sc_cmfb_0/transmission_gate_6/in VSS -14.73fF
C107 sc_cmfb_0/transmission_gate_7/in VSS 8.08fF
C108 cm VSS 31.18fF
C109 op VSS 6.58fF
C110 p1_b VSS 108.59fF
C111 on VSS -10.34fF
C112 ota_w_test_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C113 ota_w_test_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF $ **FLOATING
C114 ota_w_test_v2_without_cmfb_0/m1_18877_3928# VSS 0.05fF $ **FLOATING
C115 ota_w_test_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C116 ota_w_test_v2_without_cmfb_0/li_11121_570# VSS 8.94fF
C117 ota_w_test_v2_without_cmfb_0/li_11122_5650# VSS 2.50fF
C118 ota_w_test_v2_without_cmfb_0/li_8434_570# VSS 9.31fF
C119 bias_a VSS -334.78fF
C120 ota_w_test_v2_without_cmfb_0/li_8436_5651# VSS 6.42fF
C121 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -342.22fF
C122 bias_b VSS -357.50fF
C123 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C124 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.85fF
C125 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C126 VDD VSS 343.80fF
C127 i_bias VSS -61.96fF
C128 bias_c VSS -129.75fF
C129 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C130 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C131 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C132 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C133 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C134 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C135 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C136 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C137 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.13fF
C138 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C139 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C140 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C141 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.14fF
C142 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C143 ota_w_test_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C144 bias_d VSS -229.59fF
C145 ota_w_test_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 4.65fF
C146 ota_w_test_v2_without_cmfb_0/li_14138_570# VSS 33.60fF
C147 cmc VSS -125.24fF
C148 in VSS -28.57fF
C149 ip VSS -28.50fF
.ends

