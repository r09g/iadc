magic
tech sky130A
timestamp 1654752884
<< end >>
