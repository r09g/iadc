magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< nwell >>
rect 1089 2796 1135 2842
rect 1405 2796 1451 2842
rect 1721 2796 1767 2842
rect 2037 2796 2083 2842
rect 2353 2796 2399 2842
rect 2669 2796 2715 2842
rect 2985 2796 3031 2842
rect 3301 2796 3347 2842
rect 141 1711 187 1814
rect 3301 1757 3347 1798
rect 3140 1501 3192 1544
<< pwell >>
rect 115 167 213 231
rect 431 167 529 231
rect 747 167 845 231
rect 1063 167 1161 231
rect 1379 167 1477 231
rect 1695 167 1793 231
rect 2011 167 2109 231
rect 2327 167 2425 231
rect 2643 167 2741 231
rect 2959 167 3057 231
<< mvndiff >>
rect 141 193 187 205
rect 457 193 503 205
rect 773 193 819 205
rect 1089 193 1135 205
rect 1405 193 1451 205
rect 1721 193 1767 205
rect 2037 193 2083 205
rect 2353 193 2399 205
rect 2669 193 2715 205
rect 2985 193 3031 205
<< mvpdiff >>
rect 1089 2796 1135 2798
rect 1405 2796 1451 2798
rect 1721 2796 1767 2798
rect 2037 2796 2083 2798
rect 2353 2796 2399 2798
rect 2669 2796 2715 2798
rect 2985 2796 3031 2798
rect 3301 2796 3347 2798
<< locali >>
rect 109 2983 143 3017
rect 177 2983 215 3017
rect 249 2983 287 3017
rect 321 2983 359 3017
rect 393 2983 431 3017
rect 465 2983 503 3017
rect 537 2983 575 3017
rect 609 2983 647 3017
rect 681 2983 719 3017
rect 753 2983 791 3017
rect 825 2983 863 3017
rect 897 2983 935 3017
rect 969 2983 1007 3017
rect 1041 2983 1079 3017
rect 1113 2983 1151 3017
rect 1185 2983 1223 3017
rect 1257 2983 1295 3017
rect 1329 2983 1367 3017
rect 1401 2983 1439 3017
rect 1473 2983 1511 3017
rect 1545 2983 1583 3017
rect 1617 2983 1655 3017
rect 1689 2983 1727 3017
rect 1761 2983 1799 3017
rect 1833 2983 1871 3017
rect 1905 2983 1943 3017
rect 1977 2983 2015 3017
rect 2049 2983 2087 3017
rect 2121 2983 2159 3017
rect 2193 2983 2231 3017
rect 2265 2983 2303 3017
rect 2337 2983 2375 3017
rect 2409 2983 2447 3017
rect 2481 2983 2519 3017
rect 2553 2983 2591 3017
rect 2625 2983 2663 3017
rect 2697 2983 2735 3017
rect 2769 2983 2807 3017
rect 2841 2983 2879 3017
rect 2913 2983 2951 3017
rect 2985 2983 3023 3017
rect 3057 2983 3095 3017
rect 3129 2983 3167 3017
rect 3201 2983 3239 3017
rect 3273 2983 3311 3017
rect 3345 2983 3379 3017
rect 13 2891 47 2921
rect 13 2819 47 2857
rect 3441 2891 3475 2921
rect 3441 2819 3475 2857
rect 1095 2796 1129 2802
rect 1411 2796 1445 2802
rect 1727 2796 1761 2802
rect 2043 2796 2077 2802
rect 2359 2796 2393 2802
rect 2675 2796 2709 2802
rect 2991 2796 3025 2802
rect 3307 2796 3341 2802
rect 13 2747 47 2785
rect 13 2675 47 2713
rect 13 2603 47 2641
rect 13 2531 47 2569
rect 13 2459 47 2497
rect 13 2387 47 2425
rect 13 2315 47 2353
rect 13 2243 47 2281
rect 13 2171 47 2209
rect 13 2099 47 2137
rect 13 2027 47 2065
rect 13 1955 47 1993
rect 13 1883 47 1921
rect 13 1811 47 1849
rect 13 1739 47 1777
rect 13 1675 47 1705
rect 3441 2747 3475 2785
rect 3441 2675 3475 2713
rect 3441 2603 3475 2641
rect 3441 2531 3475 2569
rect 3441 2459 3475 2497
rect 3441 2387 3475 2425
rect 3441 2315 3475 2353
rect 3441 2243 3475 2281
rect 3441 2171 3475 2209
rect 3441 2099 3475 2137
rect 3441 2027 3475 2065
rect 3441 1955 3475 1993
rect 3441 1883 3475 1921
rect 3441 1811 3475 1849
rect 3441 1739 3475 1777
rect 3441 1675 3475 1705
rect 13 1286 47 1307
rect 13 1214 47 1252
rect 13 1142 47 1180
rect 13 1070 47 1108
rect 13 998 47 1036
rect 13 926 47 964
rect 13 854 47 892
rect 13 782 47 820
rect 13 710 47 748
rect 13 638 47 676
rect 13 566 47 604
rect 13 494 47 532
rect 13 422 47 460
rect 13 350 47 388
rect 13 278 47 316
rect 13 206 47 244
rect 3441 1286 3475 1307
rect 3441 1214 3475 1252
rect 3441 1142 3475 1180
rect 3441 1070 3475 1108
rect 3441 998 3475 1036
rect 3441 926 3475 964
rect 3441 854 3475 892
rect 3441 782 3475 820
rect 3441 710 3475 748
rect 3441 638 3475 676
rect 3441 566 3475 604
rect 3441 494 3475 532
rect 3441 422 3475 460
rect 3441 350 3475 388
rect 3441 278 3475 316
rect 3441 206 3475 244
rect 147 189 181 205
rect 463 189 497 205
rect 779 189 813 205
rect 1095 189 1129 205
rect 1411 189 1445 205
rect 1727 189 1761 205
rect 2043 189 2077 205
rect 2359 189 2393 205
rect 2675 189 2709 205
rect 2991 189 3025 205
rect 13 134 47 172
rect 13 79 47 100
rect 3441 134 3475 172
rect 3441 79 3475 100
rect 109 -17 143 17
rect 177 -17 215 17
rect 249 -17 287 17
rect 321 -17 359 17
rect 393 -17 431 17
rect 465 -17 503 17
rect 537 -17 575 17
rect 609 -17 647 17
rect 681 -17 719 17
rect 753 -17 791 17
rect 825 -17 863 17
rect 897 -17 935 17
rect 969 -17 1007 17
rect 1041 -17 1079 17
rect 1113 -17 1151 17
rect 1185 -17 1223 17
rect 1257 -17 1295 17
rect 1329 -17 1367 17
rect 1401 -17 1439 17
rect 1473 -17 1511 17
rect 1545 -17 1583 17
rect 1617 -17 1655 17
rect 1689 -17 1727 17
rect 1761 -17 1799 17
rect 1833 -17 1871 17
rect 1905 -17 1943 17
rect 1977 -17 2015 17
rect 2049 -17 2087 17
rect 2121 -17 2159 17
rect 2193 -17 2231 17
rect 2265 -17 2303 17
rect 2337 -17 2375 17
rect 2409 -17 2447 17
rect 2481 -17 2519 17
rect 2553 -17 2591 17
rect 2625 -17 2663 17
rect 2697 -17 2735 17
rect 2769 -17 2807 17
rect 2841 -17 2879 17
rect 2913 -17 2951 17
rect 2985 -17 3023 17
rect 3057 -17 3095 17
rect 3129 -17 3167 17
rect 3201 -17 3239 17
rect 3273 -17 3311 17
rect 3345 -17 3379 17
<< viali >>
rect 143 2983 177 3017
rect 215 2983 249 3017
rect 287 2983 321 3017
rect 359 2983 393 3017
rect 431 2983 465 3017
rect 503 2983 537 3017
rect 575 2983 609 3017
rect 647 2983 681 3017
rect 719 2983 753 3017
rect 791 2983 825 3017
rect 863 2983 897 3017
rect 935 2983 969 3017
rect 1007 2983 1041 3017
rect 1079 2983 1113 3017
rect 1151 2983 1185 3017
rect 1223 2983 1257 3017
rect 1295 2983 1329 3017
rect 1367 2983 1401 3017
rect 1439 2983 1473 3017
rect 1511 2983 1545 3017
rect 1583 2983 1617 3017
rect 1655 2983 1689 3017
rect 1727 2983 1761 3017
rect 1799 2983 1833 3017
rect 1871 2983 1905 3017
rect 1943 2983 1977 3017
rect 2015 2983 2049 3017
rect 2087 2983 2121 3017
rect 2159 2983 2193 3017
rect 2231 2983 2265 3017
rect 2303 2983 2337 3017
rect 2375 2983 2409 3017
rect 2447 2983 2481 3017
rect 2519 2983 2553 3017
rect 2591 2983 2625 3017
rect 2663 2983 2697 3017
rect 2735 2983 2769 3017
rect 2807 2983 2841 3017
rect 2879 2983 2913 3017
rect 2951 2983 2985 3017
rect 3023 2983 3057 3017
rect 3095 2983 3129 3017
rect 3167 2983 3201 3017
rect 3239 2983 3273 3017
rect 3311 2983 3345 3017
rect 13 2857 47 2891
rect 13 2785 47 2819
rect 3441 2857 3475 2891
rect 13 2713 47 2747
rect 13 2641 47 2675
rect 13 2569 47 2603
rect 13 2497 47 2531
rect 13 2425 47 2459
rect 13 2353 47 2387
rect 13 2281 47 2315
rect 13 2209 47 2243
rect 13 2137 47 2171
rect 13 2065 47 2099
rect 13 1993 47 2027
rect 13 1921 47 1955
rect 13 1849 47 1883
rect 13 1777 47 1811
rect 13 1705 47 1739
rect 3441 2785 3475 2819
rect 3441 2713 3475 2747
rect 3441 2641 3475 2675
rect 3441 2569 3475 2603
rect 3441 2497 3475 2531
rect 3441 2425 3475 2459
rect 3441 2353 3475 2387
rect 3441 2281 3475 2315
rect 3441 2209 3475 2243
rect 3441 2137 3475 2171
rect 3441 2065 3475 2099
rect 3441 1993 3475 2027
rect 3441 1921 3475 1955
rect 3441 1849 3475 1883
rect 3441 1777 3475 1811
rect 3441 1705 3475 1739
rect 13 1252 47 1286
rect 13 1180 47 1214
rect 13 1108 47 1142
rect 13 1036 47 1070
rect 13 964 47 998
rect 13 892 47 926
rect 13 820 47 854
rect 13 748 47 782
rect 13 676 47 710
rect 13 604 47 638
rect 13 532 47 566
rect 13 460 47 494
rect 13 388 47 422
rect 13 316 47 350
rect 13 244 47 278
rect 13 172 47 206
rect 3441 1252 3475 1286
rect 3441 1180 3475 1214
rect 3441 1108 3475 1142
rect 3441 1036 3475 1070
rect 3441 964 3475 998
rect 3441 892 3475 926
rect 3441 820 3475 854
rect 3441 748 3475 782
rect 3441 676 3475 710
rect 3441 604 3475 638
rect 3441 532 3475 566
rect 3441 460 3475 494
rect 3441 388 3475 422
rect 3441 316 3475 350
rect 3441 244 3475 278
rect 13 100 47 134
rect 3441 172 3475 206
rect 3441 100 3475 134
rect 143 -17 177 17
rect 215 -17 249 17
rect 287 -17 321 17
rect 359 -17 393 17
rect 431 -17 465 17
rect 503 -17 537 17
rect 575 -17 609 17
rect 647 -17 681 17
rect 719 -17 753 17
rect 791 -17 825 17
rect 863 -17 897 17
rect 935 -17 969 17
rect 1007 -17 1041 17
rect 1079 -17 1113 17
rect 1151 -17 1185 17
rect 1223 -17 1257 17
rect 1295 -17 1329 17
rect 1367 -17 1401 17
rect 1439 -17 1473 17
rect 1511 -17 1545 17
rect 1583 -17 1617 17
rect 1655 -17 1689 17
rect 1727 -17 1761 17
rect 1799 -17 1833 17
rect 1871 -17 1905 17
rect 1943 -17 1977 17
rect 2015 -17 2049 17
rect 2087 -17 2121 17
rect 2159 -17 2193 17
rect 2231 -17 2265 17
rect 2303 -17 2337 17
rect 2375 -17 2409 17
rect 2447 -17 2481 17
rect 2519 -17 2553 17
rect 2591 -17 2625 17
rect 2663 -17 2697 17
rect 2735 -17 2769 17
rect 2807 -17 2841 17
rect 2879 -17 2913 17
rect 2951 -17 2985 17
rect 3023 -17 3057 17
rect 3095 -17 3129 17
rect 3167 -17 3201 17
rect 3239 -17 3273 17
rect 3311 -17 3345 17
<< metal1 >>
rect 7 3017 3481 3023
rect 7 2983 143 3017
rect 177 2983 215 3017
rect 249 2983 287 3017
rect 321 2983 359 3017
rect 393 2983 431 3017
rect 465 2983 503 3017
rect 537 2983 575 3017
rect 609 2983 647 3017
rect 681 2983 719 3017
rect 753 2983 791 3017
rect 825 2983 863 3017
rect 897 2983 935 3017
rect 969 2983 1007 3017
rect 1041 2983 1079 3017
rect 1113 2983 1151 3017
rect 1185 2983 1223 3017
rect 1257 2983 1295 3017
rect 1329 2983 1367 3017
rect 1401 2983 1439 3017
rect 1473 2983 1511 3017
rect 1545 2983 1583 3017
rect 1617 2983 1655 3017
rect 1689 2983 1727 3017
rect 1761 2983 1799 3017
rect 1833 2983 1871 3017
rect 1905 2983 1943 3017
rect 1977 2983 2015 3017
rect 2049 2983 2087 3017
rect 2121 2983 2159 3017
rect 2193 2983 2231 3017
rect 2265 2983 2303 3017
rect 2337 2983 2375 3017
rect 2409 2983 2447 3017
rect 2481 2983 2519 3017
rect 2553 2983 2591 3017
rect 2625 2983 2663 3017
rect 2697 2983 2735 3017
rect 2769 2983 2807 3017
rect 2841 2983 2879 3017
rect 2913 2983 2951 3017
rect 2985 2983 3023 3017
rect 3057 2983 3095 3017
rect 3129 2983 3167 3017
rect 3201 2983 3239 3017
rect 3273 2983 3311 3017
rect 3345 2983 3481 3017
rect 7 2891 3481 2983
rect 7 2857 13 2891
rect 47 2857 3441 2891
rect 3475 2857 3481 2891
rect 7 2839 3481 2857
rect 7 2819 59 2839
rect 7 2785 13 2819
rect 47 2785 59 2819
rect 141 2789 187 2839
rect 457 2795 503 2839
rect 773 2796 819 2839
rect 1089 2796 1135 2839
rect 1405 2796 1451 2839
rect 1721 2796 1767 2839
rect 2037 2796 2083 2839
rect 2353 2796 2399 2839
rect 2669 2796 2715 2839
rect 2985 2796 3031 2839
rect 3301 2796 3347 2839
rect 3429 2819 3481 2839
rect 7 2747 59 2785
rect 7 2713 13 2747
rect 47 2713 59 2747
rect 7 2675 59 2713
rect 7 2641 13 2675
rect 47 2641 59 2675
rect 7 2603 59 2641
rect 7 2569 13 2603
rect 47 2569 59 2603
rect 7 2531 59 2569
rect 7 2497 13 2531
rect 47 2497 59 2531
rect 7 2459 59 2497
rect 7 2425 13 2459
rect 47 2425 59 2459
rect 7 2387 59 2425
rect 7 2353 13 2387
rect 47 2353 59 2387
rect 7 2315 59 2353
rect 7 2281 13 2315
rect 47 2281 59 2315
rect 7 2243 59 2281
rect 7 2209 13 2243
rect 47 2209 59 2243
rect 7 2171 59 2209
rect 7 2137 13 2171
rect 47 2137 59 2171
rect 7 2099 59 2137
rect 7 2065 13 2099
rect 47 2065 59 2099
rect 7 2027 59 2065
rect 7 1993 13 2027
rect 47 1993 59 2027
rect 7 1955 59 1993
rect 7 1921 13 1955
rect 47 1921 59 1955
rect 7 1883 59 1921
rect 7 1849 13 1883
rect 47 1849 59 1883
rect 7 1811 59 1849
rect 286 2772 358 2786
rect 286 2720 296 2772
rect 348 2720 358 2772
rect 286 2708 358 2720
rect 286 2656 296 2708
rect 348 2656 358 2708
rect 286 2644 358 2656
rect 286 2592 296 2644
rect 348 2592 358 2644
rect 286 2580 358 2592
rect 286 2528 296 2580
rect 348 2528 358 2580
rect 286 2516 358 2528
rect 286 2464 296 2516
rect 348 2464 358 2516
rect 286 2452 358 2464
rect 286 2400 296 2452
rect 348 2400 358 2452
rect 286 2388 358 2400
rect 286 2336 296 2388
rect 348 2336 358 2388
rect 286 2324 358 2336
rect 286 2272 296 2324
rect 348 2272 358 2324
rect 286 2260 358 2272
rect 286 2208 296 2260
rect 348 2208 358 2260
rect 286 2196 358 2208
rect 286 2144 296 2196
rect 348 2144 358 2196
rect 286 2132 358 2144
rect 286 2080 296 2132
rect 348 2080 358 2132
rect 286 2068 358 2080
rect 286 2016 296 2068
rect 348 2016 358 2068
rect 286 2004 358 2016
rect 286 1952 296 2004
rect 348 1952 358 2004
rect 286 1940 358 1952
rect 286 1888 296 1940
rect 348 1888 358 1940
rect 286 1876 358 1888
rect 286 1824 296 1876
rect 348 1824 358 1876
rect 7 1777 13 1811
rect 47 1777 59 1811
rect 7 1757 59 1777
rect 141 1757 187 1814
rect 286 1810 358 1824
rect 602 2772 674 2786
rect 602 2720 612 2772
rect 664 2720 674 2772
rect 602 2708 674 2720
rect 602 2656 612 2708
rect 664 2656 674 2708
rect 602 2644 674 2656
rect 602 2592 612 2644
rect 664 2592 674 2644
rect 602 2580 674 2592
rect 602 2528 612 2580
rect 664 2528 674 2580
rect 602 2516 674 2528
rect 602 2464 612 2516
rect 664 2464 674 2516
rect 602 2452 674 2464
rect 602 2400 612 2452
rect 664 2400 674 2452
rect 602 2388 674 2400
rect 602 2336 612 2388
rect 664 2336 674 2388
rect 602 2324 674 2336
rect 602 2272 612 2324
rect 664 2272 674 2324
rect 602 2260 674 2272
rect 602 2208 612 2260
rect 664 2208 674 2260
rect 602 2196 674 2208
rect 602 2144 612 2196
rect 664 2144 674 2196
rect 602 2132 674 2144
rect 602 2080 612 2132
rect 664 2080 674 2132
rect 602 2068 674 2080
rect 602 2016 612 2068
rect 664 2016 674 2068
rect 602 2004 674 2016
rect 602 1952 612 2004
rect 664 1952 674 2004
rect 602 1940 674 1952
rect 602 1888 612 1940
rect 664 1888 674 1940
rect 602 1876 674 1888
rect 602 1824 612 1876
rect 664 1824 674 1876
rect 602 1810 674 1824
rect 918 2772 990 2786
rect 918 2720 928 2772
rect 980 2720 990 2772
rect 918 2708 990 2720
rect 918 2656 928 2708
rect 980 2656 990 2708
rect 918 2644 990 2656
rect 918 2592 928 2644
rect 980 2592 990 2644
rect 918 2580 990 2592
rect 918 2528 928 2580
rect 980 2528 990 2580
rect 918 2516 990 2528
rect 918 2464 928 2516
rect 980 2464 990 2516
rect 918 2452 990 2464
rect 918 2400 928 2452
rect 980 2400 990 2452
rect 918 2388 990 2400
rect 918 2336 928 2388
rect 980 2336 990 2388
rect 918 2324 990 2336
rect 918 2272 928 2324
rect 980 2272 990 2324
rect 918 2260 990 2272
rect 918 2208 928 2260
rect 980 2208 990 2260
rect 918 2196 990 2208
rect 918 2144 928 2196
rect 980 2144 990 2196
rect 918 2132 990 2144
rect 918 2080 928 2132
rect 980 2080 990 2132
rect 918 2068 990 2080
rect 918 2016 928 2068
rect 980 2016 990 2068
rect 918 2004 990 2016
rect 918 1952 928 2004
rect 980 1952 990 2004
rect 918 1940 990 1952
rect 918 1888 928 1940
rect 980 1888 990 1940
rect 918 1876 990 1888
rect 918 1824 928 1876
rect 980 1824 990 1876
rect 918 1810 990 1824
rect 1234 2772 1306 2786
rect 1234 2720 1244 2772
rect 1296 2720 1306 2772
rect 1234 2708 1306 2720
rect 1234 2656 1244 2708
rect 1296 2656 1306 2708
rect 1234 2644 1306 2656
rect 1234 2592 1244 2644
rect 1296 2592 1306 2644
rect 1234 2580 1306 2592
rect 1234 2528 1244 2580
rect 1296 2528 1306 2580
rect 1234 2516 1306 2528
rect 1234 2464 1244 2516
rect 1296 2464 1306 2516
rect 1234 2452 1306 2464
rect 1234 2400 1244 2452
rect 1296 2400 1306 2452
rect 1234 2388 1306 2400
rect 1234 2336 1244 2388
rect 1296 2336 1306 2388
rect 1234 2324 1306 2336
rect 1234 2272 1244 2324
rect 1296 2272 1306 2324
rect 1234 2260 1306 2272
rect 1234 2208 1244 2260
rect 1296 2208 1306 2260
rect 1234 2196 1306 2208
rect 1234 2144 1244 2196
rect 1296 2144 1306 2196
rect 1234 2132 1306 2144
rect 1234 2080 1244 2132
rect 1296 2080 1306 2132
rect 1234 2068 1306 2080
rect 1234 2016 1244 2068
rect 1296 2016 1306 2068
rect 1234 2004 1306 2016
rect 1234 1952 1244 2004
rect 1296 1952 1306 2004
rect 1234 1940 1306 1952
rect 1234 1888 1244 1940
rect 1296 1888 1306 1940
rect 1234 1876 1306 1888
rect 1234 1824 1244 1876
rect 1296 1824 1306 1876
rect 1234 1810 1306 1824
rect 1550 2772 1622 2786
rect 1550 2720 1560 2772
rect 1612 2720 1622 2772
rect 1550 2708 1622 2720
rect 1550 2656 1560 2708
rect 1612 2656 1622 2708
rect 1550 2644 1622 2656
rect 1550 2592 1560 2644
rect 1612 2592 1622 2644
rect 1550 2580 1622 2592
rect 1550 2528 1560 2580
rect 1612 2528 1622 2580
rect 1550 2516 1622 2528
rect 1550 2464 1560 2516
rect 1612 2464 1622 2516
rect 1550 2452 1622 2464
rect 1550 2400 1560 2452
rect 1612 2400 1622 2452
rect 1550 2388 1622 2400
rect 1550 2336 1560 2388
rect 1612 2336 1622 2388
rect 1550 2324 1622 2336
rect 1550 2272 1560 2324
rect 1612 2272 1622 2324
rect 1550 2260 1622 2272
rect 1550 2208 1560 2260
rect 1612 2208 1622 2260
rect 1550 2196 1622 2208
rect 1550 2144 1560 2196
rect 1612 2144 1622 2196
rect 1550 2132 1622 2144
rect 1550 2080 1560 2132
rect 1612 2080 1622 2132
rect 1550 2068 1622 2080
rect 1550 2016 1560 2068
rect 1612 2016 1622 2068
rect 1550 2004 1622 2016
rect 1550 1952 1560 2004
rect 1612 1952 1622 2004
rect 1550 1940 1622 1952
rect 1550 1888 1560 1940
rect 1612 1888 1622 1940
rect 1550 1876 1622 1888
rect 1550 1824 1560 1876
rect 1612 1824 1622 1876
rect 1550 1810 1622 1824
rect 1866 2772 1938 2786
rect 1866 2720 1876 2772
rect 1928 2720 1938 2772
rect 1866 2708 1938 2720
rect 1866 2656 1876 2708
rect 1928 2656 1938 2708
rect 1866 2644 1938 2656
rect 1866 2592 1876 2644
rect 1928 2592 1938 2644
rect 1866 2580 1938 2592
rect 1866 2528 1876 2580
rect 1928 2528 1938 2580
rect 1866 2516 1938 2528
rect 1866 2464 1876 2516
rect 1928 2464 1938 2516
rect 1866 2452 1938 2464
rect 1866 2400 1876 2452
rect 1928 2400 1938 2452
rect 1866 2388 1938 2400
rect 1866 2336 1876 2388
rect 1928 2336 1938 2388
rect 1866 2324 1938 2336
rect 1866 2272 1876 2324
rect 1928 2272 1938 2324
rect 1866 2260 1938 2272
rect 1866 2208 1876 2260
rect 1928 2208 1938 2260
rect 1866 2196 1938 2208
rect 1866 2144 1876 2196
rect 1928 2144 1938 2196
rect 1866 2132 1938 2144
rect 1866 2080 1876 2132
rect 1928 2080 1938 2132
rect 1866 2068 1938 2080
rect 1866 2016 1876 2068
rect 1928 2016 1938 2068
rect 1866 2004 1938 2016
rect 1866 1952 1876 2004
rect 1928 1952 1938 2004
rect 1866 1940 1938 1952
rect 1866 1888 1876 1940
rect 1928 1888 1938 1940
rect 1866 1876 1938 1888
rect 1866 1824 1876 1876
rect 1928 1824 1938 1876
rect 1866 1810 1938 1824
rect 2182 2772 2254 2786
rect 2182 2720 2192 2772
rect 2244 2720 2254 2772
rect 2182 2708 2254 2720
rect 2182 2656 2192 2708
rect 2244 2656 2254 2708
rect 2182 2644 2254 2656
rect 2182 2592 2192 2644
rect 2244 2592 2254 2644
rect 2182 2580 2254 2592
rect 2182 2528 2192 2580
rect 2244 2528 2254 2580
rect 2182 2516 2254 2528
rect 2182 2464 2192 2516
rect 2244 2464 2254 2516
rect 2182 2452 2254 2464
rect 2182 2400 2192 2452
rect 2244 2400 2254 2452
rect 2182 2388 2254 2400
rect 2182 2336 2192 2388
rect 2244 2336 2254 2388
rect 2182 2324 2254 2336
rect 2182 2272 2192 2324
rect 2244 2272 2254 2324
rect 2182 2260 2254 2272
rect 2182 2208 2192 2260
rect 2244 2208 2254 2260
rect 2182 2196 2254 2208
rect 2182 2144 2192 2196
rect 2244 2144 2254 2196
rect 2182 2132 2254 2144
rect 2182 2080 2192 2132
rect 2244 2080 2254 2132
rect 2182 2068 2254 2080
rect 2182 2016 2192 2068
rect 2244 2016 2254 2068
rect 2182 2004 2254 2016
rect 2182 1952 2192 2004
rect 2244 1952 2254 2004
rect 2182 1940 2254 1952
rect 2182 1888 2192 1940
rect 2244 1888 2254 1940
rect 2182 1876 2254 1888
rect 2182 1824 2192 1876
rect 2244 1824 2254 1876
rect 2182 1810 2254 1824
rect 2498 2772 2570 2786
rect 2498 2720 2508 2772
rect 2560 2720 2570 2772
rect 2498 2708 2570 2720
rect 2498 2656 2508 2708
rect 2560 2656 2570 2708
rect 2498 2644 2570 2656
rect 2498 2592 2508 2644
rect 2560 2592 2570 2644
rect 2498 2580 2570 2592
rect 2498 2528 2508 2580
rect 2560 2528 2570 2580
rect 2498 2516 2570 2528
rect 2498 2464 2508 2516
rect 2560 2464 2570 2516
rect 2498 2452 2570 2464
rect 2498 2400 2508 2452
rect 2560 2400 2570 2452
rect 2498 2388 2570 2400
rect 2498 2336 2508 2388
rect 2560 2336 2570 2388
rect 2498 2324 2570 2336
rect 2498 2272 2508 2324
rect 2560 2272 2570 2324
rect 2498 2260 2570 2272
rect 2498 2208 2508 2260
rect 2560 2208 2570 2260
rect 2498 2196 2570 2208
rect 2498 2144 2508 2196
rect 2560 2144 2570 2196
rect 2498 2132 2570 2144
rect 2498 2080 2508 2132
rect 2560 2080 2570 2132
rect 2498 2068 2570 2080
rect 2498 2016 2508 2068
rect 2560 2016 2570 2068
rect 2498 2004 2570 2016
rect 2498 1952 2508 2004
rect 2560 1952 2570 2004
rect 2498 1940 2570 1952
rect 2498 1888 2508 1940
rect 2560 1888 2570 1940
rect 2498 1876 2570 1888
rect 2498 1824 2508 1876
rect 2560 1824 2570 1876
rect 2498 1810 2570 1824
rect 2814 2772 2886 2786
rect 2814 2720 2824 2772
rect 2876 2720 2886 2772
rect 2814 2708 2886 2720
rect 2814 2656 2824 2708
rect 2876 2656 2886 2708
rect 2814 2644 2886 2656
rect 2814 2592 2824 2644
rect 2876 2592 2886 2644
rect 2814 2580 2886 2592
rect 2814 2528 2824 2580
rect 2876 2528 2886 2580
rect 2814 2516 2886 2528
rect 2814 2464 2824 2516
rect 2876 2464 2886 2516
rect 2814 2452 2886 2464
rect 2814 2400 2824 2452
rect 2876 2400 2886 2452
rect 2814 2388 2886 2400
rect 2814 2336 2824 2388
rect 2876 2336 2886 2388
rect 2814 2324 2886 2336
rect 2814 2272 2824 2324
rect 2876 2272 2886 2324
rect 2814 2260 2886 2272
rect 2814 2208 2824 2260
rect 2876 2208 2886 2260
rect 2814 2196 2886 2208
rect 2814 2144 2824 2196
rect 2876 2144 2886 2196
rect 2814 2132 2886 2144
rect 2814 2080 2824 2132
rect 2876 2080 2886 2132
rect 2814 2068 2886 2080
rect 2814 2016 2824 2068
rect 2876 2016 2886 2068
rect 2814 2004 2886 2016
rect 2814 1952 2824 2004
rect 2876 1952 2886 2004
rect 2814 1940 2886 1952
rect 2814 1888 2824 1940
rect 2876 1888 2886 1940
rect 2814 1876 2886 1888
rect 2814 1824 2824 1876
rect 2876 1824 2886 1876
rect 2814 1810 2886 1824
rect 3130 2772 3202 2786
rect 3130 2720 3140 2772
rect 3192 2720 3202 2772
rect 3130 2708 3202 2720
rect 3130 2656 3140 2708
rect 3192 2656 3202 2708
rect 3130 2644 3202 2656
rect 3130 2592 3140 2644
rect 3192 2592 3202 2644
rect 3130 2580 3202 2592
rect 3130 2528 3140 2580
rect 3192 2528 3202 2580
rect 3130 2516 3202 2528
rect 3130 2464 3140 2516
rect 3192 2464 3202 2516
rect 3130 2452 3202 2464
rect 3130 2400 3140 2452
rect 3192 2400 3202 2452
rect 3130 2388 3202 2400
rect 3130 2336 3140 2388
rect 3192 2336 3202 2388
rect 3130 2324 3202 2336
rect 3130 2272 3140 2324
rect 3192 2272 3202 2324
rect 3130 2260 3202 2272
rect 3130 2208 3140 2260
rect 3192 2208 3202 2260
rect 3130 2196 3202 2208
rect 3130 2144 3140 2196
rect 3192 2144 3202 2196
rect 3130 2132 3202 2144
rect 3130 2080 3140 2132
rect 3192 2080 3202 2132
rect 3130 2068 3202 2080
rect 3130 2016 3140 2068
rect 3192 2016 3202 2068
rect 3130 2004 3202 2016
rect 3130 1952 3140 2004
rect 3192 1952 3202 2004
rect 3130 1940 3202 1952
rect 3130 1888 3140 1940
rect 3192 1888 3202 1940
rect 3130 1876 3202 1888
rect 3130 1824 3140 1876
rect 3192 1824 3202 1876
rect 3130 1810 3202 1824
rect 3429 2785 3441 2819
rect 3475 2785 3481 2819
rect 3429 2747 3481 2785
rect 3429 2713 3441 2747
rect 3475 2713 3481 2747
rect 3429 2675 3481 2713
rect 3429 2641 3441 2675
rect 3475 2641 3481 2675
rect 3429 2603 3481 2641
rect 3429 2569 3441 2603
rect 3475 2569 3481 2603
rect 3429 2531 3481 2569
rect 3429 2497 3441 2531
rect 3475 2497 3481 2531
rect 3429 2459 3481 2497
rect 3429 2425 3441 2459
rect 3475 2425 3481 2459
rect 3429 2387 3481 2425
rect 3429 2353 3441 2387
rect 3475 2353 3481 2387
rect 3429 2315 3481 2353
rect 3429 2281 3441 2315
rect 3475 2281 3481 2315
rect 3429 2243 3481 2281
rect 3429 2209 3441 2243
rect 3475 2209 3481 2243
rect 3429 2171 3481 2209
rect 3429 2137 3441 2171
rect 3475 2137 3481 2171
rect 3429 2099 3481 2137
rect 3429 2065 3441 2099
rect 3475 2065 3481 2099
rect 3429 2027 3481 2065
rect 3429 1993 3441 2027
rect 3475 1993 3481 2027
rect 3429 1955 3481 1993
rect 3429 1921 3441 1955
rect 3475 1921 3481 1955
rect 3429 1883 3481 1921
rect 3429 1849 3441 1883
rect 3475 1849 3481 1883
rect 3429 1811 3481 1849
rect 3301 1757 3347 1798
rect 3429 1777 3441 1811
rect 3475 1777 3481 1811
rect 3429 1757 3481 1777
rect 7 1739 3481 1757
rect 7 1705 13 1739
rect 47 1711 3441 1739
rect 47 1705 53 1711
rect 7 1663 53 1705
rect 3435 1705 3441 1711
rect 3475 1705 3481 1739
rect 3435 1663 3481 1705
rect -65 1518 3553 1555
rect -65 1466 296 1518
rect 348 1466 612 1518
rect 664 1466 928 1518
rect 980 1466 1244 1518
rect 1296 1466 1560 1518
rect 1612 1466 1876 1518
rect 1928 1466 2192 1518
rect 2244 1466 2508 1518
rect 2560 1466 2824 1518
rect 2876 1466 3140 1518
rect 3192 1466 3553 1518
rect -65 1427 3553 1466
rect 7 1286 53 1319
rect 7 1252 13 1286
rect 47 1271 53 1286
rect 3435 1286 3481 1319
rect 3435 1271 3441 1286
rect 47 1252 3441 1271
rect 3475 1252 3481 1286
rect 7 1225 3481 1252
rect 7 1214 53 1225
rect 7 1180 13 1214
rect 47 1180 53 1214
rect 3301 1189 3347 1225
rect 3435 1214 3481 1225
rect 7 1142 53 1180
rect 7 1108 13 1142
rect 47 1108 53 1142
rect 7 1070 53 1108
rect 7 1036 13 1070
rect 47 1036 53 1070
rect 7 998 53 1036
rect 7 964 13 998
rect 47 964 53 998
rect 7 926 53 964
rect 7 892 13 926
rect 47 892 53 926
rect 7 854 53 892
rect 7 820 13 854
rect 47 820 53 854
rect 7 782 53 820
rect 7 748 13 782
rect 47 748 53 782
rect 7 710 53 748
rect 7 676 13 710
rect 47 676 53 710
rect 7 638 53 676
rect 7 604 13 638
rect 47 604 53 638
rect 7 566 53 604
rect 7 532 13 566
rect 47 532 53 566
rect 7 494 53 532
rect 7 460 13 494
rect 47 460 53 494
rect 7 422 53 460
rect 7 388 13 422
rect 47 388 53 422
rect 7 350 53 388
rect 7 316 13 350
rect 47 316 53 350
rect 7 278 53 316
rect 7 244 13 278
rect 47 244 53 278
rect 7 206 53 244
rect 7 172 13 206
rect 47 172 53 206
rect 286 1167 358 1181
rect 286 1115 296 1167
rect 348 1115 358 1167
rect 286 1103 358 1115
rect 286 1051 296 1103
rect 348 1051 358 1103
rect 286 1039 358 1051
rect 286 987 296 1039
rect 348 987 358 1039
rect 286 975 358 987
rect 286 923 296 975
rect 348 923 358 975
rect 286 911 358 923
rect 286 859 296 911
rect 348 859 358 911
rect 286 847 358 859
rect 286 795 296 847
rect 348 795 358 847
rect 286 783 358 795
rect 286 731 296 783
rect 348 731 358 783
rect 286 719 358 731
rect 286 667 296 719
rect 348 667 358 719
rect 286 655 358 667
rect 286 603 296 655
rect 348 603 358 655
rect 286 591 358 603
rect 286 539 296 591
rect 348 539 358 591
rect 286 527 358 539
rect 286 475 296 527
rect 348 475 358 527
rect 286 463 358 475
rect 286 411 296 463
rect 348 411 358 463
rect 286 399 358 411
rect 286 347 296 399
rect 348 347 358 399
rect 286 335 358 347
rect 286 283 296 335
rect 348 283 358 335
rect 286 271 358 283
rect 286 219 296 271
rect 348 219 358 271
rect 286 205 358 219
rect 602 1167 674 1181
rect 602 1115 612 1167
rect 664 1115 674 1167
rect 602 1103 674 1115
rect 602 1051 612 1103
rect 664 1051 674 1103
rect 602 1039 674 1051
rect 602 987 612 1039
rect 664 987 674 1039
rect 602 975 674 987
rect 602 923 612 975
rect 664 923 674 975
rect 602 911 674 923
rect 602 859 612 911
rect 664 859 674 911
rect 602 847 674 859
rect 602 795 612 847
rect 664 795 674 847
rect 602 783 674 795
rect 602 731 612 783
rect 664 731 674 783
rect 602 719 674 731
rect 602 667 612 719
rect 664 667 674 719
rect 602 655 674 667
rect 602 603 612 655
rect 664 603 674 655
rect 602 591 674 603
rect 602 539 612 591
rect 664 539 674 591
rect 602 527 674 539
rect 602 475 612 527
rect 664 475 674 527
rect 602 463 674 475
rect 602 411 612 463
rect 664 411 674 463
rect 602 399 674 411
rect 602 347 612 399
rect 664 347 674 399
rect 602 335 674 347
rect 602 283 612 335
rect 664 283 674 335
rect 602 271 674 283
rect 602 219 612 271
rect 664 219 674 271
rect 602 205 674 219
rect 918 1167 990 1181
rect 918 1115 928 1167
rect 980 1115 990 1167
rect 918 1103 990 1115
rect 918 1051 928 1103
rect 980 1051 990 1103
rect 918 1039 990 1051
rect 918 987 928 1039
rect 980 987 990 1039
rect 918 975 990 987
rect 918 923 928 975
rect 980 923 990 975
rect 918 911 990 923
rect 918 859 928 911
rect 980 859 990 911
rect 918 847 990 859
rect 918 795 928 847
rect 980 795 990 847
rect 918 783 990 795
rect 918 731 928 783
rect 980 731 990 783
rect 918 719 990 731
rect 918 667 928 719
rect 980 667 990 719
rect 918 655 990 667
rect 918 603 928 655
rect 980 603 990 655
rect 918 591 990 603
rect 918 539 928 591
rect 980 539 990 591
rect 918 527 990 539
rect 918 475 928 527
rect 980 475 990 527
rect 918 463 990 475
rect 918 411 928 463
rect 980 411 990 463
rect 918 399 990 411
rect 918 347 928 399
rect 980 347 990 399
rect 918 335 990 347
rect 918 283 928 335
rect 980 283 990 335
rect 918 271 990 283
rect 918 219 928 271
rect 980 219 990 271
rect 918 205 990 219
rect 1234 1167 1306 1181
rect 1234 1115 1244 1167
rect 1296 1115 1306 1167
rect 1234 1103 1306 1115
rect 1234 1051 1244 1103
rect 1296 1051 1306 1103
rect 1234 1039 1306 1051
rect 1234 987 1244 1039
rect 1296 987 1306 1039
rect 1234 975 1306 987
rect 1234 923 1244 975
rect 1296 923 1306 975
rect 1234 911 1306 923
rect 1234 859 1244 911
rect 1296 859 1306 911
rect 1234 847 1306 859
rect 1234 795 1244 847
rect 1296 795 1306 847
rect 1234 783 1306 795
rect 1234 731 1244 783
rect 1296 731 1306 783
rect 1234 719 1306 731
rect 1234 667 1244 719
rect 1296 667 1306 719
rect 1234 655 1306 667
rect 1234 603 1244 655
rect 1296 603 1306 655
rect 1234 591 1306 603
rect 1234 539 1244 591
rect 1296 539 1306 591
rect 1234 527 1306 539
rect 1234 475 1244 527
rect 1296 475 1306 527
rect 1234 463 1306 475
rect 1234 411 1244 463
rect 1296 411 1306 463
rect 1234 399 1306 411
rect 1234 347 1244 399
rect 1296 347 1306 399
rect 1234 335 1306 347
rect 1234 283 1244 335
rect 1296 283 1306 335
rect 1234 271 1306 283
rect 1234 219 1244 271
rect 1296 219 1306 271
rect 1234 205 1306 219
rect 1550 1167 1622 1181
rect 1550 1115 1560 1167
rect 1612 1115 1622 1167
rect 1550 1103 1622 1115
rect 1550 1051 1560 1103
rect 1612 1051 1622 1103
rect 1550 1039 1622 1051
rect 1550 987 1560 1039
rect 1612 987 1622 1039
rect 1550 975 1622 987
rect 1550 923 1560 975
rect 1612 923 1622 975
rect 1550 911 1622 923
rect 1550 859 1560 911
rect 1612 859 1622 911
rect 1550 847 1622 859
rect 1550 795 1560 847
rect 1612 795 1622 847
rect 1550 783 1622 795
rect 1550 731 1560 783
rect 1612 731 1622 783
rect 1550 719 1622 731
rect 1550 667 1560 719
rect 1612 667 1622 719
rect 1550 655 1622 667
rect 1550 603 1560 655
rect 1612 603 1622 655
rect 1550 591 1622 603
rect 1550 539 1560 591
rect 1612 539 1622 591
rect 1550 527 1622 539
rect 1550 475 1560 527
rect 1612 475 1622 527
rect 1550 463 1622 475
rect 1550 411 1560 463
rect 1612 411 1622 463
rect 1550 399 1622 411
rect 1550 347 1560 399
rect 1612 347 1622 399
rect 1550 335 1622 347
rect 1550 283 1560 335
rect 1612 283 1622 335
rect 1550 271 1622 283
rect 1550 219 1560 271
rect 1612 219 1622 271
rect 1550 205 1622 219
rect 1866 1167 1938 1181
rect 1866 1115 1876 1167
rect 1928 1115 1938 1167
rect 1866 1103 1938 1115
rect 1866 1051 1876 1103
rect 1928 1051 1938 1103
rect 1866 1039 1938 1051
rect 1866 987 1876 1039
rect 1928 987 1938 1039
rect 1866 975 1938 987
rect 1866 923 1876 975
rect 1928 923 1938 975
rect 1866 911 1938 923
rect 1866 859 1876 911
rect 1928 859 1938 911
rect 1866 847 1938 859
rect 1866 795 1876 847
rect 1928 795 1938 847
rect 1866 783 1938 795
rect 1866 731 1876 783
rect 1928 731 1938 783
rect 1866 719 1938 731
rect 1866 667 1876 719
rect 1928 667 1938 719
rect 1866 655 1938 667
rect 1866 603 1876 655
rect 1928 603 1938 655
rect 1866 591 1938 603
rect 1866 539 1876 591
rect 1928 539 1938 591
rect 1866 527 1938 539
rect 1866 475 1876 527
rect 1928 475 1938 527
rect 1866 463 1938 475
rect 1866 411 1876 463
rect 1928 411 1938 463
rect 1866 399 1938 411
rect 1866 347 1876 399
rect 1928 347 1938 399
rect 1866 335 1938 347
rect 1866 283 1876 335
rect 1928 283 1938 335
rect 1866 271 1938 283
rect 1866 219 1876 271
rect 1928 219 1938 271
rect 1866 205 1938 219
rect 2182 1167 2254 1181
rect 2182 1115 2192 1167
rect 2244 1115 2254 1167
rect 2182 1103 2254 1115
rect 2182 1051 2192 1103
rect 2244 1051 2254 1103
rect 2182 1039 2254 1051
rect 2182 987 2192 1039
rect 2244 987 2254 1039
rect 2182 975 2254 987
rect 2182 923 2192 975
rect 2244 923 2254 975
rect 2182 911 2254 923
rect 2182 859 2192 911
rect 2244 859 2254 911
rect 2182 847 2254 859
rect 2182 795 2192 847
rect 2244 795 2254 847
rect 2182 783 2254 795
rect 2182 731 2192 783
rect 2244 731 2254 783
rect 2182 719 2254 731
rect 2182 667 2192 719
rect 2244 667 2254 719
rect 2182 655 2254 667
rect 2182 603 2192 655
rect 2244 603 2254 655
rect 2182 591 2254 603
rect 2182 539 2192 591
rect 2244 539 2254 591
rect 2182 527 2254 539
rect 2182 475 2192 527
rect 2244 475 2254 527
rect 2182 463 2254 475
rect 2182 411 2192 463
rect 2244 411 2254 463
rect 2182 399 2254 411
rect 2182 347 2192 399
rect 2244 347 2254 399
rect 2182 335 2254 347
rect 2182 283 2192 335
rect 2244 283 2254 335
rect 2182 271 2254 283
rect 2182 219 2192 271
rect 2244 219 2254 271
rect 2182 205 2254 219
rect 2498 1167 2570 1181
rect 2498 1115 2508 1167
rect 2560 1115 2570 1167
rect 2498 1103 2570 1115
rect 2498 1051 2508 1103
rect 2560 1051 2570 1103
rect 2498 1039 2570 1051
rect 2498 987 2508 1039
rect 2560 987 2570 1039
rect 2498 975 2570 987
rect 2498 923 2508 975
rect 2560 923 2570 975
rect 2498 911 2570 923
rect 2498 859 2508 911
rect 2560 859 2570 911
rect 2498 847 2570 859
rect 2498 795 2508 847
rect 2560 795 2570 847
rect 2498 783 2570 795
rect 2498 731 2508 783
rect 2560 731 2570 783
rect 2498 719 2570 731
rect 2498 667 2508 719
rect 2560 667 2570 719
rect 2498 655 2570 667
rect 2498 603 2508 655
rect 2560 603 2570 655
rect 2498 591 2570 603
rect 2498 539 2508 591
rect 2560 539 2570 591
rect 2498 527 2570 539
rect 2498 475 2508 527
rect 2560 475 2570 527
rect 2498 463 2570 475
rect 2498 411 2508 463
rect 2560 411 2570 463
rect 2498 399 2570 411
rect 2498 347 2508 399
rect 2560 347 2570 399
rect 2498 335 2570 347
rect 2498 283 2508 335
rect 2560 283 2570 335
rect 2498 271 2570 283
rect 2498 219 2508 271
rect 2560 219 2570 271
rect 2498 205 2570 219
rect 2814 1167 2886 1181
rect 2814 1115 2824 1167
rect 2876 1115 2886 1167
rect 2814 1103 2886 1115
rect 2814 1051 2824 1103
rect 2876 1051 2886 1103
rect 2814 1039 2886 1051
rect 2814 987 2824 1039
rect 2876 987 2886 1039
rect 2814 975 2886 987
rect 2814 923 2824 975
rect 2876 923 2886 975
rect 2814 911 2886 923
rect 2814 859 2824 911
rect 2876 859 2886 911
rect 2814 847 2886 859
rect 2814 795 2824 847
rect 2876 795 2886 847
rect 2814 783 2886 795
rect 2814 731 2824 783
rect 2876 731 2886 783
rect 2814 719 2886 731
rect 2814 667 2824 719
rect 2876 667 2886 719
rect 2814 655 2886 667
rect 2814 603 2824 655
rect 2876 603 2886 655
rect 2814 591 2886 603
rect 2814 539 2824 591
rect 2876 539 2886 591
rect 2814 527 2886 539
rect 2814 475 2824 527
rect 2876 475 2886 527
rect 2814 463 2886 475
rect 2814 411 2824 463
rect 2876 411 2886 463
rect 2814 399 2886 411
rect 2814 347 2824 399
rect 2876 347 2886 399
rect 2814 335 2886 347
rect 2814 283 2824 335
rect 2876 283 2886 335
rect 2814 271 2886 283
rect 2814 219 2824 271
rect 2876 219 2886 271
rect 2814 205 2886 219
rect 3130 1167 3202 1181
rect 3130 1115 3140 1167
rect 3192 1115 3202 1167
rect 3130 1103 3202 1115
rect 3130 1051 3140 1103
rect 3192 1051 3202 1103
rect 3130 1039 3202 1051
rect 3130 987 3140 1039
rect 3192 987 3202 1039
rect 3130 975 3202 987
rect 3130 923 3140 975
rect 3192 923 3202 975
rect 3130 911 3202 923
rect 3130 859 3140 911
rect 3192 859 3202 911
rect 3130 847 3202 859
rect 3130 795 3140 847
rect 3192 795 3202 847
rect 3130 783 3202 795
rect 3130 731 3140 783
rect 3192 731 3202 783
rect 3130 719 3202 731
rect 3130 667 3140 719
rect 3192 667 3202 719
rect 3130 655 3202 667
rect 3130 603 3140 655
rect 3192 603 3202 655
rect 3130 591 3202 603
rect 3130 539 3140 591
rect 3192 539 3202 591
rect 3130 527 3202 539
rect 3130 475 3140 527
rect 3192 475 3202 527
rect 3130 463 3202 475
rect 3130 411 3140 463
rect 3192 411 3202 463
rect 3130 399 3202 411
rect 3130 347 3140 399
rect 3192 347 3202 399
rect 3130 335 3202 347
rect 3130 283 3140 335
rect 3192 283 3202 335
rect 3130 271 3202 283
rect 3130 219 3140 271
rect 3192 219 3202 271
rect 3130 205 3202 219
rect 3435 1180 3441 1214
rect 3475 1180 3481 1214
rect 3435 1142 3481 1180
rect 3435 1108 3441 1142
rect 3475 1108 3481 1142
rect 3435 1070 3481 1108
rect 3435 1036 3441 1070
rect 3475 1036 3481 1070
rect 3435 998 3481 1036
rect 3435 964 3441 998
rect 3475 964 3481 998
rect 3435 926 3481 964
rect 3435 892 3441 926
rect 3475 892 3481 926
rect 3435 854 3481 892
rect 3435 820 3441 854
rect 3475 820 3481 854
rect 3435 782 3481 820
rect 3435 748 3441 782
rect 3475 748 3481 782
rect 3435 710 3481 748
rect 3435 676 3441 710
rect 3475 676 3481 710
rect 3435 638 3481 676
rect 3435 604 3441 638
rect 3475 604 3481 638
rect 3435 566 3481 604
rect 3435 532 3441 566
rect 3475 532 3481 566
rect 3435 494 3481 532
rect 3435 460 3441 494
rect 3475 460 3481 494
rect 3435 422 3481 460
rect 3435 388 3441 422
rect 3475 388 3481 422
rect 3435 350 3481 388
rect 3435 316 3441 350
rect 3475 316 3481 350
rect 3435 278 3481 316
rect 3435 244 3441 278
rect 3475 244 3481 278
rect 3435 206 3481 244
rect 7 161 53 172
rect 141 161 187 205
rect 457 161 503 205
rect 773 161 819 205
rect 1089 161 1135 205
rect 1405 161 1451 205
rect 1721 161 1767 205
rect 2037 161 2083 205
rect 2353 161 2399 205
rect 2669 161 2715 205
rect 2985 161 3031 205
rect 3301 161 3347 204
rect 3435 172 3441 206
rect 3475 172 3481 206
rect 3435 161 3481 172
rect 7 134 3481 161
rect 7 100 13 134
rect 47 100 3441 134
rect 3475 100 3481 134
rect 7 17 3481 100
rect 7 -17 143 17
rect 177 -17 215 17
rect 249 -17 287 17
rect 321 -17 359 17
rect 393 -17 431 17
rect 465 -17 503 17
rect 537 -17 575 17
rect 609 -17 647 17
rect 681 -17 719 17
rect 753 -17 791 17
rect 825 -17 863 17
rect 897 -17 935 17
rect 969 -17 1007 17
rect 1041 -17 1079 17
rect 1113 -17 1151 17
rect 1185 -17 1223 17
rect 1257 -17 1295 17
rect 1329 -17 1367 17
rect 1401 -17 1439 17
rect 1473 -17 1511 17
rect 1545 -17 1583 17
rect 1617 -17 1655 17
rect 1689 -17 1727 17
rect 1761 -17 1799 17
rect 1833 -17 1871 17
rect 1905 -17 1943 17
rect 1977 -17 2015 17
rect 2049 -17 2087 17
rect 2121 -17 2159 17
rect 2193 -17 2231 17
rect 2265 -17 2303 17
rect 2337 -17 2375 17
rect 2409 -17 2447 17
rect 2481 -17 2519 17
rect 2553 -17 2591 17
rect 2625 -17 2663 17
rect 2697 -17 2735 17
rect 2769 -17 2807 17
rect 2841 -17 2879 17
rect 2913 -17 2951 17
rect 2985 -17 3023 17
rect 3057 -17 3095 17
rect 3129 -17 3167 17
rect 3201 -17 3239 17
rect 3273 -17 3311 17
rect 3345 -17 3481 17
rect 7 -23 3481 -17
<< via1 >>
rect 296 2720 348 2772
rect 296 2656 348 2708
rect 296 2592 348 2644
rect 296 2528 348 2580
rect 296 2464 348 2516
rect 296 2400 348 2452
rect 296 2336 348 2388
rect 296 2272 348 2324
rect 296 2208 348 2260
rect 296 2144 348 2196
rect 296 2080 348 2132
rect 296 2016 348 2068
rect 296 1952 348 2004
rect 296 1888 348 1940
rect 296 1824 348 1876
rect 612 2720 664 2772
rect 612 2656 664 2708
rect 612 2592 664 2644
rect 612 2528 664 2580
rect 612 2464 664 2516
rect 612 2400 664 2452
rect 612 2336 664 2388
rect 612 2272 664 2324
rect 612 2208 664 2260
rect 612 2144 664 2196
rect 612 2080 664 2132
rect 612 2016 664 2068
rect 612 1952 664 2004
rect 612 1888 664 1940
rect 612 1824 664 1876
rect 928 2720 980 2772
rect 928 2656 980 2708
rect 928 2592 980 2644
rect 928 2528 980 2580
rect 928 2464 980 2516
rect 928 2400 980 2452
rect 928 2336 980 2388
rect 928 2272 980 2324
rect 928 2208 980 2260
rect 928 2144 980 2196
rect 928 2080 980 2132
rect 928 2016 980 2068
rect 928 1952 980 2004
rect 928 1888 980 1940
rect 928 1824 980 1876
rect 1244 2720 1296 2772
rect 1244 2656 1296 2708
rect 1244 2592 1296 2644
rect 1244 2528 1296 2580
rect 1244 2464 1296 2516
rect 1244 2400 1296 2452
rect 1244 2336 1296 2388
rect 1244 2272 1296 2324
rect 1244 2208 1296 2260
rect 1244 2144 1296 2196
rect 1244 2080 1296 2132
rect 1244 2016 1296 2068
rect 1244 1952 1296 2004
rect 1244 1888 1296 1940
rect 1244 1824 1296 1876
rect 1560 2720 1612 2772
rect 1560 2656 1612 2708
rect 1560 2592 1612 2644
rect 1560 2528 1612 2580
rect 1560 2464 1612 2516
rect 1560 2400 1612 2452
rect 1560 2336 1612 2388
rect 1560 2272 1612 2324
rect 1560 2208 1612 2260
rect 1560 2144 1612 2196
rect 1560 2080 1612 2132
rect 1560 2016 1612 2068
rect 1560 1952 1612 2004
rect 1560 1888 1612 1940
rect 1560 1824 1612 1876
rect 1876 2720 1928 2772
rect 1876 2656 1928 2708
rect 1876 2592 1928 2644
rect 1876 2528 1928 2580
rect 1876 2464 1928 2516
rect 1876 2400 1928 2452
rect 1876 2336 1928 2388
rect 1876 2272 1928 2324
rect 1876 2208 1928 2260
rect 1876 2144 1928 2196
rect 1876 2080 1928 2132
rect 1876 2016 1928 2068
rect 1876 1952 1928 2004
rect 1876 1888 1928 1940
rect 1876 1824 1928 1876
rect 2192 2720 2244 2772
rect 2192 2656 2244 2708
rect 2192 2592 2244 2644
rect 2192 2528 2244 2580
rect 2192 2464 2244 2516
rect 2192 2400 2244 2452
rect 2192 2336 2244 2388
rect 2192 2272 2244 2324
rect 2192 2208 2244 2260
rect 2192 2144 2244 2196
rect 2192 2080 2244 2132
rect 2192 2016 2244 2068
rect 2192 1952 2244 2004
rect 2192 1888 2244 1940
rect 2192 1824 2244 1876
rect 2508 2720 2560 2772
rect 2508 2656 2560 2708
rect 2508 2592 2560 2644
rect 2508 2528 2560 2580
rect 2508 2464 2560 2516
rect 2508 2400 2560 2452
rect 2508 2336 2560 2388
rect 2508 2272 2560 2324
rect 2508 2208 2560 2260
rect 2508 2144 2560 2196
rect 2508 2080 2560 2132
rect 2508 2016 2560 2068
rect 2508 1952 2560 2004
rect 2508 1888 2560 1940
rect 2508 1824 2560 1876
rect 2824 2720 2876 2772
rect 2824 2656 2876 2708
rect 2824 2592 2876 2644
rect 2824 2528 2876 2580
rect 2824 2464 2876 2516
rect 2824 2400 2876 2452
rect 2824 2336 2876 2388
rect 2824 2272 2876 2324
rect 2824 2208 2876 2260
rect 2824 2144 2876 2196
rect 2824 2080 2876 2132
rect 2824 2016 2876 2068
rect 2824 1952 2876 2004
rect 2824 1888 2876 1940
rect 2824 1824 2876 1876
rect 3140 2720 3192 2772
rect 3140 2656 3192 2708
rect 3140 2592 3192 2644
rect 3140 2528 3192 2580
rect 3140 2464 3192 2516
rect 3140 2400 3192 2452
rect 3140 2336 3192 2388
rect 3140 2272 3192 2324
rect 3140 2208 3192 2260
rect 3140 2144 3192 2196
rect 3140 2080 3192 2132
rect 3140 2016 3192 2068
rect 3140 1952 3192 2004
rect 3140 1888 3192 1940
rect 3140 1824 3192 1876
rect 296 1466 348 1518
rect 612 1466 664 1518
rect 928 1466 980 1518
rect 1244 1466 1296 1518
rect 1560 1466 1612 1518
rect 1876 1466 1928 1518
rect 2192 1466 2244 1518
rect 2508 1466 2560 1518
rect 2824 1466 2876 1518
rect 3140 1466 3192 1518
rect 296 1115 348 1167
rect 296 1051 348 1103
rect 296 987 348 1039
rect 296 923 348 975
rect 296 859 348 911
rect 296 795 348 847
rect 296 731 348 783
rect 296 667 348 719
rect 296 603 348 655
rect 296 539 348 591
rect 296 475 348 527
rect 296 411 348 463
rect 296 347 348 399
rect 296 283 348 335
rect 296 219 348 271
rect 612 1115 664 1167
rect 612 1051 664 1103
rect 612 987 664 1039
rect 612 923 664 975
rect 612 859 664 911
rect 612 795 664 847
rect 612 731 664 783
rect 612 667 664 719
rect 612 603 664 655
rect 612 539 664 591
rect 612 475 664 527
rect 612 411 664 463
rect 612 347 664 399
rect 612 283 664 335
rect 612 219 664 271
rect 928 1115 980 1167
rect 928 1051 980 1103
rect 928 987 980 1039
rect 928 923 980 975
rect 928 859 980 911
rect 928 795 980 847
rect 928 731 980 783
rect 928 667 980 719
rect 928 603 980 655
rect 928 539 980 591
rect 928 475 980 527
rect 928 411 980 463
rect 928 347 980 399
rect 928 283 980 335
rect 928 219 980 271
rect 1244 1115 1296 1167
rect 1244 1051 1296 1103
rect 1244 987 1296 1039
rect 1244 923 1296 975
rect 1244 859 1296 911
rect 1244 795 1296 847
rect 1244 731 1296 783
rect 1244 667 1296 719
rect 1244 603 1296 655
rect 1244 539 1296 591
rect 1244 475 1296 527
rect 1244 411 1296 463
rect 1244 347 1296 399
rect 1244 283 1296 335
rect 1244 219 1296 271
rect 1560 1115 1612 1167
rect 1560 1051 1612 1103
rect 1560 987 1612 1039
rect 1560 923 1612 975
rect 1560 859 1612 911
rect 1560 795 1612 847
rect 1560 731 1612 783
rect 1560 667 1612 719
rect 1560 603 1612 655
rect 1560 539 1612 591
rect 1560 475 1612 527
rect 1560 411 1612 463
rect 1560 347 1612 399
rect 1560 283 1612 335
rect 1560 219 1612 271
rect 1876 1115 1928 1167
rect 1876 1051 1928 1103
rect 1876 987 1928 1039
rect 1876 923 1928 975
rect 1876 859 1928 911
rect 1876 795 1928 847
rect 1876 731 1928 783
rect 1876 667 1928 719
rect 1876 603 1928 655
rect 1876 539 1928 591
rect 1876 475 1928 527
rect 1876 411 1928 463
rect 1876 347 1928 399
rect 1876 283 1928 335
rect 1876 219 1928 271
rect 2192 1115 2244 1167
rect 2192 1051 2244 1103
rect 2192 987 2244 1039
rect 2192 923 2244 975
rect 2192 859 2244 911
rect 2192 795 2244 847
rect 2192 731 2244 783
rect 2192 667 2244 719
rect 2192 603 2244 655
rect 2192 539 2244 591
rect 2192 475 2244 527
rect 2192 411 2244 463
rect 2192 347 2244 399
rect 2192 283 2244 335
rect 2192 219 2244 271
rect 2508 1115 2560 1167
rect 2508 1051 2560 1103
rect 2508 987 2560 1039
rect 2508 923 2560 975
rect 2508 859 2560 911
rect 2508 795 2560 847
rect 2508 731 2560 783
rect 2508 667 2560 719
rect 2508 603 2560 655
rect 2508 539 2560 591
rect 2508 475 2560 527
rect 2508 411 2560 463
rect 2508 347 2560 399
rect 2508 283 2560 335
rect 2508 219 2560 271
rect 2824 1115 2876 1167
rect 2824 1051 2876 1103
rect 2824 987 2876 1039
rect 2824 923 2876 975
rect 2824 859 2876 911
rect 2824 795 2876 847
rect 2824 731 2876 783
rect 2824 667 2876 719
rect 2824 603 2876 655
rect 2824 539 2876 591
rect 2824 475 2876 527
rect 2824 411 2876 463
rect 2824 347 2876 399
rect 2824 283 2876 335
rect 2824 219 2876 271
rect 3140 1115 3192 1167
rect 3140 1051 3192 1103
rect 3140 987 3192 1039
rect 3140 923 3192 975
rect 3140 859 3192 911
rect 3140 795 3192 847
rect 3140 731 3192 783
rect 3140 667 3192 719
rect 3140 603 3192 655
rect 3140 539 3192 591
rect 3140 475 3192 527
rect 3140 411 3192 463
rect 3140 347 3192 399
rect 3140 283 3192 335
rect 3140 219 3192 271
<< metal2 >>
rect 296 2772 348 2796
rect 296 2708 348 2720
rect 296 2644 348 2656
rect 296 2580 348 2592
rect 296 2516 348 2528
rect 296 2452 348 2464
rect 296 2388 348 2400
rect 296 2324 348 2336
rect 296 2260 348 2272
rect 296 2196 348 2208
rect 296 2132 348 2144
rect 296 2068 348 2080
rect 296 2004 348 2016
rect 296 1940 348 1952
rect 296 1876 348 1888
rect 296 1518 348 1824
rect 296 1167 348 1466
rect 296 1103 348 1115
rect 296 1039 348 1051
rect 296 975 348 987
rect 296 911 348 923
rect 296 847 348 859
rect 296 783 348 795
rect 296 719 348 731
rect 296 655 348 667
rect 296 591 348 603
rect 296 527 348 539
rect 296 463 348 475
rect 296 399 348 411
rect 296 335 348 347
rect 296 271 348 283
rect 296 195 348 219
rect 612 2772 664 2796
rect 612 2708 664 2720
rect 612 2644 664 2656
rect 612 2580 664 2592
rect 612 2516 664 2528
rect 612 2452 664 2464
rect 612 2388 664 2400
rect 612 2324 664 2336
rect 612 2260 664 2272
rect 612 2196 664 2208
rect 612 2132 664 2144
rect 612 2068 664 2080
rect 612 2004 664 2016
rect 612 1940 664 1952
rect 612 1876 664 1888
rect 612 1518 664 1824
rect 612 1167 664 1466
rect 612 1103 664 1115
rect 612 1039 664 1051
rect 612 975 664 987
rect 612 911 664 923
rect 612 847 664 859
rect 612 783 664 795
rect 612 719 664 731
rect 612 655 664 667
rect 612 591 664 603
rect 612 527 664 539
rect 612 463 664 475
rect 612 399 664 411
rect 612 335 664 347
rect 612 271 664 283
rect 612 195 664 219
rect 928 2772 980 2796
rect 928 2708 980 2720
rect 928 2644 980 2656
rect 928 2580 980 2592
rect 928 2516 980 2528
rect 928 2452 980 2464
rect 928 2388 980 2400
rect 928 2324 980 2336
rect 928 2260 980 2272
rect 928 2196 980 2208
rect 928 2132 980 2144
rect 928 2068 980 2080
rect 928 2004 980 2016
rect 928 1940 980 1952
rect 928 1876 980 1888
rect 928 1518 980 1824
rect 928 1167 980 1466
rect 928 1103 980 1115
rect 928 1039 980 1051
rect 928 975 980 987
rect 928 911 980 923
rect 928 847 980 859
rect 928 783 980 795
rect 928 719 980 731
rect 928 655 980 667
rect 928 591 980 603
rect 928 527 980 539
rect 928 463 980 475
rect 928 399 980 411
rect 928 335 980 347
rect 928 271 980 283
rect 928 195 980 219
rect 1244 2772 1296 2796
rect 1244 2708 1296 2720
rect 1244 2644 1296 2656
rect 1244 2580 1296 2592
rect 1244 2516 1296 2528
rect 1244 2452 1296 2464
rect 1244 2388 1296 2400
rect 1244 2324 1296 2336
rect 1244 2260 1296 2272
rect 1244 2196 1296 2208
rect 1244 2132 1296 2144
rect 1244 2068 1296 2080
rect 1244 2004 1296 2016
rect 1244 1940 1296 1952
rect 1244 1876 1296 1888
rect 1244 1518 1296 1824
rect 1244 1167 1296 1466
rect 1244 1103 1296 1115
rect 1244 1039 1296 1051
rect 1244 975 1296 987
rect 1244 911 1296 923
rect 1244 847 1296 859
rect 1244 783 1296 795
rect 1244 719 1296 731
rect 1244 655 1296 667
rect 1244 591 1296 603
rect 1244 527 1296 539
rect 1244 463 1296 475
rect 1244 399 1296 411
rect 1244 335 1296 347
rect 1244 271 1296 283
rect 1244 195 1296 219
rect 1560 2772 1612 2796
rect 1560 2708 1612 2720
rect 1560 2644 1612 2656
rect 1560 2580 1612 2592
rect 1560 2516 1612 2528
rect 1560 2452 1612 2464
rect 1560 2388 1612 2400
rect 1560 2324 1612 2336
rect 1560 2260 1612 2272
rect 1560 2196 1612 2208
rect 1560 2132 1612 2144
rect 1560 2068 1612 2080
rect 1560 2004 1612 2016
rect 1560 1940 1612 1952
rect 1560 1876 1612 1888
rect 1560 1518 1612 1824
rect 1560 1167 1612 1466
rect 1560 1103 1612 1115
rect 1560 1039 1612 1051
rect 1560 975 1612 987
rect 1560 911 1612 923
rect 1560 847 1612 859
rect 1560 783 1612 795
rect 1560 719 1612 731
rect 1560 655 1612 667
rect 1560 591 1612 603
rect 1560 527 1612 539
rect 1560 463 1612 475
rect 1560 399 1612 411
rect 1560 335 1612 347
rect 1560 271 1612 283
rect 1560 195 1612 219
rect 1876 2772 1928 2796
rect 1876 2708 1928 2720
rect 1876 2644 1928 2656
rect 1876 2580 1928 2592
rect 1876 2516 1928 2528
rect 1876 2452 1928 2464
rect 1876 2388 1928 2400
rect 1876 2324 1928 2336
rect 1876 2260 1928 2272
rect 1876 2196 1928 2208
rect 1876 2132 1928 2144
rect 1876 2068 1928 2080
rect 1876 2004 1928 2016
rect 1876 1940 1928 1952
rect 1876 1876 1928 1888
rect 1876 1518 1928 1824
rect 1876 1167 1928 1466
rect 1876 1103 1928 1115
rect 1876 1039 1928 1051
rect 1876 975 1928 987
rect 1876 911 1928 923
rect 1876 847 1928 859
rect 1876 783 1928 795
rect 1876 719 1928 731
rect 1876 655 1928 667
rect 1876 591 1928 603
rect 1876 527 1928 539
rect 1876 463 1928 475
rect 1876 399 1928 411
rect 1876 335 1928 347
rect 1876 271 1928 283
rect 1876 195 1928 219
rect 2192 2772 2244 2796
rect 2192 2708 2244 2720
rect 2192 2644 2244 2656
rect 2192 2580 2244 2592
rect 2192 2516 2244 2528
rect 2192 2452 2244 2464
rect 2192 2388 2244 2400
rect 2192 2324 2244 2336
rect 2192 2260 2244 2272
rect 2192 2196 2244 2208
rect 2192 2132 2244 2144
rect 2192 2068 2244 2080
rect 2192 2004 2244 2016
rect 2192 1940 2244 1952
rect 2192 1876 2244 1888
rect 2192 1518 2244 1824
rect 2192 1167 2244 1466
rect 2192 1103 2244 1115
rect 2192 1039 2244 1051
rect 2192 975 2244 987
rect 2192 911 2244 923
rect 2192 847 2244 859
rect 2192 783 2244 795
rect 2192 719 2244 731
rect 2192 655 2244 667
rect 2192 591 2244 603
rect 2192 527 2244 539
rect 2192 463 2244 475
rect 2192 399 2244 411
rect 2192 335 2244 347
rect 2192 271 2244 283
rect 2192 195 2244 219
rect 2508 2772 2560 2796
rect 2508 2708 2560 2720
rect 2508 2644 2560 2656
rect 2508 2580 2560 2592
rect 2508 2516 2560 2528
rect 2508 2452 2560 2464
rect 2508 2388 2560 2400
rect 2508 2324 2560 2336
rect 2508 2260 2560 2272
rect 2508 2196 2560 2208
rect 2508 2132 2560 2144
rect 2508 2068 2560 2080
rect 2508 2004 2560 2016
rect 2508 1940 2560 1952
rect 2508 1876 2560 1888
rect 2508 1518 2560 1824
rect 2508 1167 2560 1466
rect 2508 1103 2560 1115
rect 2508 1039 2560 1051
rect 2508 975 2560 987
rect 2508 911 2560 923
rect 2508 847 2560 859
rect 2508 783 2560 795
rect 2508 719 2560 731
rect 2508 655 2560 667
rect 2508 591 2560 603
rect 2508 527 2560 539
rect 2508 463 2560 475
rect 2508 399 2560 411
rect 2508 335 2560 347
rect 2508 271 2560 283
rect 2508 195 2560 219
rect 2824 2772 2876 2796
rect 2824 2708 2876 2720
rect 2824 2644 2876 2656
rect 2824 2580 2876 2592
rect 2824 2516 2876 2528
rect 2824 2452 2876 2464
rect 2824 2388 2876 2400
rect 2824 2324 2876 2336
rect 2824 2260 2876 2272
rect 2824 2196 2876 2208
rect 2824 2132 2876 2144
rect 2824 2068 2876 2080
rect 2824 2004 2876 2016
rect 2824 1940 2876 1952
rect 2824 1876 2876 1888
rect 2824 1518 2876 1824
rect 2824 1167 2876 1466
rect 2824 1103 2876 1115
rect 2824 1039 2876 1051
rect 2824 975 2876 987
rect 2824 911 2876 923
rect 2824 847 2876 859
rect 2824 783 2876 795
rect 2824 719 2876 731
rect 2824 655 2876 667
rect 2824 591 2876 603
rect 2824 527 2876 539
rect 2824 463 2876 475
rect 2824 399 2876 411
rect 2824 335 2876 347
rect 2824 271 2876 283
rect 2824 195 2876 219
rect 3140 2772 3192 2796
rect 3140 2708 3192 2720
rect 3140 2644 3192 2656
rect 3140 2580 3192 2592
rect 3140 2516 3192 2528
rect 3140 2452 3192 2464
rect 3140 2388 3192 2400
rect 3140 2324 3192 2336
rect 3140 2260 3192 2272
rect 3140 2196 3192 2208
rect 3140 2132 3192 2144
rect 3140 2068 3192 2080
rect 3140 2004 3192 2016
rect 3140 1940 3192 1952
rect 3140 1876 3192 1888
rect 3140 1518 3192 1824
rect 3140 1167 3192 1466
rect 3140 1103 3192 1115
rect 3140 1039 3192 1051
rect 3140 975 3192 987
rect 3140 911 3192 923
rect 3140 847 3192 859
rect 3140 783 3192 795
rect 3140 719 3192 731
rect 3140 655 3192 667
rect 3140 591 3192 603
rect 3140 527 3192 539
rect 3140 463 3192 475
rect 3140 399 3192 411
rect 3140 335 3192 347
rect 3140 271 3192 283
rect 3140 195 3192 219
use sky130_fd_pr__nfet_g5v0d10v5_BRTJC6  sky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0
timestamp 1654583101
transform 1 0 1744 0 1 693
box -1769 -748 1769 748
use sky130_fd_pr__pfet_g5v0d10v5_CADZ46  sky130_fd_pr__pfet_g5v0d10v5_CADZ46_0
timestamp 1654583101
transform 1 0 1744 0 1 2298
box -1809 -797 1809 797
<< labels >>
flabel metal1 s -54 1487 -54 1487 1 FreeSans 500 0 0 0 esd
port 1 nsew
flabel metal1 s 30 2927 30 2927 1 FreeSans 500 0 0 0 VDD
port 2 nsew
flabel metal1 s 30 71 30 71 1 FreeSans 500 0 0 0 VSS
port 3 nsew
<< end >>
