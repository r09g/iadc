magic
tech sky130A
magscale 1 2
timestamp 1654727055
<< nwell >>
rect -3266 -716 -1972 -66
rect -1018 -1059 -298 -738
rect -742 -1304 -298 -1059
rect 285 -1180 3100 -530
rect -3266 -2050 -1972 -1400
rect -742 -2071 -298 -1826
rect -1294 -2392 -298 -2071
rect 285 -2514 3100 -1864
rect -3266 -3428 -1972 -2778
rect -1294 -3235 -298 -2914
rect -742 -3480 -298 -3235
rect 285 -3892 3100 -3242
rect -3266 -4806 -1972 -4156
rect -742 -4568 -298 -4002
rect 285 -5270 3100 -4620
<< pwell >>
rect 1553 -68 1809 -66
rect -951 -494 -917 -460
rect -583 -494 -549 -460
rect -938 -498 -917 -494
rect -570 -498 -549 -494
rect -938 -515 -635 -498
rect -938 -525 -615 -515
rect -570 -525 -384 -498
rect -938 -680 -384 -525
rect 285 -530 3100 -68
rect -3266 -1178 -1972 -716
rect -701 -1586 -384 -1362
rect 1553 -1402 1809 -1400
rect -701 -1768 -337 -1586
rect -3266 -2512 -1972 -2050
rect 285 -1864 3100 -1402
rect -1253 -2615 -337 -2450
rect -1241 -2632 -337 -2615
rect -1122 -2636 -1101 -2632
rect -1135 -2670 -1101 -2636
rect -857 -2663 -825 -2641
rect -767 -2665 -735 -2643
rect -1122 -2674 -1101 -2670
rect -584 -2674 -550 -2632
rect -1253 -2701 -1167 -2691
rect -1122 -2701 -936 -2674
rect -701 -2701 -615 -2691
rect -607 -2701 -337 -2674
rect -1253 -2856 -337 -2701
rect 1553 -2780 1809 -2778
rect -3266 -3890 -1972 -3428
rect 285 -3242 3100 -2780
rect -701 -3693 -337 -3538
rect -701 -3703 -615 -3693
rect -607 -3720 -337 -3693
rect -584 -3724 -550 -3720
rect -584 -3758 -549 -3724
rect -570 -3762 -549 -3758
rect -701 -3789 -615 -3779
rect -570 -3789 -384 -3762
rect -702 -3944 -338 -3789
rect 1553 -4158 1809 -4156
rect 285 -4620 3100 -4158
rect -701 -4781 -337 -4626
rect -701 -4791 -615 -4781
rect -3266 -5268 -1972 -4806
rect -570 -4808 -384 -4781
rect -570 -4812 -549 -4808
rect -583 -4846 -549 -4812
<< nmos >>
rect 485 -382 515 -278
rect 581 -382 611 -278
rect 677 -382 707 -278
rect 773 -382 803 -278
rect 869 -382 899 -278
rect 965 -382 995 -278
rect 1061 -382 1091 -278
rect 1157 -382 1187 -278
rect 1253 -382 1283 -278
rect 1349 -382 1379 -278
rect 1661 -384 1691 -284
rect 2006 -382 2036 -278
rect 2102 -382 2132 -278
rect 2198 -382 2228 -278
rect 2294 -382 2324 -278
rect 2390 -382 2420 -278
rect 2486 -382 2516 -278
rect 2582 -382 2612 -278
rect 2678 -382 2708 -278
rect 2774 -382 2804 -278
rect 2870 -382 2900 -278
rect -3066 -968 -3036 -864
rect -2970 -968 -2940 -864
rect -2874 -968 -2844 -864
rect -2778 -968 -2748 -864
rect -2682 -968 -2652 -864
rect -2586 -968 -2556 -864
rect -2490 -968 -2460 -864
rect -2394 -968 -2364 -864
rect -2298 -968 -2268 -864
rect -2202 -968 -2172 -864
rect 485 -1716 515 -1612
rect 581 -1716 611 -1612
rect 677 -1716 707 -1612
rect 773 -1716 803 -1612
rect 869 -1716 899 -1612
rect 965 -1716 995 -1612
rect 1061 -1716 1091 -1612
rect 1157 -1716 1187 -1612
rect 1253 -1716 1283 -1612
rect 1349 -1716 1379 -1612
rect 1661 -1718 1691 -1618
rect 2006 -1716 2036 -1612
rect 2102 -1716 2132 -1612
rect 2198 -1716 2228 -1612
rect 2294 -1716 2324 -1612
rect 2390 -1716 2420 -1612
rect 2486 -1716 2516 -1612
rect 2582 -1716 2612 -1612
rect 2678 -1716 2708 -1612
rect 2774 -1716 2804 -1612
rect 2870 -1716 2900 -1612
rect -3066 -2302 -3036 -2198
rect -2970 -2302 -2940 -2198
rect -2874 -2302 -2844 -2198
rect -2778 -2302 -2748 -2198
rect -2682 -2302 -2652 -2198
rect -2586 -2302 -2556 -2198
rect -2490 -2302 -2460 -2198
rect -2394 -2302 -2364 -2198
rect -2298 -2302 -2268 -2198
rect -2202 -2302 -2172 -2198
rect 485 -3094 515 -2990
rect 581 -3094 611 -2990
rect 677 -3094 707 -2990
rect 773 -3094 803 -2990
rect 869 -3094 899 -2990
rect 965 -3094 995 -2990
rect 1061 -3094 1091 -2990
rect 1157 -3094 1187 -2990
rect 1253 -3094 1283 -2990
rect 1349 -3094 1379 -2990
rect 1661 -3096 1691 -2996
rect 2006 -3094 2036 -2990
rect 2102 -3094 2132 -2990
rect 2198 -3094 2228 -2990
rect 2294 -3094 2324 -2990
rect 2390 -3094 2420 -2990
rect 2486 -3094 2516 -2990
rect 2582 -3094 2612 -2990
rect 2678 -3094 2708 -2990
rect 2774 -3094 2804 -2990
rect 2870 -3094 2900 -2990
rect -3066 -3680 -3036 -3576
rect -2970 -3680 -2940 -3576
rect -2874 -3680 -2844 -3576
rect -2778 -3680 -2748 -3576
rect -2682 -3680 -2652 -3576
rect -2586 -3680 -2556 -3576
rect -2490 -3680 -2460 -3576
rect -2394 -3680 -2364 -3576
rect -2298 -3680 -2268 -3576
rect -2202 -3680 -2172 -3576
rect 485 -4472 515 -4368
rect 581 -4472 611 -4368
rect 677 -4472 707 -4368
rect 773 -4472 803 -4368
rect 869 -4472 899 -4368
rect 965 -4472 995 -4368
rect 1061 -4472 1091 -4368
rect 1157 -4472 1187 -4368
rect 1253 -4472 1283 -4368
rect 1349 -4472 1379 -4368
rect 1661 -4474 1691 -4374
rect 2006 -4472 2036 -4368
rect 2102 -4472 2132 -4368
rect 2198 -4472 2228 -4368
rect 2294 -4472 2324 -4368
rect 2390 -4472 2420 -4368
rect 2486 -4472 2516 -4368
rect 2582 -4472 2612 -4368
rect 2678 -4472 2708 -4368
rect 2774 -4472 2804 -4368
rect 2870 -4472 2900 -4368
rect -3066 -5058 -3036 -4954
rect -2970 -5058 -2940 -4954
rect -2874 -5058 -2844 -4954
rect -2778 -5058 -2748 -4954
rect -2682 -5058 -2652 -4954
rect -2586 -5058 -2556 -4954
rect -2490 -5058 -2460 -4954
rect -2394 -5058 -2364 -4954
rect -2298 -5058 -2268 -4954
rect -2202 -5058 -2172 -4954
<< scnmos >>
rect -860 -654 -830 -524
rect -492 -654 -462 -524
rect -492 -1518 -462 -1388
rect -529 -1742 -499 -1612
rect -445 -1742 -415 -1612
rect -1044 -2606 -1014 -2476
rect -529 -2606 -499 -2476
rect -445 -2606 -415 -2476
rect -1044 -2830 -1014 -2700
rect -529 -2830 -499 -2700
rect -445 -2830 -415 -2700
rect -529 -3694 -499 -3564
rect -445 -3694 -415 -3564
rect -492 -3918 -462 -3788
rect -492 -4782 -462 -4652
<< pmos >>
rect -3066 -558 -3036 -286
rect -2970 -558 -2940 -286
rect -2874 -558 -2844 -286
rect -2778 -558 -2748 -286
rect -2682 -558 -2652 -286
rect -2586 -558 -2556 -286
rect -2490 -558 -2460 -286
rect -2394 -558 -2364 -286
rect -2298 -558 -2268 -286
rect -2202 -558 -2172 -286
rect 485 -960 515 -688
rect 581 -960 611 -688
rect 677 -960 707 -688
rect 773 -960 803 -688
rect 869 -960 899 -688
rect 965 -960 995 -688
rect 1061 -960 1091 -688
rect 1157 -960 1187 -688
rect 1253 -960 1283 -688
rect 1349 -960 1379 -688
rect 2006 -960 2036 -688
rect 2102 -960 2132 -688
rect 2198 -960 2228 -688
rect 2294 -960 2324 -688
rect 2390 -960 2420 -688
rect 2486 -960 2516 -688
rect 2582 -960 2612 -688
rect 2678 -960 2708 -688
rect 2774 -960 2804 -688
rect 2870 -960 2900 -688
rect -3066 -1892 -3036 -1620
rect -2970 -1892 -2940 -1620
rect -2874 -1892 -2844 -1620
rect -2778 -1892 -2748 -1620
rect -2682 -1892 -2652 -1620
rect -2586 -1892 -2556 -1620
rect -2490 -1892 -2460 -1620
rect -2394 -1892 -2364 -1620
rect -2298 -1892 -2268 -1620
rect -2202 -1892 -2172 -1620
rect 485 -2294 515 -2022
rect 581 -2294 611 -2022
rect 677 -2294 707 -2022
rect 773 -2294 803 -2022
rect 869 -2294 899 -2022
rect 965 -2294 995 -2022
rect 1061 -2294 1091 -2022
rect 1157 -2294 1187 -2022
rect 1253 -2294 1283 -2022
rect 1349 -2294 1379 -2022
rect 2006 -2294 2036 -2022
rect 2102 -2294 2132 -2022
rect 2198 -2294 2228 -2022
rect 2294 -2294 2324 -2022
rect 2390 -2294 2420 -2022
rect 2486 -2294 2516 -2022
rect 2582 -2294 2612 -2022
rect 2678 -2294 2708 -2022
rect 2774 -2294 2804 -2022
rect 2870 -2294 2900 -2022
rect -3066 -3270 -3036 -2998
rect -2970 -3270 -2940 -2998
rect -2874 -3270 -2844 -2998
rect -2778 -3270 -2748 -2998
rect -2682 -3270 -2652 -2998
rect -2586 -3270 -2556 -2998
rect -2490 -3270 -2460 -2998
rect -2394 -3270 -2364 -2998
rect -2298 -3270 -2268 -2998
rect -2202 -3270 -2172 -2998
rect 485 -3672 515 -3400
rect 581 -3672 611 -3400
rect 677 -3672 707 -3400
rect 773 -3672 803 -3400
rect 869 -3672 899 -3400
rect 965 -3672 995 -3400
rect 1061 -3672 1091 -3400
rect 1157 -3672 1187 -3400
rect 1253 -3672 1283 -3400
rect 1349 -3672 1379 -3400
rect 2006 -3672 2036 -3400
rect 2102 -3672 2132 -3400
rect 2198 -3672 2228 -3400
rect 2294 -3672 2324 -3400
rect 2390 -3672 2420 -3400
rect 2486 -3672 2516 -3400
rect 2582 -3672 2612 -3400
rect 2678 -3672 2708 -3400
rect 2774 -3672 2804 -3400
rect 2870 -3672 2900 -3400
rect -3066 -4648 -3036 -4376
rect -2970 -4648 -2940 -4376
rect -2874 -4648 -2844 -4376
rect -2778 -4648 -2748 -4376
rect -2682 -4648 -2652 -4376
rect -2586 -4648 -2556 -4376
rect -2490 -4648 -2460 -4376
rect -2394 -4648 -2364 -4376
rect -2298 -4648 -2268 -4376
rect -2202 -4648 -2172 -4376
rect 485 -5050 515 -4778
rect 581 -5050 611 -4778
rect 677 -5050 707 -4778
rect 773 -5050 803 -4778
rect 869 -5050 899 -4778
rect 965 -5050 995 -4778
rect 1061 -5050 1091 -4778
rect 1157 -5050 1187 -4778
rect 1253 -5050 1283 -4778
rect 1349 -5050 1379 -4778
rect 2006 -5050 2036 -4778
rect 2102 -5050 2132 -4778
rect 2198 -5050 2228 -4778
rect 2294 -5050 2324 -4778
rect 2390 -5050 2420 -4778
rect 2486 -5050 2516 -4778
rect 2582 -5050 2612 -4778
rect 2678 -5050 2708 -4778
rect 2774 -5050 2804 -4778
rect 2870 -5050 2900 -4778
<< scpmoshvt >>
rect -860 -974 -830 -774
rect -492 -974 -462 -774
rect -492 -1268 -462 -1068
rect -529 -2062 -499 -1862
rect -445 -2062 -415 -1862
rect -1044 -2356 -1014 -2156
rect -529 -2356 -499 -2156
rect -445 -2356 -415 -2156
rect -1044 -3150 -1014 -2950
rect -529 -3150 -499 -2950
rect -445 -3150 -415 -2950
rect -529 -3444 -499 -3244
rect -445 -3444 -415 -3244
rect -492 -4238 -462 -4038
rect -492 -4532 -462 -4332
<< ndiff >>
rect 423 -290 485 -278
rect 423 -370 435 -290
rect 469 -370 485 -290
rect 423 -382 485 -370
rect 515 -290 581 -278
rect 515 -370 531 -290
rect 565 -370 581 -290
rect 515 -382 581 -370
rect 611 -290 677 -278
rect 611 -370 627 -290
rect 661 -370 677 -290
rect 611 -382 677 -370
rect 707 -290 773 -278
rect 707 -370 723 -290
rect 757 -370 773 -290
rect 707 -382 773 -370
rect 803 -290 869 -278
rect 803 -370 819 -290
rect 853 -370 869 -290
rect 803 -382 869 -370
rect 899 -290 965 -278
rect 899 -370 915 -290
rect 949 -370 965 -290
rect 899 -382 965 -370
rect 995 -290 1061 -278
rect 995 -370 1011 -290
rect 1045 -370 1061 -290
rect 995 -382 1061 -370
rect 1091 -290 1157 -278
rect 1091 -370 1107 -290
rect 1141 -370 1157 -290
rect 1091 -382 1157 -370
rect 1187 -290 1253 -278
rect 1187 -370 1203 -290
rect 1237 -370 1253 -290
rect 1187 -382 1253 -370
rect 1283 -290 1349 -278
rect 1283 -370 1299 -290
rect 1333 -370 1349 -290
rect 1283 -382 1349 -370
rect 1379 -290 1441 -278
rect 1379 -370 1395 -290
rect 1429 -370 1441 -290
rect 1379 -382 1441 -370
rect 1603 -296 1661 -284
rect 1603 -372 1615 -296
rect 1649 -372 1661 -296
rect 1603 -384 1661 -372
rect 1691 -296 1749 -284
rect 1691 -372 1703 -296
rect 1737 -372 1749 -296
rect 1691 -384 1749 -372
rect 1944 -290 2006 -278
rect 1944 -370 1956 -290
rect 1990 -370 2006 -290
rect 1944 -382 2006 -370
rect 2036 -290 2102 -278
rect 2036 -370 2052 -290
rect 2086 -370 2102 -290
rect 2036 -382 2102 -370
rect 2132 -290 2198 -278
rect 2132 -370 2148 -290
rect 2182 -370 2198 -290
rect 2132 -382 2198 -370
rect 2228 -290 2294 -278
rect 2228 -370 2244 -290
rect 2278 -370 2294 -290
rect 2228 -382 2294 -370
rect 2324 -290 2390 -278
rect 2324 -370 2340 -290
rect 2374 -370 2390 -290
rect 2324 -382 2390 -370
rect 2420 -290 2486 -278
rect 2420 -370 2436 -290
rect 2470 -370 2486 -290
rect 2420 -382 2486 -370
rect 2516 -290 2582 -278
rect 2516 -370 2532 -290
rect 2566 -370 2582 -290
rect 2516 -382 2582 -370
rect 2612 -290 2678 -278
rect 2612 -370 2628 -290
rect 2662 -370 2678 -290
rect 2612 -382 2678 -370
rect 2708 -290 2774 -278
rect 2708 -370 2724 -290
rect 2758 -370 2774 -290
rect 2708 -382 2774 -370
rect 2804 -290 2870 -278
rect 2804 -370 2820 -290
rect 2854 -370 2870 -290
rect 2804 -382 2870 -370
rect 2900 -290 2962 -278
rect 2900 -370 2916 -290
rect 2950 -370 2962 -290
rect 2900 -382 2962 -370
rect -912 -540 -860 -524
rect -912 -574 -904 -540
rect -870 -574 -860 -540
rect -912 -608 -860 -574
rect -912 -642 -904 -608
rect -870 -642 -860 -608
rect -912 -654 -860 -642
rect -830 -540 -778 -524
rect -830 -574 -820 -540
rect -786 -574 -778 -540
rect -544 -540 -492 -524
rect -830 -608 -778 -574
rect -830 -642 -820 -608
rect -786 -642 -778 -608
rect -830 -654 -778 -642
rect -544 -574 -536 -540
rect -502 -574 -492 -540
rect -544 -608 -492 -574
rect -544 -642 -536 -608
rect -502 -642 -492 -608
rect -544 -654 -492 -642
rect -462 -540 -410 -524
rect -462 -574 -452 -540
rect -418 -574 -410 -540
rect -462 -608 -410 -574
rect -462 -642 -452 -608
rect -418 -642 -410 -608
rect -462 -654 -410 -642
rect -3128 -876 -3066 -864
rect -3128 -956 -3116 -876
rect -3082 -956 -3066 -876
rect -3128 -968 -3066 -956
rect -3036 -876 -2970 -864
rect -3036 -956 -3020 -876
rect -2986 -956 -2970 -876
rect -3036 -968 -2970 -956
rect -2940 -876 -2874 -864
rect -2940 -956 -2924 -876
rect -2890 -956 -2874 -876
rect -2940 -968 -2874 -956
rect -2844 -876 -2778 -864
rect -2844 -956 -2828 -876
rect -2794 -956 -2778 -876
rect -2844 -968 -2778 -956
rect -2748 -876 -2682 -864
rect -2748 -956 -2732 -876
rect -2698 -956 -2682 -876
rect -2748 -968 -2682 -956
rect -2652 -876 -2586 -864
rect -2652 -956 -2636 -876
rect -2602 -956 -2586 -876
rect -2652 -968 -2586 -956
rect -2556 -876 -2490 -864
rect -2556 -956 -2540 -876
rect -2506 -956 -2490 -876
rect -2556 -968 -2490 -956
rect -2460 -876 -2394 -864
rect -2460 -956 -2444 -876
rect -2410 -956 -2394 -876
rect -2460 -968 -2394 -956
rect -2364 -876 -2298 -864
rect -2364 -956 -2348 -876
rect -2314 -956 -2298 -876
rect -2364 -968 -2298 -956
rect -2268 -876 -2202 -864
rect -2268 -956 -2252 -876
rect -2218 -956 -2202 -876
rect -2268 -968 -2202 -956
rect -2172 -876 -2110 -864
rect -2172 -956 -2156 -876
rect -2122 -956 -2110 -876
rect -2172 -968 -2110 -956
rect -544 -1400 -492 -1388
rect -544 -1434 -536 -1400
rect -502 -1434 -492 -1400
rect -544 -1468 -492 -1434
rect -544 -1502 -536 -1468
rect -502 -1502 -492 -1468
rect -544 -1518 -492 -1502
rect -462 -1400 -410 -1388
rect -462 -1434 -452 -1400
rect -418 -1434 -410 -1400
rect -462 -1468 -410 -1434
rect -462 -1502 -452 -1468
rect -418 -1502 -410 -1468
rect -462 -1518 -410 -1502
rect -581 -1624 -529 -1612
rect -581 -1658 -573 -1624
rect -539 -1658 -529 -1624
rect -581 -1692 -529 -1658
rect -581 -1726 -573 -1692
rect -539 -1726 -529 -1692
rect -581 -1742 -529 -1726
rect -499 -1742 -445 -1612
rect -415 -1624 -363 -1612
rect -415 -1658 -405 -1624
rect -371 -1658 -363 -1624
rect -415 -1692 -363 -1658
rect -415 -1726 -405 -1692
rect -371 -1726 -363 -1692
rect -415 -1742 -363 -1726
rect 423 -1624 485 -1612
rect 423 -1704 435 -1624
rect 469 -1704 485 -1624
rect 423 -1716 485 -1704
rect 515 -1624 581 -1612
rect 515 -1704 531 -1624
rect 565 -1704 581 -1624
rect 515 -1716 581 -1704
rect 611 -1624 677 -1612
rect 611 -1704 627 -1624
rect 661 -1704 677 -1624
rect 611 -1716 677 -1704
rect 707 -1624 773 -1612
rect 707 -1704 723 -1624
rect 757 -1704 773 -1624
rect 707 -1716 773 -1704
rect 803 -1624 869 -1612
rect 803 -1704 819 -1624
rect 853 -1704 869 -1624
rect 803 -1716 869 -1704
rect 899 -1624 965 -1612
rect 899 -1704 915 -1624
rect 949 -1704 965 -1624
rect 899 -1716 965 -1704
rect 995 -1624 1061 -1612
rect 995 -1704 1011 -1624
rect 1045 -1704 1061 -1624
rect 995 -1716 1061 -1704
rect 1091 -1624 1157 -1612
rect 1091 -1704 1107 -1624
rect 1141 -1704 1157 -1624
rect 1091 -1716 1157 -1704
rect 1187 -1624 1253 -1612
rect 1187 -1704 1203 -1624
rect 1237 -1704 1253 -1624
rect 1187 -1716 1253 -1704
rect 1283 -1624 1349 -1612
rect 1283 -1704 1299 -1624
rect 1333 -1704 1349 -1624
rect 1283 -1716 1349 -1704
rect 1379 -1624 1441 -1612
rect 1379 -1704 1395 -1624
rect 1429 -1704 1441 -1624
rect 1379 -1716 1441 -1704
rect 1603 -1630 1661 -1618
rect 1603 -1706 1615 -1630
rect 1649 -1706 1661 -1630
rect 1603 -1718 1661 -1706
rect 1691 -1630 1749 -1618
rect 1691 -1706 1703 -1630
rect 1737 -1706 1749 -1630
rect 1691 -1718 1749 -1706
rect 1944 -1624 2006 -1612
rect 1944 -1704 1956 -1624
rect 1990 -1704 2006 -1624
rect 1944 -1716 2006 -1704
rect 2036 -1624 2102 -1612
rect 2036 -1704 2052 -1624
rect 2086 -1704 2102 -1624
rect 2036 -1716 2102 -1704
rect 2132 -1624 2198 -1612
rect 2132 -1704 2148 -1624
rect 2182 -1704 2198 -1624
rect 2132 -1716 2198 -1704
rect 2228 -1624 2294 -1612
rect 2228 -1704 2244 -1624
rect 2278 -1704 2294 -1624
rect 2228 -1716 2294 -1704
rect 2324 -1624 2390 -1612
rect 2324 -1704 2340 -1624
rect 2374 -1704 2390 -1624
rect 2324 -1716 2390 -1704
rect 2420 -1624 2486 -1612
rect 2420 -1704 2436 -1624
rect 2470 -1704 2486 -1624
rect 2420 -1716 2486 -1704
rect 2516 -1624 2582 -1612
rect 2516 -1704 2532 -1624
rect 2566 -1704 2582 -1624
rect 2516 -1716 2582 -1704
rect 2612 -1624 2678 -1612
rect 2612 -1704 2628 -1624
rect 2662 -1704 2678 -1624
rect 2612 -1716 2678 -1704
rect 2708 -1624 2774 -1612
rect 2708 -1704 2724 -1624
rect 2758 -1704 2774 -1624
rect 2708 -1716 2774 -1704
rect 2804 -1624 2870 -1612
rect 2804 -1704 2820 -1624
rect 2854 -1704 2870 -1624
rect 2804 -1716 2870 -1704
rect 2900 -1624 2962 -1612
rect 2900 -1704 2916 -1624
rect 2950 -1704 2962 -1624
rect 2900 -1716 2962 -1704
rect -3128 -2210 -3066 -2198
rect -3128 -2290 -3116 -2210
rect -3082 -2290 -3066 -2210
rect -3128 -2302 -3066 -2290
rect -3036 -2210 -2970 -2198
rect -3036 -2290 -3020 -2210
rect -2986 -2290 -2970 -2210
rect -3036 -2302 -2970 -2290
rect -2940 -2210 -2874 -2198
rect -2940 -2290 -2924 -2210
rect -2890 -2290 -2874 -2210
rect -2940 -2302 -2874 -2290
rect -2844 -2210 -2778 -2198
rect -2844 -2290 -2828 -2210
rect -2794 -2290 -2778 -2210
rect -2844 -2302 -2778 -2290
rect -2748 -2210 -2682 -2198
rect -2748 -2290 -2732 -2210
rect -2698 -2290 -2682 -2210
rect -2748 -2302 -2682 -2290
rect -2652 -2210 -2586 -2198
rect -2652 -2290 -2636 -2210
rect -2602 -2290 -2586 -2210
rect -2652 -2302 -2586 -2290
rect -2556 -2210 -2490 -2198
rect -2556 -2290 -2540 -2210
rect -2506 -2290 -2490 -2210
rect -2556 -2302 -2490 -2290
rect -2460 -2210 -2394 -2198
rect -2460 -2290 -2444 -2210
rect -2410 -2290 -2394 -2210
rect -2460 -2302 -2394 -2290
rect -2364 -2210 -2298 -2198
rect -2364 -2290 -2348 -2210
rect -2314 -2290 -2298 -2210
rect -2364 -2302 -2298 -2290
rect -2268 -2210 -2202 -2198
rect -2268 -2290 -2252 -2210
rect -2218 -2290 -2202 -2210
rect -2268 -2302 -2202 -2290
rect -2172 -2210 -2110 -2198
rect -2172 -2290 -2156 -2210
rect -2122 -2290 -2110 -2210
rect -2172 -2302 -2110 -2290
rect -1096 -2488 -1044 -2476
rect -1096 -2522 -1088 -2488
rect -1054 -2522 -1044 -2488
rect -1096 -2556 -1044 -2522
rect -1096 -2590 -1088 -2556
rect -1054 -2590 -1044 -2556
rect -1096 -2606 -1044 -2590
rect -1014 -2488 -962 -2476
rect -1014 -2522 -1004 -2488
rect -970 -2522 -962 -2488
rect -1014 -2556 -962 -2522
rect -1014 -2590 -1004 -2556
rect -970 -2590 -962 -2556
rect -581 -2492 -529 -2476
rect -581 -2526 -573 -2492
rect -539 -2526 -529 -2492
rect -581 -2560 -529 -2526
rect -1014 -2606 -962 -2590
rect -581 -2594 -573 -2560
rect -539 -2594 -529 -2560
rect -581 -2606 -529 -2594
rect -499 -2606 -445 -2476
rect -415 -2492 -363 -2476
rect -415 -2526 -405 -2492
rect -371 -2526 -363 -2492
rect -415 -2560 -363 -2526
rect -415 -2594 -405 -2560
rect -371 -2594 -363 -2560
rect -415 -2606 -363 -2594
rect -1096 -2716 -1044 -2700
rect -1096 -2750 -1088 -2716
rect -1054 -2750 -1044 -2716
rect -1096 -2784 -1044 -2750
rect -1096 -2818 -1088 -2784
rect -1054 -2818 -1044 -2784
rect -1096 -2830 -1044 -2818
rect -1014 -2716 -962 -2700
rect -1014 -2750 -1004 -2716
rect -970 -2750 -962 -2716
rect -581 -2712 -529 -2700
rect -1014 -2784 -962 -2750
rect -1014 -2818 -1004 -2784
rect -970 -2818 -962 -2784
rect -1014 -2830 -962 -2818
rect -581 -2746 -573 -2712
rect -539 -2746 -529 -2712
rect -581 -2780 -529 -2746
rect -581 -2814 -573 -2780
rect -539 -2814 -529 -2780
rect -581 -2830 -529 -2814
rect -499 -2830 -445 -2700
rect -415 -2712 -363 -2700
rect -415 -2746 -405 -2712
rect -371 -2746 -363 -2712
rect -415 -2780 -363 -2746
rect -415 -2814 -405 -2780
rect -371 -2814 -363 -2780
rect -415 -2830 -363 -2814
rect 423 -3002 485 -2990
rect 423 -3082 435 -3002
rect 469 -3082 485 -3002
rect 423 -3094 485 -3082
rect 515 -3002 581 -2990
rect 515 -3082 531 -3002
rect 565 -3082 581 -3002
rect 515 -3094 581 -3082
rect 611 -3002 677 -2990
rect 611 -3082 627 -3002
rect 661 -3082 677 -3002
rect 611 -3094 677 -3082
rect 707 -3002 773 -2990
rect 707 -3082 723 -3002
rect 757 -3082 773 -3002
rect 707 -3094 773 -3082
rect 803 -3002 869 -2990
rect 803 -3082 819 -3002
rect 853 -3082 869 -3002
rect 803 -3094 869 -3082
rect 899 -3002 965 -2990
rect 899 -3082 915 -3002
rect 949 -3082 965 -3002
rect 899 -3094 965 -3082
rect 995 -3002 1061 -2990
rect 995 -3082 1011 -3002
rect 1045 -3082 1061 -3002
rect 995 -3094 1061 -3082
rect 1091 -3002 1157 -2990
rect 1091 -3082 1107 -3002
rect 1141 -3082 1157 -3002
rect 1091 -3094 1157 -3082
rect 1187 -3002 1253 -2990
rect 1187 -3082 1203 -3002
rect 1237 -3082 1253 -3002
rect 1187 -3094 1253 -3082
rect 1283 -3002 1349 -2990
rect 1283 -3082 1299 -3002
rect 1333 -3082 1349 -3002
rect 1283 -3094 1349 -3082
rect 1379 -3002 1441 -2990
rect 1379 -3082 1395 -3002
rect 1429 -3082 1441 -3002
rect 1379 -3094 1441 -3082
rect 1603 -3008 1661 -2996
rect 1603 -3084 1615 -3008
rect 1649 -3084 1661 -3008
rect 1603 -3096 1661 -3084
rect 1691 -3008 1749 -2996
rect 1691 -3084 1703 -3008
rect 1737 -3084 1749 -3008
rect 1691 -3096 1749 -3084
rect 1944 -3002 2006 -2990
rect 1944 -3082 1956 -3002
rect 1990 -3082 2006 -3002
rect 1944 -3094 2006 -3082
rect 2036 -3002 2102 -2990
rect 2036 -3082 2052 -3002
rect 2086 -3082 2102 -3002
rect 2036 -3094 2102 -3082
rect 2132 -3002 2198 -2990
rect 2132 -3082 2148 -3002
rect 2182 -3082 2198 -3002
rect 2132 -3094 2198 -3082
rect 2228 -3002 2294 -2990
rect 2228 -3082 2244 -3002
rect 2278 -3082 2294 -3002
rect 2228 -3094 2294 -3082
rect 2324 -3002 2390 -2990
rect 2324 -3082 2340 -3002
rect 2374 -3082 2390 -3002
rect 2324 -3094 2390 -3082
rect 2420 -3002 2486 -2990
rect 2420 -3082 2436 -3002
rect 2470 -3082 2486 -3002
rect 2420 -3094 2486 -3082
rect 2516 -3002 2582 -2990
rect 2516 -3082 2532 -3002
rect 2566 -3082 2582 -3002
rect 2516 -3094 2582 -3082
rect 2612 -3002 2678 -2990
rect 2612 -3082 2628 -3002
rect 2662 -3082 2678 -3002
rect 2612 -3094 2678 -3082
rect 2708 -3002 2774 -2990
rect 2708 -3082 2724 -3002
rect 2758 -3082 2774 -3002
rect 2708 -3094 2774 -3082
rect 2804 -3002 2870 -2990
rect 2804 -3082 2820 -3002
rect 2854 -3082 2870 -3002
rect 2804 -3094 2870 -3082
rect 2900 -3002 2962 -2990
rect 2900 -3082 2916 -3002
rect 2950 -3082 2962 -3002
rect 2900 -3094 2962 -3082
rect -3128 -3588 -3066 -3576
rect -3128 -3668 -3116 -3588
rect -3082 -3668 -3066 -3588
rect -3128 -3680 -3066 -3668
rect -3036 -3588 -2970 -3576
rect -3036 -3668 -3020 -3588
rect -2986 -3668 -2970 -3588
rect -3036 -3680 -2970 -3668
rect -2940 -3588 -2874 -3576
rect -2940 -3668 -2924 -3588
rect -2890 -3668 -2874 -3588
rect -2940 -3680 -2874 -3668
rect -2844 -3588 -2778 -3576
rect -2844 -3668 -2828 -3588
rect -2794 -3668 -2778 -3588
rect -2844 -3680 -2778 -3668
rect -2748 -3588 -2682 -3576
rect -2748 -3668 -2732 -3588
rect -2698 -3668 -2682 -3588
rect -2748 -3680 -2682 -3668
rect -2652 -3588 -2586 -3576
rect -2652 -3668 -2636 -3588
rect -2602 -3668 -2586 -3588
rect -2652 -3680 -2586 -3668
rect -2556 -3588 -2490 -3576
rect -2556 -3668 -2540 -3588
rect -2506 -3668 -2490 -3588
rect -2556 -3680 -2490 -3668
rect -2460 -3588 -2394 -3576
rect -2460 -3668 -2444 -3588
rect -2410 -3668 -2394 -3588
rect -2460 -3680 -2394 -3668
rect -2364 -3588 -2298 -3576
rect -2364 -3668 -2348 -3588
rect -2314 -3668 -2298 -3588
rect -2364 -3680 -2298 -3668
rect -2268 -3588 -2202 -3576
rect -2268 -3668 -2252 -3588
rect -2218 -3668 -2202 -3588
rect -2268 -3680 -2202 -3668
rect -2172 -3588 -2110 -3576
rect -2172 -3668 -2156 -3588
rect -2122 -3668 -2110 -3588
rect -2172 -3680 -2110 -3668
rect -581 -3580 -529 -3564
rect -581 -3614 -573 -3580
rect -539 -3614 -529 -3580
rect -581 -3648 -529 -3614
rect -581 -3682 -573 -3648
rect -539 -3682 -529 -3648
rect -581 -3694 -529 -3682
rect -499 -3694 -445 -3564
rect -415 -3580 -363 -3564
rect -415 -3614 -405 -3580
rect -371 -3614 -363 -3580
rect -415 -3648 -363 -3614
rect -415 -3682 -405 -3648
rect -371 -3682 -363 -3648
rect -415 -3694 -363 -3682
rect -544 -3804 -492 -3788
rect -544 -3838 -536 -3804
rect -502 -3838 -492 -3804
rect -544 -3872 -492 -3838
rect -544 -3906 -536 -3872
rect -502 -3906 -492 -3872
rect -544 -3918 -492 -3906
rect -462 -3804 -410 -3788
rect -462 -3838 -452 -3804
rect -418 -3838 -410 -3804
rect -462 -3872 -410 -3838
rect -462 -3906 -452 -3872
rect -418 -3906 -410 -3872
rect -462 -3918 -410 -3906
rect 423 -4380 485 -4368
rect 423 -4460 435 -4380
rect 469 -4460 485 -4380
rect 423 -4472 485 -4460
rect 515 -4380 581 -4368
rect 515 -4460 531 -4380
rect 565 -4460 581 -4380
rect 515 -4472 581 -4460
rect 611 -4380 677 -4368
rect 611 -4460 627 -4380
rect 661 -4460 677 -4380
rect 611 -4472 677 -4460
rect 707 -4380 773 -4368
rect 707 -4460 723 -4380
rect 757 -4460 773 -4380
rect 707 -4472 773 -4460
rect 803 -4380 869 -4368
rect 803 -4460 819 -4380
rect 853 -4460 869 -4380
rect 803 -4472 869 -4460
rect 899 -4380 965 -4368
rect 899 -4460 915 -4380
rect 949 -4460 965 -4380
rect 899 -4472 965 -4460
rect 995 -4380 1061 -4368
rect 995 -4460 1011 -4380
rect 1045 -4460 1061 -4380
rect 995 -4472 1061 -4460
rect 1091 -4380 1157 -4368
rect 1091 -4460 1107 -4380
rect 1141 -4460 1157 -4380
rect 1091 -4472 1157 -4460
rect 1187 -4380 1253 -4368
rect 1187 -4460 1203 -4380
rect 1237 -4460 1253 -4380
rect 1187 -4472 1253 -4460
rect 1283 -4380 1349 -4368
rect 1283 -4460 1299 -4380
rect 1333 -4460 1349 -4380
rect 1283 -4472 1349 -4460
rect 1379 -4380 1441 -4368
rect 1379 -4460 1395 -4380
rect 1429 -4460 1441 -4380
rect 1379 -4472 1441 -4460
rect 1603 -4386 1661 -4374
rect 1603 -4462 1615 -4386
rect 1649 -4462 1661 -4386
rect 1603 -4474 1661 -4462
rect 1691 -4386 1749 -4374
rect 1691 -4462 1703 -4386
rect 1737 -4462 1749 -4386
rect 1691 -4474 1749 -4462
rect 1944 -4380 2006 -4368
rect 1944 -4460 1956 -4380
rect 1990 -4460 2006 -4380
rect 1944 -4472 2006 -4460
rect 2036 -4380 2102 -4368
rect 2036 -4460 2052 -4380
rect 2086 -4460 2102 -4380
rect 2036 -4472 2102 -4460
rect 2132 -4380 2198 -4368
rect 2132 -4460 2148 -4380
rect 2182 -4460 2198 -4380
rect 2132 -4472 2198 -4460
rect 2228 -4380 2294 -4368
rect 2228 -4460 2244 -4380
rect 2278 -4460 2294 -4380
rect 2228 -4472 2294 -4460
rect 2324 -4380 2390 -4368
rect 2324 -4460 2340 -4380
rect 2374 -4460 2390 -4380
rect 2324 -4472 2390 -4460
rect 2420 -4380 2486 -4368
rect 2420 -4460 2436 -4380
rect 2470 -4460 2486 -4380
rect 2420 -4472 2486 -4460
rect 2516 -4380 2582 -4368
rect 2516 -4460 2532 -4380
rect 2566 -4460 2582 -4380
rect 2516 -4472 2582 -4460
rect 2612 -4380 2678 -4368
rect 2612 -4460 2628 -4380
rect 2662 -4460 2678 -4380
rect 2612 -4472 2678 -4460
rect 2708 -4380 2774 -4368
rect 2708 -4460 2724 -4380
rect 2758 -4460 2774 -4380
rect 2708 -4472 2774 -4460
rect 2804 -4380 2870 -4368
rect 2804 -4460 2820 -4380
rect 2854 -4460 2870 -4380
rect 2804 -4472 2870 -4460
rect 2900 -4380 2962 -4368
rect 2900 -4460 2916 -4380
rect 2950 -4460 2962 -4380
rect 2900 -4472 2962 -4460
rect -544 -4664 -492 -4652
rect -544 -4698 -536 -4664
rect -502 -4698 -492 -4664
rect -544 -4732 -492 -4698
rect -544 -4766 -536 -4732
rect -502 -4766 -492 -4732
rect -544 -4782 -492 -4766
rect -462 -4664 -410 -4652
rect -462 -4698 -452 -4664
rect -418 -4698 -410 -4664
rect -462 -4732 -410 -4698
rect -462 -4766 -452 -4732
rect -418 -4766 -410 -4732
rect -462 -4782 -410 -4766
rect -3128 -4966 -3066 -4954
rect -3128 -5046 -3116 -4966
rect -3082 -5046 -3066 -4966
rect -3128 -5058 -3066 -5046
rect -3036 -4966 -2970 -4954
rect -3036 -5046 -3020 -4966
rect -2986 -5046 -2970 -4966
rect -3036 -5058 -2970 -5046
rect -2940 -4966 -2874 -4954
rect -2940 -5046 -2924 -4966
rect -2890 -5046 -2874 -4966
rect -2940 -5058 -2874 -5046
rect -2844 -4966 -2778 -4954
rect -2844 -5046 -2828 -4966
rect -2794 -5046 -2778 -4966
rect -2844 -5058 -2778 -5046
rect -2748 -4966 -2682 -4954
rect -2748 -5046 -2732 -4966
rect -2698 -5046 -2682 -4966
rect -2748 -5058 -2682 -5046
rect -2652 -4966 -2586 -4954
rect -2652 -5046 -2636 -4966
rect -2602 -5046 -2586 -4966
rect -2652 -5058 -2586 -5046
rect -2556 -4966 -2490 -4954
rect -2556 -5046 -2540 -4966
rect -2506 -5046 -2490 -4966
rect -2556 -5058 -2490 -5046
rect -2460 -4966 -2394 -4954
rect -2460 -5046 -2444 -4966
rect -2410 -5046 -2394 -4966
rect -2460 -5058 -2394 -5046
rect -2364 -4966 -2298 -4954
rect -2364 -5046 -2348 -4966
rect -2314 -5046 -2298 -4966
rect -2364 -5058 -2298 -5046
rect -2268 -4966 -2202 -4954
rect -2268 -5046 -2252 -4966
rect -2218 -5046 -2202 -4966
rect -2268 -5058 -2202 -5046
rect -2172 -4966 -2110 -4954
rect -2172 -5046 -2156 -4966
rect -2122 -5046 -2110 -4966
rect -2172 -5058 -2110 -5046
<< pdiff >>
rect -3128 -298 -3066 -286
rect -3128 -546 -3116 -298
rect -3082 -546 -3066 -298
rect -3128 -558 -3066 -546
rect -3036 -298 -2970 -286
rect -3036 -546 -3020 -298
rect -2986 -546 -2970 -298
rect -3036 -558 -2970 -546
rect -2940 -298 -2874 -286
rect -2940 -546 -2924 -298
rect -2890 -546 -2874 -298
rect -2940 -558 -2874 -546
rect -2844 -298 -2778 -286
rect -2844 -546 -2828 -298
rect -2794 -546 -2778 -298
rect -2844 -558 -2778 -546
rect -2748 -298 -2682 -286
rect -2748 -546 -2732 -298
rect -2698 -546 -2682 -298
rect -2748 -558 -2682 -546
rect -2652 -298 -2586 -286
rect -2652 -546 -2636 -298
rect -2602 -546 -2586 -298
rect -2652 -558 -2586 -546
rect -2556 -298 -2490 -286
rect -2556 -546 -2540 -298
rect -2506 -546 -2490 -298
rect -2556 -558 -2490 -546
rect -2460 -298 -2394 -286
rect -2460 -546 -2444 -298
rect -2410 -546 -2394 -298
rect -2460 -558 -2394 -546
rect -2364 -298 -2298 -286
rect -2364 -546 -2348 -298
rect -2314 -546 -2298 -298
rect -2364 -558 -2298 -546
rect -2268 -298 -2202 -286
rect -2268 -546 -2252 -298
rect -2218 -546 -2202 -298
rect -2268 -558 -2202 -546
rect -2172 -298 -2110 -286
rect -2172 -546 -2156 -298
rect -2122 -546 -2110 -298
rect -2172 -558 -2110 -546
rect -912 -792 -860 -774
rect -912 -826 -904 -792
rect -870 -826 -860 -792
rect -912 -860 -860 -826
rect -912 -894 -904 -860
rect -870 -894 -860 -860
rect -912 -928 -860 -894
rect -912 -962 -904 -928
rect -870 -962 -860 -928
rect -912 -974 -860 -962
rect -830 -792 -778 -774
rect -830 -826 -820 -792
rect -786 -826 -778 -792
rect -830 -860 -778 -826
rect -830 -894 -820 -860
rect -786 -894 -778 -860
rect -830 -928 -778 -894
rect -830 -962 -820 -928
rect -786 -962 -778 -928
rect -544 -792 -492 -774
rect -544 -826 -536 -792
rect -502 -826 -492 -792
rect -544 -860 -492 -826
rect -544 -894 -536 -860
rect -502 -894 -492 -860
rect -544 -928 -492 -894
rect -830 -974 -778 -962
rect -544 -962 -536 -928
rect -502 -962 -492 -928
rect -544 -974 -492 -962
rect -462 -792 -410 -774
rect -462 -826 -452 -792
rect -418 -826 -410 -792
rect -462 -860 -410 -826
rect -462 -894 -452 -860
rect -418 -894 -410 -860
rect -462 -928 -410 -894
rect -462 -962 -452 -928
rect -418 -962 -410 -928
rect -462 -974 -410 -962
rect 423 -700 485 -688
rect 423 -948 435 -700
rect 469 -948 485 -700
rect 423 -960 485 -948
rect 515 -700 581 -688
rect 515 -948 531 -700
rect 565 -948 581 -700
rect 515 -960 581 -948
rect 611 -700 677 -688
rect 611 -948 627 -700
rect 661 -948 677 -700
rect 611 -960 677 -948
rect 707 -700 773 -688
rect 707 -948 723 -700
rect 757 -948 773 -700
rect 707 -960 773 -948
rect 803 -700 869 -688
rect 803 -948 819 -700
rect 853 -948 869 -700
rect 803 -960 869 -948
rect 899 -700 965 -688
rect 899 -948 915 -700
rect 949 -948 965 -700
rect 899 -960 965 -948
rect 995 -700 1061 -688
rect 995 -948 1011 -700
rect 1045 -948 1061 -700
rect 995 -960 1061 -948
rect 1091 -700 1157 -688
rect 1091 -948 1107 -700
rect 1141 -948 1157 -700
rect 1091 -960 1157 -948
rect 1187 -700 1253 -688
rect 1187 -948 1203 -700
rect 1237 -948 1253 -700
rect 1187 -960 1253 -948
rect 1283 -700 1349 -688
rect 1283 -948 1299 -700
rect 1333 -948 1349 -700
rect 1283 -960 1349 -948
rect 1379 -700 1441 -688
rect 1379 -948 1395 -700
rect 1429 -948 1441 -700
rect 1379 -960 1441 -948
rect -544 -1080 -492 -1068
rect -544 -1114 -536 -1080
rect -502 -1114 -492 -1080
rect -544 -1148 -492 -1114
rect -544 -1182 -536 -1148
rect -502 -1182 -492 -1148
rect -544 -1216 -492 -1182
rect -544 -1250 -536 -1216
rect -502 -1250 -492 -1216
rect -544 -1268 -492 -1250
rect -462 -1080 -410 -1068
rect -462 -1114 -452 -1080
rect -418 -1114 -410 -1080
rect -462 -1148 -410 -1114
rect 1944 -700 2006 -688
rect 1944 -948 1956 -700
rect 1990 -948 2006 -700
rect 1944 -960 2006 -948
rect 2036 -700 2102 -688
rect 2036 -948 2052 -700
rect 2086 -948 2102 -700
rect 2036 -960 2102 -948
rect 2132 -700 2198 -688
rect 2132 -948 2148 -700
rect 2182 -948 2198 -700
rect 2132 -960 2198 -948
rect 2228 -700 2294 -688
rect 2228 -948 2244 -700
rect 2278 -948 2294 -700
rect 2228 -960 2294 -948
rect 2324 -700 2390 -688
rect 2324 -948 2340 -700
rect 2374 -948 2390 -700
rect 2324 -960 2390 -948
rect 2420 -700 2486 -688
rect 2420 -948 2436 -700
rect 2470 -948 2486 -700
rect 2420 -960 2486 -948
rect 2516 -700 2582 -688
rect 2516 -948 2532 -700
rect 2566 -948 2582 -700
rect 2516 -960 2582 -948
rect 2612 -700 2678 -688
rect 2612 -948 2628 -700
rect 2662 -948 2678 -700
rect 2612 -960 2678 -948
rect 2708 -700 2774 -688
rect 2708 -948 2724 -700
rect 2758 -948 2774 -700
rect 2708 -960 2774 -948
rect 2804 -700 2870 -688
rect 2804 -948 2820 -700
rect 2854 -948 2870 -700
rect 2804 -960 2870 -948
rect 2900 -700 2962 -688
rect 2900 -948 2916 -700
rect 2950 -948 2962 -700
rect 2900 -960 2962 -948
rect -462 -1182 -452 -1148
rect -418 -1182 -410 -1148
rect -462 -1216 -410 -1182
rect -462 -1250 -452 -1216
rect -418 -1250 -410 -1216
rect -462 -1268 -410 -1250
rect -3128 -1632 -3066 -1620
rect -3128 -1880 -3116 -1632
rect -3082 -1880 -3066 -1632
rect -3128 -1892 -3066 -1880
rect -3036 -1632 -2970 -1620
rect -3036 -1880 -3020 -1632
rect -2986 -1880 -2970 -1632
rect -3036 -1892 -2970 -1880
rect -2940 -1632 -2874 -1620
rect -2940 -1880 -2924 -1632
rect -2890 -1880 -2874 -1632
rect -2940 -1892 -2874 -1880
rect -2844 -1632 -2778 -1620
rect -2844 -1880 -2828 -1632
rect -2794 -1880 -2778 -1632
rect -2844 -1892 -2778 -1880
rect -2748 -1632 -2682 -1620
rect -2748 -1880 -2732 -1632
rect -2698 -1880 -2682 -1632
rect -2748 -1892 -2682 -1880
rect -2652 -1632 -2586 -1620
rect -2652 -1880 -2636 -1632
rect -2602 -1880 -2586 -1632
rect -2652 -1892 -2586 -1880
rect -2556 -1632 -2490 -1620
rect -2556 -1880 -2540 -1632
rect -2506 -1880 -2490 -1632
rect -2556 -1892 -2490 -1880
rect -2460 -1632 -2394 -1620
rect -2460 -1880 -2444 -1632
rect -2410 -1880 -2394 -1632
rect -2460 -1892 -2394 -1880
rect -2364 -1632 -2298 -1620
rect -2364 -1880 -2348 -1632
rect -2314 -1880 -2298 -1632
rect -2364 -1892 -2298 -1880
rect -2268 -1632 -2202 -1620
rect -2268 -1880 -2252 -1632
rect -2218 -1880 -2202 -1632
rect -2268 -1892 -2202 -1880
rect -2172 -1632 -2110 -1620
rect -2172 -1880 -2156 -1632
rect -2122 -1880 -2110 -1632
rect -2172 -1892 -2110 -1880
rect -581 -1880 -529 -1862
rect -581 -1914 -573 -1880
rect -539 -1914 -529 -1880
rect -581 -1948 -529 -1914
rect -581 -1982 -573 -1948
rect -539 -1982 -529 -1948
rect -581 -2016 -529 -1982
rect -581 -2050 -573 -2016
rect -539 -2050 -529 -2016
rect -581 -2062 -529 -2050
rect -499 -1880 -445 -1862
rect -499 -1914 -489 -1880
rect -455 -1914 -445 -1880
rect -499 -1948 -445 -1914
rect -499 -1982 -489 -1948
rect -455 -1982 -445 -1948
rect -499 -2016 -445 -1982
rect -499 -2050 -489 -2016
rect -455 -2050 -445 -2016
rect -499 -2062 -445 -2050
rect -415 -1880 -363 -1862
rect -415 -1914 -405 -1880
rect -371 -1914 -363 -1880
rect -415 -1948 -363 -1914
rect -415 -1982 -405 -1948
rect -371 -1982 -363 -1948
rect -415 -2016 -363 -1982
rect -415 -2050 -405 -2016
rect -371 -2050 -363 -2016
rect -415 -2062 -363 -2050
rect -1096 -2168 -1044 -2156
rect -1096 -2202 -1088 -2168
rect -1054 -2202 -1044 -2168
rect -1096 -2236 -1044 -2202
rect -1096 -2270 -1088 -2236
rect -1054 -2270 -1044 -2236
rect -1096 -2304 -1044 -2270
rect -1096 -2338 -1088 -2304
rect -1054 -2338 -1044 -2304
rect -1096 -2356 -1044 -2338
rect -1014 -2168 -962 -2156
rect -1014 -2202 -1004 -2168
rect -970 -2202 -962 -2168
rect -581 -2168 -529 -2156
rect -1014 -2236 -962 -2202
rect -1014 -2270 -1004 -2236
rect -970 -2270 -962 -2236
rect -1014 -2304 -962 -2270
rect -1014 -2338 -1004 -2304
rect -970 -2338 -962 -2304
rect -1014 -2356 -962 -2338
rect -581 -2202 -573 -2168
rect -539 -2202 -529 -2168
rect -581 -2236 -529 -2202
rect -581 -2270 -573 -2236
rect -539 -2270 -529 -2236
rect -581 -2304 -529 -2270
rect -581 -2338 -573 -2304
rect -539 -2338 -529 -2304
rect -581 -2356 -529 -2338
rect -499 -2168 -445 -2156
rect -499 -2202 -489 -2168
rect -455 -2202 -445 -2168
rect -499 -2236 -445 -2202
rect -499 -2270 -489 -2236
rect -455 -2270 -445 -2236
rect -499 -2304 -445 -2270
rect -499 -2338 -489 -2304
rect -455 -2338 -445 -2304
rect -499 -2356 -445 -2338
rect -415 -2168 -363 -2156
rect -415 -2202 -405 -2168
rect -371 -2202 -363 -2168
rect -415 -2236 -363 -2202
rect -415 -2270 -405 -2236
rect -371 -2270 -363 -2236
rect -415 -2304 -363 -2270
rect -415 -2338 -405 -2304
rect -371 -2338 -363 -2304
rect -415 -2356 -363 -2338
rect 423 -2034 485 -2022
rect 423 -2282 435 -2034
rect 469 -2282 485 -2034
rect 423 -2294 485 -2282
rect 515 -2034 581 -2022
rect 515 -2282 531 -2034
rect 565 -2282 581 -2034
rect 515 -2294 581 -2282
rect 611 -2034 677 -2022
rect 611 -2282 627 -2034
rect 661 -2282 677 -2034
rect 611 -2294 677 -2282
rect 707 -2034 773 -2022
rect 707 -2282 723 -2034
rect 757 -2282 773 -2034
rect 707 -2294 773 -2282
rect 803 -2034 869 -2022
rect 803 -2282 819 -2034
rect 853 -2282 869 -2034
rect 803 -2294 869 -2282
rect 899 -2034 965 -2022
rect 899 -2282 915 -2034
rect 949 -2282 965 -2034
rect 899 -2294 965 -2282
rect 995 -2034 1061 -2022
rect 995 -2282 1011 -2034
rect 1045 -2282 1061 -2034
rect 995 -2294 1061 -2282
rect 1091 -2034 1157 -2022
rect 1091 -2282 1107 -2034
rect 1141 -2282 1157 -2034
rect 1091 -2294 1157 -2282
rect 1187 -2034 1253 -2022
rect 1187 -2282 1203 -2034
rect 1237 -2282 1253 -2034
rect 1187 -2294 1253 -2282
rect 1283 -2034 1349 -2022
rect 1283 -2282 1299 -2034
rect 1333 -2282 1349 -2034
rect 1283 -2294 1349 -2282
rect 1379 -2034 1441 -2022
rect 1379 -2282 1395 -2034
rect 1429 -2282 1441 -2034
rect 1379 -2294 1441 -2282
rect 1944 -2034 2006 -2022
rect 1944 -2282 1956 -2034
rect 1990 -2282 2006 -2034
rect 1944 -2294 2006 -2282
rect 2036 -2034 2102 -2022
rect 2036 -2282 2052 -2034
rect 2086 -2282 2102 -2034
rect 2036 -2294 2102 -2282
rect 2132 -2034 2198 -2022
rect 2132 -2282 2148 -2034
rect 2182 -2282 2198 -2034
rect 2132 -2294 2198 -2282
rect 2228 -2034 2294 -2022
rect 2228 -2282 2244 -2034
rect 2278 -2282 2294 -2034
rect 2228 -2294 2294 -2282
rect 2324 -2034 2390 -2022
rect 2324 -2282 2340 -2034
rect 2374 -2282 2390 -2034
rect 2324 -2294 2390 -2282
rect 2420 -2034 2486 -2022
rect 2420 -2282 2436 -2034
rect 2470 -2282 2486 -2034
rect 2420 -2294 2486 -2282
rect 2516 -2034 2582 -2022
rect 2516 -2282 2532 -2034
rect 2566 -2282 2582 -2034
rect 2516 -2294 2582 -2282
rect 2612 -2034 2678 -2022
rect 2612 -2282 2628 -2034
rect 2662 -2282 2678 -2034
rect 2612 -2294 2678 -2282
rect 2708 -2034 2774 -2022
rect 2708 -2282 2724 -2034
rect 2758 -2282 2774 -2034
rect 2708 -2294 2774 -2282
rect 2804 -2034 2870 -2022
rect 2804 -2282 2820 -2034
rect 2854 -2282 2870 -2034
rect 2804 -2294 2870 -2282
rect 2900 -2034 2962 -2022
rect 2900 -2282 2916 -2034
rect 2950 -2282 2962 -2034
rect 2900 -2294 2962 -2282
rect -3128 -3010 -3066 -2998
rect -3128 -3258 -3116 -3010
rect -3082 -3258 -3066 -3010
rect -3128 -3270 -3066 -3258
rect -3036 -3010 -2970 -2998
rect -3036 -3258 -3020 -3010
rect -2986 -3258 -2970 -3010
rect -3036 -3270 -2970 -3258
rect -2940 -3010 -2874 -2998
rect -2940 -3258 -2924 -3010
rect -2890 -3258 -2874 -3010
rect -2940 -3270 -2874 -3258
rect -2844 -3010 -2778 -2998
rect -2844 -3258 -2828 -3010
rect -2794 -3258 -2778 -3010
rect -2844 -3270 -2778 -3258
rect -2748 -3010 -2682 -2998
rect -2748 -3258 -2732 -3010
rect -2698 -3258 -2682 -3010
rect -2748 -3270 -2682 -3258
rect -2652 -3010 -2586 -2998
rect -2652 -3258 -2636 -3010
rect -2602 -3258 -2586 -3010
rect -2652 -3270 -2586 -3258
rect -2556 -3010 -2490 -2998
rect -2556 -3258 -2540 -3010
rect -2506 -3258 -2490 -3010
rect -2556 -3270 -2490 -3258
rect -2460 -3010 -2394 -2998
rect -2460 -3258 -2444 -3010
rect -2410 -3258 -2394 -3010
rect -2460 -3270 -2394 -3258
rect -2364 -3010 -2298 -2998
rect -2364 -3258 -2348 -3010
rect -2314 -3258 -2298 -3010
rect -2364 -3270 -2298 -3258
rect -2268 -3010 -2202 -2998
rect -2268 -3258 -2252 -3010
rect -2218 -3258 -2202 -3010
rect -2268 -3270 -2202 -3258
rect -2172 -3010 -2110 -2998
rect -2172 -3258 -2156 -3010
rect -2122 -3258 -2110 -3010
rect -2172 -3270 -2110 -3258
rect -1096 -2968 -1044 -2950
rect -1096 -3002 -1088 -2968
rect -1054 -3002 -1044 -2968
rect -1096 -3036 -1044 -3002
rect -1096 -3070 -1088 -3036
rect -1054 -3070 -1044 -3036
rect -1096 -3104 -1044 -3070
rect -1096 -3138 -1088 -3104
rect -1054 -3138 -1044 -3104
rect -1096 -3150 -1044 -3138
rect -1014 -2968 -962 -2950
rect -1014 -3002 -1004 -2968
rect -970 -3002 -962 -2968
rect -1014 -3036 -962 -3002
rect -1014 -3070 -1004 -3036
rect -970 -3070 -962 -3036
rect -1014 -3104 -962 -3070
rect -1014 -3138 -1004 -3104
rect -970 -3138 -962 -3104
rect -581 -2968 -529 -2950
rect -581 -3002 -573 -2968
rect -539 -3002 -529 -2968
rect -581 -3036 -529 -3002
rect -581 -3070 -573 -3036
rect -539 -3070 -529 -3036
rect -581 -3104 -529 -3070
rect -1014 -3150 -962 -3138
rect -581 -3138 -573 -3104
rect -539 -3138 -529 -3104
rect -581 -3150 -529 -3138
rect -499 -2968 -445 -2950
rect -499 -3002 -489 -2968
rect -455 -3002 -445 -2968
rect -499 -3036 -445 -3002
rect -499 -3070 -489 -3036
rect -455 -3070 -445 -3036
rect -499 -3104 -445 -3070
rect -499 -3138 -489 -3104
rect -455 -3138 -445 -3104
rect -499 -3150 -445 -3138
rect -415 -2968 -363 -2950
rect -415 -3002 -405 -2968
rect -371 -3002 -363 -2968
rect -415 -3036 -363 -3002
rect -415 -3070 -405 -3036
rect -371 -3070 -363 -3036
rect -415 -3104 -363 -3070
rect -415 -3138 -405 -3104
rect -371 -3138 -363 -3104
rect -415 -3150 -363 -3138
rect -581 -3256 -529 -3244
rect -581 -3290 -573 -3256
rect -539 -3290 -529 -3256
rect -581 -3324 -529 -3290
rect -581 -3358 -573 -3324
rect -539 -3358 -529 -3324
rect -581 -3392 -529 -3358
rect -581 -3426 -573 -3392
rect -539 -3426 -529 -3392
rect -581 -3444 -529 -3426
rect -499 -3256 -445 -3244
rect -499 -3290 -489 -3256
rect -455 -3290 -445 -3256
rect -499 -3324 -445 -3290
rect -499 -3358 -489 -3324
rect -455 -3358 -445 -3324
rect -499 -3392 -445 -3358
rect -499 -3426 -489 -3392
rect -455 -3426 -445 -3392
rect -499 -3444 -445 -3426
rect -415 -3256 -363 -3244
rect -415 -3290 -405 -3256
rect -371 -3290 -363 -3256
rect -415 -3324 -363 -3290
rect -415 -3358 -405 -3324
rect -371 -3358 -363 -3324
rect -415 -3392 -363 -3358
rect -415 -3426 -405 -3392
rect -371 -3426 -363 -3392
rect -415 -3444 -363 -3426
rect 423 -3412 485 -3400
rect 423 -3660 435 -3412
rect 469 -3660 485 -3412
rect 423 -3672 485 -3660
rect 515 -3412 581 -3400
rect 515 -3660 531 -3412
rect 565 -3660 581 -3412
rect 515 -3672 581 -3660
rect 611 -3412 677 -3400
rect 611 -3660 627 -3412
rect 661 -3660 677 -3412
rect 611 -3672 677 -3660
rect 707 -3412 773 -3400
rect 707 -3660 723 -3412
rect 757 -3660 773 -3412
rect 707 -3672 773 -3660
rect 803 -3412 869 -3400
rect 803 -3660 819 -3412
rect 853 -3660 869 -3412
rect 803 -3672 869 -3660
rect 899 -3412 965 -3400
rect 899 -3660 915 -3412
rect 949 -3660 965 -3412
rect 899 -3672 965 -3660
rect 995 -3412 1061 -3400
rect 995 -3660 1011 -3412
rect 1045 -3660 1061 -3412
rect 995 -3672 1061 -3660
rect 1091 -3412 1157 -3400
rect 1091 -3660 1107 -3412
rect 1141 -3660 1157 -3412
rect 1091 -3672 1157 -3660
rect 1187 -3412 1253 -3400
rect 1187 -3660 1203 -3412
rect 1237 -3660 1253 -3412
rect 1187 -3672 1253 -3660
rect 1283 -3412 1349 -3400
rect 1283 -3660 1299 -3412
rect 1333 -3660 1349 -3412
rect 1283 -3672 1349 -3660
rect 1379 -3412 1441 -3400
rect 1379 -3660 1395 -3412
rect 1429 -3660 1441 -3412
rect 1379 -3672 1441 -3660
rect 1944 -3412 2006 -3400
rect 1944 -3660 1956 -3412
rect 1990 -3660 2006 -3412
rect 1944 -3672 2006 -3660
rect 2036 -3412 2102 -3400
rect 2036 -3660 2052 -3412
rect 2086 -3660 2102 -3412
rect 2036 -3672 2102 -3660
rect 2132 -3412 2198 -3400
rect 2132 -3660 2148 -3412
rect 2182 -3660 2198 -3412
rect 2132 -3672 2198 -3660
rect 2228 -3412 2294 -3400
rect 2228 -3660 2244 -3412
rect 2278 -3660 2294 -3412
rect 2228 -3672 2294 -3660
rect 2324 -3412 2390 -3400
rect 2324 -3660 2340 -3412
rect 2374 -3660 2390 -3412
rect 2324 -3672 2390 -3660
rect 2420 -3412 2486 -3400
rect 2420 -3660 2436 -3412
rect 2470 -3660 2486 -3412
rect 2420 -3672 2486 -3660
rect 2516 -3412 2582 -3400
rect 2516 -3660 2532 -3412
rect 2566 -3660 2582 -3412
rect 2516 -3672 2582 -3660
rect 2612 -3412 2678 -3400
rect 2612 -3660 2628 -3412
rect 2662 -3660 2678 -3412
rect 2612 -3672 2678 -3660
rect 2708 -3412 2774 -3400
rect 2708 -3660 2724 -3412
rect 2758 -3660 2774 -3412
rect 2708 -3672 2774 -3660
rect 2804 -3412 2870 -3400
rect 2804 -3660 2820 -3412
rect 2854 -3660 2870 -3412
rect 2804 -3672 2870 -3660
rect 2900 -3412 2962 -3400
rect 2900 -3660 2916 -3412
rect 2950 -3660 2962 -3412
rect 2900 -3672 2962 -3660
rect -544 -4056 -492 -4038
rect -544 -4090 -536 -4056
rect -502 -4090 -492 -4056
rect -544 -4124 -492 -4090
rect -544 -4158 -536 -4124
rect -502 -4158 -492 -4124
rect -544 -4192 -492 -4158
rect -544 -4226 -536 -4192
rect -502 -4226 -492 -4192
rect -544 -4238 -492 -4226
rect -462 -4056 -410 -4038
rect -462 -4090 -452 -4056
rect -418 -4090 -410 -4056
rect -462 -4124 -410 -4090
rect -462 -4158 -452 -4124
rect -418 -4158 -410 -4124
rect -462 -4192 -410 -4158
rect -462 -4226 -452 -4192
rect -418 -4226 -410 -4192
rect -462 -4238 -410 -4226
rect -3128 -4388 -3066 -4376
rect -3128 -4636 -3116 -4388
rect -3082 -4636 -3066 -4388
rect -3128 -4648 -3066 -4636
rect -3036 -4388 -2970 -4376
rect -3036 -4636 -3020 -4388
rect -2986 -4636 -2970 -4388
rect -3036 -4648 -2970 -4636
rect -2940 -4388 -2874 -4376
rect -2940 -4636 -2924 -4388
rect -2890 -4636 -2874 -4388
rect -2940 -4648 -2874 -4636
rect -2844 -4388 -2778 -4376
rect -2844 -4636 -2828 -4388
rect -2794 -4636 -2778 -4388
rect -2844 -4648 -2778 -4636
rect -2748 -4388 -2682 -4376
rect -2748 -4636 -2732 -4388
rect -2698 -4636 -2682 -4388
rect -2748 -4648 -2682 -4636
rect -2652 -4388 -2586 -4376
rect -2652 -4636 -2636 -4388
rect -2602 -4636 -2586 -4388
rect -2652 -4648 -2586 -4636
rect -2556 -4388 -2490 -4376
rect -2556 -4636 -2540 -4388
rect -2506 -4636 -2490 -4388
rect -2556 -4648 -2490 -4636
rect -2460 -4388 -2394 -4376
rect -2460 -4636 -2444 -4388
rect -2410 -4636 -2394 -4388
rect -2460 -4648 -2394 -4636
rect -2364 -4388 -2298 -4376
rect -2364 -4636 -2348 -4388
rect -2314 -4636 -2298 -4388
rect -2364 -4648 -2298 -4636
rect -2268 -4388 -2202 -4376
rect -2268 -4636 -2252 -4388
rect -2218 -4636 -2202 -4388
rect -2268 -4648 -2202 -4636
rect -2172 -4388 -2110 -4376
rect -2172 -4636 -2156 -4388
rect -2122 -4636 -2110 -4388
rect -2172 -4648 -2110 -4636
rect -544 -4344 -492 -4332
rect -544 -4378 -536 -4344
rect -502 -4378 -492 -4344
rect -544 -4412 -492 -4378
rect -544 -4446 -536 -4412
rect -502 -4446 -492 -4412
rect -544 -4480 -492 -4446
rect -544 -4514 -536 -4480
rect -502 -4514 -492 -4480
rect -544 -4532 -492 -4514
rect -462 -4344 -410 -4332
rect -462 -4378 -452 -4344
rect -418 -4378 -410 -4344
rect -462 -4412 -410 -4378
rect -462 -4446 -452 -4412
rect -418 -4446 -410 -4412
rect -462 -4480 -410 -4446
rect -462 -4514 -452 -4480
rect -418 -4514 -410 -4480
rect -462 -4532 -410 -4514
rect 423 -4790 485 -4778
rect 423 -5038 435 -4790
rect 469 -5038 485 -4790
rect 423 -5050 485 -5038
rect 515 -4790 581 -4778
rect 515 -5038 531 -4790
rect 565 -5038 581 -4790
rect 515 -5050 581 -5038
rect 611 -4790 677 -4778
rect 611 -5038 627 -4790
rect 661 -5038 677 -4790
rect 611 -5050 677 -5038
rect 707 -4790 773 -4778
rect 707 -5038 723 -4790
rect 757 -5038 773 -4790
rect 707 -5050 773 -5038
rect 803 -4790 869 -4778
rect 803 -5038 819 -4790
rect 853 -5038 869 -4790
rect 803 -5050 869 -5038
rect 899 -4790 965 -4778
rect 899 -5038 915 -4790
rect 949 -5038 965 -4790
rect 899 -5050 965 -5038
rect 995 -4790 1061 -4778
rect 995 -5038 1011 -4790
rect 1045 -5038 1061 -4790
rect 995 -5050 1061 -5038
rect 1091 -4790 1157 -4778
rect 1091 -5038 1107 -4790
rect 1141 -5038 1157 -4790
rect 1091 -5050 1157 -5038
rect 1187 -4790 1253 -4778
rect 1187 -5038 1203 -4790
rect 1237 -5038 1253 -4790
rect 1187 -5050 1253 -5038
rect 1283 -4790 1349 -4778
rect 1283 -5038 1299 -4790
rect 1333 -5038 1349 -4790
rect 1283 -5050 1349 -5038
rect 1379 -4790 1441 -4778
rect 1379 -5038 1395 -4790
rect 1429 -5038 1441 -4790
rect 1379 -5050 1441 -5038
rect 1944 -4790 2006 -4778
rect 1944 -5038 1956 -4790
rect 1990 -5038 2006 -4790
rect 1944 -5050 2006 -5038
rect 2036 -4790 2102 -4778
rect 2036 -5038 2052 -4790
rect 2086 -5038 2102 -4790
rect 2036 -5050 2102 -5038
rect 2132 -4790 2198 -4778
rect 2132 -5038 2148 -4790
rect 2182 -5038 2198 -4790
rect 2132 -5050 2198 -5038
rect 2228 -4790 2294 -4778
rect 2228 -5038 2244 -4790
rect 2278 -5038 2294 -4790
rect 2228 -5050 2294 -5038
rect 2324 -4790 2390 -4778
rect 2324 -5038 2340 -4790
rect 2374 -5038 2390 -4790
rect 2324 -5050 2390 -5038
rect 2420 -4790 2486 -4778
rect 2420 -5038 2436 -4790
rect 2470 -5038 2486 -4790
rect 2420 -5050 2486 -5038
rect 2516 -4790 2582 -4778
rect 2516 -5038 2532 -4790
rect 2566 -5038 2582 -4790
rect 2516 -5050 2582 -5038
rect 2612 -4790 2678 -4778
rect 2612 -5038 2628 -4790
rect 2662 -5038 2678 -4790
rect 2612 -5050 2678 -5038
rect 2708 -4790 2774 -4778
rect 2708 -5038 2724 -4790
rect 2758 -5038 2774 -4790
rect 2708 -5050 2774 -5038
rect 2804 -4790 2870 -4778
rect 2804 -5038 2820 -4790
rect 2854 -5038 2870 -4790
rect 2804 -5050 2870 -5038
rect 2900 -4790 2962 -4778
rect 2900 -5038 2916 -4790
rect 2950 -5038 2962 -4790
rect 2900 -5050 2962 -5038
<< ndiffc >>
rect 435 -370 469 -290
rect 531 -370 565 -290
rect 627 -370 661 -290
rect 723 -370 757 -290
rect 819 -370 853 -290
rect 915 -370 949 -290
rect 1011 -370 1045 -290
rect 1107 -370 1141 -290
rect 1203 -370 1237 -290
rect 1299 -370 1333 -290
rect 1395 -370 1429 -290
rect 1615 -372 1649 -296
rect 1703 -372 1737 -296
rect 1956 -370 1990 -290
rect 2052 -370 2086 -290
rect 2148 -370 2182 -290
rect 2244 -370 2278 -290
rect 2340 -370 2374 -290
rect 2436 -370 2470 -290
rect 2532 -370 2566 -290
rect 2628 -370 2662 -290
rect 2724 -370 2758 -290
rect 2820 -370 2854 -290
rect 2916 -370 2950 -290
rect -904 -574 -870 -540
rect -904 -642 -870 -608
rect -820 -574 -786 -540
rect -820 -642 -786 -608
rect -536 -574 -502 -540
rect -536 -642 -502 -608
rect -452 -574 -418 -540
rect -452 -642 -418 -608
rect -3116 -956 -3082 -876
rect -3020 -956 -2986 -876
rect -2924 -956 -2890 -876
rect -2828 -956 -2794 -876
rect -2732 -956 -2698 -876
rect -2636 -956 -2602 -876
rect -2540 -956 -2506 -876
rect -2444 -956 -2410 -876
rect -2348 -956 -2314 -876
rect -2252 -956 -2218 -876
rect -2156 -956 -2122 -876
rect -536 -1434 -502 -1400
rect -536 -1502 -502 -1468
rect -452 -1434 -418 -1400
rect -452 -1502 -418 -1468
rect -573 -1658 -539 -1624
rect -573 -1726 -539 -1692
rect -405 -1658 -371 -1624
rect -405 -1726 -371 -1692
rect 435 -1704 469 -1624
rect 531 -1704 565 -1624
rect 627 -1704 661 -1624
rect 723 -1704 757 -1624
rect 819 -1704 853 -1624
rect 915 -1704 949 -1624
rect 1011 -1704 1045 -1624
rect 1107 -1704 1141 -1624
rect 1203 -1704 1237 -1624
rect 1299 -1704 1333 -1624
rect 1395 -1704 1429 -1624
rect 1615 -1706 1649 -1630
rect 1703 -1706 1737 -1630
rect 1956 -1704 1990 -1624
rect 2052 -1704 2086 -1624
rect 2148 -1704 2182 -1624
rect 2244 -1704 2278 -1624
rect 2340 -1704 2374 -1624
rect 2436 -1704 2470 -1624
rect 2532 -1704 2566 -1624
rect 2628 -1704 2662 -1624
rect 2724 -1704 2758 -1624
rect 2820 -1704 2854 -1624
rect 2916 -1704 2950 -1624
rect -3116 -2290 -3082 -2210
rect -3020 -2290 -2986 -2210
rect -2924 -2290 -2890 -2210
rect -2828 -2290 -2794 -2210
rect -2732 -2290 -2698 -2210
rect -2636 -2290 -2602 -2210
rect -2540 -2290 -2506 -2210
rect -2444 -2290 -2410 -2210
rect -2348 -2290 -2314 -2210
rect -2252 -2290 -2218 -2210
rect -2156 -2290 -2122 -2210
rect -1088 -2522 -1054 -2488
rect -1088 -2590 -1054 -2556
rect -1004 -2522 -970 -2488
rect -1004 -2590 -970 -2556
rect -573 -2526 -539 -2492
rect -573 -2594 -539 -2560
rect -405 -2526 -371 -2492
rect -405 -2594 -371 -2560
rect -1088 -2750 -1054 -2716
rect -1088 -2818 -1054 -2784
rect -1004 -2750 -970 -2716
rect -1004 -2818 -970 -2784
rect -573 -2746 -539 -2712
rect -573 -2814 -539 -2780
rect -405 -2746 -371 -2712
rect -405 -2814 -371 -2780
rect 435 -3082 469 -3002
rect 531 -3082 565 -3002
rect 627 -3082 661 -3002
rect 723 -3082 757 -3002
rect 819 -3082 853 -3002
rect 915 -3082 949 -3002
rect 1011 -3082 1045 -3002
rect 1107 -3082 1141 -3002
rect 1203 -3082 1237 -3002
rect 1299 -3082 1333 -3002
rect 1395 -3082 1429 -3002
rect 1615 -3084 1649 -3008
rect 1703 -3084 1737 -3008
rect 1956 -3082 1990 -3002
rect 2052 -3082 2086 -3002
rect 2148 -3082 2182 -3002
rect 2244 -3082 2278 -3002
rect 2340 -3082 2374 -3002
rect 2436 -3082 2470 -3002
rect 2532 -3082 2566 -3002
rect 2628 -3082 2662 -3002
rect 2724 -3082 2758 -3002
rect 2820 -3082 2854 -3002
rect 2916 -3082 2950 -3002
rect -3116 -3668 -3082 -3588
rect -3020 -3668 -2986 -3588
rect -2924 -3668 -2890 -3588
rect -2828 -3668 -2794 -3588
rect -2732 -3668 -2698 -3588
rect -2636 -3668 -2602 -3588
rect -2540 -3668 -2506 -3588
rect -2444 -3668 -2410 -3588
rect -2348 -3668 -2314 -3588
rect -2252 -3668 -2218 -3588
rect -2156 -3668 -2122 -3588
rect -573 -3614 -539 -3580
rect -573 -3682 -539 -3648
rect -405 -3614 -371 -3580
rect -405 -3682 -371 -3648
rect -536 -3838 -502 -3804
rect -536 -3906 -502 -3872
rect -452 -3838 -418 -3804
rect -452 -3906 -418 -3872
rect 435 -4460 469 -4380
rect 531 -4460 565 -4380
rect 627 -4460 661 -4380
rect 723 -4460 757 -4380
rect 819 -4460 853 -4380
rect 915 -4460 949 -4380
rect 1011 -4460 1045 -4380
rect 1107 -4460 1141 -4380
rect 1203 -4460 1237 -4380
rect 1299 -4460 1333 -4380
rect 1395 -4460 1429 -4380
rect 1615 -4462 1649 -4386
rect 1703 -4462 1737 -4386
rect 1956 -4460 1990 -4380
rect 2052 -4460 2086 -4380
rect 2148 -4460 2182 -4380
rect 2244 -4460 2278 -4380
rect 2340 -4460 2374 -4380
rect 2436 -4460 2470 -4380
rect 2532 -4460 2566 -4380
rect 2628 -4460 2662 -4380
rect 2724 -4460 2758 -4380
rect 2820 -4460 2854 -4380
rect 2916 -4460 2950 -4380
rect -536 -4698 -502 -4664
rect -536 -4766 -502 -4732
rect -452 -4698 -418 -4664
rect -452 -4766 -418 -4732
rect -3116 -5046 -3082 -4966
rect -3020 -5046 -2986 -4966
rect -2924 -5046 -2890 -4966
rect -2828 -5046 -2794 -4966
rect -2732 -5046 -2698 -4966
rect -2636 -5046 -2602 -4966
rect -2540 -5046 -2506 -4966
rect -2444 -5046 -2410 -4966
rect -2348 -5046 -2314 -4966
rect -2252 -5046 -2218 -4966
rect -2156 -5046 -2122 -4966
<< pdiffc >>
rect -3116 -546 -3082 -298
rect -3020 -546 -2986 -298
rect -2924 -546 -2890 -298
rect -2828 -546 -2794 -298
rect -2732 -546 -2698 -298
rect -2636 -546 -2602 -298
rect -2540 -546 -2506 -298
rect -2444 -546 -2410 -298
rect -2348 -546 -2314 -298
rect -2252 -546 -2218 -298
rect -2156 -546 -2122 -298
rect -904 -826 -870 -792
rect -904 -894 -870 -860
rect -904 -962 -870 -928
rect -820 -826 -786 -792
rect -820 -894 -786 -860
rect -820 -962 -786 -928
rect -536 -826 -502 -792
rect -536 -894 -502 -860
rect -536 -962 -502 -928
rect -452 -826 -418 -792
rect -452 -894 -418 -860
rect -452 -962 -418 -928
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect -536 -1114 -502 -1080
rect -536 -1182 -502 -1148
rect -536 -1250 -502 -1216
rect -452 -1114 -418 -1080
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect -452 -1182 -418 -1148
rect -452 -1250 -418 -1216
rect -3116 -1880 -3082 -1632
rect -3020 -1880 -2986 -1632
rect -2924 -1880 -2890 -1632
rect -2828 -1880 -2794 -1632
rect -2732 -1880 -2698 -1632
rect -2636 -1880 -2602 -1632
rect -2540 -1880 -2506 -1632
rect -2444 -1880 -2410 -1632
rect -2348 -1880 -2314 -1632
rect -2252 -1880 -2218 -1632
rect -2156 -1880 -2122 -1632
rect -573 -1914 -539 -1880
rect -573 -1982 -539 -1948
rect -573 -2050 -539 -2016
rect -489 -1914 -455 -1880
rect -489 -1982 -455 -1948
rect -489 -2050 -455 -2016
rect -405 -1914 -371 -1880
rect -405 -1982 -371 -1948
rect -405 -2050 -371 -2016
rect -1088 -2202 -1054 -2168
rect -1088 -2270 -1054 -2236
rect -1088 -2338 -1054 -2304
rect -1004 -2202 -970 -2168
rect -1004 -2270 -970 -2236
rect -1004 -2338 -970 -2304
rect -573 -2202 -539 -2168
rect -573 -2270 -539 -2236
rect -573 -2338 -539 -2304
rect -489 -2202 -455 -2168
rect -489 -2270 -455 -2236
rect -489 -2338 -455 -2304
rect -405 -2202 -371 -2168
rect -405 -2270 -371 -2236
rect -405 -2338 -371 -2304
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
rect -3116 -3258 -3082 -3010
rect -3020 -3258 -2986 -3010
rect -2924 -3258 -2890 -3010
rect -2828 -3258 -2794 -3010
rect -2732 -3258 -2698 -3010
rect -2636 -3258 -2602 -3010
rect -2540 -3258 -2506 -3010
rect -2444 -3258 -2410 -3010
rect -2348 -3258 -2314 -3010
rect -2252 -3258 -2218 -3010
rect -2156 -3258 -2122 -3010
rect -1088 -3002 -1054 -2968
rect -1088 -3070 -1054 -3036
rect -1088 -3138 -1054 -3104
rect -1004 -3002 -970 -2968
rect -1004 -3070 -970 -3036
rect -1004 -3138 -970 -3104
rect -573 -3002 -539 -2968
rect -573 -3070 -539 -3036
rect -573 -3138 -539 -3104
rect -489 -3002 -455 -2968
rect -489 -3070 -455 -3036
rect -489 -3138 -455 -3104
rect -405 -3002 -371 -2968
rect -405 -3070 -371 -3036
rect -405 -3138 -371 -3104
rect -573 -3290 -539 -3256
rect -573 -3358 -539 -3324
rect -573 -3426 -539 -3392
rect -489 -3290 -455 -3256
rect -489 -3358 -455 -3324
rect -489 -3426 -455 -3392
rect -405 -3290 -371 -3256
rect -405 -3358 -371 -3324
rect -405 -3426 -371 -3392
rect 435 -3660 469 -3412
rect 531 -3660 565 -3412
rect 627 -3660 661 -3412
rect 723 -3660 757 -3412
rect 819 -3660 853 -3412
rect 915 -3660 949 -3412
rect 1011 -3660 1045 -3412
rect 1107 -3660 1141 -3412
rect 1203 -3660 1237 -3412
rect 1299 -3660 1333 -3412
rect 1395 -3660 1429 -3412
rect 1956 -3660 1990 -3412
rect 2052 -3660 2086 -3412
rect 2148 -3660 2182 -3412
rect 2244 -3660 2278 -3412
rect 2340 -3660 2374 -3412
rect 2436 -3660 2470 -3412
rect 2532 -3660 2566 -3412
rect 2628 -3660 2662 -3412
rect 2724 -3660 2758 -3412
rect 2820 -3660 2854 -3412
rect 2916 -3660 2950 -3412
rect -536 -4090 -502 -4056
rect -536 -4158 -502 -4124
rect -536 -4226 -502 -4192
rect -452 -4090 -418 -4056
rect -452 -4158 -418 -4124
rect -452 -4226 -418 -4192
rect -3116 -4636 -3082 -4388
rect -3020 -4636 -2986 -4388
rect -2924 -4636 -2890 -4388
rect -2828 -4636 -2794 -4388
rect -2732 -4636 -2698 -4388
rect -2636 -4636 -2602 -4388
rect -2540 -4636 -2506 -4388
rect -2444 -4636 -2410 -4388
rect -2348 -4636 -2314 -4388
rect -2252 -4636 -2218 -4388
rect -2156 -4636 -2122 -4388
rect -536 -4378 -502 -4344
rect -536 -4446 -502 -4412
rect -536 -4514 -502 -4480
rect -452 -4378 -418 -4344
rect -452 -4446 -418 -4412
rect -452 -4514 -418 -4480
rect 435 -5038 469 -4790
rect 531 -5038 565 -4790
rect 627 -5038 661 -4790
rect 723 -5038 757 -4790
rect 819 -5038 853 -4790
rect 915 -5038 949 -4790
rect 1011 -5038 1045 -4790
rect 1107 -5038 1141 -4790
rect 1203 -5038 1237 -4790
rect 1299 -5038 1333 -4790
rect 1395 -5038 1429 -4790
rect 1956 -5038 1990 -4790
rect 2052 -5038 2086 -4790
rect 2148 -5038 2182 -4790
rect 2244 -5038 2278 -4790
rect 2340 -5038 2374 -4790
rect 2436 -5038 2470 -4790
rect 2532 -5038 2566 -4790
rect 2628 -5038 2662 -4790
rect 2724 -5038 2758 -4790
rect 2820 -5038 2854 -4790
rect 2916 -5038 2950 -4790
<< psubdiff >>
rect 321 -138 417 -104
rect 1447 -138 1543 -104
rect 321 -200 355 -138
rect 1509 -200 1543 -138
rect 321 -460 355 -398
rect 1842 -138 1938 -104
rect 2968 -138 3064 -104
rect 1842 -200 1876 -138
rect 1509 -460 1543 -398
rect 3030 -200 3064 -138
rect 321 -494 417 -460
rect 1447 -494 1543 -460
rect 1842 -460 1876 -398
rect 3030 -460 3064 -398
rect 1842 -494 1938 -460
rect 2968 -494 3064 -460
rect -675 -588 -641 -541
rect -675 -646 -641 -622
rect -3230 -786 -3134 -752
rect -2104 -786 -2008 -752
rect -3230 -848 -3196 -786
rect -2042 -848 -2008 -786
rect -3230 -1108 -3196 -1046
rect -2042 -1108 -2008 -1046
rect -3230 -1142 -3134 -1108
rect -2104 -1142 -2008 -1108
rect -675 -1420 -641 -1396
rect -675 -1501 -641 -1454
rect 321 -1472 417 -1438
rect 1447 -1472 1543 -1438
rect 321 -1534 355 -1472
rect -675 -1676 -641 -1629
rect -675 -1734 -641 -1710
rect 1509 -1534 1543 -1472
rect 321 -1794 355 -1732
rect 1842 -1472 1938 -1438
rect 2968 -1472 3064 -1438
rect 1842 -1534 1876 -1472
rect 1509 -1794 1543 -1732
rect 3030 -1534 3064 -1472
rect 321 -1828 417 -1794
rect 1447 -1828 1543 -1794
rect 1842 -1794 1876 -1732
rect 3030 -1794 3064 -1732
rect 1842 -1828 1938 -1794
rect 2968 -1828 3064 -1794
rect -3230 -2120 -3134 -2086
rect -2104 -2120 -2008 -2086
rect -3230 -2182 -3196 -2120
rect -2042 -2182 -2008 -2120
rect -3230 -2442 -3196 -2380
rect -2042 -2442 -2008 -2380
rect -3230 -2476 -3134 -2442
rect -2104 -2476 -2008 -2442
rect -1227 -2508 -1193 -2484
rect -1227 -2589 -1193 -2542
rect -675 -2508 -641 -2484
rect -675 -2589 -641 -2542
rect -1227 -2764 -1193 -2717
rect -1227 -2822 -1193 -2798
rect -675 -2764 -641 -2717
rect -675 -2822 -641 -2798
rect 321 -2850 417 -2816
rect 1447 -2850 1543 -2816
rect 321 -2912 355 -2850
rect 1509 -2912 1543 -2850
rect 321 -3172 355 -3110
rect 1842 -2850 1938 -2816
rect 2968 -2850 3064 -2816
rect 1842 -2912 1876 -2850
rect 1509 -3172 1543 -3110
rect 3030 -2912 3064 -2850
rect 321 -3206 417 -3172
rect 1447 -3206 1543 -3172
rect 1842 -3172 1876 -3110
rect 3030 -3172 3064 -3110
rect 1842 -3206 1938 -3172
rect 2968 -3206 3064 -3172
rect -3230 -3498 -3134 -3464
rect -2104 -3498 -2008 -3464
rect -3230 -3560 -3196 -3498
rect -2042 -3560 -2008 -3498
rect -3230 -3820 -3196 -3758
rect -675 -3596 -641 -3572
rect -675 -3677 -641 -3630
rect -2042 -3820 -2008 -3758
rect -3230 -3854 -3134 -3820
rect -2104 -3854 -2008 -3820
rect -675 -3852 -641 -3805
rect -675 -3910 -641 -3886
rect 321 -4228 417 -4194
rect 1447 -4228 1543 -4194
rect 321 -4290 355 -4228
rect 1509 -4290 1543 -4228
rect 321 -4550 355 -4488
rect 1842 -4228 1938 -4194
rect 2968 -4228 3064 -4194
rect 1842 -4290 1876 -4228
rect 1509 -4550 1543 -4488
rect 3030 -4290 3064 -4228
rect 321 -4584 417 -4550
rect 1447 -4584 1543 -4550
rect 1842 -4550 1876 -4488
rect 3030 -4550 3064 -4488
rect 1842 -4584 1938 -4550
rect 2968 -4584 3064 -4550
rect -675 -4684 -641 -4660
rect -675 -4765 -641 -4718
rect -3230 -4876 -3134 -4842
rect -2104 -4876 -2008 -4842
rect -3230 -4938 -3196 -4876
rect -2042 -4938 -2008 -4876
rect -3230 -5198 -3196 -5136
rect -2042 -5198 -2008 -5136
rect -3230 -5232 -3134 -5198
rect -2104 -5232 -2008 -5198
<< nsubdiff >>
rect -3230 -136 -3134 -102
rect -2104 -136 -2008 -102
rect -3230 -198 -3196 -136
rect -2042 -198 -2008 -136
rect -3230 -646 -3196 -584
rect -2042 -646 -2008 -584
rect -3230 -680 -3134 -646
rect -2104 -680 -2008 -646
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect 1509 -662 1543 -600
rect -675 -806 -641 -782
rect -675 -899 -641 -840
rect -675 -957 -641 -933
rect -675 -1109 -641 -1085
rect -675 -1202 -641 -1143
rect -675 -1260 -641 -1236
rect 321 -1110 355 -1048
rect 1509 -1110 1543 -1048
rect 321 -1144 417 -1110
rect 1447 -1144 1543 -1110
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1842 -1110 1876 -1048
rect 3030 -1110 3064 -1048
rect 1842 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect -3230 -1470 -3134 -1436
rect -2104 -1470 -2008 -1436
rect -3230 -1532 -3196 -1470
rect -2042 -1532 -2008 -1470
rect -3230 -1980 -3196 -1918
rect -2042 -1980 -2008 -1918
rect -3230 -2014 -3134 -1980
rect -2104 -2014 -2008 -1980
rect -675 -1894 -641 -1870
rect -675 -1987 -641 -1928
rect -675 -2045 -641 -2021
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect -1227 -2197 -1193 -2173
rect -1227 -2290 -1193 -2231
rect -1227 -2348 -1193 -2324
rect -675 -2197 -641 -2173
rect -675 -2290 -641 -2231
rect -675 -2348 -641 -2324
rect 321 -2444 355 -2382
rect 1509 -2444 1543 -2382
rect 321 -2478 417 -2444
rect 1447 -2478 1543 -2444
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1842 -2444 1876 -2382
rect 3030 -2444 3064 -2382
rect 1842 -2478 1938 -2444
rect 2968 -2478 3064 -2444
rect -3230 -2848 -3134 -2814
rect -2104 -2848 -2008 -2814
rect -3230 -2910 -3196 -2848
rect -2042 -2910 -2008 -2848
rect -1227 -2982 -1193 -2958
rect -1227 -3075 -1193 -3016
rect -1227 -3133 -1193 -3109
rect -675 -2982 -641 -2958
rect -675 -3075 -641 -3016
rect -675 -3133 -641 -3109
rect -3230 -3358 -3196 -3296
rect -2042 -3358 -2008 -3296
rect -3230 -3392 -3134 -3358
rect -2104 -3392 -2008 -3358
rect -675 -3285 -641 -3261
rect -675 -3378 -641 -3319
rect -675 -3436 -641 -3412
rect 321 -3312 417 -3278
rect 1447 -3312 1543 -3278
rect 321 -3374 355 -3312
rect 1509 -3374 1543 -3312
rect 321 -3822 355 -3760
rect 1509 -3822 1543 -3760
rect 321 -3856 417 -3822
rect 1447 -3856 1543 -3822
rect 1842 -3312 1938 -3278
rect 2968 -3312 3064 -3278
rect 1842 -3374 1876 -3312
rect 3030 -3374 3064 -3312
rect 1842 -3822 1876 -3760
rect 3030 -3822 3064 -3760
rect 1842 -3856 1938 -3822
rect 2968 -3856 3064 -3822
rect -675 -4070 -641 -4046
rect -675 -4163 -641 -4104
rect -3230 -4226 -3134 -4192
rect -2104 -4226 -2008 -4192
rect -675 -4221 -641 -4197
rect -3230 -4288 -3196 -4226
rect -2042 -4288 -2008 -4226
rect -675 -4373 -641 -4349
rect -675 -4466 -641 -4407
rect -675 -4524 -641 -4500
rect -3230 -4736 -3196 -4674
rect -2042 -4736 -2008 -4674
rect -3230 -4770 -3134 -4736
rect -2104 -4770 -2008 -4736
rect 321 -4690 417 -4656
rect 1447 -4690 1543 -4656
rect 321 -4752 355 -4690
rect 1509 -4752 1543 -4690
rect 321 -5200 355 -5138
rect 1509 -5200 1543 -5138
rect 321 -5234 417 -5200
rect 1447 -5234 1543 -5200
rect 1842 -4690 1938 -4656
rect 2968 -4690 3064 -4656
rect 1842 -4752 1876 -4690
rect 3030 -4752 3064 -4690
rect 1842 -5200 1876 -5138
rect 3030 -5200 3064 -5138
rect 1842 -5234 1938 -5200
rect 2968 -5234 3064 -5200
<< psubdiffcont >>
rect 417 -138 1447 -104
rect 321 -398 355 -200
rect 1509 -398 1543 -200
rect 1938 -138 2968 -104
rect 1842 -398 1876 -200
rect 417 -494 1447 -460
rect 3030 -398 3064 -200
rect 1938 -494 2968 -460
rect -675 -622 -641 -588
rect -3134 -786 -2104 -752
rect -3230 -1046 -3196 -848
rect -2042 -1046 -2008 -848
rect -3134 -1142 -2104 -1108
rect -675 -1454 -641 -1420
rect 417 -1472 1447 -1438
rect -675 -1710 -641 -1676
rect 321 -1732 355 -1534
rect 1509 -1732 1543 -1534
rect 1938 -1472 2968 -1438
rect 1842 -1732 1876 -1534
rect 417 -1828 1447 -1794
rect 3030 -1732 3064 -1534
rect 1938 -1828 2968 -1794
rect -3134 -2120 -2104 -2086
rect -3230 -2380 -3196 -2182
rect -2042 -2380 -2008 -2182
rect -3134 -2476 -2104 -2442
rect -1227 -2542 -1193 -2508
rect -675 -2542 -641 -2508
rect -1227 -2798 -1193 -2764
rect -675 -2798 -641 -2764
rect 417 -2850 1447 -2816
rect 321 -3110 355 -2912
rect 1509 -3110 1543 -2912
rect 1938 -2850 2968 -2816
rect 1842 -3110 1876 -2912
rect 417 -3206 1447 -3172
rect 3030 -3110 3064 -2912
rect 1938 -3206 2968 -3172
rect -3134 -3498 -2104 -3464
rect -3230 -3758 -3196 -3560
rect -2042 -3758 -2008 -3560
rect -675 -3630 -641 -3596
rect -3134 -3854 -2104 -3820
rect -675 -3886 -641 -3852
rect 417 -4228 1447 -4194
rect 321 -4488 355 -4290
rect 1509 -4488 1543 -4290
rect 1938 -4228 2968 -4194
rect 1842 -4488 1876 -4290
rect 417 -4584 1447 -4550
rect 3030 -4488 3064 -4290
rect 1938 -4584 2968 -4550
rect -675 -4718 -641 -4684
rect -3134 -4876 -2104 -4842
rect -3230 -5136 -3196 -4938
rect -2042 -5136 -2008 -4938
rect -3134 -5232 -2104 -5198
<< nsubdiffcont >>
rect -3134 -136 -2104 -102
rect -3230 -584 -3196 -198
rect -2042 -584 -2008 -198
rect -3134 -680 -2104 -646
rect 417 -600 1447 -566
rect -675 -840 -641 -806
rect -675 -933 -641 -899
rect 321 -1048 355 -662
rect -675 -1143 -641 -1109
rect -675 -1236 -641 -1202
rect 1509 -1048 1543 -662
rect 417 -1144 1447 -1110
rect 1938 -600 2968 -566
rect 1842 -1048 1876 -662
rect 3030 -1048 3064 -662
rect 1938 -1144 2968 -1110
rect -3134 -1470 -2104 -1436
rect -3230 -1918 -3196 -1532
rect -2042 -1918 -2008 -1532
rect -3134 -2014 -2104 -1980
rect -675 -1928 -641 -1894
rect -675 -2021 -641 -1987
rect 417 -1934 1447 -1900
rect -1227 -2231 -1193 -2197
rect -1227 -2324 -1193 -2290
rect -675 -2231 -641 -2197
rect -675 -2324 -641 -2290
rect 321 -2382 355 -1996
rect 1509 -2382 1543 -1996
rect 417 -2478 1447 -2444
rect 1938 -1934 2968 -1900
rect 1842 -2382 1876 -1996
rect 3030 -2382 3064 -1996
rect 1938 -2478 2968 -2444
rect -3134 -2848 -2104 -2814
rect -3230 -3296 -3196 -2910
rect -2042 -3296 -2008 -2910
rect -1227 -3016 -1193 -2982
rect -1227 -3109 -1193 -3075
rect -675 -3016 -641 -2982
rect -675 -3109 -641 -3075
rect -3134 -3392 -2104 -3358
rect -675 -3319 -641 -3285
rect -675 -3412 -641 -3378
rect 417 -3312 1447 -3278
rect 321 -3760 355 -3374
rect 1509 -3760 1543 -3374
rect 417 -3856 1447 -3822
rect 1938 -3312 2968 -3278
rect 1842 -3760 1876 -3374
rect 3030 -3760 3064 -3374
rect 1938 -3856 2968 -3822
rect -675 -4104 -641 -4070
rect -3134 -4226 -2104 -4192
rect -675 -4197 -641 -4163
rect -3230 -4674 -3196 -4288
rect -2042 -4674 -2008 -4288
rect -675 -4407 -641 -4373
rect -675 -4500 -641 -4466
rect -3134 -4770 -2104 -4736
rect 417 -4690 1447 -4656
rect 321 -5138 355 -4752
rect 1509 -5138 1543 -4752
rect 417 -5234 1447 -5200
rect 1938 -4690 2968 -4656
rect 1842 -5138 1876 -4752
rect 3030 -5138 3064 -4752
rect 1938 -5234 2968 -5200
<< poly >>
rect -3132 -204 -2106 -188
rect -3132 -238 -3116 -204
rect -3082 -238 -2924 -204
rect -2890 -238 -2732 -204
rect -2698 -238 -2540 -204
rect -2506 -238 -2348 -204
rect -2314 -238 -2156 -204
rect -2122 -238 -2106 -204
rect -3132 -254 -2106 -238
rect -3066 -286 -3036 -254
rect -2970 -286 -2940 -254
rect -2874 -286 -2844 -254
rect -2778 -286 -2748 -254
rect -2682 -286 -2652 -254
rect -2586 -286 -2556 -254
rect -2490 -286 -2460 -254
rect -2394 -286 -2364 -254
rect -2298 -286 -2268 -254
rect -2202 -286 -2172 -254
rect -3066 -584 -3036 -558
rect -2970 -584 -2940 -558
rect -2874 -584 -2844 -558
rect -2778 -584 -2748 -558
rect -2682 -584 -2652 -558
rect -2586 -584 -2556 -558
rect -2490 -584 -2460 -558
rect -2394 -584 -2364 -558
rect -2298 -584 -2268 -558
rect -2202 -584 -2172 -558
rect 419 -197 1445 -181
rect 419 -231 435 -197
rect 469 -231 627 -197
rect 661 -231 819 -197
rect 853 -231 1011 -197
rect 1045 -231 1203 -197
rect 1237 -231 1395 -197
rect 1429 -231 1445 -197
rect 419 -247 1445 -231
rect 485 -278 515 -247
rect 581 -278 611 -247
rect 677 -278 707 -247
rect 773 -278 803 -247
rect 869 -278 899 -247
rect 965 -278 995 -247
rect 1061 -278 1091 -247
rect 1157 -278 1187 -247
rect 1253 -278 1283 -247
rect 1349 -278 1379 -247
rect 485 -408 515 -382
rect 581 -408 611 -382
rect 677 -408 707 -382
rect 773 -408 803 -382
rect 869 -408 899 -382
rect 965 -408 995 -382
rect 1061 -408 1091 -382
rect 1157 -408 1187 -382
rect 1253 -408 1283 -382
rect 1349 -408 1379 -382
rect 1661 -284 1691 -258
rect 1661 -406 1691 -384
rect 1940 -197 2966 -181
rect 1940 -231 1956 -197
rect 1990 -231 2148 -197
rect 2182 -231 2340 -197
rect 2374 -231 2532 -197
rect 2566 -231 2724 -197
rect 2758 -231 2916 -197
rect 2950 -231 2966 -197
rect 1940 -247 2966 -231
rect 2006 -278 2036 -247
rect 2102 -278 2132 -247
rect 2198 -278 2228 -247
rect 2294 -278 2324 -247
rect 2390 -278 2420 -247
rect 2486 -278 2516 -247
rect 2582 -278 2612 -247
rect 2678 -278 2708 -247
rect 2774 -278 2804 -247
rect 2870 -278 2900 -247
rect 1643 -422 1709 -406
rect 1643 -456 1659 -422
rect 1693 -456 1709 -422
rect 1643 -472 1709 -456
rect 2006 -408 2036 -382
rect 2102 -408 2132 -382
rect 2198 -408 2228 -382
rect 2294 -408 2324 -382
rect 2390 -408 2420 -382
rect 2486 -408 2516 -382
rect 2582 -408 2612 -382
rect 2678 -408 2708 -382
rect 2774 -408 2804 -382
rect 2870 -408 2900 -382
rect -860 -524 -830 -498
rect -492 -524 -462 -498
rect -860 -676 -830 -654
rect -492 -676 -462 -654
rect -916 -692 -830 -676
rect -916 -726 -900 -692
rect -866 -726 -830 -692
rect -916 -742 -830 -726
rect -548 -692 -462 -676
rect -548 -726 -532 -692
rect -498 -726 -462 -692
rect -548 -742 -462 -726
rect -860 -774 -830 -742
rect -492 -774 -462 -742
rect -3066 -864 -3036 -838
rect -2970 -864 -2940 -838
rect -2874 -864 -2844 -838
rect -2778 -864 -2748 -838
rect -2682 -864 -2652 -838
rect -2586 -864 -2556 -838
rect -2490 -864 -2460 -838
rect -2394 -864 -2364 -838
rect -2298 -864 -2268 -838
rect -2202 -864 -2172 -838
rect -3066 -999 -3036 -968
rect -2970 -999 -2940 -968
rect -2874 -999 -2844 -968
rect -2778 -999 -2748 -968
rect -2682 -999 -2652 -968
rect -2586 -999 -2556 -968
rect -2490 -999 -2460 -968
rect -2394 -999 -2364 -968
rect -2298 -999 -2268 -968
rect -2202 -999 -2172 -968
rect -3132 -1015 -2106 -999
rect -3132 -1049 -3116 -1015
rect -3082 -1049 -2924 -1015
rect -2890 -1049 -2732 -1015
rect -2698 -1049 -2540 -1015
rect -2506 -1049 -2348 -1015
rect -2314 -1049 -2156 -1015
rect -2122 -1049 -2106 -1015
rect -3132 -1065 -2106 -1049
rect -860 -1000 -830 -974
rect -492 -1000 -462 -974
rect -492 -1068 -462 -1042
rect 485 -688 515 -662
rect 581 -688 611 -662
rect 677 -688 707 -662
rect 773 -688 803 -662
rect 869 -688 899 -662
rect 965 -688 995 -662
rect 1061 -688 1091 -662
rect 1157 -688 1187 -662
rect 1253 -688 1283 -662
rect 1349 -688 1379 -662
rect 485 -992 515 -960
rect 581 -992 611 -960
rect 677 -992 707 -960
rect 773 -992 803 -960
rect 869 -992 899 -960
rect 965 -992 995 -960
rect 1061 -992 1091 -960
rect 1157 -992 1187 -960
rect 1253 -992 1283 -960
rect 1349 -992 1379 -960
rect 419 -1008 1445 -992
rect 419 -1042 435 -1008
rect 469 -1042 627 -1008
rect 661 -1042 819 -1008
rect 853 -1042 1011 -1008
rect 1045 -1042 1203 -1008
rect 1237 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 419 -1058 1445 -1042
rect 2006 -688 2036 -662
rect 2102 -688 2132 -662
rect 2198 -688 2228 -662
rect 2294 -688 2324 -662
rect 2390 -688 2420 -662
rect 2486 -688 2516 -662
rect 2582 -688 2612 -662
rect 2678 -688 2708 -662
rect 2774 -688 2804 -662
rect 2870 -688 2900 -662
rect 2006 -992 2036 -960
rect 2102 -992 2132 -960
rect 2198 -992 2228 -960
rect 2294 -992 2324 -960
rect 2390 -992 2420 -960
rect 2486 -992 2516 -960
rect 2582 -992 2612 -960
rect 2678 -992 2708 -960
rect 2774 -992 2804 -960
rect 2870 -992 2900 -960
rect 1940 -1008 2966 -992
rect 1940 -1042 1956 -1008
rect 1990 -1042 2148 -1008
rect 2182 -1042 2340 -1008
rect 2374 -1042 2532 -1008
rect 2566 -1042 2724 -1008
rect 2758 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1940 -1058 2966 -1042
rect -492 -1300 -462 -1268
rect -548 -1316 -462 -1300
rect -548 -1350 -532 -1316
rect -498 -1350 -462 -1316
rect -548 -1366 -462 -1350
rect -492 -1388 -462 -1366
rect -3132 -1538 -2106 -1522
rect -3132 -1572 -3116 -1538
rect -3082 -1572 -2924 -1538
rect -2890 -1572 -2732 -1538
rect -2698 -1572 -2540 -1538
rect -2506 -1572 -2348 -1538
rect -2314 -1572 -2156 -1538
rect -2122 -1572 -2106 -1538
rect -3132 -1588 -2106 -1572
rect -3066 -1620 -3036 -1588
rect -2970 -1620 -2940 -1588
rect -2874 -1620 -2844 -1588
rect -2778 -1620 -2748 -1588
rect -2682 -1620 -2652 -1588
rect -2586 -1620 -2556 -1588
rect -2490 -1620 -2460 -1588
rect -2394 -1620 -2364 -1588
rect -2298 -1620 -2268 -1588
rect -2202 -1620 -2172 -1588
rect -3066 -1918 -3036 -1892
rect -2970 -1918 -2940 -1892
rect -2874 -1918 -2844 -1892
rect -2778 -1918 -2748 -1892
rect -2682 -1918 -2652 -1892
rect -2586 -1918 -2556 -1892
rect -2490 -1918 -2460 -1892
rect -2394 -1918 -2364 -1892
rect -2298 -1918 -2268 -1892
rect -2202 -1918 -2172 -1892
rect -492 -1544 -462 -1518
rect -529 -1612 -499 -1586
rect -445 -1612 -415 -1586
rect 419 -1531 1445 -1515
rect 419 -1565 435 -1531
rect 469 -1565 627 -1531
rect 661 -1565 819 -1531
rect 853 -1565 1011 -1531
rect 1045 -1565 1203 -1531
rect 1237 -1565 1395 -1531
rect 1429 -1565 1445 -1531
rect 419 -1581 1445 -1565
rect 485 -1612 515 -1581
rect 581 -1612 611 -1581
rect 677 -1612 707 -1581
rect 773 -1612 803 -1581
rect 869 -1612 899 -1581
rect 965 -1612 995 -1581
rect 1061 -1612 1091 -1581
rect 1157 -1612 1187 -1581
rect 1253 -1612 1283 -1581
rect 1349 -1612 1379 -1581
rect -529 -1764 -499 -1742
rect -591 -1780 -499 -1764
rect -591 -1814 -576 -1780
rect -542 -1814 -499 -1780
rect -591 -1830 -499 -1814
rect -529 -1862 -499 -1830
rect -445 -1764 -415 -1742
rect -445 -1780 -357 -1764
rect -445 -1814 -408 -1780
rect -374 -1814 -357 -1780
rect -445 -1830 -357 -1814
rect 485 -1742 515 -1716
rect 581 -1742 611 -1716
rect 677 -1742 707 -1716
rect 773 -1742 803 -1716
rect 869 -1742 899 -1716
rect 965 -1742 995 -1716
rect 1061 -1742 1091 -1716
rect 1157 -1742 1187 -1716
rect 1253 -1742 1283 -1716
rect 1349 -1742 1379 -1716
rect 1661 -1618 1691 -1592
rect 1661 -1740 1691 -1718
rect 1940 -1531 2966 -1515
rect 1940 -1565 1956 -1531
rect 1990 -1565 2148 -1531
rect 2182 -1565 2340 -1531
rect 2374 -1565 2532 -1531
rect 2566 -1565 2724 -1531
rect 2758 -1565 2916 -1531
rect 2950 -1565 2966 -1531
rect 1940 -1581 2966 -1565
rect 2006 -1612 2036 -1581
rect 2102 -1612 2132 -1581
rect 2198 -1612 2228 -1581
rect 2294 -1612 2324 -1581
rect 2390 -1612 2420 -1581
rect 2486 -1612 2516 -1581
rect 2582 -1612 2612 -1581
rect 2678 -1612 2708 -1581
rect 2774 -1612 2804 -1581
rect 2870 -1612 2900 -1581
rect 1643 -1756 1709 -1740
rect 1643 -1790 1659 -1756
rect 1693 -1790 1709 -1756
rect 1643 -1806 1709 -1790
rect 2006 -1742 2036 -1716
rect 2102 -1742 2132 -1716
rect 2198 -1742 2228 -1716
rect 2294 -1742 2324 -1716
rect 2390 -1742 2420 -1716
rect 2486 -1742 2516 -1716
rect 2582 -1742 2612 -1716
rect 2678 -1742 2708 -1716
rect 2774 -1742 2804 -1716
rect 2870 -1742 2900 -1716
rect -445 -1862 -415 -1830
rect -529 -2088 -499 -2062
rect -445 -2088 -415 -2062
rect -3066 -2198 -3036 -2172
rect -2970 -2198 -2940 -2172
rect -2874 -2198 -2844 -2172
rect -2778 -2198 -2748 -2172
rect -2682 -2198 -2652 -2172
rect -2586 -2198 -2556 -2172
rect -2490 -2198 -2460 -2172
rect -2394 -2198 -2364 -2172
rect -2298 -2198 -2268 -2172
rect -2202 -2198 -2172 -2172
rect -1044 -2156 -1014 -2130
rect -529 -2156 -499 -2130
rect -445 -2156 -415 -2130
rect -3066 -2333 -3036 -2302
rect -2970 -2333 -2940 -2302
rect -2874 -2333 -2844 -2302
rect -2778 -2333 -2748 -2302
rect -2682 -2333 -2652 -2302
rect -2586 -2333 -2556 -2302
rect -2490 -2333 -2460 -2302
rect -2394 -2333 -2364 -2302
rect -2298 -2333 -2268 -2302
rect -2202 -2333 -2172 -2302
rect -3132 -2349 -2106 -2333
rect -3132 -2383 -3116 -2349
rect -3082 -2383 -2924 -2349
rect -2890 -2383 -2732 -2349
rect -2698 -2383 -2540 -2349
rect -2506 -2383 -2348 -2349
rect -2314 -2383 -2156 -2349
rect -2122 -2383 -2106 -2349
rect -3132 -2399 -2106 -2383
rect -1044 -2388 -1014 -2356
rect -529 -2388 -499 -2356
rect -1100 -2404 -1014 -2388
rect -1100 -2438 -1084 -2404
rect -1050 -2438 -1014 -2404
rect -1100 -2454 -1014 -2438
rect -591 -2404 -499 -2388
rect -591 -2438 -576 -2404
rect -542 -2438 -499 -2404
rect -591 -2454 -499 -2438
rect -1044 -2476 -1014 -2454
rect -529 -2476 -499 -2454
rect -445 -2388 -415 -2356
rect 485 -2022 515 -1996
rect 581 -2022 611 -1996
rect 677 -2022 707 -1996
rect 773 -2022 803 -1996
rect 869 -2022 899 -1996
rect 965 -2022 995 -1996
rect 1061 -2022 1091 -1996
rect 1157 -2022 1187 -1996
rect 1253 -2022 1283 -1996
rect 1349 -2022 1379 -1996
rect 485 -2326 515 -2294
rect 581 -2326 611 -2294
rect 677 -2326 707 -2294
rect 773 -2326 803 -2294
rect 869 -2326 899 -2294
rect 965 -2326 995 -2294
rect 1061 -2326 1091 -2294
rect 1157 -2326 1187 -2294
rect 1253 -2326 1283 -2294
rect 1349 -2326 1379 -2294
rect -445 -2404 -357 -2388
rect -445 -2438 -408 -2404
rect -374 -2438 -357 -2404
rect -445 -2454 -357 -2438
rect 419 -2342 1445 -2326
rect 419 -2376 435 -2342
rect 469 -2376 627 -2342
rect 661 -2376 819 -2342
rect 853 -2376 1011 -2342
rect 1045 -2376 1203 -2342
rect 1237 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 419 -2392 1445 -2376
rect -445 -2476 -415 -2454
rect 2006 -2022 2036 -1996
rect 2102 -2022 2132 -1996
rect 2198 -2022 2228 -1996
rect 2294 -2022 2324 -1996
rect 2390 -2022 2420 -1996
rect 2486 -2022 2516 -1996
rect 2582 -2022 2612 -1996
rect 2678 -2022 2708 -1996
rect 2774 -2022 2804 -1996
rect 2870 -2022 2900 -1996
rect 2006 -2326 2036 -2294
rect 2102 -2326 2132 -2294
rect 2198 -2326 2228 -2294
rect 2294 -2326 2324 -2294
rect 2390 -2326 2420 -2294
rect 2486 -2326 2516 -2294
rect 2582 -2326 2612 -2294
rect 2678 -2326 2708 -2294
rect 2774 -2326 2804 -2294
rect 2870 -2326 2900 -2294
rect 1940 -2342 2966 -2326
rect 1940 -2376 1956 -2342
rect 1990 -2376 2148 -2342
rect 2182 -2376 2340 -2342
rect 2374 -2376 2532 -2342
rect 2566 -2376 2724 -2342
rect 2758 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1940 -2392 2966 -2376
rect -1044 -2632 -1014 -2606
rect -529 -2632 -499 -2606
rect -445 -2632 -415 -2606
rect -1044 -2700 -1014 -2674
rect -529 -2700 -499 -2674
rect -445 -2700 -415 -2674
rect -3132 -2916 -2106 -2900
rect -3132 -2950 -3116 -2916
rect -3082 -2950 -2924 -2916
rect -2890 -2950 -2732 -2916
rect -2698 -2950 -2540 -2916
rect -2506 -2950 -2348 -2916
rect -2314 -2950 -2156 -2916
rect -2122 -2950 -2106 -2916
rect -3132 -2966 -2106 -2950
rect -1044 -2852 -1014 -2830
rect -529 -2852 -499 -2830
rect -3066 -2998 -3036 -2966
rect -2970 -2998 -2940 -2966
rect -2874 -2998 -2844 -2966
rect -2778 -2998 -2748 -2966
rect -2682 -2998 -2652 -2966
rect -2586 -2998 -2556 -2966
rect -2490 -2998 -2460 -2966
rect -2394 -2998 -2364 -2966
rect -2298 -2998 -2268 -2966
rect -2202 -2998 -2172 -2966
rect -3066 -3296 -3036 -3270
rect -2970 -3296 -2940 -3270
rect -2874 -3296 -2844 -3270
rect -2778 -3296 -2748 -3270
rect -2682 -3296 -2652 -3270
rect -2586 -3296 -2556 -3270
rect -2490 -3296 -2460 -3270
rect -2394 -3296 -2364 -3270
rect -2298 -3296 -2268 -3270
rect -2202 -3296 -2172 -3270
rect -1100 -2868 -1014 -2852
rect -1100 -2902 -1084 -2868
rect -1050 -2902 -1014 -2868
rect -1100 -2918 -1014 -2902
rect -591 -2868 -499 -2852
rect -591 -2902 -576 -2868
rect -542 -2902 -499 -2868
rect -591 -2918 -499 -2902
rect -1044 -2950 -1014 -2918
rect -529 -2950 -499 -2918
rect -445 -2852 -415 -2830
rect -445 -2868 -357 -2852
rect -445 -2902 -408 -2868
rect -374 -2902 -357 -2868
rect -445 -2918 -357 -2902
rect -445 -2950 -415 -2918
rect 419 -2909 1445 -2893
rect 419 -2943 435 -2909
rect 469 -2943 627 -2909
rect 661 -2943 819 -2909
rect 853 -2943 1011 -2909
rect 1045 -2943 1203 -2909
rect 1237 -2943 1395 -2909
rect 1429 -2943 1445 -2909
rect 419 -2959 1445 -2943
rect 485 -2990 515 -2959
rect 581 -2990 611 -2959
rect 677 -2990 707 -2959
rect 773 -2990 803 -2959
rect 869 -2990 899 -2959
rect 965 -2990 995 -2959
rect 1061 -2990 1091 -2959
rect 1157 -2990 1187 -2959
rect 1253 -2990 1283 -2959
rect 1349 -2990 1379 -2959
rect -1044 -3176 -1014 -3150
rect -529 -3176 -499 -3150
rect -445 -3176 -415 -3150
rect 485 -3120 515 -3094
rect 581 -3120 611 -3094
rect 677 -3120 707 -3094
rect 773 -3120 803 -3094
rect 869 -3120 899 -3094
rect 965 -3120 995 -3094
rect 1061 -3120 1091 -3094
rect 1157 -3120 1187 -3094
rect 1253 -3120 1283 -3094
rect 1349 -3120 1379 -3094
rect 1661 -2996 1691 -2970
rect 1661 -3118 1691 -3096
rect 1940 -2909 2966 -2893
rect 1940 -2943 1956 -2909
rect 1990 -2943 2148 -2909
rect 2182 -2943 2340 -2909
rect 2374 -2943 2532 -2909
rect 2566 -2943 2724 -2909
rect 2758 -2943 2916 -2909
rect 2950 -2943 2966 -2909
rect 1940 -2959 2966 -2943
rect 2006 -2990 2036 -2959
rect 2102 -2990 2132 -2959
rect 2198 -2990 2228 -2959
rect 2294 -2990 2324 -2959
rect 2390 -2990 2420 -2959
rect 2486 -2990 2516 -2959
rect 2582 -2990 2612 -2959
rect 2678 -2990 2708 -2959
rect 2774 -2990 2804 -2959
rect 2870 -2990 2900 -2959
rect 1643 -3134 1709 -3118
rect 1643 -3168 1659 -3134
rect 1693 -3168 1709 -3134
rect 1643 -3184 1709 -3168
rect 2006 -3120 2036 -3094
rect 2102 -3120 2132 -3094
rect 2198 -3120 2228 -3094
rect 2294 -3120 2324 -3094
rect 2390 -3120 2420 -3094
rect 2486 -3120 2516 -3094
rect 2582 -3120 2612 -3094
rect 2678 -3120 2708 -3094
rect 2774 -3120 2804 -3094
rect 2870 -3120 2900 -3094
rect -529 -3244 -499 -3218
rect -445 -3244 -415 -3218
rect -529 -3476 -499 -3444
rect -3066 -3576 -3036 -3550
rect -2970 -3576 -2940 -3550
rect -2874 -3576 -2844 -3550
rect -2778 -3576 -2748 -3550
rect -2682 -3576 -2652 -3550
rect -2586 -3576 -2556 -3550
rect -2490 -3576 -2460 -3550
rect -2394 -3576 -2364 -3550
rect -2298 -3576 -2268 -3550
rect -2202 -3576 -2172 -3550
rect -591 -3492 -499 -3476
rect -591 -3526 -576 -3492
rect -542 -3526 -499 -3492
rect -591 -3542 -499 -3526
rect -3066 -3711 -3036 -3680
rect -2970 -3711 -2940 -3680
rect -2874 -3711 -2844 -3680
rect -2778 -3711 -2748 -3680
rect -2682 -3711 -2652 -3680
rect -2586 -3711 -2556 -3680
rect -2490 -3711 -2460 -3680
rect -2394 -3711 -2364 -3680
rect -2298 -3711 -2268 -3680
rect -2202 -3711 -2172 -3680
rect -3132 -3727 -2106 -3711
rect -3132 -3761 -3116 -3727
rect -3082 -3761 -2924 -3727
rect -2890 -3761 -2732 -3727
rect -2698 -3761 -2540 -3727
rect -2506 -3761 -2348 -3727
rect -2314 -3761 -2156 -3727
rect -2122 -3761 -2106 -3727
rect -3132 -3777 -2106 -3761
rect -529 -3564 -499 -3542
rect -445 -3476 -415 -3444
rect -445 -3492 -357 -3476
rect -445 -3526 -408 -3492
rect -374 -3526 -357 -3492
rect -445 -3542 -357 -3526
rect -445 -3564 -415 -3542
rect -529 -3720 -499 -3694
rect -445 -3720 -415 -3694
rect 485 -3400 515 -3374
rect 581 -3400 611 -3374
rect 677 -3400 707 -3374
rect 773 -3400 803 -3374
rect 869 -3400 899 -3374
rect 965 -3400 995 -3374
rect 1061 -3400 1091 -3374
rect 1157 -3400 1187 -3374
rect 1253 -3400 1283 -3374
rect 1349 -3400 1379 -3374
rect 485 -3704 515 -3672
rect 581 -3704 611 -3672
rect 677 -3704 707 -3672
rect 773 -3704 803 -3672
rect 869 -3704 899 -3672
rect 965 -3704 995 -3672
rect 1061 -3704 1091 -3672
rect 1157 -3704 1187 -3672
rect 1253 -3704 1283 -3672
rect 1349 -3704 1379 -3672
rect -492 -3788 -462 -3762
rect 419 -3720 1445 -3704
rect 419 -3754 435 -3720
rect 469 -3754 627 -3720
rect 661 -3754 819 -3720
rect 853 -3754 1011 -3720
rect 1045 -3754 1203 -3720
rect 1237 -3754 1395 -3720
rect 1429 -3754 1445 -3720
rect 419 -3770 1445 -3754
rect 2006 -3400 2036 -3374
rect 2102 -3400 2132 -3374
rect 2198 -3400 2228 -3374
rect 2294 -3400 2324 -3374
rect 2390 -3400 2420 -3374
rect 2486 -3400 2516 -3374
rect 2582 -3400 2612 -3374
rect 2678 -3400 2708 -3374
rect 2774 -3400 2804 -3374
rect 2870 -3400 2900 -3374
rect 2006 -3704 2036 -3672
rect 2102 -3704 2132 -3672
rect 2198 -3704 2228 -3672
rect 2294 -3704 2324 -3672
rect 2390 -3704 2420 -3672
rect 2486 -3704 2516 -3672
rect 2582 -3704 2612 -3672
rect 2678 -3704 2708 -3672
rect 2774 -3704 2804 -3672
rect 2870 -3704 2900 -3672
rect 1940 -3720 2966 -3704
rect 1940 -3754 1956 -3720
rect 1990 -3754 2148 -3720
rect 2182 -3754 2340 -3720
rect 2374 -3754 2532 -3720
rect 2566 -3754 2724 -3720
rect 2758 -3754 2916 -3720
rect 2950 -3754 2966 -3720
rect 1940 -3770 2966 -3754
rect -492 -3940 -462 -3918
rect -548 -3956 -462 -3940
rect -548 -3990 -532 -3956
rect -498 -3990 -462 -3956
rect -548 -4006 -462 -3990
rect -492 -4038 -462 -4006
rect -3132 -4294 -2106 -4278
rect -3132 -4328 -3116 -4294
rect -3082 -4328 -2924 -4294
rect -2890 -4328 -2732 -4294
rect -2698 -4328 -2540 -4294
rect -2506 -4328 -2348 -4294
rect -2314 -4328 -2156 -4294
rect -2122 -4328 -2106 -4294
rect -3132 -4344 -2106 -4328
rect -492 -4264 -462 -4238
rect -3066 -4376 -3036 -4344
rect -2970 -4376 -2940 -4344
rect -2874 -4376 -2844 -4344
rect -2778 -4376 -2748 -4344
rect -2682 -4376 -2652 -4344
rect -2586 -4376 -2556 -4344
rect -2490 -4376 -2460 -4344
rect -2394 -4376 -2364 -4344
rect -2298 -4376 -2268 -4344
rect -2202 -4376 -2172 -4344
rect -3066 -4674 -3036 -4648
rect -2970 -4674 -2940 -4648
rect -2874 -4674 -2844 -4648
rect -2778 -4674 -2748 -4648
rect -2682 -4674 -2652 -4648
rect -2586 -4674 -2556 -4648
rect -2490 -4674 -2460 -4648
rect -2394 -4674 -2364 -4648
rect -2298 -4674 -2268 -4648
rect -2202 -4674 -2172 -4648
rect -492 -4332 -462 -4306
rect 419 -4287 1445 -4271
rect 419 -4321 435 -4287
rect 469 -4321 627 -4287
rect 661 -4321 819 -4287
rect 853 -4321 1011 -4287
rect 1045 -4321 1203 -4287
rect 1237 -4321 1395 -4287
rect 1429 -4321 1445 -4287
rect 419 -4337 1445 -4321
rect 485 -4368 515 -4337
rect 581 -4368 611 -4337
rect 677 -4368 707 -4337
rect 773 -4368 803 -4337
rect 869 -4368 899 -4337
rect 965 -4368 995 -4337
rect 1061 -4368 1091 -4337
rect 1157 -4368 1187 -4337
rect 1253 -4368 1283 -4337
rect 1349 -4368 1379 -4337
rect -492 -4564 -462 -4532
rect -548 -4580 -462 -4564
rect -548 -4614 -532 -4580
rect -498 -4614 -462 -4580
rect 485 -4498 515 -4472
rect 581 -4498 611 -4472
rect 677 -4498 707 -4472
rect 773 -4498 803 -4472
rect 869 -4498 899 -4472
rect 965 -4498 995 -4472
rect 1061 -4498 1091 -4472
rect 1157 -4498 1187 -4472
rect 1253 -4498 1283 -4472
rect 1349 -4498 1379 -4472
rect 1661 -4374 1691 -4348
rect 1661 -4496 1691 -4474
rect 1940 -4287 2966 -4271
rect 1940 -4321 1956 -4287
rect 1990 -4321 2148 -4287
rect 2182 -4321 2340 -4287
rect 2374 -4321 2532 -4287
rect 2566 -4321 2724 -4287
rect 2758 -4321 2916 -4287
rect 2950 -4321 2966 -4287
rect 1940 -4337 2966 -4321
rect 2006 -4368 2036 -4337
rect 2102 -4368 2132 -4337
rect 2198 -4368 2228 -4337
rect 2294 -4368 2324 -4337
rect 2390 -4368 2420 -4337
rect 2486 -4368 2516 -4337
rect 2582 -4368 2612 -4337
rect 2678 -4368 2708 -4337
rect 2774 -4368 2804 -4337
rect 2870 -4368 2900 -4337
rect 1643 -4512 1709 -4496
rect 1643 -4546 1659 -4512
rect 1693 -4546 1709 -4512
rect 1643 -4562 1709 -4546
rect 2006 -4498 2036 -4472
rect 2102 -4498 2132 -4472
rect 2198 -4498 2228 -4472
rect 2294 -4498 2324 -4472
rect 2390 -4498 2420 -4472
rect 2486 -4498 2516 -4472
rect 2582 -4498 2612 -4472
rect 2678 -4498 2708 -4472
rect 2774 -4498 2804 -4472
rect 2870 -4498 2900 -4472
rect -548 -4630 -462 -4614
rect -492 -4652 -462 -4630
rect -492 -4808 -462 -4782
rect -3066 -4954 -3036 -4928
rect -2970 -4954 -2940 -4928
rect -2874 -4954 -2844 -4928
rect -2778 -4954 -2748 -4928
rect -2682 -4954 -2652 -4928
rect -2586 -4954 -2556 -4928
rect -2490 -4954 -2460 -4928
rect -2394 -4954 -2364 -4928
rect -2298 -4954 -2268 -4928
rect -2202 -4954 -2172 -4928
rect -3066 -5089 -3036 -5058
rect -2970 -5089 -2940 -5058
rect -2874 -5089 -2844 -5058
rect -2778 -5089 -2748 -5058
rect -2682 -5089 -2652 -5058
rect -2586 -5089 -2556 -5058
rect -2490 -5089 -2460 -5058
rect -2394 -5089 -2364 -5058
rect -2298 -5089 -2268 -5058
rect -2202 -5089 -2172 -5058
rect -3132 -5105 -2106 -5089
rect -3132 -5139 -3116 -5105
rect -3082 -5139 -2924 -5105
rect -2890 -5139 -2732 -5105
rect -2698 -5139 -2540 -5105
rect -2506 -5139 -2348 -5105
rect -2314 -5139 -2156 -5105
rect -2122 -5139 -2106 -5105
rect -3132 -5155 -2106 -5139
rect 485 -4778 515 -4752
rect 581 -4778 611 -4752
rect 677 -4778 707 -4752
rect 773 -4778 803 -4752
rect 869 -4778 899 -4752
rect 965 -4778 995 -4752
rect 1061 -4778 1091 -4752
rect 1157 -4778 1187 -4752
rect 1253 -4778 1283 -4752
rect 1349 -4778 1379 -4752
rect 485 -5082 515 -5050
rect 581 -5082 611 -5050
rect 677 -5082 707 -5050
rect 773 -5082 803 -5050
rect 869 -5082 899 -5050
rect 965 -5082 995 -5050
rect 1061 -5082 1091 -5050
rect 1157 -5082 1187 -5050
rect 1253 -5082 1283 -5050
rect 1349 -5082 1379 -5050
rect 419 -5098 1445 -5082
rect 419 -5132 435 -5098
rect 469 -5132 627 -5098
rect 661 -5132 819 -5098
rect 853 -5132 1011 -5098
rect 1045 -5132 1203 -5098
rect 1237 -5132 1395 -5098
rect 1429 -5132 1445 -5098
rect 419 -5148 1445 -5132
rect 2006 -4778 2036 -4752
rect 2102 -4778 2132 -4752
rect 2198 -4778 2228 -4752
rect 2294 -4778 2324 -4752
rect 2390 -4778 2420 -4752
rect 2486 -4778 2516 -4752
rect 2582 -4778 2612 -4752
rect 2678 -4778 2708 -4752
rect 2774 -4778 2804 -4752
rect 2870 -4778 2900 -4752
rect 2006 -5082 2036 -5050
rect 2102 -5082 2132 -5050
rect 2198 -5082 2228 -5050
rect 2294 -5082 2324 -5050
rect 2390 -5082 2420 -5050
rect 2486 -5082 2516 -5050
rect 2582 -5082 2612 -5050
rect 2678 -5082 2708 -5050
rect 2774 -5082 2804 -5050
rect 2870 -5082 2900 -5050
rect 1940 -5098 2966 -5082
rect 1940 -5132 1956 -5098
rect 1990 -5132 2148 -5098
rect 2182 -5132 2340 -5098
rect 2374 -5132 2532 -5098
rect 2566 -5132 2724 -5098
rect 2758 -5132 2916 -5098
rect 2950 -5132 2966 -5098
rect 1940 -5148 2966 -5132
<< polycont >>
rect -3116 -238 -3082 -204
rect -2924 -238 -2890 -204
rect -2732 -238 -2698 -204
rect -2540 -238 -2506 -204
rect -2348 -238 -2314 -204
rect -2156 -238 -2122 -204
rect 435 -231 469 -197
rect 627 -231 661 -197
rect 819 -231 853 -197
rect 1011 -231 1045 -197
rect 1203 -231 1237 -197
rect 1395 -231 1429 -197
rect 1956 -231 1990 -197
rect 2148 -231 2182 -197
rect 2340 -231 2374 -197
rect 2532 -231 2566 -197
rect 2724 -231 2758 -197
rect 2916 -231 2950 -197
rect 1659 -456 1693 -422
rect -900 -726 -866 -692
rect -532 -726 -498 -692
rect -3116 -1049 -3082 -1015
rect -2924 -1049 -2890 -1015
rect -2732 -1049 -2698 -1015
rect -2540 -1049 -2506 -1015
rect -2348 -1049 -2314 -1015
rect -2156 -1049 -2122 -1015
rect 435 -1042 469 -1008
rect 627 -1042 661 -1008
rect 819 -1042 853 -1008
rect 1011 -1042 1045 -1008
rect 1203 -1042 1237 -1008
rect 1395 -1042 1429 -1008
rect 1956 -1042 1990 -1008
rect 2148 -1042 2182 -1008
rect 2340 -1042 2374 -1008
rect 2532 -1042 2566 -1008
rect 2724 -1042 2758 -1008
rect 2916 -1042 2950 -1008
rect -532 -1350 -498 -1316
rect -3116 -1572 -3082 -1538
rect -2924 -1572 -2890 -1538
rect -2732 -1572 -2698 -1538
rect -2540 -1572 -2506 -1538
rect -2348 -1572 -2314 -1538
rect -2156 -1572 -2122 -1538
rect 435 -1565 469 -1531
rect 627 -1565 661 -1531
rect 819 -1565 853 -1531
rect 1011 -1565 1045 -1531
rect 1203 -1565 1237 -1531
rect 1395 -1565 1429 -1531
rect -576 -1814 -542 -1780
rect -408 -1814 -374 -1780
rect 1956 -1565 1990 -1531
rect 2148 -1565 2182 -1531
rect 2340 -1565 2374 -1531
rect 2532 -1565 2566 -1531
rect 2724 -1565 2758 -1531
rect 2916 -1565 2950 -1531
rect 1659 -1790 1693 -1756
rect -3116 -2383 -3082 -2349
rect -2924 -2383 -2890 -2349
rect -2732 -2383 -2698 -2349
rect -2540 -2383 -2506 -2349
rect -2348 -2383 -2314 -2349
rect -2156 -2383 -2122 -2349
rect -1084 -2438 -1050 -2404
rect -576 -2438 -542 -2404
rect -408 -2438 -374 -2404
rect 435 -2376 469 -2342
rect 627 -2376 661 -2342
rect 819 -2376 853 -2342
rect 1011 -2376 1045 -2342
rect 1203 -2376 1237 -2342
rect 1395 -2376 1429 -2342
rect 1956 -2376 1990 -2342
rect 2148 -2376 2182 -2342
rect 2340 -2376 2374 -2342
rect 2532 -2376 2566 -2342
rect 2724 -2376 2758 -2342
rect 2916 -2376 2950 -2342
rect -3116 -2950 -3082 -2916
rect -2924 -2950 -2890 -2916
rect -2732 -2950 -2698 -2916
rect -2540 -2950 -2506 -2916
rect -2348 -2950 -2314 -2916
rect -2156 -2950 -2122 -2916
rect -1084 -2902 -1050 -2868
rect -576 -2902 -542 -2868
rect -408 -2902 -374 -2868
rect 435 -2943 469 -2909
rect 627 -2943 661 -2909
rect 819 -2943 853 -2909
rect 1011 -2943 1045 -2909
rect 1203 -2943 1237 -2909
rect 1395 -2943 1429 -2909
rect 1956 -2943 1990 -2909
rect 2148 -2943 2182 -2909
rect 2340 -2943 2374 -2909
rect 2532 -2943 2566 -2909
rect 2724 -2943 2758 -2909
rect 2916 -2943 2950 -2909
rect 1659 -3168 1693 -3134
rect -576 -3526 -542 -3492
rect -3116 -3761 -3082 -3727
rect -2924 -3761 -2890 -3727
rect -2732 -3761 -2698 -3727
rect -2540 -3761 -2506 -3727
rect -2348 -3761 -2314 -3727
rect -2156 -3761 -2122 -3727
rect -408 -3526 -374 -3492
rect 435 -3754 469 -3720
rect 627 -3754 661 -3720
rect 819 -3754 853 -3720
rect 1011 -3754 1045 -3720
rect 1203 -3754 1237 -3720
rect 1395 -3754 1429 -3720
rect 1956 -3754 1990 -3720
rect 2148 -3754 2182 -3720
rect 2340 -3754 2374 -3720
rect 2532 -3754 2566 -3720
rect 2724 -3754 2758 -3720
rect 2916 -3754 2950 -3720
rect -532 -3990 -498 -3956
rect -3116 -4328 -3082 -4294
rect -2924 -4328 -2890 -4294
rect -2732 -4328 -2698 -4294
rect -2540 -4328 -2506 -4294
rect -2348 -4328 -2314 -4294
rect -2156 -4328 -2122 -4294
rect 435 -4321 469 -4287
rect 627 -4321 661 -4287
rect 819 -4321 853 -4287
rect 1011 -4321 1045 -4287
rect 1203 -4321 1237 -4287
rect 1395 -4321 1429 -4287
rect -532 -4614 -498 -4580
rect 1956 -4321 1990 -4287
rect 2148 -4321 2182 -4287
rect 2340 -4321 2374 -4287
rect 2532 -4321 2566 -4287
rect 2724 -4321 2758 -4287
rect 2916 -4321 2950 -4287
rect 1659 -4546 1693 -4512
rect -3116 -5139 -3082 -5105
rect -2924 -5139 -2890 -5105
rect -2732 -5139 -2698 -5105
rect -2540 -5139 -2506 -5105
rect -2348 -5139 -2314 -5105
rect -2156 -5139 -2122 -5105
rect 435 -5132 469 -5098
rect 627 -5132 661 -5098
rect 819 -5132 853 -5098
rect 1011 -5132 1045 -5098
rect 1203 -5132 1237 -5098
rect 1395 -5132 1429 -5098
rect 1956 -5132 1990 -5098
rect 2148 -5132 2182 -5098
rect 2340 -5132 2374 -5098
rect 2532 -5132 2566 -5098
rect 2724 -5132 2758 -5098
rect 2916 -5132 2950 -5098
<< locali >>
rect -3843 224 3659 352
rect -3230 -136 -3134 -102
rect -2104 -118 -2008 -102
rect -1670 -118 -1542 224
rect -2104 -136 -1542 -118
rect -3230 -198 -3196 -136
rect -2042 -182 -1542 -136
rect -3132 -201 -2106 -196
rect -3132 -204 -2348 -201
rect -2314 -204 -2106 -201
rect -3132 -238 -3116 -204
rect -3082 -238 -2924 -204
rect -2890 -238 -2732 -204
rect -2698 -238 -2540 -204
rect -2506 -238 -2348 -204
rect -2314 -238 -2156 -204
rect -2122 -238 -2106 -204
rect -3132 -246 -2106 -238
rect -2042 -198 -2008 -182
rect -3116 -298 -3082 -282
rect -3116 -562 -3082 -546
rect -3020 -298 -2986 -282
rect -3020 -562 -2986 -546
rect -2924 -298 -2890 -282
rect -2924 -562 -2890 -546
rect -2828 -298 -2794 -282
rect -2828 -562 -2794 -546
rect -2732 -298 -2698 -282
rect -2732 -562 -2698 -546
rect -2636 -298 -2602 -282
rect -2636 -562 -2602 -546
rect -2540 -298 -2506 -282
rect -2540 -562 -2506 -546
rect -2444 -298 -2410 -282
rect -2444 -562 -2410 -546
rect -2348 -298 -2314 -282
rect -2348 -562 -2314 -546
rect -2252 -298 -2218 -282
rect -2252 -562 -2218 -546
rect -2156 -298 -2122 -282
rect -2156 -562 -2122 -546
rect -3230 -646 -3196 -584
rect -2042 -646 -2008 -584
rect -3230 -680 -3134 -646
rect -2104 -680 -2008 -646
rect -3230 -786 -3134 -752
rect -2104 -786 -2008 -752
rect -3230 -848 -3196 -786
rect -3564 -1046 -3230 -1024
rect -2042 -848 -2008 -786
rect -3116 -876 -3082 -860
rect -3116 -972 -3082 -956
rect -3020 -876 -2986 -860
rect -3020 -972 -2986 -956
rect -2924 -876 -2890 -860
rect -2924 -972 -2890 -956
rect -2828 -876 -2794 -860
rect -2828 -972 -2794 -956
rect -2732 -876 -2698 -860
rect -2732 -972 -2698 -956
rect -2636 -876 -2602 -860
rect -2636 -972 -2602 -956
rect -2540 -876 -2506 -860
rect -2540 -972 -2506 -956
rect -2444 -876 -2410 -860
rect -2444 -972 -2410 -956
rect -2348 -876 -2314 -860
rect -2348 -972 -2314 -956
rect -2252 -876 -2218 -860
rect -2252 -972 -2218 -956
rect -2156 -876 -2122 -860
rect -2156 -972 -2122 -956
rect -3564 -1088 -3196 -1046
rect -3132 -1015 -2106 -1007
rect -3132 -1049 -3116 -1015
rect -3082 -1049 -2924 -1015
rect -2890 -1049 -2732 -1015
rect -2698 -1049 -2540 -1015
rect -2506 -1049 -2348 -1015
rect -2314 -1019 -2156 -1015
rect -2122 -1016 -2106 -1015
rect -2311 -1049 -2156 -1019
rect -3132 -1053 -2345 -1049
rect -2311 -1050 -2155 -1049
rect -2121 -1050 -2106 -1016
rect -2311 -1053 -2106 -1050
rect -3132 -1057 -2106 -1053
rect -3564 -2383 -3500 -1088
rect -3230 -1108 -3196 -1088
rect -2042 -1108 -2008 -1046
rect -3230 -1142 -3134 -1108
rect -2104 -1142 -2008 -1108
rect -1670 -989 -1542 -182
rect -165 -102 1647 -5
rect -165 -104 1889 -102
rect -165 -133 417 -104
rect -165 -444 -37 -133
rect -355 -460 -37 -444
rect -980 -494 -951 -460
rect -917 -494 -859 -460
rect -825 -494 -767 -460
rect -733 -494 -675 -460
rect -641 -494 -583 -460
rect -549 -494 -491 -460
rect -457 -494 -399 -460
rect -365 -494 -37 -460
rect 321 -138 417 -133
rect 1447 -138 1938 -104
rect 2968 -138 3064 -104
rect 321 -200 355 -138
rect 1509 -170 1876 -138
rect 419 -197 1445 -189
rect 419 -231 435 -197
rect 469 -231 627 -197
rect 661 -231 819 -197
rect 853 -231 1011 -197
rect 1045 -231 1203 -197
rect 1237 -231 1395 -197
rect 1429 -231 1445 -197
rect 419 -239 1445 -231
rect 1509 -200 1543 -170
rect 435 -290 469 -274
rect 435 -386 469 -370
rect 531 -290 565 -274
rect 531 -386 565 -370
rect 627 -290 661 -274
rect 627 -386 661 -370
rect 723 -290 757 -274
rect 723 -386 757 -370
rect 819 -290 853 -274
rect 819 -386 853 -370
rect 915 -290 949 -274
rect 915 -386 949 -370
rect 1011 -290 1045 -274
rect 1011 -386 1045 -370
rect 1107 -290 1141 -274
rect 1107 -386 1141 -370
rect 1203 -290 1237 -274
rect 1203 -386 1237 -370
rect 1299 -290 1333 -274
rect 1299 -386 1333 -370
rect 1395 -290 1429 -274
rect 1395 -386 1429 -370
rect 1842 -200 1876 -170
rect 321 -460 355 -398
rect 1615 -296 1649 -280
rect 1615 -388 1649 -372
rect 1703 -296 1737 -280
rect 1703 -388 1737 -372
rect 1509 -460 1543 -398
rect 1940 -197 2966 -189
rect 1940 -231 1956 -197
rect 1990 -231 2148 -197
rect 2182 -231 2340 -197
rect 2374 -231 2532 -197
rect 2566 -231 2724 -197
rect 2758 -231 2916 -197
rect 2950 -231 2966 -197
rect 1940 -239 2966 -231
rect 3030 -200 3064 -138
rect 1956 -290 1990 -274
rect 1956 -386 1990 -370
rect 2052 -290 2086 -274
rect 2052 -386 2086 -370
rect 2148 -290 2182 -274
rect 2148 -386 2182 -370
rect 2244 -290 2278 -274
rect 2244 -386 2278 -370
rect 2340 -290 2374 -274
rect 2340 -386 2374 -370
rect 2436 -290 2470 -274
rect 2436 -386 2470 -370
rect 2532 -290 2566 -274
rect 2532 -386 2566 -370
rect 2628 -290 2662 -274
rect 2628 -386 2662 -370
rect 2724 -290 2758 -274
rect 2724 -386 2758 -370
rect 2820 -290 2854 -274
rect 2820 -386 2854 -370
rect 2916 -290 2950 -274
rect 2916 -386 2950 -370
rect 1643 -456 1659 -422
rect 1693 -456 1709 -422
rect 321 -494 417 -460
rect 1447 -494 1543 -460
rect 1842 -460 1876 -398
rect 3030 -460 3064 -398
rect 1842 -494 1938 -460
rect 2968 -494 3064 -460
rect -916 -540 -870 -494
rect -916 -574 -904 -540
rect -916 -608 -870 -574
rect -916 -642 -904 -608
rect -916 -658 -870 -642
rect -836 -540 -770 -528
rect -836 -574 -820 -540
rect -786 -574 -770 -540
rect -836 -603 -770 -574
rect -836 -637 -822 -603
rect -788 -608 -770 -603
rect -836 -642 -820 -637
rect -786 -642 -770 -608
rect -687 -588 -629 -494
rect -687 -622 -675 -588
rect -641 -622 -629 -588
rect -687 -639 -629 -622
rect -548 -540 -502 -494
rect -355 -508 -37 -494
rect -548 -574 -536 -540
rect -548 -608 -502 -574
rect -836 -654 -770 -642
rect -916 -698 -900 -692
rect -916 -732 -905 -698
rect -866 -726 -850 -692
rect -871 -732 -850 -726
rect -916 -740 -850 -732
rect -816 -774 -770 -654
rect -548 -642 -536 -608
rect -548 -658 -502 -642
rect -468 -540 -402 -528
rect -468 -574 -452 -540
rect -418 -574 -402 -540
rect -468 -594 -402 -574
rect -468 -642 -452 -594
rect -418 -642 -402 -594
rect -468 -654 -402 -642
rect -548 -700 -532 -692
rect -548 -734 -538 -700
rect -498 -726 -482 -692
rect -504 -734 -482 -726
rect -548 -740 -482 -734
rect -912 -792 -870 -776
rect -912 -826 -904 -792
rect -912 -860 -870 -826
rect -912 -894 -904 -860
rect -912 -928 -870 -894
rect -912 -962 -904 -928
rect -912 -989 -870 -962
rect -836 -792 -770 -774
rect -836 -826 -820 -792
rect -786 -826 -770 -792
rect -836 -860 -770 -826
rect -836 -894 -820 -860
rect -786 -894 -770 -860
rect -836 -928 -770 -894
rect -836 -962 -820 -928
rect -786 -962 -770 -928
rect -836 -970 -770 -962
rect -687 -806 -629 -771
rect -448 -774 -402 -654
rect -687 -840 -675 -806
rect -641 -840 -629 -806
rect -687 -899 -629 -840
rect -687 -933 -675 -899
rect -641 -933 -629 -899
rect -1670 -1004 -870 -989
rect -687 -1004 -629 -933
rect -544 -792 -502 -776
rect -544 -826 -536 -792
rect -544 -860 -502 -826
rect -544 -894 -536 -860
rect -544 -928 -502 -894
rect -544 -962 -536 -928
rect -544 -1004 -502 -962
rect -468 -792 -402 -774
rect -468 -826 -452 -792
rect -418 -826 -402 -792
rect -468 -860 -402 -826
rect -468 -894 -452 -860
rect -418 -894 -402 -860
rect -468 -928 -402 -894
rect -468 -962 -452 -928
rect -418 -962 -402 -928
rect -468 -970 -402 -962
rect -1670 -1038 -951 -1004
rect -917 -1038 -859 -1004
rect -825 -1038 -767 -1004
rect -733 -1038 -675 -1004
rect -641 -1038 -583 -1004
rect -549 -1038 -491 -1004
rect -457 -1038 -399 -1004
rect -365 -1038 -336 -1004
rect -1670 -1053 -891 -1038
rect -3230 -1470 -3134 -1436
rect -2104 -1443 -2008 -1436
rect -1670 -1443 -1542 -1053
rect -687 -1109 -629 -1038
rect -687 -1143 -675 -1109
rect -641 -1143 -629 -1109
rect -687 -1202 -629 -1143
rect -687 -1236 -675 -1202
rect -641 -1236 -629 -1202
rect -687 -1271 -629 -1236
rect -544 -1080 -502 -1038
rect -544 -1114 -536 -1080
rect -544 -1148 -502 -1114
rect -544 -1182 -536 -1148
rect -544 -1216 -502 -1182
rect -544 -1250 -536 -1216
rect -544 -1266 -502 -1250
rect -468 -1080 -402 -1072
rect -468 -1114 -452 -1080
rect -418 -1114 -402 -1080
rect -468 -1148 -402 -1114
rect -468 -1182 -452 -1148
rect -418 -1182 -402 -1148
rect -468 -1197 -402 -1182
rect -468 -1231 -453 -1197
rect -419 -1216 -402 -1197
rect -468 -1250 -452 -1231
rect -418 -1250 -402 -1216
rect -468 -1268 -402 -1250
rect -548 -1312 -482 -1302
rect -548 -1346 -534 -1312
rect -500 -1316 -482 -1312
rect -548 -1350 -532 -1346
rect -498 -1350 -482 -1316
rect -548 -1400 -502 -1384
rect -448 -1388 -402 -1268
rect -2104 -1470 -1542 -1443
rect -3230 -1532 -3196 -1470
rect -2042 -1507 -1542 -1470
rect -3132 -1538 -2106 -1530
rect -3132 -1572 -3116 -1538
rect -3082 -1572 -2924 -1538
rect -2890 -1572 -2732 -1538
rect -2698 -1572 -2540 -1538
rect -2506 -1572 -2348 -1538
rect -2314 -1572 -2156 -1538
rect -2122 -1572 -2106 -1538
rect -3132 -1580 -2106 -1572
rect -2042 -1532 -2008 -1507
rect -3116 -1632 -3082 -1616
rect -3116 -1896 -3082 -1880
rect -3020 -1632 -2986 -1616
rect -3020 -1896 -2986 -1880
rect -2924 -1632 -2890 -1616
rect -2924 -1896 -2890 -1880
rect -2828 -1632 -2794 -1616
rect -2828 -1896 -2794 -1880
rect -2732 -1632 -2698 -1616
rect -2732 -1896 -2698 -1880
rect -2636 -1632 -2602 -1616
rect -2636 -1896 -2602 -1880
rect -2540 -1632 -2506 -1616
rect -2540 -1896 -2506 -1880
rect -2444 -1632 -2410 -1616
rect -2444 -1896 -2410 -1880
rect -2348 -1632 -2314 -1616
rect -2348 -1896 -2314 -1880
rect -2252 -1632 -2218 -1616
rect -2252 -1896 -2218 -1880
rect -2156 -1632 -2122 -1616
rect -2156 -1896 -2122 -1880
rect -3230 -1980 -3196 -1918
rect -2042 -1980 -2008 -1918
rect -3230 -2014 -3134 -1980
rect -2104 -2014 -2008 -1980
rect -1670 -2082 -1542 -1507
rect -687 -1420 -629 -1403
rect -687 -1454 -675 -1420
rect -641 -1454 -629 -1420
rect -687 -1548 -629 -1454
rect -548 -1434 -536 -1400
rect -548 -1468 -502 -1434
rect -548 -1502 -536 -1468
rect -548 -1548 -502 -1502
rect -468 -1400 -402 -1388
rect -468 -1434 -452 -1400
rect -418 -1434 -402 -1400
rect -468 -1468 -402 -1434
rect -468 -1502 -452 -1468
rect -418 -1502 -402 -1468
rect -468 -1514 -402 -1502
rect -165 -1334 -37 -508
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect 1509 -662 1543 -600
rect 435 -700 469 -684
rect 435 -964 469 -948
rect 531 -700 565 -684
rect 531 -964 565 -948
rect 627 -700 661 -684
rect 627 -964 661 -948
rect 723 -700 757 -684
rect 723 -964 757 -948
rect 819 -700 853 -684
rect 819 -964 853 -948
rect 915 -700 949 -684
rect 915 -964 949 -948
rect 1011 -700 1045 -684
rect 1011 -964 1045 -948
rect 1107 -700 1141 -684
rect 1107 -964 1141 -948
rect 1203 -700 1237 -684
rect 1203 -964 1237 -948
rect 1299 -700 1333 -684
rect 1299 -964 1333 -948
rect 1395 -700 1429 -684
rect 1395 -964 1429 -948
rect 321 -1110 355 -1048
rect 419 -1008 1445 -1000
rect 419 -1042 435 -1008
rect 469 -1042 627 -1008
rect 661 -1042 819 -1008
rect 853 -1042 1011 -1008
rect 1045 -1042 1203 -1008
rect 1237 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 419 -1050 1445 -1042
rect 1509 -1076 1543 -1048
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1956 -700 1990 -684
rect 1956 -964 1990 -948
rect 2052 -700 2086 -684
rect 2052 -964 2086 -948
rect 2148 -700 2182 -684
rect 2148 -964 2182 -948
rect 2244 -700 2278 -684
rect 2244 -964 2278 -948
rect 2340 -700 2374 -684
rect 2340 -964 2374 -948
rect 2436 -700 2470 -684
rect 2436 -964 2470 -948
rect 2532 -700 2566 -684
rect 2532 -964 2566 -948
rect 2628 -700 2662 -684
rect 2628 -964 2662 -948
rect 2724 -700 2758 -684
rect 2724 -964 2758 -948
rect 2820 -700 2854 -684
rect 2820 -964 2854 -948
rect 2916 -700 2950 -684
rect 2916 -964 2950 -948
rect 1842 -1076 1876 -1048
rect 1940 -1008 2966 -1000
rect 1940 -1042 1956 -1008
rect 1990 -1042 2148 -1008
rect 2182 -1042 2340 -1008
rect 2374 -1042 2532 -1008
rect 2566 -1042 2724 -1008
rect 2758 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1940 -1050 2966 -1042
rect 3030 -1069 3064 -1048
rect 3329 -1069 3457 224
rect 1509 -1110 1882 -1076
rect 3030 -1110 3457 -1069
rect 321 -1144 417 -1110
rect 1447 -1144 1938 -1110
rect 2968 -1144 3457 -1110
rect 1677 -1249 3457 -1144
rect -165 -1436 1650 -1334
rect -165 -1438 1889 -1436
rect -165 -1472 417 -1438
rect 1447 -1472 1938 -1438
rect 2968 -1472 3064 -1438
rect -165 -1503 355 -1472
rect -165 -1548 -37 -1503
rect -704 -1582 -675 -1548
rect -641 -1582 -583 -1548
rect -549 -1582 -491 -1548
rect -457 -1582 -399 -1548
rect -365 -1582 -37 -1548
rect -687 -1676 -629 -1582
rect -687 -1710 -675 -1676
rect -641 -1710 -629 -1676
rect -687 -1727 -629 -1710
rect -595 -1624 -533 -1582
rect -595 -1658 -573 -1624
rect -539 -1658 -533 -1624
rect -595 -1692 -533 -1658
rect -595 -1726 -573 -1692
rect -539 -1726 -533 -1692
rect -595 -1742 -533 -1726
rect -492 -1624 -353 -1616
rect -492 -1658 -405 -1624
rect -371 -1658 -353 -1624
rect -492 -1676 -353 -1658
rect -492 -1710 -469 -1676
rect -435 -1692 -353 -1676
rect -435 -1710 -405 -1692
rect -492 -1726 -405 -1710
rect -371 -1726 -353 -1692
rect -492 -1742 -353 -1726
rect -593 -1780 -526 -1776
rect -593 -1784 -576 -1780
rect -593 -1818 -582 -1784
rect -542 -1814 -526 -1780
rect -548 -1818 -526 -1814
rect -593 -1830 -526 -1818
rect -687 -1894 -629 -1859
rect -492 -1862 -458 -1742
rect -424 -1819 -408 -1780
rect -374 -1819 -357 -1780
rect -424 -1830 -357 -1819
rect -687 -1928 -675 -1894
rect -641 -1928 -629 -1894
rect -687 -1987 -629 -1928
rect -687 -2021 -675 -1987
rect -641 -2021 -629 -1987
rect -3230 -2120 -3134 -2086
rect -2104 -2120 -2008 -2086
rect -3230 -2182 -3196 -2120
rect -2042 -2182 -2008 -2120
rect -3116 -2210 -3082 -2194
rect -3116 -2306 -3082 -2290
rect -3020 -2210 -2986 -2194
rect -3020 -2306 -2986 -2290
rect -2924 -2210 -2890 -2194
rect -2924 -2306 -2890 -2290
rect -2828 -2210 -2794 -2194
rect -2828 -2306 -2794 -2290
rect -2732 -2210 -2698 -2194
rect -2732 -2306 -2698 -2290
rect -2636 -2210 -2602 -2194
rect -2636 -2306 -2602 -2290
rect -2540 -2210 -2506 -2194
rect -2540 -2306 -2506 -2290
rect -2444 -2210 -2410 -2194
rect -2444 -2306 -2410 -2290
rect -2348 -2210 -2314 -2194
rect -2348 -2306 -2314 -2290
rect -2252 -2210 -2218 -2194
rect -2252 -2306 -2218 -2290
rect -2156 -2210 -2122 -2194
rect -2156 -2306 -2122 -2290
rect -3230 -2383 -3196 -2380
rect -3564 -2442 -3196 -2383
rect -3132 -2349 -2106 -2341
rect -3132 -2383 -3116 -2349
rect -3082 -2383 -2924 -2349
rect -2890 -2383 -2732 -2349
rect -2698 -2383 -2540 -2349
rect -2506 -2383 -2348 -2349
rect -2314 -2383 -2156 -2349
rect -2122 -2383 -2106 -2349
rect -3132 -2391 -2106 -2383
rect -2042 -2442 -2008 -2380
rect -3564 -2447 -3134 -2442
rect -3564 -3782 -3500 -2447
rect -3230 -2476 -3134 -2447
rect -2104 -2476 -2008 -2442
rect -1670 -2092 -1220 -2082
rect -687 -2092 -629 -2021
rect -595 -1880 -539 -1864
rect -595 -1914 -573 -1880
rect -595 -1948 -539 -1914
rect -595 -1982 -573 -1948
rect -595 -2016 -539 -1982
rect -595 -2050 -573 -2016
rect -595 -2092 -539 -2050
rect -505 -1880 -439 -1862
rect -505 -1914 -489 -1880
rect -455 -1914 -439 -1880
rect -505 -1948 -439 -1914
rect -505 -1982 -489 -1948
rect -455 -1982 -439 -1948
rect -505 -2016 -439 -1982
rect -505 -2050 -489 -2016
rect -455 -2050 -439 -2016
rect -505 -2058 -439 -2050
rect -405 -1880 -353 -1864
rect -371 -1914 -353 -1880
rect -405 -1948 -353 -1914
rect -371 -1982 -353 -1948
rect -405 -2016 -353 -1982
rect -371 -2050 -353 -2016
rect -405 -2092 -353 -2050
rect -1670 -2126 -1227 -2092
rect -1193 -2126 -1135 -2092
rect -1101 -2126 -1043 -2092
rect -1009 -2126 -951 -2092
rect -917 -2126 -859 -2092
rect -825 -2126 -767 -2092
rect -733 -2126 -675 -2092
rect -641 -2126 -583 -2092
rect -549 -2126 -491 -2092
rect -457 -2126 -399 -2092
rect -365 -2126 -336 -2092
rect -1670 -2146 -1181 -2126
rect -3230 -2848 -3134 -2814
rect -2104 -2841 -2008 -2814
rect -1670 -2841 -1542 -2146
rect -1239 -2197 -1181 -2146
rect -1239 -2231 -1227 -2197
rect -1193 -2231 -1181 -2197
rect -1239 -2290 -1181 -2231
rect -1239 -2324 -1227 -2290
rect -1193 -2324 -1181 -2290
rect -1239 -2359 -1181 -2324
rect -1096 -2168 -1054 -2126
rect -1096 -2202 -1088 -2168
rect -1096 -2236 -1054 -2202
rect -1096 -2270 -1088 -2236
rect -1096 -2304 -1054 -2270
rect -1096 -2338 -1088 -2304
rect -1096 -2354 -1054 -2338
rect -1020 -2168 -954 -2160
rect -1020 -2202 -1004 -2168
rect -970 -2202 -954 -2168
rect -1020 -2236 -954 -2202
rect -1020 -2270 -1004 -2236
rect -970 -2270 -954 -2236
rect -1020 -2304 -954 -2270
rect -1020 -2338 -1004 -2304
rect -970 -2338 -954 -2304
rect -1020 -2356 -954 -2338
rect -1100 -2398 -1034 -2390
rect -1100 -2432 -1091 -2398
rect -1057 -2404 -1034 -2398
rect -1100 -2438 -1084 -2432
rect -1050 -2438 -1034 -2404
rect -1100 -2488 -1054 -2472
rect -1000 -2476 -954 -2356
rect -687 -2197 -629 -2126
rect -687 -2231 -675 -2197
rect -641 -2231 -629 -2197
rect -687 -2290 -629 -2231
rect -687 -2324 -675 -2290
rect -641 -2324 -629 -2290
rect -687 -2359 -629 -2324
rect -595 -2168 -539 -2126
rect -595 -2202 -573 -2168
rect -595 -2236 -539 -2202
rect -595 -2270 -573 -2236
rect -595 -2304 -539 -2270
rect -595 -2338 -573 -2304
rect -595 -2354 -539 -2338
rect -505 -2168 -439 -2160
rect -505 -2202 -489 -2168
rect -455 -2202 -439 -2168
rect -505 -2236 -439 -2202
rect -505 -2338 -489 -2236
rect -455 -2338 -439 -2236
rect -505 -2356 -439 -2338
rect -405 -2168 -353 -2126
rect -371 -2202 -353 -2168
rect -405 -2236 -353 -2202
rect -371 -2270 -353 -2236
rect -405 -2304 -353 -2270
rect -371 -2338 -353 -2304
rect -405 -2354 -353 -2338
rect -593 -2398 -526 -2388
rect -593 -2432 -583 -2398
rect -549 -2404 -526 -2398
rect -593 -2438 -576 -2432
rect -542 -2438 -526 -2404
rect -593 -2442 -526 -2438
rect -492 -2476 -458 -2356
rect -424 -2395 -357 -2388
rect -424 -2404 -402 -2395
rect -424 -2438 -408 -2404
rect -368 -2429 -357 -2395
rect -374 -2438 -357 -2429
rect -1239 -2508 -1181 -2491
rect -1239 -2542 -1227 -2508
rect -1193 -2542 -1181 -2508
rect -1239 -2636 -1181 -2542
rect -1100 -2522 -1088 -2488
rect -1100 -2556 -1054 -2522
rect -1100 -2590 -1088 -2556
rect -1100 -2636 -1054 -2590
rect -1020 -2488 -954 -2476
rect -1020 -2522 -1004 -2488
rect -970 -2522 -954 -2488
rect -1020 -2556 -954 -2522
rect -1020 -2590 -1004 -2556
rect -970 -2590 -954 -2556
rect -1020 -2602 -954 -2590
rect -687 -2508 -629 -2491
rect -687 -2542 -675 -2508
rect -641 -2542 -629 -2508
rect -687 -2636 -629 -2542
rect -595 -2492 -533 -2476
rect -595 -2526 -573 -2492
rect -539 -2526 -533 -2492
rect -595 -2560 -533 -2526
rect -595 -2594 -573 -2560
rect -539 -2594 -533 -2560
rect -595 -2636 -533 -2594
rect -492 -2492 -353 -2476
rect -492 -2526 -405 -2492
rect -371 -2526 -353 -2492
rect -492 -2560 -353 -2526
rect -492 -2594 -405 -2560
rect -371 -2594 -353 -2560
rect -492 -2602 -353 -2594
rect -165 -2636 -37 -1582
rect 321 -1534 355 -1503
rect 1509 -1504 1876 -1472
rect 419 -1531 1445 -1523
rect 419 -1565 435 -1531
rect 469 -1565 627 -1531
rect 661 -1565 819 -1531
rect 853 -1565 1011 -1531
rect 1045 -1565 1203 -1531
rect 1237 -1565 1395 -1531
rect 1429 -1565 1445 -1531
rect 419 -1573 1445 -1565
rect 1509 -1534 1543 -1504
rect 435 -1624 469 -1608
rect 435 -1720 469 -1704
rect 531 -1624 565 -1608
rect 531 -1720 565 -1704
rect 627 -1624 661 -1608
rect 627 -1720 661 -1704
rect 723 -1624 757 -1608
rect 723 -1720 757 -1704
rect 819 -1624 853 -1608
rect 819 -1720 853 -1704
rect 915 -1624 949 -1608
rect 915 -1720 949 -1704
rect 1011 -1624 1045 -1608
rect 1011 -1720 1045 -1704
rect 1107 -1624 1141 -1608
rect 1107 -1720 1141 -1704
rect 1203 -1624 1237 -1608
rect 1203 -1720 1237 -1704
rect 1299 -1624 1333 -1608
rect 1299 -1720 1333 -1704
rect 1395 -1624 1429 -1608
rect 1395 -1720 1429 -1704
rect 1842 -1534 1876 -1504
rect 321 -1794 355 -1732
rect 1615 -1630 1649 -1614
rect 1615 -1722 1649 -1706
rect 1703 -1630 1737 -1614
rect 1703 -1722 1737 -1706
rect 1509 -1794 1543 -1732
rect 1940 -1531 2966 -1523
rect 1940 -1565 1956 -1531
rect 1990 -1565 2148 -1531
rect 2182 -1565 2340 -1531
rect 2374 -1565 2532 -1531
rect 2566 -1565 2724 -1531
rect 2758 -1565 2916 -1531
rect 2950 -1565 2966 -1531
rect 1940 -1573 2966 -1565
rect 3030 -1534 3064 -1472
rect 1956 -1624 1990 -1608
rect 1956 -1720 1990 -1704
rect 2052 -1624 2086 -1608
rect 2052 -1720 2086 -1704
rect 2148 -1624 2182 -1608
rect 2148 -1720 2182 -1704
rect 2244 -1624 2278 -1608
rect 2244 -1720 2278 -1704
rect 2340 -1624 2374 -1608
rect 2340 -1720 2374 -1704
rect 2436 -1624 2470 -1608
rect 2436 -1720 2470 -1704
rect 2532 -1624 2566 -1608
rect 2532 -1720 2566 -1704
rect 2628 -1624 2662 -1608
rect 2628 -1720 2662 -1704
rect 2724 -1624 2758 -1608
rect 2724 -1720 2758 -1704
rect 2820 -1624 2854 -1608
rect 2820 -1720 2854 -1704
rect 2916 -1624 2950 -1608
rect 2916 -1720 2950 -1704
rect 1643 -1790 1659 -1756
rect 1693 -1790 1709 -1756
rect 321 -1828 417 -1794
rect 1447 -1828 1543 -1794
rect 1842 -1794 1876 -1732
rect 3030 -1794 3064 -1732
rect 1842 -1828 1938 -1794
rect 2968 -1828 3064 -1794
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect 435 -2034 469 -2018
rect 435 -2298 469 -2282
rect 531 -2034 565 -2018
rect 531 -2298 565 -2282
rect 627 -2034 661 -2018
rect 627 -2298 661 -2282
rect 723 -2034 757 -2018
rect 723 -2298 757 -2282
rect 819 -2034 853 -2018
rect 819 -2298 853 -2282
rect 915 -2034 949 -2018
rect 915 -2298 949 -2282
rect 1011 -2034 1045 -2018
rect 1011 -2298 1045 -2282
rect 1107 -2034 1141 -2018
rect 1107 -2298 1141 -2282
rect 1203 -2034 1237 -2018
rect 1203 -2298 1237 -2282
rect 1299 -2034 1333 -2018
rect 1299 -2298 1333 -2282
rect 1395 -2034 1429 -2018
rect 1395 -2298 1429 -2282
rect 321 -2444 355 -2382
rect 419 -2342 1445 -2334
rect 419 -2376 435 -2342
rect 469 -2376 627 -2342
rect 661 -2376 819 -2342
rect 853 -2376 1011 -2342
rect 1045 -2376 1203 -2342
rect 1237 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 419 -2384 1445 -2376
rect 1509 -2410 1543 -2382
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1956 -2034 1990 -2018
rect 1956 -2298 1990 -2282
rect 2052 -2034 2086 -2018
rect 2052 -2298 2086 -2282
rect 2148 -2034 2182 -2018
rect 2148 -2298 2182 -2282
rect 2244 -2034 2278 -2018
rect 2244 -2298 2278 -2282
rect 2340 -2034 2374 -2018
rect 2340 -2298 2374 -2282
rect 2436 -2034 2470 -2018
rect 2436 -2298 2470 -2282
rect 2532 -2034 2566 -2018
rect 2532 -2298 2566 -2282
rect 2628 -2034 2662 -2018
rect 2628 -2298 2662 -2282
rect 2724 -2034 2758 -2018
rect 2724 -2298 2758 -2282
rect 2820 -2034 2854 -2018
rect 2820 -2298 2854 -2282
rect 2916 -2034 2950 -2018
rect 2916 -2298 2950 -2282
rect 1842 -2410 1876 -2382
rect 1940 -2342 2966 -2334
rect 1940 -2376 1956 -2342
rect 1990 -2376 2148 -2342
rect 2182 -2376 2340 -2342
rect 2374 -2376 2532 -2342
rect 2566 -2376 2724 -2342
rect 2758 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1940 -2384 2966 -2376
rect 3030 -2396 3064 -2382
rect 3329 -2396 3457 -1249
rect 1509 -2444 1882 -2410
rect 3030 -2444 3457 -2396
rect 321 -2478 417 -2444
rect 1447 -2478 1938 -2444
rect 2968 -2478 3457 -2444
rect 1686 -2575 3457 -2478
rect -1256 -2670 -1227 -2636
rect -1193 -2670 -1135 -2636
rect -1101 -2670 -1043 -2636
rect -1009 -2670 -951 -2636
rect -917 -2670 -859 -2636
rect -825 -2670 -767 -2636
rect -733 -2670 -675 -2636
rect -641 -2670 -583 -2636
rect -549 -2670 -491 -2636
rect -457 -2670 -399 -2636
rect -365 -2670 -37 -2636
rect -1239 -2764 -1181 -2670
rect -1239 -2798 -1227 -2764
rect -1193 -2798 -1181 -2764
rect -1239 -2815 -1181 -2798
rect -1100 -2716 -1054 -2670
rect -1100 -2750 -1088 -2716
rect -1100 -2784 -1054 -2750
rect -1100 -2818 -1088 -2784
rect -1100 -2834 -1054 -2818
rect -1020 -2716 -954 -2704
rect -1020 -2750 -1004 -2716
rect -970 -2750 -954 -2716
rect -1020 -2784 -954 -2750
rect -1020 -2818 -1004 -2784
rect -970 -2818 -954 -2784
rect -687 -2764 -629 -2670
rect -687 -2798 -675 -2764
rect -641 -2798 -629 -2764
rect -687 -2815 -629 -2798
rect -595 -2712 -533 -2670
rect -595 -2746 -573 -2712
rect -539 -2746 -533 -2712
rect -595 -2780 -533 -2746
rect -595 -2814 -573 -2780
rect -539 -2814 -533 -2780
rect -1020 -2830 -954 -2818
rect -595 -2830 -533 -2814
rect -492 -2712 -353 -2704
rect -492 -2746 -405 -2712
rect -371 -2746 -353 -2712
rect -492 -2780 -353 -2746
rect -492 -2814 -405 -2780
rect -371 -2814 -353 -2780
rect -492 -2830 -353 -2814
rect -165 -2713 -37 -2670
rect -165 -2814 1647 -2713
rect -165 -2816 1889 -2814
rect -2104 -2848 -1542 -2841
rect -3230 -2910 -3196 -2848
rect -2042 -2905 -1542 -2848
rect -3132 -2916 -2106 -2908
rect -3132 -2950 -3116 -2916
rect -3082 -2950 -2924 -2916
rect -2890 -2950 -2732 -2916
rect -2698 -2950 -2540 -2916
rect -2506 -2950 -2348 -2916
rect -2314 -2950 -2156 -2916
rect -2122 -2950 -2106 -2916
rect -3132 -2958 -2106 -2950
rect -2042 -2910 -2008 -2905
rect -3116 -3010 -3082 -2994
rect -3116 -3274 -3082 -3258
rect -3020 -3010 -2986 -2994
rect -3020 -3274 -2986 -3258
rect -2924 -3010 -2890 -2994
rect -2924 -3274 -2890 -3258
rect -2828 -3010 -2794 -2994
rect -2828 -3274 -2794 -3258
rect -2732 -3010 -2698 -2994
rect -2732 -3274 -2698 -3258
rect -2636 -3010 -2602 -2994
rect -2636 -3274 -2602 -3258
rect -2540 -3010 -2506 -2994
rect -2540 -3274 -2506 -3258
rect -2444 -3010 -2410 -2994
rect -2444 -3274 -2410 -3258
rect -2348 -3010 -2314 -2994
rect -2348 -3274 -2314 -3258
rect -2252 -3010 -2218 -2994
rect -2252 -3274 -2218 -3258
rect -2156 -3010 -2122 -2994
rect -2156 -3274 -2122 -3258
rect -3230 -3358 -3196 -3296
rect -2042 -3358 -2008 -3296
rect -3230 -3392 -3134 -3358
rect -2104 -3392 -2008 -3358
rect -1670 -3164 -1542 -2905
rect -1100 -2874 -1084 -2868
rect -1100 -2908 -1089 -2874
rect -1050 -2902 -1034 -2868
rect -1055 -2908 -1034 -2902
rect -1100 -2916 -1034 -2908
rect -1000 -2874 -954 -2830
rect -1000 -2908 -994 -2874
rect -960 -2908 -954 -2874
rect -1239 -2982 -1181 -2947
rect -1000 -2950 -954 -2908
rect -593 -2868 -526 -2864
rect -593 -2902 -576 -2868
rect -542 -2874 -526 -2868
rect -593 -2908 -574 -2902
rect -540 -2908 -526 -2874
rect -593 -2918 -526 -2908
rect -1239 -3016 -1227 -2982
rect -1193 -3016 -1181 -2982
rect -1239 -3075 -1181 -3016
rect -1239 -3109 -1227 -3075
rect -1193 -3109 -1181 -3075
rect -1239 -3164 -1181 -3109
rect -1670 -3180 -1181 -3164
rect -1096 -2968 -1054 -2952
rect -1096 -3002 -1088 -2968
rect -1096 -3036 -1054 -3002
rect -1096 -3070 -1088 -3036
rect -1096 -3104 -1054 -3070
rect -1096 -3138 -1088 -3104
rect -1096 -3180 -1054 -3138
rect -1020 -2968 -954 -2950
rect -1020 -3002 -1004 -2968
rect -970 -3002 -954 -2968
rect -1020 -3036 -954 -3002
rect -1020 -3070 -1004 -3036
rect -970 -3070 -954 -3036
rect -1020 -3104 -954 -3070
rect -1020 -3138 -1004 -3104
rect -970 -3138 -954 -3104
rect -1020 -3146 -954 -3138
rect -687 -2982 -629 -2947
rect -492 -2950 -458 -2830
rect -165 -2850 417 -2816
rect 1447 -2850 1938 -2816
rect 2968 -2850 3064 -2816
rect -424 -2902 -408 -2868
rect -374 -2875 -357 -2868
rect -424 -2909 -401 -2902
rect -367 -2909 -357 -2875
rect -424 -2918 -357 -2909
rect -165 -2882 355 -2850
rect -687 -3016 -675 -2982
rect -641 -3016 -629 -2982
rect -687 -3075 -629 -3016
rect -687 -3109 -675 -3075
rect -641 -3109 -629 -3075
rect -687 -3180 -629 -3109
rect -595 -2968 -539 -2952
rect -595 -3002 -573 -2968
rect -595 -3036 -539 -3002
rect -595 -3070 -573 -3036
rect -595 -3104 -539 -3070
rect -595 -3138 -573 -3104
rect -595 -3180 -539 -3138
rect -505 -2968 -439 -2950
rect -505 -3002 -489 -2968
rect -455 -3002 -439 -2968
rect -505 -3036 -439 -3002
rect -505 -3070 -490 -3036
rect -455 -3070 -439 -3036
rect -505 -3104 -439 -3070
rect -505 -3138 -489 -3104
rect -455 -3138 -439 -3104
rect -505 -3146 -439 -3138
rect -405 -2968 -353 -2952
rect -371 -3002 -353 -2968
rect -405 -3036 -353 -3002
rect -371 -3070 -353 -3036
rect -405 -3104 -353 -3070
rect -371 -3138 -353 -3104
rect -405 -3180 -353 -3138
rect -1670 -3214 -1227 -3180
rect -1193 -3214 -1135 -3180
rect -1101 -3214 -1043 -3180
rect -1009 -3214 -951 -3180
rect -917 -3214 -859 -3180
rect -825 -3214 -767 -3180
rect -733 -3214 -675 -3180
rect -641 -3214 -583 -3180
rect -549 -3214 -491 -3180
rect -457 -3214 -399 -3180
rect -365 -3214 -336 -3180
rect -1670 -3228 -1203 -3214
rect -3230 -3498 -3134 -3464
rect -2104 -3498 -2008 -3464
rect -3230 -3560 -3196 -3498
rect -2042 -3560 -2008 -3498
rect -3116 -3588 -3082 -3572
rect -3116 -3684 -3082 -3668
rect -3020 -3588 -2986 -3572
rect -3020 -3684 -2986 -3668
rect -2924 -3588 -2890 -3572
rect -2924 -3684 -2890 -3668
rect -2828 -3588 -2794 -3572
rect -2828 -3684 -2794 -3668
rect -2732 -3588 -2698 -3572
rect -2732 -3684 -2698 -3668
rect -2636 -3588 -2602 -3572
rect -2636 -3684 -2602 -3668
rect -2540 -3588 -2506 -3572
rect -2540 -3684 -2506 -3668
rect -2444 -3588 -2410 -3572
rect -2444 -3684 -2410 -3668
rect -2348 -3588 -2314 -3572
rect -2348 -3684 -2314 -3668
rect -2252 -3588 -2218 -3572
rect -2252 -3684 -2218 -3668
rect -2156 -3588 -2122 -3572
rect -2156 -3684 -2122 -3668
rect -3230 -3782 -3196 -3758
rect -3132 -3727 -2106 -3719
rect -3132 -3761 -3116 -3727
rect -3082 -3761 -2924 -3727
rect -2890 -3761 -2732 -3727
rect -2698 -3761 -2540 -3727
rect -2506 -3761 -2348 -3727
rect -2314 -3761 -2156 -3727
rect -2122 -3761 -2106 -3727
rect -3132 -3769 -2106 -3761
rect -3564 -3820 -3196 -3782
rect -2042 -3820 -2008 -3758
rect -3564 -3846 -3134 -3820
rect -3564 -5168 -3500 -3846
rect -3230 -3854 -3134 -3846
rect -2104 -3854 -2008 -3820
rect -3230 -4226 -3134 -4192
rect -2104 -4226 -2008 -4192
rect -3230 -4288 -3196 -4226
rect -2042 -4239 -2008 -4226
rect -1670 -4239 -1542 -3228
rect -687 -3285 -629 -3214
rect -687 -3319 -675 -3285
rect -641 -3319 -629 -3285
rect -687 -3378 -629 -3319
rect -687 -3412 -675 -3378
rect -641 -3412 -629 -3378
rect -687 -3447 -629 -3412
rect -595 -3256 -539 -3214
rect -595 -3290 -573 -3256
rect -595 -3324 -539 -3290
rect -595 -3358 -573 -3324
rect -595 -3392 -539 -3358
rect -595 -3426 -573 -3392
rect -595 -3442 -539 -3426
rect -505 -3256 -439 -3248
rect -505 -3290 -489 -3256
rect -455 -3290 -439 -3256
rect -505 -3324 -439 -3290
rect -505 -3358 -489 -3324
rect -455 -3358 -439 -3324
rect -505 -3392 -439 -3358
rect -505 -3426 -489 -3392
rect -455 -3426 -439 -3392
rect -505 -3444 -439 -3426
rect -405 -3256 -353 -3214
rect -371 -3290 -353 -3256
rect -405 -3324 -353 -3290
rect -371 -3358 -353 -3324
rect -405 -3392 -353 -3358
rect -371 -3426 -353 -3392
rect -405 -3442 -353 -3426
rect -593 -3492 -526 -3476
rect -593 -3526 -576 -3492
rect -542 -3526 -526 -3492
rect -593 -3530 -526 -3526
rect -492 -3564 -458 -3444
rect -424 -3487 -357 -3476
rect -424 -3492 -405 -3487
rect -424 -3526 -408 -3492
rect -371 -3521 -357 -3487
rect -374 -3526 -357 -3521
rect -687 -3596 -629 -3579
rect -687 -3630 -675 -3596
rect -641 -3630 -629 -3596
rect -687 -3724 -629 -3630
rect -595 -3580 -533 -3564
rect -595 -3614 -573 -3580
rect -539 -3614 -533 -3580
rect -595 -3648 -533 -3614
rect -595 -3682 -573 -3648
rect -539 -3682 -533 -3648
rect -595 -3724 -533 -3682
rect -492 -3580 -353 -3564
rect -492 -3590 -405 -3580
rect -458 -3614 -405 -3590
rect -371 -3614 -353 -3580
rect -458 -3624 -353 -3614
rect -492 -3648 -353 -3624
rect -492 -3682 -405 -3648
rect -371 -3682 -353 -3648
rect -492 -3690 -353 -3682
rect -165 -3724 -37 -2882
rect 321 -2912 355 -2882
rect 1509 -2882 1876 -2850
rect 419 -2909 1445 -2901
rect 419 -2943 435 -2909
rect 469 -2943 627 -2909
rect 661 -2943 819 -2909
rect 853 -2943 1011 -2909
rect 1045 -2943 1203 -2909
rect 1237 -2943 1395 -2909
rect 1429 -2943 1445 -2909
rect 419 -2951 1445 -2943
rect 1509 -2912 1543 -2882
rect 435 -3002 469 -2986
rect 435 -3098 469 -3082
rect 531 -3002 565 -2986
rect 531 -3098 565 -3082
rect 627 -3002 661 -2986
rect 627 -3098 661 -3082
rect 723 -3002 757 -2986
rect 723 -3098 757 -3082
rect 819 -3002 853 -2986
rect 819 -3098 853 -3082
rect 915 -3002 949 -2986
rect 915 -3098 949 -3082
rect 1011 -3002 1045 -2986
rect 1011 -3098 1045 -3082
rect 1107 -3002 1141 -2986
rect 1107 -3098 1141 -3082
rect 1203 -3002 1237 -2986
rect 1203 -3098 1237 -3082
rect 1299 -3002 1333 -2986
rect 1299 -3098 1333 -3082
rect 1395 -3002 1429 -2986
rect 1395 -3098 1429 -3082
rect 1842 -2912 1876 -2882
rect 321 -3172 355 -3110
rect 1615 -3008 1649 -2992
rect 1615 -3100 1649 -3084
rect 1703 -3008 1737 -2992
rect 1703 -3100 1737 -3084
rect 1509 -3172 1543 -3110
rect 1940 -2909 2966 -2901
rect 1940 -2943 1956 -2909
rect 1990 -2943 2148 -2909
rect 2182 -2943 2340 -2909
rect 2374 -2943 2532 -2909
rect 2566 -2943 2724 -2909
rect 2758 -2943 2916 -2909
rect 2950 -2943 2966 -2909
rect 1940 -2951 2966 -2943
rect 3030 -2912 3064 -2850
rect 1956 -3002 1990 -2986
rect 1956 -3098 1990 -3082
rect 2052 -3002 2086 -2986
rect 2052 -3098 2086 -3082
rect 2148 -3002 2182 -2986
rect 2148 -3098 2182 -3082
rect 2244 -3002 2278 -2986
rect 2244 -3098 2278 -3082
rect 2340 -3002 2374 -2986
rect 2340 -3098 2374 -3082
rect 2436 -3002 2470 -2986
rect 2436 -3098 2470 -3082
rect 2532 -3002 2566 -2986
rect 2532 -3098 2566 -3082
rect 2628 -3002 2662 -2986
rect 2628 -3098 2662 -3082
rect 2724 -3002 2758 -2986
rect 2724 -3098 2758 -3082
rect 2820 -3002 2854 -2986
rect 2820 -3098 2854 -3082
rect 2916 -3002 2950 -2986
rect 2916 -3098 2950 -3082
rect 1643 -3168 1659 -3134
rect 1693 -3168 1709 -3134
rect 321 -3206 417 -3172
rect 1447 -3206 1543 -3172
rect 1842 -3172 1876 -3110
rect 3030 -3172 3064 -3110
rect 1842 -3206 1938 -3172
rect 2968 -3206 3064 -3172
rect -704 -3758 -675 -3724
rect -641 -3758 -583 -3724
rect -549 -3758 -491 -3724
rect -457 -3758 -399 -3724
rect -365 -3758 -37 -3724
rect -687 -3852 -629 -3758
rect -687 -3886 -675 -3852
rect -641 -3886 -629 -3852
rect -687 -3903 -629 -3886
rect -548 -3804 -502 -3758
rect -548 -3838 -536 -3804
rect -548 -3872 -502 -3838
rect -548 -3906 -536 -3872
rect -548 -3922 -502 -3906
rect -468 -3804 -402 -3792
rect -468 -3838 -452 -3804
rect -418 -3838 -402 -3804
rect -468 -3872 -402 -3838
rect -468 -3906 -452 -3872
rect -418 -3906 -402 -3872
rect -468 -3918 -402 -3906
rect -548 -3961 -532 -3956
rect -548 -3995 -539 -3961
rect -498 -3990 -482 -3956
rect -505 -3995 -482 -3990
rect -548 -4004 -482 -3995
rect -2042 -4258 -1542 -4239
rect -687 -4070 -629 -4035
rect -448 -4038 -402 -3918
rect -687 -4104 -675 -4070
rect -641 -4104 -629 -4070
rect -687 -4163 -629 -4104
rect -687 -4197 -675 -4163
rect -641 -4197 -629 -4163
rect -687 -4258 -629 -4197
rect -2042 -4268 -629 -4258
rect -544 -4056 -502 -4040
rect -544 -4090 -536 -4056
rect -544 -4124 -502 -4090
rect -544 -4158 -536 -4124
rect -544 -4192 -502 -4158
rect -544 -4226 -536 -4192
rect -544 -4268 -502 -4226
rect -468 -4056 -402 -4038
rect -468 -4090 -452 -4056
rect -418 -4090 -402 -4056
rect -468 -4120 -402 -4090
rect -468 -4154 -453 -4120
rect -419 -4124 -402 -4120
rect -468 -4158 -452 -4154
rect -418 -4158 -402 -4124
rect -468 -4192 -402 -4158
rect -468 -4226 -452 -4192
rect -418 -4226 -402 -4192
rect -468 -4234 -402 -4226
rect -165 -4083 -37 -3758
rect 321 -3312 417 -3278
rect 1447 -3312 1543 -3278
rect 321 -3374 355 -3312
rect 1509 -3374 1543 -3312
rect 435 -3412 469 -3396
rect 435 -3676 469 -3660
rect 531 -3412 565 -3396
rect 531 -3676 565 -3660
rect 627 -3412 661 -3396
rect 627 -3676 661 -3660
rect 723 -3412 757 -3396
rect 723 -3676 757 -3660
rect 819 -3412 853 -3396
rect 819 -3676 853 -3660
rect 915 -3412 949 -3396
rect 915 -3676 949 -3660
rect 1011 -3412 1045 -3396
rect 1011 -3676 1045 -3660
rect 1107 -3412 1141 -3396
rect 1107 -3676 1141 -3660
rect 1203 -3412 1237 -3396
rect 1203 -3676 1237 -3660
rect 1299 -3412 1333 -3396
rect 1299 -3676 1333 -3660
rect 1395 -3412 1429 -3396
rect 1395 -3676 1429 -3660
rect 321 -3822 355 -3760
rect 419 -3720 1445 -3712
rect 419 -3754 435 -3720
rect 469 -3754 627 -3720
rect 661 -3754 819 -3720
rect 853 -3754 1011 -3720
rect 1045 -3754 1203 -3720
rect 1237 -3754 1395 -3720
rect 1429 -3754 1445 -3720
rect 419 -3762 1445 -3754
rect 1509 -3788 1543 -3760
rect 1842 -3312 1938 -3278
rect 2968 -3312 3064 -3278
rect 1842 -3374 1876 -3312
rect 3030 -3374 3064 -3312
rect 1956 -3412 1990 -3396
rect 1956 -3676 1990 -3660
rect 2052 -3412 2086 -3396
rect 2052 -3676 2086 -3660
rect 2148 -3412 2182 -3396
rect 2148 -3676 2182 -3660
rect 2244 -3412 2278 -3396
rect 2244 -3676 2278 -3660
rect 2340 -3412 2374 -3396
rect 2340 -3676 2374 -3660
rect 2436 -3412 2470 -3396
rect 2436 -3676 2470 -3660
rect 2532 -3412 2566 -3396
rect 2532 -3676 2566 -3660
rect 2628 -3412 2662 -3396
rect 2628 -3676 2662 -3660
rect 2724 -3412 2758 -3396
rect 2724 -3676 2758 -3660
rect 2820 -3412 2854 -3396
rect 2820 -3676 2854 -3660
rect 2916 -3412 2950 -3396
rect 2916 -3676 2950 -3660
rect 1842 -3788 1876 -3760
rect 1940 -3720 2966 -3712
rect 1940 -3754 1956 -3720
rect 1990 -3754 2148 -3720
rect 2182 -3754 2340 -3720
rect 2374 -3754 2532 -3720
rect 2566 -3754 2724 -3720
rect 2758 -3754 2916 -3720
rect 2950 -3754 2966 -3720
rect 1940 -3762 2966 -3754
rect 3030 -3779 3064 -3760
rect 3329 -3779 3457 -2575
rect 1509 -3822 1882 -3788
rect 3030 -3822 3457 -3779
rect 321 -3856 417 -3822
rect 1447 -3856 1938 -3822
rect 2968 -3856 3457 -3822
rect 1686 -3959 3457 -3856
rect -165 -4192 1661 -4083
rect -165 -4194 1889 -4192
rect -165 -4228 417 -4194
rect 1447 -4228 1938 -4194
rect 2968 -4228 3064 -4194
rect -165 -4264 355 -4228
rect -3132 -4294 -2106 -4286
rect -3132 -4328 -3116 -4294
rect -3082 -4328 -2924 -4294
rect -2890 -4328 -2732 -4294
rect -2698 -4328 -2540 -4294
rect -2506 -4328 -2348 -4294
rect -2314 -4328 -2156 -4294
rect -2122 -4328 -2106 -4294
rect -3132 -4336 -2106 -4328
rect -2042 -4288 -675 -4268
rect -3116 -4388 -3082 -4372
rect -3116 -4652 -3082 -4636
rect -3020 -4388 -2986 -4372
rect -3020 -4652 -2986 -4636
rect -2924 -4388 -2890 -4372
rect -2924 -4652 -2890 -4636
rect -2828 -4388 -2794 -4372
rect -2828 -4652 -2794 -4636
rect -2732 -4388 -2698 -4372
rect -2732 -4652 -2698 -4636
rect -2636 -4388 -2602 -4372
rect -2636 -4652 -2602 -4636
rect -2540 -4388 -2506 -4372
rect -2540 -4652 -2506 -4636
rect -2444 -4388 -2410 -4372
rect -2444 -4652 -2410 -4636
rect -2348 -4388 -2314 -4372
rect -2348 -4652 -2314 -4636
rect -2252 -4388 -2218 -4372
rect -2252 -4652 -2218 -4636
rect -2156 -4388 -2122 -4372
rect -2156 -4652 -2122 -4636
rect -3230 -4736 -3196 -4674
rect -2008 -4302 -675 -4288
rect -641 -4302 -583 -4268
rect -549 -4302 -491 -4268
rect -457 -4302 -399 -4268
rect -365 -4302 -336 -4268
rect -2008 -4303 -629 -4302
rect -1670 -4322 -629 -4303
rect -1670 -4324 -1542 -4322
rect -687 -4373 -629 -4322
rect -687 -4407 -675 -4373
rect -641 -4407 -629 -4373
rect -687 -4466 -629 -4407
rect -687 -4500 -675 -4466
rect -641 -4500 -629 -4466
rect -687 -4535 -629 -4500
rect -544 -4344 -502 -4302
rect -544 -4378 -536 -4344
rect -544 -4412 -502 -4378
rect -544 -4446 -536 -4412
rect -544 -4480 -502 -4446
rect -544 -4514 -536 -4480
rect -544 -4530 -502 -4514
rect -468 -4344 -402 -4336
rect -468 -4378 -452 -4344
rect -418 -4378 -402 -4344
rect -468 -4412 -402 -4378
rect -468 -4452 -452 -4412
rect -418 -4452 -402 -4412
rect -468 -4480 -402 -4452
rect -468 -4514 -452 -4480
rect -418 -4514 -402 -4480
rect -468 -4532 -402 -4514
rect -548 -4574 -482 -4566
rect -548 -4608 -540 -4574
rect -506 -4580 -482 -4574
rect -548 -4614 -532 -4608
rect -498 -4614 -482 -4580
rect -548 -4664 -502 -4648
rect -448 -4652 -402 -4532
rect -2042 -4736 -2008 -4674
rect -3230 -4770 -3134 -4736
rect -2104 -4770 -2008 -4736
rect -687 -4684 -629 -4667
rect -687 -4718 -675 -4684
rect -641 -4718 -629 -4684
rect -687 -4812 -629 -4718
rect -548 -4698 -536 -4664
rect -548 -4732 -502 -4698
rect -548 -4766 -536 -4732
rect -548 -4812 -502 -4766
rect -468 -4664 -402 -4652
rect -468 -4698 -452 -4664
rect -418 -4698 -402 -4664
rect -468 -4732 -402 -4698
rect -468 -4766 -452 -4732
rect -418 -4766 -402 -4732
rect -468 -4778 -402 -4766
rect -165 -4812 -37 -4264
rect 321 -4290 355 -4264
rect 1509 -4260 1876 -4228
rect 419 -4287 1445 -4279
rect 419 -4321 435 -4287
rect 469 -4321 627 -4287
rect 661 -4321 819 -4287
rect 853 -4321 1011 -4287
rect 1045 -4321 1203 -4287
rect 1237 -4321 1395 -4287
rect 1429 -4321 1445 -4287
rect 419 -4329 1445 -4321
rect 1509 -4290 1543 -4260
rect 435 -4380 469 -4364
rect 435 -4476 469 -4460
rect 531 -4380 565 -4364
rect 531 -4476 565 -4460
rect 627 -4380 661 -4364
rect 627 -4476 661 -4460
rect 723 -4380 757 -4364
rect 723 -4476 757 -4460
rect 819 -4380 853 -4364
rect 819 -4476 853 -4460
rect 915 -4380 949 -4364
rect 915 -4476 949 -4460
rect 1011 -4380 1045 -4364
rect 1011 -4476 1045 -4460
rect 1107 -4380 1141 -4364
rect 1107 -4476 1141 -4460
rect 1203 -4380 1237 -4364
rect 1203 -4476 1237 -4460
rect 1299 -4380 1333 -4364
rect 1299 -4476 1333 -4460
rect 1395 -4380 1429 -4364
rect 1395 -4476 1429 -4460
rect 1842 -4290 1876 -4260
rect 321 -4550 355 -4488
rect 1615 -4386 1649 -4370
rect 1615 -4478 1649 -4462
rect 1703 -4386 1737 -4370
rect 1703 -4478 1737 -4462
rect 1509 -4550 1543 -4488
rect 1940 -4287 2966 -4279
rect 1940 -4321 1956 -4287
rect 1990 -4321 2148 -4287
rect 2182 -4321 2340 -4287
rect 2374 -4321 2532 -4287
rect 2566 -4321 2724 -4287
rect 2758 -4321 2916 -4287
rect 2950 -4321 2966 -4287
rect 1940 -4329 2966 -4321
rect 3030 -4290 3064 -4228
rect 1956 -4380 1990 -4364
rect 1956 -4476 1990 -4460
rect 2052 -4380 2086 -4364
rect 2052 -4476 2086 -4460
rect 2148 -4380 2182 -4364
rect 2148 -4476 2182 -4460
rect 2244 -4380 2278 -4364
rect 2244 -4476 2278 -4460
rect 2340 -4380 2374 -4364
rect 2340 -4476 2374 -4460
rect 2436 -4380 2470 -4364
rect 2436 -4476 2470 -4460
rect 2532 -4380 2566 -4364
rect 2532 -4476 2566 -4460
rect 2628 -4380 2662 -4364
rect 2628 -4476 2662 -4460
rect 2724 -4380 2758 -4364
rect 2724 -4476 2758 -4460
rect 2820 -4380 2854 -4364
rect 2820 -4476 2854 -4460
rect 2916 -4380 2950 -4364
rect 2916 -4476 2950 -4460
rect 1643 -4546 1659 -4512
rect 1693 -4546 1709 -4512
rect 321 -4584 417 -4550
rect 1447 -4584 1543 -4550
rect 1842 -4550 1876 -4488
rect 3030 -4550 3064 -4488
rect 1842 -4584 1938 -4550
rect 2968 -4584 3064 -4550
rect -3230 -4876 -3134 -4842
rect -2104 -4876 -2008 -4842
rect -704 -4846 -675 -4812
rect -641 -4846 -583 -4812
rect -549 -4846 -491 -4812
rect -457 -4846 -399 -4812
rect -365 -4846 -37 -4812
rect -3230 -4938 -3196 -4876
rect -2042 -4938 -2008 -4876
rect -3116 -4966 -3082 -4950
rect -3116 -5062 -3082 -5046
rect -3020 -4966 -2986 -4950
rect -3020 -5062 -2986 -5046
rect -2924 -4966 -2890 -4950
rect -2924 -5062 -2890 -5046
rect -2828 -4966 -2794 -4950
rect -2828 -5062 -2794 -5046
rect -2732 -4966 -2698 -4950
rect -2732 -5062 -2698 -5046
rect -2636 -4966 -2602 -4950
rect -2636 -5062 -2602 -5046
rect -2540 -4966 -2506 -4950
rect -2540 -5062 -2506 -5046
rect -2444 -4966 -2410 -4950
rect -2444 -5062 -2410 -5046
rect -2348 -4966 -2314 -4950
rect -2348 -5062 -2314 -5046
rect -2252 -4966 -2218 -4950
rect -2252 -5062 -2218 -5046
rect -2156 -4966 -2122 -4950
rect -2156 -5062 -2122 -5046
rect -3230 -5168 -3196 -5136
rect -3132 -5105 -2106 -5097
rect -3132 -5139 -3116 -5105
rect -3082 -5139 -2924 -5105
rect -2890 -5139 -2732 -5105
rect -2698 -5139 -2540 -5105
rect -2506 -5139 -2348 -5105
rect -2314 -5139 -2156 -5105
rect -2122 -5139 -2106 -5105
rect -3132 -5147 -2106 -5139
rect -3564 -5198 -3196 -5168
rect -2042 -5198 -2008 -5136
rect -3564 -5232 -3134 -5198
rect -2104 -5232 -2008 -5198
rect -3564 -5564 -3500 -5232
rect -165 -5564 -37 -4846
rect 321 -4690 417 -4656
rect 1447 -4690 1543 -4656
rect 321 -4752 355 -4690
rect 1509 -4752 1543 -4690
rect 435 -4790 469 -4774
rect 435 -5054 469 -5038
rect 531 -4790 565 -4774
rect 531 -5054 565 -5038
rect 627 -4790 661 -4774
rect 627 -5054 661 -5038
rect 723 -4790 757 -4774
rect 723 -5054 757 -5038
rect 819 -4790 853 -4774
rect 819 -5054 853 -5038
rect 915 -4790 949 -4774
rect 915 -5054 949 -5038
rect 1011 -4790 1045 -4774
rect 1011 -5054 1045 -5038
rect 1107 -4790 1141 -4774
rect 1107 -5054 1141 -5038
rect 1203 -4790 1237 -4774
rect 1203 -5054 1237 -5038
rect 1299 -4790 1333 -4774
rect 1299 -5054 1333 -5038
rect 1395 -4790 1429 -4774
rect 1395 -5054 1429 -5038
rect 321 -5200 355 -5138
rect 419 -5098 1445 -5090
rect 419 -5132 435 -5098
rect 469 -5132 627 -5098
rect 661 -5132 819 -5098
rect 853 -5132 1011 -5098
rect 1045 -5132 1203 -5098
rect 1237 -5132 1395 -5098
rect 1429 -5132 1445 -5098
rect 419 -5140 1445 -5132
rect 1509 -5166 1543 -5138
rect 1842 -4690 1938 -4656
rect 2968 -4690 3064 -4656
rect 1842 -4752 1876 -4690
rect 3030 -4752 3064 -4690
rect 1956 -4790 1990 -4774
rect 1956 -5054 1990 -5038
rect 2052 -4790 2086 -4774
rect 2052 -5054 2086 -5038
rect 2148 -4790 2182 -4774
rect 2148 -5054 2182 -5038
rect 2244 -4790 2278 -4774
rect 2244 -5054 2278 -5038
rect 2340 -4790 2374 -4774
rect 2340 -5054 2374 -5038
rect 2436 -4790 2470 -4774
rect 2436 -5054 2470 -5038
rect 2532 -4790 2566 -4774
rect 2532 -5054 2566 -5038
rect 2628 -4790 2662 -4774
rect 2628 -5054 2662 -5038
rect 2724 -4790 2758 -4774
rect 2724 -5054 2758 -5038
rect 2820 -4790 2854 -4774
rect 2820 -5054 2854 -5038
rect 2916 -4790 2950 -4774
rect 2916 -5054 2950 -5038
rect 1842 -5166 1876 -5138
rect 1940 -5098 2966 -5090
rect 1940 -5132 1956 -5098
rect 1990 -5132 2148 -5098
rect 2182 -5132 2340 -5098
rect 2374 -5132 2532 -5098
rect 2566 -5132 2724 -5098
rect 2758 -5132 2916 -5098
rect 2950 -5132 2966 -5098
rect 1940 -5140 2966 -5132
rect 1509 -5200 1882 -5166
rect 3030 -5200 3064 -5138
rect 321 -5234 417 -5200
rect 1447 -5234 1938 -5200
rect 2968 -5227 3064 -5200
rect 3329 -5227 3457 -3959
rect 2968 -5234 3457 -5227
rect 1661 -5355 3457 -5234
rect -3827 -5692 3675 -5564
<< viali >>
rect -2348 -204 -2314 -201
rect -2348 -235 -2314 -204
rect -2156 -238 -2122 -204
rect -3116 -546 -3082 -298
rect -3020 -546 -2986 -298
rect -2924 -546 -2890 -298
rect -2828 -546 -2794 -298
rect -2732 -546 -2698 -298
rect -2636 -546 -2602 -298
rect -2540 -546 -2506 -298
rect -2444 -546 -2410 -298
rect -2348 -546 -2314 -298
rect -2252 -546 -2218 -298
rect -2156 -546 -2122 -298
rect -3116 -956 -3082 -876
rect -3020 -956 -2986 -876
rect -2924 -956 -2890 -876
rect -2828 -956 -2794 -876
rect -2732 -956 -2698 -876
rect -2636 -956 -2602 -876
rect -2540 -956 -2506 -876
rect -2444 -956 -2410 -876
rect -2348 -956 -2314 -876
rect -2252 -956 -2218 -876
rect -2156 -956 -2122 -876
rect -2345 -1049 -2314 -1019
rect -2314 -1049 -2311 -1019
rect -2155 -1049 -2122 -1016
rect -2122 -1049 -2121 -1016
rect -2345 -1053 -2311 -1049
rect -2155 -1050 -2121 -1049
rect -951 -494 -917 -460
rect -859 -494 -825 -460
rect -767 -494 -733 -460
rect -675 -494 -641 -460
rect -583 -494 -549 -460
rect -491 -494 -457 -460
rect -399 -494 -365 -460
rect 435 -231 469 -197
rect 1395 -231 1429 -197
rect 435 -370 469 -290
rect 531 -370 565 -290
rect 627 -370 661 -290
rect 723 -370 757 -290
rect 819 -370 853 -290
rect 915 -370 949 -290
rect 1011 -370 1045 -290
rect 1107 -370 1141 -290
rect 1203 -370 1237 -290
rect 1299 -370 1333 -290
rect 1395 -370 1429 -290
rect 1509 -385 1543 -285
rect 1615 -372 1649 -296
rect 1703 -372 1737 -296
rect 1956 -231 1990 -197
rect 2916 -231 2950 -197
rect 1956 -370 1990 -290
rect 2052 -370 2086 -290
rect 2148 -370 2182 -290
rect 2244 -370 2278 -290
rect 2340 -370 2374 -290
rect 2436 -370 2470 -290
rect 2532 -370 2566 -290
rect 2628 -370 2662 -290
rect 2724 -370 2758 -290
rect 2820 -370 2854 -290
rect 2916 -370 2950 -290
rect 1659 -456 1693 -422
rect -822 -608 -788 -603
rect -822 -637 -820 -608
rect -820 -637 -788 -608
rect -905 -726 -900 -698
rect -900 -726 -871 -698
rect -905 -732 -871 -726
rect -452 -608 -418 -594
rect -452 -628 -418 -608
rect -538 -726 -532 -700
rect -532 -726 -504 -700
rect -538 -734 -504 -726
rect -951 -1038 -917 -1004
rect -859 -1038 -825 -1004
rect -767 -1038 -733 -1004
rect -675 -1038 -641 -1004
rect -583 -1038 -549 -1004
rect -491 -1038 -457 -1004
rect -399 -1038 -365 -1004
rect -453 -1216 -419 -1197
rect -453 -1231 -452 -1216
rect -452 -1231 -419 -1216
rect -534 -1316 -500 -1312
rect -534 -1346 -532 -1316
rect -532 -1346 -500 -1316
rect -2348 -1572 -2314 -1538
rect -2156 -1572 -2122 -1538
rect -3116 -1880 -3082 -1632
rect -3020 -1880 -2986 -1632
rect -2924 -1880 -2890 -1632
rect -2828 -1880 -2794 -1632
rect -2732 -1880 -2698 -1632
rect -2636 -1880 -2602 -1632
rect -2540 -1880 -2506 -1632
rect -2444 -1880 -2410 -1632
rect -2348 -1880 -2314 -1632
rect -2252 -1880 -2218 -1632
rect -2156 -1880 -2122 -1632
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect 435 -1042 469 -1008
rect 1395 -1042 1429 -1008
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect 1956 -1042 1990 -1008
rect 2916 -1042 2950 -1008
rect -675 -1582 -641 -1548
rect -583 -1582 -549 -1548
rect -491 -1582 -457 -1548
rect -399 -1582 -365 -1548
rect -469 -1710 -435 -1676
rect -582 -1814 -576 -1784
rect -576 -1814 -548 -1784
rect -582 -1818 -548 -1814
rect -408 -1814 -374 -1785
rect -408 -1819 -374 -1814
rect -3116 -2290 -3082 -2210
rect -3020 -2290 -2986 -2210
rect -2924 -2290 -2890 -2210
rect -2828 -2290 -2794 -2210
rect -2732 -2290 -2698 -2210
rect -2636 -2290 -2602 -2210
rect -2540 -2290 -2506 -2210
rect -2444 -2290 -2410 -2210
rect -2348 -2290 -2314 -2210
rect -2252 -2290 -2218 -2210
rect -2156 -2290 -2122 -2210
rect -2348 -2383 -2314 -2349
rect -2156 -2383 -2122 -2349
rect -1227 -2126 -1193 -2092
rect -1135 -2126 -1101 -2092
rect -1043 -2126 -1009 -2092
rect -951 -2126 -917 -2092
rect -859 -2126 -825 -2092
rect -767 -2126 -733 -2092
rect -675 -2126 -641 -2092
rect -583 -2126 -549 -2092
rect -491 -2126 -457 -2092
rect -399 -2126 -365 -2092
rect -1004 -2270 -970 -2236
rect -1091 -2404 -1057 -2398
rect -1091 -2432 -1084 -2404
rect -1084 -2432 -1057 -2404
rect -489 -2304 -455 -2270
rect -583 -2404 -549 -2398
rect -583 -2432 -576 -2404
rect -576 -2432 -549 -2404
rect -402 -2404 -368 -2395
rect -402 -2429 -374 -2404
rect -374 -2429 -368 -2404
rect 435 -1565 469 -1531
rect 1395 -1565 1429 -1531
rect 435 -1704 469 -1624
rect 531 -1704 565 -1624
rect 627 -1704 661 -1624
rect 723 -1704 757 -1624
rect 819 -1704 853 -1624
rect 915 -1704 949 -1624
rect 1011 -1704 1045 -1624
rect 1107 -1704 1141 -1624
rect 1203 -1704 1237 -1624
rect 1299 -1704 1333 -1624
rect 1395 -1704 1429 -1624
rect 1509 -1719 1543 -1619
rect 1615 -1706 1649 -1630
rect 1703 -1706 1737 -1630
rect 1956 -1565 1990 -1531
rect 2916 -1565 2950 -1531
rect 1956 -1704 1990 -1624
rect 2052 -1704 2086 -1624
rect 2148 -1704 2182 -1624
rect 2244 -1704 2278 -1624
rect 2340 -1704 2374 -1624
rect 2436 -1704 2470 -1624
rect 2532 -1704 2566 -1624
rect 2628 -1704 2662 -1624
rect 2724 -1704 2758 -1624
rect 2820 -1704 2854 -1624
rect 2916 -1704 2950 -1624
rect 1659 -1790 1693 -1756
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 435 -2376 469 -2342
rect 1395 -2376 1429 -2342
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
rect 1956 -2376 1990 -2342
rect 2916 -2376 2950 -2342
rect -1227 -2670 -1193 -2636
rect -1135 -2670 -1101 -2636
rect -1043 -2670 -1009 -2636
rect -951 -2670 -917 -2636
rect -859 -2670 -825 -2636
rect -767 -2670 -733 -2636
rect -675 -2670 -641 -2636
rect -583 -2670 -549 -2636
rect -491 -2670 -457 -2636
rect -399 -2670 -365 -2636
rect -2348 -2950 -2314 -2916
rect -2156 -2950 -2122 -2916
rect -3116 -3258 -3082 -3010
rect -3020 -3258 -2986 -3010
rect -2924 -3258 -2890 -3010
rect -2828 -3258 -2794 -3010
rect -2732 -3258 -2698 -3010
rect -2636 -3258 -2602 -3010
rect -2540 -3258 -2506 -3010
rect -2444 -3258 -2410 -3010
rect -2348 -3258 -2314 -3010
rect -2252 -3258 -2218 -3010
rect -2156 -3258 -2122 -3010
rect -1089 -2902 -1084 -2874
rect -1084 -2902 -1055 -2874
rect -1089 -2908 -1055 -2902
rect -994 -2908 -960 -2874
rect -574 -2902 -542 -2874
rect -542 -2902 -540 -2874
rect -574 -2908 -540 -2902
rect -401 -2902 -374 -2875
rect -374 -2902 -367 -2875
rect -401 -2909 -367 -2902
rect -490 -3070 -489 -3036
rect -489 -3070 -456 -3036
rect -1227 -3214 -1193 -3180
rect -1135 -3214 -1101 -3180
rect -1043 -3214 -1009 -3180
rect -951 -3214 -917 -3180
rect -859 -3214 -825 -3180
rect -767 -3214 -733 -3180
rect -675 -3214 -641 -3180
rect -583 -3214 -549 -3180
rect -491 -3214 -457 -3180
rect -399 -3214 -365 -3180
rect -3116 -3668 -3082 -3588
rect -3020 -3668 -2986 -3588
rect -2924 -3668 -2890 -3588
rect -2828 -3668 -2794 -3588
rect -2732 -3668 -2698 -3588
rect -2636 -3668 -2602 -3588
rect -2540 -3668 -2506 -3588
rect -2444 -3668 -2410 -3588
rect -2348 -3668 -2314 -3588
rect -2252 -3668 -2218 -3588
rect -2156 -3668 -2122 -3588
rect -2348 -3761 -2314 -3727
rect -2156 -3761 -2122 -3727
rect -576 -3526 -542 -3492
rect -405 -3492 -371 -3487
rect -405 -3521 -374 -3492
rect -374 -3521 -371 -3492
rect -492 -3624 -458 -3590
rect 435 -2943 469 -2909
rect 1395 -2943 1429 -2909
rect 435 -3082 469 -3002
rect 531 -3082 565 -3002
rect 627 -3082 661 -3002
rect 723 -3082 757 -3002
rect 819 -3082 853 -3002
rect 915 -3082 949 -3002
rect 1011 -3082 1045 -3002
rect 1107 -3082 1141 -3002
rect 1203 -3082 1237 -3002
rect 1299 -3082 1333 -3002
rect 1395 -3082 1429 -3002
rect 1509 -3097 1543 -2997
rect 1615 -3084 1649 -3008
rect 1703 -3084 1737 -3008
rect 1956 -2943 1990 -2909
rect 2916 -2943 2950 -2909
rect 1956 -3082 1990 -3002
rect 2052 -3082 2086 -3002
rect 2148 -3082 2182 -3002
rect 2244 -3082 2278 -3002
rect 2340 -3082 2374 -3002
rect 2436 -3082 2470 -3002
rect 2532 -3082 2566 -3002
rect 2628 -3082 2662 -3002
rect 2724 -3082 2758 -3002
rect 2820 -3082 2854 -3002
rect 2916 -3082 2950 -3002
rect 1659 -3168 1693 -3134
rect -675 -3758 -641 -3724
rect -583 -3758 -549 -3724
rect -491 -3758 -457 -3724
rect -399 -3758 -365 -3724
rect -539 -3990 -532 -3961
rect -532 -3990 -505 -3961
rect -539 -3995 -505 -3990
rect -453 -4124 -419 -4120
rect -453 -4154 -452 -4124
rect -452 -4154 -419 -4124
rect 435 -3660 469 -3412
rect 531 -3660 565 -3412
rect 627 -3660 661 -3412
rect 723 -3660 757 -3412
rect 819 -3660 853 -3412
rect 915 -3660 949 -3412
rect 1011 -3660 1045 -3412
rect 1107 -3660 1141 -3412
rect 1203 -3660 1237 -3412
rect 1299 -3660 1333 -3412
rect 1395 -3660 1429 -3412
rect 435 -3754 469 -3720
rect 1395 -3754 1429 -3720
rect 1956 -3660 1990 -3412
rect 2052 -3660 2086 -3412
rect 2148 -3660 2182 -3412
rect 2244 -3660 2278 -3412
rect 2340 -3660 2374 -3412
rect 2436 -3660 2470 -3412
rect 2532 -3660 2566 -3412
rect 2628 -3660 2662 -3412
rect 2724 -3660 2758 -3412
rect 2820 -3660 2854 -3412
rect 2916 -3660 2950 -3412
rect 1956 -3754 1990 -3720
rect 2916 -3754 2950 -3720
rect -2348 -4328 -2314 -4294
rect -2156 -4328 -2122 -4294
rect -3116 -4636 -3082 -4388
rect -3020 -4636 -2986 -4388
rect -2924 -4636 -2890 -4388
rect -2828 -4636 -2794 -4388
rect -2732 -4636 -2698 -4388
rect -2636 -4636 -2602 -4388
rect -2540 -4636 -2506 -4388
rect -2444 -4636 -2410 -4388
rect -2348 -4636 -2314 -4388
rect -2252 -4636 -2218 -4388
rect -2156 -4636 -2122 -4388
rect -675 -4302 -641 -4268
rect -583 -4302 -549 -4268
rect -491 -4302 -457 -4268
rect -399 -4302 -365 -4268
rect -452 -4446 -418 -4418
rect -452 -4452 -418 -4446
rect -540 -4580 -506 -4574
rect -540 -4608 -532 -4580
rect -532 -4608 -506 -4580
rect 435 -4321 469 -4287
rect 1395 -4321 1429 -4287
rect 435 -4460 469 -4380
rect 531 -4460 565 -4380
rect 627 -4460 661 -4380
rect 723 -4460 757 -4380
rect 819 -4460 853 -4380
rect 915 -4460 949 -4380
rect 1011 -4460 1045 -4380
rect 1107 -4460 1141 -4380
rect 1203 -4460 1237 -4380
rect 1299 -4460 1333 -4380
rect 1395 -4460 1429 -4380
rect 1509 -4475 1543 -4375
rect 1615 -4462 1649 -4386
rect 1703 -4462 1737 -4386
rect 1956 -4321 1990 -4287
rect 2916 -4321 2950 -4287
rect 1956 -4460 1990 -4380
rect 2052 -4460 2086 -4380
rect 2148 -4460 2182 -4380
rect 2244 -4460 2278 -4380
rect 2340 -4460 2374 -4380
rect 2436 -4460 2470 -4380
rect 2532 -4460 2566 -4380
rect 2628 -4460 2662 -4380
rect 2724 -4460 2758 -4380
rect 2820 -4460 2854 -4380
rect 2916 -4460 2950 -4380
rect 1659 -4546 1693 -4512
rect -675 -4846 -641 -4812
rect -583 -4846 -549 -4812
rect -491 -4846 -457 -4812
rect -399 -4846 -365 -4812
rect -3116 -5046 -3082 -4966
rect -3020 -5046 -2986 -4966
rect -2924 -5046 -2890 -4966
rect -2828 -5046 -2794 -4966
rect -2732 -5046 -2698 -4966
rect -2636 -5046 -2602 -4966
rect -2540 -5046 -2506 -4966
rect -2444 -5046 -2410 -4966
rect -2348 -5046 -2314 -4966
rect -2252 -5046 -2218 -4966
rect -2156 -5046 -2122 -4966
rect -2348 -5139 -2314 -5105
rect -2156 -5139 -2122 -5105
rect 435 -5038 469 -4790
rect 531 -5038 565 -4790
rect 627 -5038 661 -4790
rect 723 -5038 757 -4790
rect 819 -5038 853 -4790
rect 915 -5038 949 -4790
rect 1011 -5038 1045 -4790
rect 1107 -5038 1141 -4790
rect 1203 -5038 1237 -4790
rect 1299 -5038 1333 -4790
rect 1395 -5038 1429 -4790
rect 435 -5132 469 -5098
rect 1395 -5132 1429 -5098
rect 1956 -5038 1990 -4790
rect 2052 -5038 2086 -4790
rect 2148 -5038 2182 -4790
rect 2244 -5038 2278 -4790
rect 2340 -5038 2374 -4790
rect 2436 -5038 2470 -4790
rect 2532 -5038 2566 -4790
rect 2628 -5038 2662 -4790
rect 2724 -5038 2758 -4790
rect 2820 -5038 2854 -4790
rect 2916 -5038 2950 -4790
rect 1956 -5132 1990 -5098
rect 2916 -5132 2950 -5098
<< metal1 >>
rect -3266 -136 -2218 -102
rect -1597 -121 -1587 -69
rect -1535 -121 -914 -69
rect -862 -121 -852 -69
rect -3266 -690 -3232 -136
rect -3020 -286 -2986 -136
rect -2828 -286 -2794 -136
rect -2636 -286 -2602 -136
rect -2444 -286 -2410 -136
rect -2367 -247 -2357 -195
rect -2305 -247 -2295 -195
rect -2252 -286 -2218 -136
rect 285 -136 1333 -102
rect -2173 -246 -2163 -194
rect -2111 -246 -2101 -194
rect -1952 -246 -1942 -194
rect -1890 -246 -1416 -194
rect -1364 -246 -1354 -194
rect -3122 -298 -3076 -286
rect -3122 -546 -3116 -298
rect -3082 -546 -3076 -298
rect -3122 -558 -3076 -546
rect -3026 -298 -2980 -286
rect -3026 -546 -3020 -298
rect -2986 -546 -2980 -298
rect -3026 -558 -2980 -546
rect -2930 -298 -2884 -286
rect -2930 -546 -2924 -298
rect -2890 -546 -2884 -298
rect -2930 -558 -2884 -546
rect -2834 -298 -2788 -286
rect -2834 -546 -2828 -298
rect -2794 -546 -2788 -298
rect -2834 -558 -2788 -546
rect -2738 -298 -2692 -286
rect -2738 -546 -2732 -298
rect -2698 -546 -2692 -298
rect -2738 -558 -2692 -546
rect -2642 -298 -2596 -286
rect -2642 -546 -2636 -298
rect -2602 -546 -2596 -298
rect -2642 -558 -2596 -546
rect -2546 -298 -2500 -286
rect -2546 -546 -2540 -298
rect -2506 -546 -2500 -298
rect -2546 -558 -2500 -546
rect -2450 -298 -2404 -286
rect -2450 -546 -2444 -298
rect -2410 -546 -2404 -298
rect -2450 -558 -2404 -546
rect -2354 -298 -2308 -286
rect -2354 -546 -2348 -298
rect -2314 -546 -2308 -298
rect -2354 -558 -2308 -546
rect -2258 -298 -2212 -286
rect -2258 -546 -2252 -298
rect -2218 -546 -2212 -298
rect -2258 -558 -2212 -546
rect -2162 -298 -2116 -286
rect -2162 -546 -2156 -298
rect -2122 -546 -2116 -298
rect -980 -460 -336 -429
rect -980 -494 -951 -460
rect -917 -494 -859 -460
rect -825 -494 -767 -460
rect -733 -494 -675 -460
rect -641 -494 -583 -460
rect -549 -494 -491 -460
rect -457 -494 -399 -460
rect -365 -494 -336 -460
rect -980 -525 -336 -494
rect 285 -503 319 -136
rect 415 -238 425 -186
rect 477 -238 487 -186
rect 531 -278 565 -136
rect 723 -278 757 -136
rect 915 -278 949 -136
rect 1107 -278 1141 -136
rect 1299 -278 1333 -136
rect 1806 -136 2854 -102
rect 1377 -240 1387 -188
rect 1439 -240 1449 -188
rect 429 -290 475 -278
rect 429 -370 435 -290
rect 469 -370 475 -290
rect 429 -382 475 -370
rect 525 -290 571 -278
rect 525 -370 531 -290
rect 565 -370 571 -290
rect 525 -382 571 -370
rect 621 -290 667 -278
rect 621 -370 627 -290
rect 661 -370 667 -290
rect 621 -382 667 -370
rect 717 -290 763 -278
rect 717 -370 723 -290
rect 757 -370 763 -290
rect 717 -382 763 -370
rect 813 -290 859 -278
rect 813 -370 819 -290
rect 853 -370 859 -290
rect 813 -382 859 -370
rect 909 -290 955 -278
rect 909 -370 915 -290
rect 949 -370 955 -290
rect 909 -382 955 -370
rect 1005 -290 1051 -278
rect 1005 -370 1011 -290
rect 1045 -370 1051 -290
rect 1005 -382 1051 -370
rect 1101 -290 1147 -278
rect 1101 -370 1107 -290
rect 1141 -370 1147 -290
rect 1101 -382 1147 -370
rect 1197 -290 1243 -278
rect 1197 -370 1203 -290
rect 1237 -370 1243 -290
rect 1197 -382 1243 -370
rect 1293 -290 1339 -278
rect 1293 -370 1299 -290
rect 1333 -370 1339 -290
rect 1293 -382 1339 -370
rect 1389 -290 1435 -278
rect 1389 -370 1395 -290
rect 1429 -370 1435 -290
rect 1389 -382 1435 -370
rect 1503 -285 1549 -273
rect 1609 -285 1655 -284
rect 215 -513 319 -503
rect -2162 -558 -2116 -546
rect -80 -547 319 -513
rect -3461 -742 -3232 -690
rect -3266 -1110 -3232 -742
rect -3116 -699 -3082 -558
rect -2924 -699 -2890 -558
rect -2732 -699 -2698 -558
rect -2540 -699 -2506 -558
rect -2348 -699 -2314 -558
rect -2156 -699 -2122 -558
rect -1426 -645 -1416 -593
rect -1364 -597 -1354 -593
rect -1364 -603 -776 -597
rect -1364 -637 -822 -603
rect -788 -637 -776 -603
rect -471 -636 -461 -584
rect -409 -636 -399 -584
rect -1364 -643 -776 -637
rect -1364 -645 -1354 -643
rect -3116 -733 -1797 -699
rect -3116 -864 -3082 -733
rect -2924 -864 -2890 -733
rect -2732 -864 -2698 -733
rect -2540 -864 -2506 -733
rect -2348 -864 -2314 -733
rect -2156 -864 -2122 -733
rect -3122 -876 -3076 -864
rect -3122 -956 -3116 -876
rect -3082 -956 -3076 -876
rect -3122 -968 -3076 -956
rect -3026 -876 -2980 -864
rect -3026 -956 -3020 -876
rect -2986 -956 -2980 -876
rect -3026 -968 -2980 -956
rect -2930 -876 -2884 -864
rect -2930 -956 -2924 -876
rect -2890 -956 -2884 -876
rect -2930 -968 -2884 -956
rect -2834 -876 -2788 -864
rect -2834 -956 -2828 -876
rect -2794 -956 -2788 -876
rect -2834 -968 -2788 -956
rect -2738 -876 -2692 -864
rect -2738 -956 -2732 -876
rect -2698 -956 -2692 -876
rect -2738 -968 -2692 -956
rect -2642 -876 -2596 -864
rect -2642 -956 -2636 -876
rect -2602 -956 -2596 -876
rect -2642 -968 -2596 -956
rect -2546 -876 -2500 -864
rect -2546 -956 -2540 -876
rect -2506 -956 -2500 -876
rect -2546 -968 -2500 -956
rect -2450 -876 -2404 -864
rect -2450 -956 -2444 -876
rect -2410 -956 -2404 -876
rect -2450 -968 -2404 -956
rect -2354 -876 -2308 -864
rect -2354 -956 -2348 -876
rect -2314 -956 -2308 -876
rect -2354 -968 -2308 -956
rect -2258 -876 -2212 -864
rect -2258 -956 -2252 -876
rect -2218 -956 -2212 -876
rect -2258 -968 -2212 -956
rect -2162 -876 -2116 -864
rect -2162 -956 -2156 -876
rect -2122 -956 -2116 -876
rect -1831 -870 -1797 -733
rect -924 -742 -914 -690
rect -862 -742 -852 -690
rect -559 -746 -549 -694
rect -497 -746 -487 -694
rect -80 -870 -46 -547
rect 215 -555 319 -547
rect -1831 -904 -46 -870
rect -2162 -968 -2116 -956
rect -3020 -1110 -2986 -968
rect -2828 -1110 -2794 -968
rect -2636 -1110 -2602 -968
rect -2444 -1110 -2410 -968
rect -2367 -1060 -2357 -1008
rect -2305 -1060 -2295 -1008
rect -2252 -1110 -2218 -968
rect -980 -1004 -336 -973
rect -2176 -1058 -2166 -1006
rect -2114 -1058 -2104 -1006
rect -980 -1038 -951 -1004
rect -917 -1038 -859 -1004
rect -825 -1038 -767 -1004
rect -733 -1038 -675 -1004
rect -641 -1038 -583 -1004
rect -549 -1038 -491 -1004
rect -457 -1038 -399 -1004
rect -365 -1038 -336 -1004
rect -980 -1069 -336 -1038
rect -3266 -1144 -2218 -1110
rect 285 -1110 319 -555
rect 435 -513 469 -382
rect 627 -513 661 -382
rect 819 -513 853 -382
rect 1011 -513 1045 -382
rect 1203 -513 1237 -382
rect 1395 -513 1429 -382
rect 1503 -385 1509 -285
rect 1543 -296 1655 -285
rect 1543 -372 1615 -296
rect 1649 -372 1655 -296
rect 1543 -384 1655 -372
rect 1697 -285 1743 -284
rect 1806 -285 1840 -136
rect 1938 -240 1948 -188
rect 2000 -240 2010 -188
rect 2052 -278 2086 -136
rect 2244 -278 2278 -136
rect 2436 -278 2470 -136
rect 2628 -278 2662 -136
rect 2820 -278 2854 -136
rect 2898 -240 2908 -188
rect 2960 -240 2970 -188
rect 1697 -296 1840 -285
rect 1697 -372 1703 -296
rect 1737 -372 1840 -296
rect 1697 -384 1840 -372
rect 1950 -290 1996 -278
rect 1950 -370 1956 -290
rect 1990 -370 1996 -290
rect 1950 -382 1996 -370
rect 2046 -290 2092 -278
rect 2046 -370 2052 -290
rect 2086 -370 2092 -290
rect 2046 -382 2092 -370
rect 2142 -290 2188 -278
rect 2142 -370 2148 -290
rect 2182 -370 2188 -290
rect 2142 -382 2188 -370
rect 2238 -290 2284 -278
rect 2238 -370 2244 -290
rect 2278 -370 2284 -290
rect 2238 -382 2284 -370
rect 2334 -290 2380 -278
rect 2334 -370 2340 -290
rect 2374 -370 2380 -290
rect 2334 -382 2380 -370
rect 2430 -290 2476 -278
rect 2430 -370 2436 -290
rect 2470 -370 2476 -290
rect 2430 -382 2476 -370
rect 2526 -290 2572 -278
rect 2526 -370 2532 -290
rect 2566 -370 2572 -290
rect 2526 -382 2572 -370
rect 2622 -290 2668 -278
rect 2622 -370 2628 -290
rect 2662 -370 2668 -290
rect 2622 -382 2668 -370
rect 2718 -290 2764 -278
rect 2718 -370 2724 -290
rect 2758 -370 2764 -290
rect 2718 -382 2764 -370
rect 2814 -290 2860 -278
rect 2814 -370 2820 -290
rect 2854 -370 2860 -290
rect 2814 -382 2860 -370
rect 2910 -290 2956 -278
rect 2910 -370 2916 -290
rect 2950 -370 2956 -290
rect 2910 -382 2956 -370
rect 1543 -385 1649 -384
rect 1703 -385 1840 -384
rect 1503 -397 1549 -385
rect 1647 -422 1705 -416
rect 1647 -423 1659 -422
rect 1693 -423 1705 -422
rect 1640 -475 1650 -423
rect 1702 -475 1712 -423
rect 1806 -513 1840 -385
rect 435 -547 1840 -513
rect 435 -688 469 -547
rect 627 -688 661 -547
rect 819 -688 853 -547
rect 1011 -688 1045 -547
rect 1203 -688 1237 -547
rect 1395 -688 1429 -547
rect 429 -700 475 -688
rect 429 -948 435 -700
rect 469 -948 475 -700
rect 429 -960 475 -948
rect 525 -700 571 -688
rect 525 -948 531 -700
rect 565 -948 571 -700
rect 525 -960 571 -948
rect 621 -700 667 -688
rect 621 -948 627 -700
rect 661 -948 667 -700
rect 621 -960 667 -948
rect 717 -700 763 -688
rect 717 -948 723 -700
rect 757 -948 763 -700
rect 717 -960 763 -948
rect 813 -700 859 -688
rect 813 -948 819 -700
rect 853 -948 859 -700
rect 813 -960 859 -948
rect 909 -700 955 -688
rect 909 -948 915 -700
rect 949 -948 955 -700
rect 909 -960 955 -948
rect 1005 -700 1051 -688
rect 1005 -948 1011 -700
rect 1045 -948 1051 -700
rect 1005 -960 1051 -948
rect 1101 -700 1147 -688
rect 1101 -948 1107 -700
rect 1141 -948 1147 -700
rect 1101 -960 1147 -948
rect 1197 -700 1243 -688
rect 1197 -948 1203 -700
rect 1237 -948 1243 -700
rect 1197 -960 1243 -948
rect 1293 -700 1339 -688
rect 1293 -948 1299 -700
rect 1333 -948 1339 -700
rect 1293 -960 1339 -948
rect 1389 -700 1435 -688
rect 1389 -948 1395 -700
rect 1429 -948 1435 -700
rect 1389 -960 1435 -948
rect 416 -1051 426 -999
rect 478 -1051 488 -999
rect 531 -1110 565 -960
rect 723 -1110 757 -960
rect 915 -1110 949 -960
rect 1107 -1110 1141 -960
rect 1299 -1110 1333 -960
rect 1375 -1052 1385 -1000
rect 1437 -1052 1447 -1000
rect 285 -1144 1333 -1110
rect 1806 -1110 1840 -547
rect 1956 -513 1990 -382
rect 2148 -513 2182 -382
rect 2340 -513 2374 -382
rect 2532 -513 2566 -382
rect 2724 -513 2758 -382
rect 2916 -513 2950 -382
rect 3048 -513 3317 -504
rect 1956 -547 3317 -513
rect 1956 -688 1990 -547
rect 2148 -688 2182 -547
rect 2340 -688 2374 -547
rect 2532 -688 2566 -547
rect 2724 -688 2758 -547
rect 2916 -688 2950 -547
rect 3048 -556 3317 -547
rect 1950 -700 1996 -688
rect 1950 -948 1956 -700
rect 1990 -948 1996 -700
rect 1950 -960 1996 -948
rect 2046 -700 2092 -688
rect 2046 -948 2052 -700
rect 2086 -948 2092 -700
rect 2046 -960 2092 -948
rect 2142 -700 2188 -688
rect 2142 -948 2148 -700
rect 2182 -948 2188 -700
rect 2142 -960 2188 -948
rect 2238 -700 2284 -688
rect 2238 -948 2244 -700
rect 2278 -948 2284 -700
rect 2238 -960 2284 -948
rect 2334 -700 2380 -688
rect 2334 -948 2340 -700
rect 2374 -948 2380 -700
rect 2334 -960 2380 -948
rect 2430 -700 2476 -688
rect 2430 -948 2436 -700
rect 2470 -948 2476 -700
rect 2430 -960 2476 -948
rect 2526 -700 2572 -688
rect 2526 -948 2532 -700
rect 2566 -948 2572 -700
rect 2526 -960 2572 -948
rect 2622 -700 2668 -688
rect 2622 -948 2628 -700
rect 2662 -948 2668 -700
rect 2622 -960 2668 -948
rect 2718 -700 2764 -688
rect 2718 -948 2724 -700
rect 2758 -948 2764 -700
rect 2718 -960 2764 -948
rect 2814 -700 2860 -688
rect 2814 -948 2820 -700
rect 2854 -948 2860 -700
rect 2814 -960 2860 -948
rect 2910 -700 2956 -688
rect 2910 -948 2916 -700
rect 2950 -948 2956 -700
rect 2910 -960 2956 -948
rect 1936 -1052 1946 -1000
rect 1998 -1052 2008 -1000
rect 2052 -1110 2086 -960
rect 2244 -1110 2278 -960
rect 2436 -1110 2470 -960
rect 2628 -1110 2662 -960
rect 2820 -1110 2854 -960
rect 2896 -1052 2906 -1000
rect 2958 -1052 2968 -1000
rect 1806 -1144 2854 -1110
rect 88 -1191 98 -1188
rect -465 -1197 98 -1191
rect -465 -1231 -453 -1197
rect -419 -1231 98 -1197
rect -465 -1237 98 -1231
rect 88 -1240 98 -1237
rect 150 -1240 160 -1188
rect -549 -1312 -287 -1303
rect -549 -1346 -534 -1312
rect -500 -1346 -287 -1312
rect -549 -1355 -287 -1346
rect -235 -1355 -225 -1303
rect -3266 -1470 -2218 -1436
rect -3266 -2023 -3232 -1470
rect -3020 -1620 -2986 -1470
rect -2828 -1620 -2794 -1470
rect -2636 -1620 -2602 -1470
rect -2444 -1620 -2410 -1470
rect -2367 -1580 -2357 -1528
rect -2305 -1580 -2295 -1528
rect -2252 -1620 -2218 -1470
rect -1852 -1446 -50 -1412
rect -2175 -1581 -2165 -1529
rect -2113 -1581 -2103 -1529
rect -3122 -1632 -3076 -1620
rect -3122 -1880 -3116 -1632
rect -3082 -1880 -3076 -1632
rect -3122 -1892 -3076 -1880
rect -3026 -1632 -2980 -1620
rect -3026 -1880 -3020 -1632
rect -2986 -1880 -2980 -1632
rect -3026 -1892 -2980 -1880
rect -2930 -1632 -2884 -1620
rect -2930 -1880 -2924 -1632
rect -2890 -1880 -2884 -1632
rect -2930 -1892 -2884 -1880
rect -2834 -1632 -2788 -1620
rect -2834 -1880 -2828 -1632
rect -2794 -1880 -2788 -1632
rect -2834 -1892 -2788 -1880
rect -2738 -1632 -2692 -1620
rect -2738 -1880 -2732 -1632
rect -2698 -1880 -2692 -1632
rect -2738 -1892 -2692 -1880
rect -2642 -1632 -2596 -1620
rect -2642 -1880 -2636 -1632
rect -2602 -1880 -2596 -1632
rect -2642 -1892 -2596 -1880
rect -2546 -1632 -2500 -1620
rect -2546 -1880 -2540 -1632
rect -2506 -1880 -2500 -1632
rect -2546 -1892 -2500 -1880
rect -2450 -1632 -2404 -1620
rect -2450 -1880 -2444 -1632
rect -2410 -1880 -2404 -1632
rect -2450 -1892 -2404 -1880
rect -2354 -1632 -2308 -1620
rect -2354 -1880 -2348 -1632
rect -2314 -1880 -2308 -1632
rect -2354 -1892 -2308 -1880
rect -2258 -1632 -2212 -1620
rect -2258 -1880 -2252 -1632
rect -2218 -1880 -2212 -1632
rect -2258 -1892 -2212 -1880
rect -2162 -1632 -2116 -1620
rect -2162 -1880 -2156 -1632
rect -2122 -1880 -2116 -1632
rect -2162 -1892 -2116 -1880
rect -3461 -2075 -3232 -2023
rect -3266 -2444 -3232 -2075
rect -3116 -2033 -3082 -1892
rect -2924 -2033 -2890 -1892
rect -2732 -2033 -2698 -1892
rect -2540 -2033 -2506 -1892
rect -2348 -2033 -2314 -1892
rect -2156 -2033 -2122 -1892
rect -1852 -2033 -1818 -1446
rect -1734 -1580 -1724 -1528
rect -1672 -1580 -1416 -1528
rect -1364 -1580 -1354 -1528
rect -704 -1548 -336 -1517
rect -704 -1582 -675 -1548
rect -641 -1582 -583 -1548
rect -549 -1582 -491 -1548
rect -457 -1582 -399 -1548
rect -365 -1582 -336 -1548
rect -704 -1613 -336 -1582
rect -488 -1721 -478 -1669
rect -426 -1721 -416 -1669
rect -602 -1828 -592 -1776
rect -540 -1828 -530 -1776
rect -426 -1831 -416 -1779
rect -364 -1831 -354 -1779
rect -84 -1847 -50 -1446
rect 285 -1470 1333 -1436
rect 285 -1837 319 -1470
rect 415 -1572 425 -1520
rect 477 -1572 487 -1520
rect 531 -1612 565 -1470
rect 723 -1612 757 -1470
rect 915 -1612 949 -1470
rect 1107 -1612 1141 -1470
rect 1299 -1612 1333 -1470
rect 1806 -1470 2854 -1436
rect 1377 -1574 1387 -1522
rect 1439 -1574 1449 -1522
rect 429 -1624 475 -1612
rect 429 -1704 435 -1624
rect 469 -1704 475 -1624
rect 429 -1716 475 -1704
rect 525 -1624 571 -1612
rect 525 -1704 531 -1624
rect 565 -1704 571 -1624
rect 525 -1716 571 -1704
rect 621 -1624 667 -1612
rect 621 -1704 627 -1624
rect 661 -1704 667 -1624
rect 621 -1716 667 -1704
rect 717 -1624 763 -1612
rect 717 -1704 723 -1624
rect 757 -1704 763 -1624
rect 717 -1716 763 -1704
rect 813 -1624 859 -1612
rect 813 -1704 819 -1624
rect 853 -1704 859 -1624
rect 813 -1716 859 -1704
rect 909 -1624 955 -1612
rect 909 -1704 915 -1624
rect 949 -1704 955 -1624
rect 909 -1716 955 -1704
rect 1005 -1624 1051 -1612
rect 1005 -1704 1011 -1624
rect 1045 -1704 1051 -1624
rect 1005 -1716 1051 -1704
rect 1101 -1624 1147 -1612
rect 1101 -1704 1107 -1624
rect 1141 -1704 1147 -1624
rect 1101 -1716 1147 -1704
rect 1197 -1624 1243 -1612
rect 1197 -1704 1203 -1624
rect 1237 -1704 1243 -1624
rect 1197 -1716 1243 -1704
rect 1293 -1624 1339 -1612
rect 1293 -1704 1299 -1624
rect 1333 -1704 1339 -1624
rect 1293 -1716 1339 -1704
rect 1389 -1624 1435 -1612
rect 1389 -1704 1395 -1624
rect 1429 -1704 1435 -1624
rect 1389 -1716 1435 -1704
rect 1503 -1619 1549 -1607
rect 1609 -1619 1655 -1618
rect 215 -1847 319 -1837
rect -84 -1881 319 -1847
rect 215 -1889 319 -1881
rect -882 -1971 -872 -1919
rect -820 -1971 -416 -1919
rect -364 -1971 -354 -1919
rect -3116 -2067 -1818 -2033
rect -3116 -2198 -3082 -2067
rect -2924 -2198 -2890 -2067
rect -2732 -2198 -2698 -2067
rect -2540 -2198 -2506 -2067
rect -2348 -2198 -2314 -2067
rect -2156 -2198 -2122 -2067
rect -1256 -2092 -336 -2061
rect -1256 -2126 -1227 -2092
rect -1193 -2126 -1135 -2092
rect -1101 -2126 -1043 -2092
rect -1009 -2126 -951 -2092
rect -917 -2126 -859 -2092
rect -825 -2126 -767 -2092
rect -733 -2126 -675 -2092
rect -641 -2126 -583 -2092
rect -549 -2126 -491 -2092
rect -457 -2126 -399 -2092
rect -365 -2126 -336 -2092
rect -1256 -2157 -336 -2126
rect -3122 -2210 -3076 -2198
rect -3122 -2290 -3116 -2210
rect -3082 -2290 -3076 -2210
rect -3122 -2302 -3076 -2290
rect -3026 -2210 -2980 -2198
rect -3026 -2290 -3020 -2210
rect -2986 -2290 -2980 -2210
rect -3026 -2302 -2980 -2290
rect -2930 -2210 -2884 -2198
rect -2930 -2290 -2924 -2210
rect -2890 -2290 -2884 -2210
rect -2930 -2302 -2884 -2290
rect -2834 -2210 -2788 -2198
rect -2834 -2290 -2828 -2210
rect -2794 -2290 -2788 -2210
rect -2834 -2302 -2788 -2290
rect -2738 -2210 -2692 -2198
rect -2738 -2290 -2732 -2210
rect -2698 -2290 -2692 -2210
rect -2738 -2302 -2692 -2290
rect -2642 -2210 -2596 -2198
rect -2642 -2290 -2636 -2210
rect -2602 -2290 -2596 -2210
rect -2642 -2302 -2596 -2290
rect -2546 -2210 -2500 -2198
rect -2546 -2290 -2540 -2210
rect -2506 -2290 -2500 -2210
rect -2546 -2302 -2500 -2290
rect -2450 -2210 -2404 -2198
rect -2450 -2290 -2444 -2210
rect -2410 -2290 -2404 -2210
rect -2450 -2302 -2404 -2290
rect -2354 -2210 -2308 -2198
rect -2354 -2290 -2348 -2210
rect -2314 -2290 -2308 -2210
rect -2354 -2302 -2308 -2290
rect -2258 -2210 -2212 -2198
rect -2258 -2290 -2252 -2210
rect -2218 -2290 -2212 -2210
rect -2258 -2302 -2212 -2290
rect -2162 -2210 -2116 -2198
rect -2162 -2290 -2156 -2210
rect -2122 -2290 -2116 -2210
rect -602 -2230 -592 -2225
rect -1016 -2236 -592 -2230
rect -1016 -2270 -1004 -2236
rect -970 -2270 -592 -2236
rect -1016 -2276 -592 -2270
rect -602 -2277 -592 -2276
rect -540 -2277 -530 -2225
rect -297 -2264 -287 -2261
rect -501 -2270 -287 -2264
rect -2162 -2302 -2116 -2290
rect -3020 -2444 -2986 -2302
rect -2828 -2444 -2794 -2302
rect -2636 -2444 -2602 -2302
rect -2444 -2444 -2410 -2302
rect -2366 -2393 -2356 -2341
rect -2304 -2393 -2294 -2341
rect -2252 -2444 -2218 -2302
rect -501 -2304 -489 -2270
rect -455 -2304 -287 -2270
rect -501 -2310 -287 -2304
rect -297 -2313 -287 -2310
rect -235 -2313 -225 -2261
rect -2174 -2392 -2164 -2340
rect -2112 -2392 -2102 -2340
rect -1111 -2440 -1101 -2388
rect -1049 -2440 -762 -2388
rect -710 -2440 -700 -2388
rect -602 -2442 -592 -2390
rect -540 -2442 -530 -2390
rect -422 -2437 -412 -2385
rect -360 -2437 -350 -2385
rect -3266 -2478 -2218 -2444
rect 285 -2444 319 -1889
rect 435 -1847 469 -1716
rect 627 -1847 661 -1716
rect 819 -1847 853 -1716
rect 1011 -1847 1045 -1716
rect 1203 -1847 1237 -1716
rect 1395 -1847 1429 -1716
rect 1503 -1719 1509 -1619
rect 1543 -1630 1655 -1619
rect 1543 -1706 1615 -1630
rect 1649 -1706 1655 -1630
rect 1543 -1718 1655 -1706
rect 1697 -1619 1743 -1618
rect 1806 -1619 1840 -1470
rect 1938 -1574 1948 -1522
rect 2000 -1574 2010 -1522
rect 2052 -1612 2086 -1470
rect 2244 -1612 2278 -1470
rect 2436 -1612 2470 -1470
rect 2628 -1612 2662 -1470
rect 2820 -1612 2854 -1470
rect 2898 -1574 2908 -1522
rect 2960 -1574 2970 -1522
rect 1697 -1630 1840 -1619
rect 1697 -1706 1703 -1630
rect 1737 -1706 1840 -1630
rect 1697 -1718 1840 -1706
rect 1950 -1624 1996 -1612
rect 1950 -1704 1956 -1624
rect 1990 -1704 1996 -1624
rect 1950 -1716 1996 -1704
rect 2046 -1624 2092 -1612
rect 2046 -1704 2052 -1624
rect 2086 -1704 2092 -1624
rect 2046 -1716 2092 -1704
rect 2142 -1624 2188 -1612
rect 2142 -1704 2148 -1624
rect 2182 -1704 2188 -1624
rect 2142 -1716 2188 -1704
rect 2238 -1624 2284 -1612
rect 2238 -1704 2244 -1624
rect 2278 -1704 2284 -1624
rect 2238 -1716 2284 -1704
rect 2334 -1624 2380 -1612
rect 2334 -1704 2340 -1624
rect 2374 -1704 2380 -1624
rect 2334 -1716 2380 -1704
rect 2430 -1624 2476 -1612
rect 2430 -1704 2436 -1624
rect 2470 -1704 2476 -1624
rect 2430 -1716 2476 -1704
rect 2526 -1624 2572 -1612
rect 2526 -1704 2532 -1624
rect 2566 -1704 2572 -1624
rect 2526 -1716 2572 -1704
rect 2622 -1624 2668 -1612
rect 2622 -1704 2628 -1624
rect 2662 -1704 2668 -1624
rect 2622 -1716 2668 -1704
rect 2718 -1624 2764 -1612
rect 2718 -1704 2724 -1624
rect 2758 -1704 2764 -1624
rect 2718 -1716 2764 -1704
rect 2814 -1624 2860 -1612
rect 2814 -1704 2820 -1624
rect 2854 -1704 2860 -1624
rect 2814 -1716 2860 -1704
rect 2910 -1624 2956 -1612
rect 2910 -1704 2916 -1624
rect 2950 -1704 2956 -1624
rect 2910 -1716 2956 -1704
rect 1543 -1719 1649 -1718
rect 1703 -1719 1840 -1718
rect 1503 -1731 1549 -1719
rect 1647 -1756 1705 -1750
rect 1647 -1757 1659 -1756
rect 1693 -1757 1705 -1756
rect 1640 -1809 1650 -1757
rect 1702 -1809 1712 -1757
rect 1806 -1847 1840 -1719
rect 435 -1881 1840 -1847
rect 435 -2022 469 -1881
rect 627 -2022 661 -1881
rect 819 -2022 853 -1881
rect 1011 -2022 1045 -1881
rect 1203 -2022 1237 -1881
rect 1395 -2022 1429 -1881
rect 429 -2034 475 -2022
rect 429 -2282 435 -2034
rect 469 -2282 475 -2034
rect 429 -2294 475 -2282
rect 525 -2034 571 -2022
rect 525 -2282 531 -2034
rect 565 -2282 571 -2034
rect 525 -2294 571 -2282
rect 621 -2034 667 -2022
rect 621 -2282 627 -2034
rect 661 -2282 667 -2034
rect 621 -2294 667 -2282
rect 717 -2034 763 -2022
rect 717 -2282 723 -2034
rect 757 -2282 763 -2034
rect 717 -2294 763 -2282
rect 813 -2034 859 -2022
rect 813 -2282 819 -2034
rect 853 -2282 859 -2034
rect 813 -2294 859 -2282
rect 909 -2034 955 -2022
rect 909 -2282 915 -2034
rect 949 -2282 955 -2034
rect 909 -2294 955 -2282
rect 1005 -2034 1051 -2022
rect 1005 -2282 1011 -2034
rect 1045 -2282 1051 -2034
rect 1005 -2294 1051 -2282
rect 1101 -2034 1147 -2022
rect 1101 -2282 1107 -2034
rect 1141 -2282 1147 -2034
rect 1101 -2294 1147 -2282
rect 1197 -2034 1243 -2022
rect 1197 -2282 1203 -2034
rect 1237 -2282 1243 -2034
rect 1197 -2294 1243 -2282
rect 1293 -2034 1339 -2022
rect 1293 -2282 1299 -2034
rect 1333 -2282 1339 -2034
rect 1293 -2294 1339 -2282
rect 1389 -2034 1435 -2022
rect 1389 -2282 1395 -2034
rect 1429 -2282 1435 -2034
rect 1389 -2294 1435 -2282
rect 416 -2385 426 -2333
rect 478 -2385 488 -2333
rect 531 -2444 565 -2294
rect 723 -2444 757 -2294
rect 915 -2444 949 -2294
rect 1107 -2444 1141 -2294
rect 1299 -2444 1333 -2294
rect 1375 -2386 1385 -2334
rect 1437 -2386 1447 -2334
rect 285 -2478 1333 -2444
rect 1806 -2444 1840 -1881
rect 1956 -1847 1990 -1716
rect 2148 -1847 2182 -1716
rect 2340 -1847 2374 -1716
rect 2532 -1847 2566 -1716
rect 2724 -1847 2758 -1716
rect 2916 -1847 2950 -1716
rect 3265 -1839 3317 -556
rect 3047 -1847 3317 -1839
rect 1956 -1881 3317 -1847
rect 1956 -2022 1990 -1881
rect 2148 -2022 2182 -1881
rect 2340 -2022 2374 -1881
rect 2532 -2022 2566 -1881
rect 2724 -2022 2758 -1881
rect 2916 -2022 2950 -1881
rect 3047 -1891 3317 -1881
rect 1950 -2034 1996 -2022
rect 1950 -2282 1956 -2034
rect 1990 -2282 1996 -2034
rect 1950 -2294 1996 -2282
rect 2046 -2034 2092 -2022
rect 2046 -2282 2052 -2034
rect 2086 -2282 2092 -2034
rect 2046 -2294 2092 -2282
rect 2142 -2034 2188 -2022
rect 2142 -2282 2148 -2034
rect 2182 -2282 2188 -2034
rect 2142 -2294 2188 -2282
rect 2238 -2034 2284 -2022
rect 2238 -2282 2244 -2034
rect 2278 -2282 2284 -2034
rect 2238 -2294 2284 -2282
rect 2334 -2034 2380 -2022
rect 2334 -2282 2340 -2034
rect 2374 -2282 2380 -2034
rect 2334 -2294 2380 -2282
rect 2430 -2034 2476 -2022
rect 2430 -2282 2436 -2034
rect 2470 -2282 2476 -2034
rect 2430 -2294 2476 -2282
rect 2526 -2034 2572 -2022
rect 2526 -2282 2532 -2034
rect 2566 -2282 2572 -2034
rect 2526 -2294 2572 -2282
rect 2622 -2034 2668 -2022
rect 2622 -2282 2628 -2034
rect 2662 -2282 2668 -2034
rect 2622 -2294 2668 -2282
rect 2718 -2034 2764 -2022
rect 2718 -2282 2724 -2034
rect 2758 -2282 2764 -2034
rect 2718 -2294 2764 -2282
rect 2814 -2034 2860 -2022
rect 2814 -2282 2820 -2034
rect 2854 -2282 2860 -2034
rect 2814 -2294 2860 -2282
rect 2910 -2034 2956 -2022
rect 2910 -2282 2916 -2034
rect 2950 -2282 2956 -2034
rect 2910 -2294 2956 -2282
rect 1936 -2386 1946 -2334
rect 1998 -2386 2008 -2334
rect 2052 -2444 2086 -2294
rect 2244 -2444 2278 -2294
rect 2436 -2444 2470 -2294
rect 2628 -2444 2662 -2294
rect 2820 -2444 2854 -2294
rect 2896 -2386 2906 -2334
rect 2958 -2386 2968 -2334
rect 1806 -2478 2854 -2444
rect -1250 -2543 -1240 -2491
rect -1188 -2543 -412 -2491
rect -360 -2543 -350 -2491
rect -1256 -2636 -336 -2605
rect -1256 -2670 -1227 -2636
rect -1193 -2670 -1135 -2636
rect -1101 -2670 -1043 -2636
rect -1009 -2670 -951 -2636
rect -917 -2670 -859 -2636
rect -825 -2670 -767 -2636
rect -733 -2670 -675 -2636
rect -641 -2670 -583 -2636
rect -549 -2670 -491 -2636
rect -457 -2670 -399 -2636
rect -365 -2670 -336 -2636
rect -1256 -2701 -336 -2670
rect 3265 -2617 3317 -1891
rect 3265 -2626 3454 -2617
rect 3265 -2660 3456 -2626
rect 3265 -2669 3454 -2660
rect -3266 -2848 -2218 -2814
rect -772 -2827 -762 -2775
rect -710 -2827 -412 -2775
rect -360 -2827 -350 -2775
rect -3266 -3403 -3232 -2848
rect -3020 -2998 -2986 -2848
rect -2828 -2998 -2794 -2848
rect -2636 -2998 -2602 -2848
rect -2444 -2998 -2410 -2848
rect -2367 -2958 -2357 -2906
rect -2305 -2958 -2295 -2906
rect -2252 -2998 -2218 -2848
rect 285 -2848 1333 -2814
rect -2175 -2959 -2165 -2907
rect -2113 -2959 -2103 -2907
rect -1936 -2958 -1926 -2906
rect -1874 -2958 -1416 -2906
rect -1364 -2958 -1354 -2906
rect -1108 -2917 -1098 -2865
rect -1046 -2917 -1036 -2865
rect -1002 -2868 -872 -2864
rect -1006 -2874 -872 -2868
rect -1006 -2908 -994 -2874
rect -960 -2908 -872 -2874
rect -1006 -2914 -872 -2908
rect -1002 -2916 -872 -2914
rect -820 -2874 -527 -2864
rect -820 -2908 -574 -2874
rect -540 -2908 -527 -2874
rect -820 -2916 -527 -2908
rect -1002 -2918 -527 -2916
rect -422 -2918 -412 -2866
rect -360 -2918 -350 -2866
rect -3122 -3010 -3076 -2998
rect -3122 -3258 -3116 -3010
rect -3082 -3258 -3076 -3010
rect -3122 -3270 -3076 -3258
rect -3026 -3010 -2980 -2998
rect -3026 -3258 -3020 -3010
rect -2986 -3258 -2980 -3010
rect -3026 -3270 -2980 -3258
rect -2930 -3010 -2884 -2998
rect -2930 -3258 -2924 -3010
rect -2890 -3258 -2884 -3010
rect -2930 -3270 -2884 -3258
rect -2834 -3010 -2788 -2998
rect -2834 -3258 -2828 -3010
rect -2794 -3258 -2788 -3010
rect -2834 -3270 -2788 -3258
rect -2738 -3010 -2692 -2998
rect -2738 -3258 -2732 -3010
rect -2698 -3258 -2692 -3010
rect -2738 -3270 -2692 -3258
rect -2642 -3010 -2596 -2998
rect -2642 -3258 -2636 -3010
rect -2602 -3258 -2596 -3010
rect -2642 -3270 -2596 -3258
rect -2546 -3010 -2500 -2998
rect -2546 -3258 -2540 -3010
rect -2506 -3258 -2500 -3010
rect -2546 -3270 -2500 -3258
rect -2450 -3010 -2404 -2998
rect -2450 -3258 -2444 -3010
rect -2410 -3258 -2404 -3010
rect -2450 -3270 -2404 -3258
rect -2354 -3010 -2308 -2998
rect -2354 -3258 -2348 -3010
rect -2314 -3258 -2308 -3010
rect -2354 -3270 -2308 -3258
rect -2258 -3010 -2212 -2998
rect -2258 -3258 -2252 -3010
rect -2218 -3258 -2212 -3010
rect -2258 -3270 -2212 -3258
rect -2162 -3010 -2116 -2998
rect -2162 -3258 -2156 -3010
rect -2122 -3258 -2116 -3010
rect -246 -3030 -236 -3026
rect -502 -3036 -236 -3030
rect -502 -3070 -490 -3036
rect -456 -3070 -236 -3036
rect -502 -3076 -236 -3070
rect -246 -3078 -236 -3076
rect -184 -3078 -174 -3026
rect -1256 -3180 -336 -3149
rect -1256 -3214 -1227 -3180
rect -1193 -3214 -1135 -3180
rect -1101 -3214 -1043 -3180
rect -1009 -3214 -951 -3180
rect -917 -3214 -859 -3180
rect -825 -3214 -767 -3180
rect -733 -3214 -675 -3180
rect -641 -3214 -583 -3180
rect -549 -3214 -491 -3180
rect -457 -3214 -399 -3180
rect -365 -3214 -336 -3180
rect -1256 -3245 -336 -3214
rect 285 -3215 319 -2848
rect 415 -2950 425 -2898
rect 477 -2950 487 -2898
rect 531 -2990 565 -2848
rect 723 -2990 757 -2848
rect 915 -2990 949 -2848
rect 1107 -2990 1141 -2848
rect 1299 -2990 1333 -2848
rect 1806 -2848 2854 -2814
rect 1377 -2952 1387 -2900
rect 1439 -2952 1449 -2900
rect 429 -3002 475 -2990
rect 429 -3082 435 -3002
rect 469 -3082 475 -3002
rect 429 -3094 475 -3082
rect 525 -3002 571 -2990
rect 525 -3082 531 -3002
rect 565 -3082 571 -3002
rect 525 -3094 571 -3082
rect 621 -3002 667 -2990
rect 621 -3082 627 -3002
rect 661 -3082 667 -3002
rect 621 -3094 667 -3082
rect 717 -3002 763 -2990
rect 717 -3082 723 -3002
rect 757 -3082 763 -3002
rect 717 -3094 763 -3082
rect 813 -3002 859 -2990
rect 813 -3082 819 -3002
rect 853 -3082 859 -3002
rect 813 -3094 859 -3082
rect 909 -3002 955 -2990
rect 909 -3082 915 -3002
rect 949 -3082 955 -3002
rect 909 -3094 955 -3082
rect 1005 -3002 1051 -2990
rect 1005 -3082 1011 -3002
rect 1045 -3082 1051 -3002
rect 1005 -3094 1051 -3082
rect 1101 -3002 1147 -2990
rect 1101 -3082 1107 -3002
rect 1141 -3082 1147 -3002
rect 1101 -3094 1147 -3082
rect 1197 -3002 1243 -2990
rect 1197 -3082 1203 -3002
rect 1237 -3082 1243 -3002
rect 1197 -3094 1243 -3082
rect 1293 -3002 1339 -2990
rect 1293 -3082 1299 -3002
rect 1333 -3082 1339 -3002
rect 1293 -3094 1339 -3082
rect 1389 -3002 1435 -2990
rect 1389 -3082 1395 -3002
rect 1429 -3082 1435 -3002
rect 1389 -3094 1435 -3082
rect 1503 -2997 1549 -2985
rect 1609 -2997 1655 -2996
rect 215 -3225 319 -3215
rect -2162 -3270 -2116 -3258
rect -44 -3259 319 -3225
rect -3461 -3455 -3232 -3403
rect -3266 -3822 -3232 -3455
rect -3116 -3411 -3082 -3270
rect -2924 -3411 -2890 -3270
rect -2732 -3411 -2698 -3270
rect -2540 -3411 -2506 -3270
rect -2348 -3411 -2314 -3270
rect -2156 -3411 -2122 -3270
rect -44 -3308 -10 -3259
rect 215 -3267 319 -3259
rect -1812 -3342 -10 -3308
rect -1812 -3411 -1778 -3342
rect -3116 -3445 -1778 -3411
rect -773 -3445 -762 -3393
rect -710 -3445 -414 -3393
rect -362 -3445 -352 -3393
rect -3116 -3576 -3082 -3445
rect -2924 -3576 -2890 -3445
rect -2732 -3576 -2698 -3445
rect -2540 -3576 -2506 -3445
rect -2348 -3576 -2314 -3445
rect -2156 -3576 -2122 -3445
rect -1251 -3539 -1241 -3485
rect -1187 -3492 -528 -3485
rect -1187 -3526 -576 -3492
rect -542 -3526 -528 -3492
rect -424 -3526 -414 -3474
rect -362 -3526 -352 -3474
rect -1187 -3539 -528 -3526
rect -417 -3527 -359 -3526
rect -3122 -3588 -3076 -3576
rect -3122 -3668 -3116 -3588
rect -3082 -3668 -3076 -3588
rect -3122 -3680 -3076 -3668
rect -3026 -3588 -2980 -3576
rect -3026 -3668 -3020 -3588
rect -2986 -3668 -2980 -3588
rect -3026 -3680 -2980 -3668
rect -2930 -3588 -2884 -3576
rect -2930 -3668 -2924 -3588
rect -2890 -3668 -2884 -3588
rect -2930 -3680 -2884 -3668
rect -2834 -3588 -2788 -3576
rect -2834 -3668 -2828 -3588
rect -2794 -3668 -2788 -3588
rect -2834 -3680 -2788 -3668
rect -2738 -3588 -2692 -3576
rect -2738 -3668 -2732 -3588
rect -2698 -3668 -2692 -3588
rect -2738 -3680 -2692 -3668
rect -2642 -3588 -2596 -3576
rect -2642 -3668 -2636 -3588
rect -2602 -3668 -2596 -3588
rect -2642 -3680 -2596 -3668
rect -2546 -3588 -2500 -3576
rect -2546 -3668 -2540 -3588
rect -2506 -3668 -2500 -3588
rect -2546 -3680 -2500 -3668
rect -2450 -3588 -2404 -3576
rect -2450 -3668 -2444 -3588
rect -2410 -3668 -2404 -3588
rect -2450 -3680 -2404 -3668
rect -2354 -3588 -2308 -3576
rect -2354 -3668 -2348 -3588
rect -2314 -3668 -2308 -3588
rect -2354 -3680 -2308 -3668
rect -2258 -3588 -2212 -3576
rect -2258 -3668 -2252 -3588
rect -2218 -3668 -2212 -3588
rect -2258 -3680 -2212 -3668
rect -2162 -3588 -2116 -3576
rect -2162 -3668 -2156 -3588
rect -2122 -3668 -2116 -3588
rect -510 -3632 -500 -3580
rect -448 -3632 -438 -3580
rect -2162 -3680 -2116 -3668
rect -3020 -3822 -2986 -3680
rect -2828 -3822 -2794 -3680
rect -2636 -3822 -2602 -3680
rect -2444 -3822 -2410 -3680
rect -2366 -3767 -2356 -3715
rect -2304 -3767 -2294 -3715
rect -2252 -3822 -2218 -3680
rect -2174 -3769 -2164 -3717
rect -2112 -3769 -2102 -3717
rect -704 -3724 -336 -3693
rect -704 -3758 -675 -3724
rect -641 -3758 -583 -3724
rect -549 -3758 -491 -3724
rect -457 -3758 -399 -3724
rect -365 -3758 -336 -3724
rect -704 -3789 -336 -3758
rect -245 -3764 -235 -3712
rect -183 -3764 140 -3712
rect 192 -3764 202 -3712
rect -3266 -3856 -2218 -3822
rect 285 -3822 319 -3267
rect 435 -3225 469 -3094
rect 627 -3225 661 -3094
rect 819 -3225 853 -3094
rect 1011 -3225 1045 -3094
rect 1203 -3225 1237 -3094
rect 1395 -3225 1429 -3094
rect 1503 -3097 1509 -2997
rect 1543 -3008 1655 -2997
rect 1543 -3084 1615 -3008
rect 1649 -3084 1655 -3008
rect 1543 -3096 1655 -3084
rect 1697 -2997 1743 -2996
rect 1806 -2997 1840 -2848
rect 1938 -2952 1948 -2900
rect 2000 -2952 2010 -2900
rect 2052 -2990 2086 -2848
rect 2244 -2990 2278 -2848
rect 2436 -2990 2470 -2848
rect 2628 -2990 2662 -2848
rect 2820 -2990 2854 -2848
rect 2898 -2952 2908 -2900
rect 2960 -2952 2970 -2900
rect 1697 -3008 1840 -2997
rect 1697 -3084 1703 -3008
rect 1737 -3084 1840 -3008
rect 1697 -3096 1840 -3084
rect 1950 -3002 1996 -2990
rect 1950 -3082 1956 -3002
rect 1990 -3082 1996 -3002
rect 1950 -3094 1996 -3082
rect 2046 -3002 2092 -2990
rect 2046 -3082 2052 -3002
rect 2086 -3082 2092 -3002
rect 2046 -3094 2092 -3082
rect 2142 -3002 2188 -2990
rect 2142 -3082 2148 -3002
rect 2182 -3082 2188 -3002
rect 2142 -3094 2188 -3082
rect 2238 -3002 2284 -2990
rect 2238 -3082 2244 -3002
rect 2278 -3082 2284 -3002
rect 2238 -3094 2284 -3082
rect 2334 -3002 2380 -2990
rect 2334 -3082 2340 -3002
rect 2374 -3082 2380 -3002
rect 2334 -3094 2380 -3082
rect 2430 -3002 2476 -2990
rect 2430 -3082 2436 -3002
rect 2470 -3082 2476 -3002
rect 2430 -3094 2476 -3082
rect 2526 -3002 2572 -2990
rect 2526 -3082 2532 -3002
rect 2566 -3082 2572 -3002
rect 2526 -3094 2572 -3082
rect 2622 -3002 2668 -2990
rect 2622 -3082 2628 -3002
rect 2662 -3082 2668 -3002
rect 2622 -3094 2668 -3082
rect 2718 -3002 2764 -2990
rect 2718 -3082 2724 -3002
rect 2758 -3082 2764 -3002
rect 2718 -3094 2764 -3082
rect 2814 -3002 2860 -2990
rect 2814 -3082 2820 -3002
rect 2854 -3082 2860 -3002
rect 2814 -3094 2860 -3082
rect 2910 -3002 2956 -2990
rect 2910 -3082 2916 -3002
rect 2950 -3082 2956 -3002
rect 2910 -3094 2956 -3082
rect 1543 -3097 1649 -3096
rect 1703 -3097 1840 -3096
rect 1503 -3109 1549 -3097
rect 1647 -3134 1705 -3128
rect 1647 -3135 1659 -3134
rect 1693 -3135 1705 -3134
rect 1640 -3187 1650 -3135
rect 1702 -3187 1712 -3135
rect 1806 -3225 1840 -3097
rect 435 -3259 1840 -3225
rect 435 -3400 469 -3259
rect 627 -3400 661 -3259
rect 819 -3400 853 -3259
rect 1011 -3400 1045 -3259
rect 1203 -3400 1237 -3259
rect 1395 -3400 1429 -3259
rect 429 -3412 475 -3400
rect 429 -3660 435 -3412
rect 469 -3660 475 -3412
rect 429 -3672 475 -3660
rect 525 -3412 571 -3400
rect 525 -3660 531 -3412
rect 565 -3660 571 -3412
rect 525 -3672 571 -3660
rect 621 -3412 667 -3400
rect 621 -3660 627 -3412
rect 661 -3660 667 -3412
rect 621 -3672 667 -3660
rect 717 -3412 763 -3400
rect 717 -3660 723 -3412
rect 757 -3660 763 -3412
rect 717 -3672 763 -3660
rect 813 -3412 859 -3400
rect 813 -3660 819 -3412
rect 853 -3660 859 -3412
rect 813 -3672 859 -3660
rect 909 -3412 955 -3400
rect 909 -3660 915 -3412
rect 949 -3660 955 -3412
rect 909 -3672 955 -3660
rect 1005 -3412 1051 -3400
rect 1005 -3660 1011 -3412
rect 1045 -3660 1051 -3412
rect 1005 -3672 1051 -3660
rect 1101 -3412 1147 -3400
rect 1101 -3660 1107 -3412
rect 1141 -3660 1147 -3412
rect 1101 -3672 1147 -3660
rect 1197 -3412 1243 -3400
rect 1197 -3660 1203 -3412
rect 1237 -3660 1243 -3412
rect 1197 -3672 1243 -3660
rect 1293 -3412 1339 -3400
rect 1293 -3660 1299 -3412
rect 1333 -3660 1339 -3412
rect 1293 -3672 1339 -3660
rect 1389 -3412 1435 -3400
rect 1389 -3660 1395 -3412
rect 1429 -3660 1435 -3412
rect 1389 -3672 1435 -3660
rect 416 -3763 426 -3711
rect 478 -3763 488 -3711
rect 531 -3822 565 -3672
rect 723 -3822 757 -3672
rect 915 -3822 949 -3672
rect 1107 -3822 1141 -3672
rect 1299 -3822 1333 -3672
rect 1375 -3764 1385 -3712
rect 1437 -3764 1447 -3712
rect 285 -3856 1333 -3822
rect 1806 -3822 1840 -3259
rect 1956 -3225 1990 -3094
rect 2148 -3225 2182 -3094
rect 2340 -3225 2374 -3094
rect 2532 -3225 2566 -3094
rect 2724 -3225 2758 -3094
rect 2916 -3225 2950 -3094
rect 3265 -3216 3317 -2669
rect 3040 -3225 3317 -3216
rect 1956 -3259 3317 -3225
rect 1956 -3400 1990 -3259
rect 2148 -3400 2182 -3259
rect 2340 -3400 2374 -3259
rect 2532 -3400 2566 -3259
rect 2724 -3400 2758 -3259
rect 2916 -3400 2950 -3259
rect 3040 -3268 3317 -3259
rect 1950 -3412 1996 -3400
rect 1950 -3660 1956 -3412
rect 1990 -3660 1996 -3412
rect 1950 -3672 1996 -3660
rect 2046 -3412 2092 -3400
rect 2046 -3660 2052 -3412
rect 2086 -3660 2092 -3412
rect 2046 -3672 2092 -3660
rect 2142 -3412 2188 -3400
rect 2142 -3660 2148 -3412
rect 2182 -3660 2188 -3412
rect 2142 -3672 2188 -3660
rect 2238 -3412 2284 -3400
rect 2238 -3660 2244 -3412
rect 2278 -3660 2284 -3412
rect 2238 -3672 2284 -3660
rect 2334 -3412 2380 -3400
rect 2334 -3660 2340 -3412
rect 2374 -3660 2380 -3412
rect 2334 -3672 2380 -3660
rect 2430 -3412 2476 -3400
rect 2430 -3660 2436 -3412
rect 2470 -3660 2476 -3412
rect 2430 -3672 2476 -3660
rect 2526 -3412 2572 -3400
rect 2526 -3660 2532 -3412
rect 2566 -3660 2572 -3412
rect 2526 -3672 2572 -3660
rect 2622 -3412 2668 -3400
rect 2622 -3660 2628 -3412
rect 2662 -3660 2668 -3412
rect 2622 -3672 2668 -3660
rect 2718 -3412 2764 -3400
rect 2718 -3660 2724 -3412
rect 2758 -3660 2764 -3412
rect 2718 -3672 2764 -3660
rect 2814 -3412 2860 -3400
rect 2814 -3660 2820 -3412
rect 2854 -3660 2860 -3412
rect 2814 -3672 2860 -3660
rect 2910 -3412 2956 -3400
rect 2910 -3660 2916 -3412
rect 2950 -3660 2956 -3412
rect 2910 -3672 2956 -3660
rect 1936 -3764 1946 -3712
rect 1998 -3764 2008 -3712
rect 2052 -3822 2086 -3672
rect 2244 -3822 2278 -3672
rect 2436 -3822 2470 -3672
rect 2628 -3822 2662 -3672
rect 2820 -3822 2854 -3672
rect 2896 -3764 2906 -3712
rect 2958 -3764 2968 -3712
rect 1806 -3856 2854 -3822
rect -579 -3961 -236 -3951
rect -579 -3995 -539 -3961
rect -505 -3995 -236 -3961
rect -579 -4003 -236 -3995
rect -184 -4003 -173 -3951
rect -91 -4114 -81 -4111
rect -465 -4120 -81 -4114
rect -465 -4154 -453 -4120
rect -419 -4154 -81 -4120
rect -465 -4160 -81 -4154
rect -91 -4163 -81 -4160
rect -29 -4163 -19 -4111
rect -3266 -4226 -2218 -4192
rect -3266 -4780 -3232 -4226
rect -3020 -4376 -2986 -4226
rect -2828 -4376 -2794 -4226
rect -2636 -4376 -2602 -4226
rect -2444 -4376 -2410 -4226
rect -2367 -4336 -2357 -4284
rect -2305 -4336 -2295 -4284
rect -2252 -4376 -2218 -4226
rect 285 -4226 1333 -4192
rect -704 -4268 -336 -4237
rect -2174 -4336 -2164 -4284
rect -2112 -4336 -2102 -4284
rect -1953 -4336 -1943 -4284
rect -1891 -4336 -1416 -4284
rect -1364 -4336 -1354 -4284
rect -704 -4302 -675 -4268
rect -641 -4302 -583 -4268
rect -549 -4302 -491 -4268
rect -457 -4302 -399 -4268
rect -365 -4302 -336 -4268
rect -704 -4333 -336 -4302
rect -3122 -4388 -3076 -4376
rect -3122 -4636 -3116 -4388
rect -3082 -4636 -3076 -4388
rect -3122 -4648 -3076 -4636
rect -3026 -4388 -2980 -4376
rect -3026 -4636 -3020 -4388
rect -2986 -4636 -2980 -4388
rect -3026 -4648 -2980 -4636
rect -2930 -4388 -2884 -4376
rect -2930 -4636 -2924 -4388
rect -2890 -4636 -2884 -4388
rect -2930 -4648 -2884 -4636
rect -2834 -4388 -2788 -4376
rect -2834 -4636 -2828 -4388
rect -2794 -4636 -2788 -4388
rect -2834 -4648 -2788 -4636
rect -2738 -4388 -2692 -4376
rect -2738 -4636 -2732 -4388
rect -2698 -4636 -2692 -4388
rect -2738 -4648 -2692 -4636
rect -2642 -4388 -2596 -4376
rect -2642 -4636 -2636 -4388
rect -2602 -4636 -2596 -4388
rect -2642 -4648 -2596 -4636
rect -2546 -4388 -2500 -4376
rect -2546 -4636 -2540 -4388
rect -2506 -4636 -2500 -4388
rect -2546 -4648 -2500 -4636
rect -2450 -4388 -2404 -4376
rect -2450 -4636 -2444 -4388
rect -2410 -4636 -2404 -4388
rect -2450 -4648 -2404 -4636
rect -2354 -4388 -2308 -4376
rect -2354 -4636 -2348 -4388
rect -2314 -4636 -2308 -4388
rect -2354 -4648 -2308 -4636
rect -2258 -4388 -2212 -4376
rect -2258 -4636 -2252 -4388
rect -2218 -4636 -2212 -4388
rect -2258 -4648 -2212 -4636
rect -2162 -4388 -2116 -4376
rect -2162 -4636 -2156 -4388
rect -2122 -4636 -2116 -4388
rect 82 -4412 92 -4409
rect -464 -4418 92 -4412
rect -464 -4452 -452 -4418
rect -418 -4452 92 -4418
rect -464 -4458 92 -4452
rect 82 -4461 92 -4458
rect 144 -4461 154 -4409
rect -558 -4617 -548 -4565
rect -496 -4617 -486 -4565
rect 285 -4593 319 -4226
rect 415 -4328 425 -4276
rect 477 -4328 487 -4276
rect 531 -4368 565 -4226
rect 723 -4368 757 -4226
rect 915 -4368 949 -4226
rect 1107 -4368 1141 -4226
rect 1299 -4368 1333 -4226
rect 1806 -4226 2854 -4192
rect 1377 -4330 1387 -4278
rect 1439 -4330 1449 -4278
rect 429 -4380 475 -4368
rect 429 -4460 435 -4380
rect 469 -4460 475 -4380
rect 429 -4472 475 -4460
rect 525 -4380 571 -4368
rect 525 -4460 531 -4380
rect 565 -4460 571 -4380
rect 525 -4472 571 -4460
rect 621 -4380 667 -4368
rect 621 -4460 627 -4380
rect 661 -4460 667 -4380
rect 621 -4472 667 -4460
rect 717 -4380 763 -4368
rect 717 -4460 723 -4380
rect 757 -4460 763 -4380
rect 717 -4472 763 -4460
rect 813 -4380 859 -4368
rect 813 -4460 819 -4380
rect 853 -4460 859 -4380
rect 813 -4472 859 -4460
rect 909 -4380 955 -4368
rect 909 -4460 915 -4380
rect 949 -4460 955 -4380
rect 909 -4472 955 -4460
rect 1005 -4380 1051 -4368
rect 1005 -4460 1011 -4380
rect 1045 -4460 1051 -4380
rect 1005 -4472 1051 -4460
rect 1101 -4380 1147 -4368
rect 1101 -4460 1107 -4380
rect 1141 -4460 1147 -4380
rect 1101 -4472 1147 -4460
rect 1197 -4380 1243 -4368
rect 1197 -4460 1203 -4380
rect 1237 -4460 1243 -4380
rect 1197 -4472 1243 -4460
rect 1293 -4380 1339 -4368
rect 1293 -4460 1299 -4380
rect 1333 -4460 1339 -4380
rect 1293 -4472 1339 -4460
rect 1389 -4380 1435 -4368
rect 1389 -4460 1395 -4380
rect 1429 -4460 1435 -4380
rect 1389 -4472 1435 -4460
rect 1503 -4375 1549 -4363
rect 1609 -4375 1655 -4374
rect 215 -4603 319 -4593
rect -2162 -4648 -2116 -4636
rect -48 -4637 319 -4603
rect -3461 -4832 -3232 -4780
rect -3266 -5200 -3232 -4832
rect -3116 -4789 -3082 -4648
rect -2924 -4789 -2890 -4648
rect -2732 -4789 -2698 -4648
rect -2540 -4789 -2506 -4648
rect -2348 -4789 -2314 -4648
rect -2156 -4789 -2122 -4648
rect -48 -4674 -14 -4637
rect 215 -4645 319 -4637
rect -1808 -4708 -14 -4674
rect -1808 -4789 -1774 -4708
rect -3116 -4823 -1774 -4789
rect -704 -4812 -336 -4781
rect -3116 -4954 -3082 -4823
rect -2924 -4954 -2890 -4823
rect -2732 -4954 -2698 -4823
rect -2540 -4954 -2506 -4823
rect -2348 -4954 -2314 -4823
rect -2156 -4954 -2122 -4823
rect -704 -4846 -675 -4812
rect -641 -4846 -583 -4812
rect -549 -4846 -491 -4812
rect -457 -4846 -399 -4812
rect -365 -4846 -336 -4812
rect -704 -4877 -336 -4846
rect -3122 -4966 -3076 -4954
rect -3122 -5046 -3116 -4966
rect -3082 -5046 -3076 -4966
rect -3122 -5058 -3076 -5046
rect -3026 -4966 -2980 -4954
rect -3026 -5046 -3020 -4966
rect -2986 -5046 -2980 -4966
rect -3026 -5058 -2980 -5046
rect -2930 -4966 -2884 -4954
rect -2930 -5046 -2924 -4966
rect -2890 -5046 -2884 -4966
rect -2930 -5058 -2884 -5046
rect -2834 -4966 -2788 -4954
rect -2834 -5046 -2828 -4966
rect -2794 -5046 -2788 -4966
rect -2834 -5058 -2788 -5046
rect -2738 -4966 -2692 -4954
rect -2738 -5046 -2732 -4966
rect -2698 -5046 -2692 -4966
rect -2738 -5058 -2692 -5046
rect -2642 -4966 -2596 -4954
rect -2642 -5046 -2636 -4966
rect -2602 -5046 -2596 -4966
rect -2642 -5058 -2596 -5046
rect -2546 -4966 -2500 -4954
rect -2546 -5046 -2540 -4966
rect -2506 -5046 -2500 -4966
rect -2546 -5058 -2500 -5046
rect -2450 -4966 -2404 -4954
rect -2450 -5046 -2444 -4966
rect -2410 -5046 -2404 -4966
rect -2450 -5058 -2404 -5046
rect -2354 -4966 -2308 -4954
rect -2354 -5046 -2348 -4966
rect -2314 -5046 -2308 -4966
rect -2354 -5058 -2308 -5046
rect -2258 -4966 -2212 -4954
rect -2258 -5046 -2252 -4966
rect -2218 -5046 -2212 -4966
rect -2258 -5058 -2212 -5046
rect -2162 -4966 -2116 -4954
rect -2162 -5046 -2156 -4966
rect -2122 -5046 -2116 -4966
rect -2162 -5058 -2116 -5046
rect -3020 -5200 -2986 -5058
rect -2828 -5200 -2794 -5058
rect -2636 -5200 -2602 -5058
rect -2444 -5200 -2410 -5058
rect -2368 -5149 -2358 -5097
rect -2306 -5149 -2296 -5097
rect -2252 -5200 -2218 -5058
rect -2173 -5149 -2163 -5097
rect -2111 -5149 -2101 -5097
rect -3266 -5234 -2218 -5200
rect 285 -5200 319 -4645
rect 435 -4603 469 -4472
rect 627 -4603 661 -4472
rect 819 -4603 853 -4472
rect 1011 -4603 1045 -4472
rect 1203 -4603 1237 -4472
rect 1395 -4603 1429 -4472
rect 1503 -4475 1509 -4375
rect 1543 -4386 1655 -4375
rect 1543 -4462 1615 -4386
rect 1649 -4462 1655 -4386
rect 1543 -4474 1655 -4462
rect 1697 -4375 1743 -4374
rect 1806 -4375 1840 -4226
rect 1938 -4330 1948 -4278
rect 2000 -4330 2010 -4278
rect 2052 -4368 2086 -4226
rect 2244 -4368 2278 -4226
rect 2436 -4368 2470 -4226
rect 2628 -4368 2662 -4226
rect 2820 -4368 2854 -4226
rect 2898 -4330 2908 -4278
rect 2960 -4330 2970 -4278
rect 1697 -4386 1840 -4375
rect 1697 -4462 1703 -4386
rect 1737 -4462 1840 -4386
rect 1697 -4474 1840 -4462
rect 1950 -4380 1996 -4368
rect 1950 -4460 1956 -4380
rect 1990 -4460 1996 -4380
rect 1950 -4472 1996 -4460
rect 2046 -4380 2092 -4368
rect 2046 -4460 2052 -4380
rect 2086 -4460 2092 -4380
rect 2046 -4472 2092 -4460
rect 2142 -4380 2188 -4368
rect 2142 -4460 2148 -4380
rect 2182 -4460 2188 -4380
rect 2142 -4472 2188 -4460
rect 2238 -4380 2284 -4368
rect 2238 -4460 2244 -4380
rect 2278 -4460 2284 -4380
rect 2238 -4472 2284 -4460
rect 2334 -4380 2380 -4368
rect 2334 -4460 2340 -4380
rect 2374 -4460 2380 -4380
rect 2334 -4472 2380 -4460
rect 2430 -4380 2476 -4368
rect 2430 -4460 2436 -4380
rect 2470 -4460 2476 -4380
rect 2430 -4472 2476 -4460
rect 2526 -4380 2572 -4368
rect 2526 -4460 2532 -4380
rect 2566 -4460 2572 -4380
rect 2526 -4472 2572 -4460
rect 2622 -4380 2668 -4368
rect 2622 -4460 2628 -4380
rect 2662 -4460 2668 -4380
rect 2622 -4472 2668 -4460
rect 2718 -4380 2764 -4368
rect 2718 -4460 2724 -4380
rect 2758 -4460 2764 -4380
rect 2718 -4472 2764 -4460
rect 2814 -4380 2860 -4368
rect 2814 -4460 2820 -4380
rect 2854 -4460 2860 -4380
rect 2814 -4472 2860 -4460
rect 2910 -4380 2956 -4368
rect 2910 -4460 2916 -4380
rect 2950 -4460 2956 -4380
rect 2910 -4472 2956 -4460
rect 1543 -4475 1649 -4474
rect 1703 -4475 1840 -4474
rect 1503 -4487 1549 -4475
rect 1647 -4512 1705 -4506
rect 1647 -4513 1659 -4512
rect 1693 -4513 1705 -4512
rect 1640 -4565 1650 -4513
rect 1702 -4565 1712 -4513
rect 1806 -4603 1840 -4475
rect 435 -4637 1840 -4603
rect 435 -4778 469 -4637
rect 627 -4778 661 -4637
rect 819 -4778 853 -4637
rect 1011 -4778 1045 -4637
rect 1203 -4778 1237 -4637
rect 1395 -4778 1429 -4637
rect 429 -4790 475 -4778
rect 429 -5038 435 -4790
rect 469 -5038 475 -4790
rect 429 -5050 475 -5038
rect 525 -4790 571 -4778
rect 525 -5038 531 -4790
rect 565 -5038 571 -4790
rect 525 -5050 571 -5038
rect 621 -4790 667 -4778
rect 621 -5038 627 -4790
rect 661 -5038 667 -4790
rect 621 -5050 667 -5038
rect 717 -4790 763 -4778
rect 717 -5038 723 -4790
rect 757 -5038 763 -4790
rect 717 -5050 763 -5038
rect 813 -4790 859 -4778
rect 813 -5038 819 -4790
rect 853 -5038 859 -4790
rect 813 -5050 859 -5038
rect 909 -4790 955 -4778
rect 909 -5038 915 -4790
rect 949 -5038 955 -4790
rect 909 -5050 955 -5038
rect 1005 -4790 1051 -4778
rect 1005 -5038 1011 -4790
rect 1045 -5038 1051 -4790
rect 1005 -5050 1051 -5038
rect 1101 -4790 1147 -4778
rect 1101 -5038 1107 -4790
rect 1141 -5038 1147 -4790
rect 1101 -5050 1147 -5038
rect 1197 -4790 1243 -4778
rect 1197 -5038 1203 -4790
rect 1237 -5038 1243 -4790
rect 1197 -5050 1243 -5038
rect 1293 -4790 1339 -4778
rect 1293 -5038 1299 -4790
rect 1333 -5038 1339 -4790
rect 1293 -5050 1339 -5038
rect 1389 -4790 1435 -4778
rect 1389 -5038 1395 -4790
rect 1429 -5038 1435 -4790
rect 1389 -5050 1435 -5038
rect 416 -5141 426 -5089
rect 478 -5141 488 -5089
rect 531 -5200 565 -5050
rect 723 -5200 757 -5050
rect 915 -5200 949 -5050
rect 1107 -5200 1141 -5050
rect 1299 -5200 1333 -5050
rect 1375 -5142 1385 -5090
rect 1437 -5142 1447 -5090
rect 285 -5234 1333 -5200
rect 1806 -5200 1840 -4637
rect 1956 -4603 1990 -4472
rect 2148 -4603 2182 -4472
rect 2340 -4603 2374 -4472
rect 2532 -4603 2566 -4472
rect 2724 -4603 2758 -4472
rect 2916 -4603 2950 -4472
rect 3265 -4595 3317 -3268
rect 3043 -4603 3317 -4595
rect 1956 -4637 3317 -4603
rect 1956 -4778 1990 -4637
rect 2148 -4778 2182 -4637
rect 2340 -4778 2374 -4637
rect 2532 -4778 2566 -4637
rect 2724 -4778 2758 -4637
rect 2916 -4778 2950 -4637
rect 3043 -4647 3317 -4637
rect 1950 -4790 1996 -4778
rect 1950 -5038 1956 -4790
rect 1990 -5038 1996 -4790
rect 1950 -5050 1996 -5038
rect 2046 -4790 2092 -4778
rect 2046 -5038 2052 -4790
rect 2086 -5038 2092 -4790
rect 2046 -5050 2092 -5038
rect 2142 -4790 2188 -4778
rect 2142 -5038 2148 -4790
rect 2182 -5038 2188 -4790
rect 2142 -5050 2188 -5038
rect 2238 -4790 2284 -4778
rect 2238 -5038 2244 -4790
rect 2278 -5038 2284 -4790
rect 2238 -5050 2284 -5038
rect 2334 -4790 2380 -4778
rect 2334 -5038 2340 -4790
rect 2374 -5038 2380 -4790
rect 2334 -5050 2380 -5038
rect 2430 -4790 2476 -4778
rect 2430 -5038 2436 -4790
rect 2470 -5038 2476 -4790
rect 2430 -5050 2476 -5038
rect 2526 -4790 2572 -4778
rect 2526 -5038 2532 -4790
rect 2566 -5038 2572 -4790
rect 2526 -5050 2572 -5038
rect 2622 -4790 2668 -4778
rect 2622 -5038 2628 -4790
rect 2662 -5038 2668 -4790
rect 2622 -5050 2668 -5038
rect 2718 -4790 2764 -4778
rect 2718 -5038 2724 -4790
rect 2758 -5038 2764 -4790
rect 2718 -5050 2764 -5038
rect 2814 -4790 2860 -4778
rect 2814 -5038 2820 -4790
rect 2854 -5038 2860 -4790
rect 2814 -5050 2860 -5038
rect 2910 -4790 2956 -4778
rect 2910 -5038 2916 -4790
rect 2950 -5038 2956 -4790
rect 2910 -5050 2956 -5038
rect 1936 -5142 1946 -5090
rect 1998 -5142 2008 -5090
rect 2052 -5200 2086 -5050
rect 2244 -5200 2278 -5050
rect 2436 -5200 2470 -5050
rect 2628 -5200 2662 -5050
rect 2820 -5200 2854 -5050
rect 2896 -5142 2906 -5090
rect 2958 -5142 2968 -5090
rect 1806 -5234 2854 -5200
<< via1 >>
rect -1587 -121 -1535 -69
rect -914 -121 -862 -69
rect -2357 -201 -2305 -195
rect -2357 -235 -2348 -201
rect -2348 -235 -2314 -201
rect -2314 -235 -2305 -201
rect -2357 -247 -2305 -235
rect -2163 -204 -2111 -194
rect -2163 -238 -2156 -204
rect -2156 -238 -2122 -204
rect -2122 -238 -2111 -204
rect -2163 -246 -2111 -238
rect -1942 -246 -1890 -194
rect -1416 -246 -1364 -194
rect 425 -197 477 -186
rect 425 -231 435 -197
rect 435 -231 469 -197
rect 469 -231 477 -197
rect 425 -238 477 -231
rect 1387 -197 1439 -188
rect 1387 -231 1395 -197
rect 1395 -231 1429 -197
rect 1429 -231 1439 -197
rect 1387 -240 1439 -231
rect -1416 -645 -1364 -593
rect -461 -594 -409 -584
rect -461 -628 -452 -594
rect -452 -628 -418 -594
rect -418 -628 -409 -594
rect -461 -636 -409 -628
rect -914 -698 -862 -690
rect -914 -732 -905 -698
rect -905 -732 -871 -698
rect -871 -732 -862 -698
rect -914 -742 -862 -732
rect -549 -700 -497 -694
rect -549 -734 -538 -700
rect -538 -734 -504 -700
rect -504 -734 -497 -700
rect -549 -746 -497 -734
rect -2357 -1019 -2305 -1008
rect -2357 -1053 -2345 -1019
rect -2345 -1053 -2311 -1019
rect -2311 -1053 -2305 -1019
rect -2357 -1060 -2305 -1053
rect -2166 -1016 -2114 -1006
rect -2166 -1050 -2155 -1016
rect -2155 -1050 -2121 -1016
rect -2121 -1050 -2114 -1016
rect -2166 -1058 -2114 -1050
rect 1948 -197 2000 -188
rect 1948 -231 1956 -197
rect 1956 -231 1990 -197
rect 1990 -231 2000 -197
rect 1948 -240 2000 -231
rect 2908 -197 2960 -188
rect 2908 -231 2916 -197
rect 2916 -231 2950 -197
rect 2950 -231 2960 -197
rect 2908 -240 2960 -231
rect 1650 -456 1659 -423
rect 1659 -456 1693 -423
rect 1693 -456 1702 -423
rect 1650 -475 1702 -456
rect 426 -1008 478 -999
rect 426 -1042 435 -1008
rect 435 -1042 469 -1008
rect 469 -1042 478 -1008
rect 426 -1051 478 -1042
rect 1385 -1008 1437 -1000
rect 1385 -1042 1395 -1008
rect 1395 -1042 1429 -1008
rect 1429 -1042 1437 -1008
rect 1385 -1052 1437 -1042
rect 1946 -1008 1998 -1000
rect 1946 -1042 1956 -1008
rect 1956 -1042 1990 -1008
rect 1990 -1042 1998 -1008
rect 1946 -1052 1998 -1042
rect 2906 -1008 2958 -1000
rect 2906 -1042 2916 -1008
rect 2916 -1042 2950 -1008
rect 2950 -1042 2958 -1008
rect 2906 -1052 2958 -1042
rect 98 -1240 150 -1188
rect -287 -1355 -235 -1303
rect -2357 -1538 -2305 -1528
rect -2357 -1572 -2348 -1538
rect -2348 -1572 -2314 -1538
rect -2314 -1572 -2305 -1538
rect -2357 -1580 -2305 -1572
rect -2165 -1538 -2113 -1529
rect -2165 -1572 -2156 -1538
rect -2156 -1572 -2122 -1538
rect -2122 -1572 -2113 -1538
rect -2165 -1581 -2113 -1572
rect -1724 -1580 -1672 -1528
rect -1416 -1580 -1364 -1528
rect -478 -1676 -426 -1669
rect -478 -1710 -469 -1676
rect -469 -1710 -435 -1676
rect -435 -1710 -426 -1676
rect -478 -1721 -426 -1710
rect -592 -1784 -540 -1776
rect -592 -1818 -582 -1784
rect -582 -1818 -548 -1784
rect -548 -1818 -540 -1784
rect -592 -1828 -540 -1818
rect -416 -1785 -364 -1779
rect -416 -1819 -408 -1785
rect -408 -1819 -374 -1785
rect -374 -1819 -364 -1785
rect -416 -1831 -364 -1819
rect 425 -1531 477 -1520
rect 425 -1565 435 -1531
rect 435 -1565 469 -1531
rect 469 -1565 477 -1531
rect 425 -1572 477 -1565
rect 1387 -1531 1439 -1522
rect 1387 -1565 1395 -1531
rect 1395 -1565 1429 -1531
rect 1429 -1565 1439 -1531
rect 1387 -1574 1439 -1565
rect -872 -1971 -820 -1919
rect -416 -1971 -364 -1919
rect -592 -2277 -540 -2225
rect -2356 -2349 -2304 -2341
rect -2356 -2383 -2348 -2349
rect -2348 -2383 -2314 -2349
rect -2314 -2383 -2304 -2349
rect -2356 -2393 -2304 -2383
rect -287 -2313 -235 -2261
rect -2164 -2349 -2112 -2340
rect -2164 -2383 -2156 -2349
rect -2156 -2383 -2122 -2349
rect -2122 -2383 -2112 -2349
rect -2164 -2392 -2112 -2383
rect -1101 -2398 -1049 -2388
rect -1101 -2432 -1091 -2398
rect -1091 -2432 -1057 -2398
rect -1057 -2432 -1049 -2398
rect -1101 -2440 -1049 -2432
rect -762 -2440 -710 -2388
rect -592 -2398 -540 -2390
rect -592 -2432 -583 -2398
rect -583 -2432 -549 -2398
rect -549 -2432 -540 -2398
rect -592 -2442 -540 -2432
rect -412 -2395 -360 -2385
rect -412 -2429 -402 -2395
rect -402 -2429 -368 -2395
rect -368 -2429 -360 -2395
rect -412 -2437 -360 -2429
rect 1948 -1531 2000 -1522
rect 1948 -1565 1956 -1531
rect 1956 -1565 1990 -1531
rect 1990 -1565 2000 -1531
rect 1948 -1574 2000 -1565
rect 2908 -1531 2960 -1522
rect 2908 -1565 2916 -1531
rect 2916 -1565 2950 -1531
rect 2950 -1565 2960 -1531
rect 2908 -1574 2960 -1565
rect 1650 -1790 1659 -1757
rect 1659 -1790 1693 -1757
rect 1693 -1790 1702 -1757
rect 1650 -1809 1702 -1790
rect 426 -2342 478 -2333
rect 426 -2376 435 -2342
rect 435 -2376 469 -2342
rect 469 -2376 478 -2342
rect 426 -2385 478 -2376
rect 1385 -2342 1437 -2334
rect 1385 -2376 1395 -2342
rect 1395 -2376 1429 -2342
rect 1429 -2376 1437 -2342
rect 1385 -2386 1437 -2376
rect 1946 -2342 1998 -2334
rect 1946 -2376 1956 -2342
rect 1956 -2376 1990 -2342
rect 1990 -2376 1998 -2342
rect 1946 -2386 1998 -2376
rect 2906 -2342 2958 -2334
rect 2906 -2376 2916 -2342
rect 2916 -2376 2950 -2342
rect 2950 -2376 2958 -2342
rect 2906 -2386 2958 -2376
rect -1240 -2543 -1188 -2491
rect -412 -2543 -360 -2491
rect -762 -2827 -710 -2775
rect -412 -2827 -360 -2775
rect -2357 -2916 -2305 -2906
rect -2357 -2950 -2348 -2916
rect -2348 -2950 -2314 -2916
rect -2314 -2950 -2305 -2916
rect -2357 -2958 -2305 -2950
rect -2165 -2916 -2113 -2907
rect -2165 -2950 -2156 -2916
rect -2156 -2950 -2122 -2916
rect -2122 -2950 -2113 -2916
rect -2165 -2959 -2113 -2950
rect -1926 -2958 -1874 -2906
rect -1416 -2958 -1364 -2906
rect -1098 -2874 -1046 -2865
rect -1098 -2908 -1089 -2874
rect -1089 -2908 -1055 -2874
rect -1055 -2908 -1046 -2874
rect -1098 -2917 -1046 -2908
rect -872 -2916 -820 -2864
rect -412 -2875 -360 -2866
rect -412 -2909 -401 -2875
rect -401 -2909 -367 -2875
rect -367 -2909 -360 -2875
rect -412 -2918 -360 -2909
rect -236 -3078 -184 -3026
rect 425 -2909 477 -2898
rect 425 -2943 435 -2909
rect 435 -2943 469 -2909
rect 469 -2943 477 -2909
rect 425 -2950 477 -2943
rect 1387 -2909 1439 -2900
rect 1387 -2943 1395 -2909
rect 1395 -2943 1429 -2909
rect 1429 -2943 1439 -2909
rect 1387 -2952 1439 -2943
rect -762 -3445 -710 -3393
rect -414 -3445 -362 -3393
rect -1241 -3539 -1187 -3485
rect -414 -3487 -362 -3474
rect -414 -3521 -405 -3487
rect -405 -3521 -371 -3487
rect -371 -3521 -362 -3487
rect -414 -3526 -362 -3521
rect -500 -3590 -448 -3580
rect -500 -3624 -492 -3590
rect -492 -3624 -458 -3590
rect -458 -3624 -448 -3590
rect -500 -3632 -448 -3624
rect -2356 -3727 -2304 -3715
rect -2356 -3761 -2348 -3727
rect -2348 -3761 -2314 -3727
rect -2314 -3761 -2304 -3727
rect -2356 -3767 -2304 -3761
rect -2164 -3727 -2112 -3717
rect -2164 -3761 -2156 -3727
rect -2156 -3761 -2122 -3727
rect -2122 -3761 -2112 -3727
rect -2164 -3769 -2112 -3761
rect -235 -3764 -183 -3712
rect 140 -3764 192 -3712
rect 1948 -2909 2000 -2900
rect 1948 -2943 1956 -2909
rect 1956 -2943 1990 -2909
rect 1990 -2943 2000 -2909
rect 1948 -2952 2000 -2943
rect 2908 -2909 2960 -2900
rect 2908 -2943 2916 -2909
rect 2916 -2943 2950 -2909
rect 2950 -2943 2960 -2909
rect 2908 -2952 2960 -2943
rect 1650 -3168 1659 -3135
rect 1659 -3168 1693 -3135
rect 1693 -3168 1702 -3135
rect 1650 -3187 1702 -3168
rect 426 -3720 478 -3711
rect 426 -3754 435 -3720
rect 435 -3754 469 -3720
rect 469 -3754 478 -3720
rect 426 -3763 478 -3754
rect 1385 -3720 1437 -3712
rect 1385 -3754 1395 -3720
rect 1395 -3754 1429 -3720
rect 1429 -3754 1437 -3720
rect 1385 -3764 1437 -3754
rect 1946 -3720 1998 -3712
rect 1946 -3754 1956 -3720
rect 1956 -3754 1990 -3720
rect 1990 -3754 1998 -3720
rect 1946 -3764 1998 -3754
rect 2906 -3720 2958 -3712
rect 2906 -3754 2916 -3720
rect 2916 -3754 2950 -3720
rect 2950 -3754 2958 -3720
rect 2906 -3764 2958 -3754
rect -236 -4003 -184 -3951
rect -81 -4163 -29 -4111
rect -2357 -4294 -2305 -4284
rect -2357 -4328 -2348 -4294
rect -2348 -4328 -2314 -4294
rect -2314 -4328 -2305 -4294
rect -2357 -4336 -2305 -4328
rect -2164 -4294 -2112 -4284
rect -2164 -4328 -2156 -4294
rect -2156 -4328 -2122 -4294
rect -2122 -4328 -2112 -4294
rect -2164 -4336 -2112 -4328
rect -1943 -4336 -1891 -4284
rect -1416 -4336 -1364 -4284
rect 92 -4461 144 -4409
rect -548 -4574 -496 -4565
rect -548 -4608 -540 -4574
rect -540 -4608 -506 -4574
rect -506 -4608 -496 -4574
rect -548 -4617 -496 -4608
rect 425 -4287 477 -4276
rect 425 -4321 435 -4287
rect 435 -4321 469 -4287
rect 469 -4321 477 -4287
rect 425 -4328 477 -4321
rect 1387 -4287 1439 -4278
rect 1387 -4321 1395 -4287
rect 1395 -4321 1429 -4287
rect 1429 -4321 1439 -4287
rect 1387 -4330 1439 -4321
rect -2358 -5105 -2306 -5097
rect -2358 -5139 -2348 -5105
rect -2348 -5139 -2314 -5105
rect -2314 -5139 -2306 -5105
rect -2358 -5149 -2306 -5139
rect -2163 -5105 -2111 -5097
rect -2163 -5139 -2156 -5105
rect -2156 -5139 -2122 -5105
rect -2122 -5139 -2111 -5105
rect -2163 -5149 -2111 -5139
rect 1948 -4287 2000 -4278
rect 1948 -4321 1956 -4287
rect 1956 -4321 1990 -4287
rect 1990 -4321 2000 -4287
rect 1948 -4330 2000 -4321
rect 2908 -4287 2960 -4278
rect 2908 -4321 2916 -4287
rect 2916 -4321 2950 -4287
rect 2950 -4321 2960 -4287
rect 2908 -4330 2960 -4321
rect 1650 -4546 1659 -4513
rect 1659 -4546 1693 -4513
rect 1693 -4546 1702 -4513
rect 1650 -4565 1702 -4546
rect 426 -5098 478 -5089
rect 426 -5132 435 -5098
rect 435 -5132 469 -5098
rect 469 -5132 478 -5098
rect 426 -5141 478 -5132
rect 1385 -5098 1437 -5090
rect 1385 -5132 1395 -5098
rect 1395 -5132 1429 -5098
rect 1429 -5132 1437 -5098
rect 1385 -5142 1437 -5132
rect 1946 -5098 1998 -5090
rect 1946 -5132 1956 -5098
rect 1956 -5132 1990 -5098
rect 1990 -5132 1998 -5098
rect 1946 -5142 1998 -5132
rect 2906 -5098 2958 -5090
rect 2906 -5132 2916 -5098
rect 2916 -5132 2950 -5098
rect 2950 -5132 2958 -5098
rect 2906 -5142 2958 -5132
<< metal2 >>
rect -1587 -69 -1535 148
rect -2357 -194 -2305 -185
rect -2163 -194 -2111 -184
rect -1942 -194 -1890 -184
rect -2357 -195 -2163 -194
rect -2305 -246 -2163 -195
rect -2111 -246 -1942 -194
rect -2357 -257 -2305 -247
rect -2163 -256 -2111 -246
rect -1942 -256 -1890 -246
rect -2357 -1001 -2305 -998
rect -2166 -1001 -2114 -996
rect -1587 -1001 -1535 -121
rect -2357 -1006 -1535 -1001
rect -2357 -1008 -2166 -1006
rect -2305 -1053 -2166 -1008
rect -2357 -1070 -2305 -1060
rect -2114 -1053 -1535 -1006
rect -2166 -1068 -2114 -1058
rect -2357 -1528 -2305 -1518
rect -2165 -1528 -2113 -1519
rect -1724 -1528 -1672 -1518
rect -2365 -1580 -2357 -1528
rect -2305 -1529 -1724 -1528
rect -2305 -1580 -2165 -1529
rect -2357 -1590 -2305 -1580
rect -2113 -1580 -1724 -1529
rect -2165 -1591 -2113 -1581
rect -1724 -1590 -1672 -1580
rect -2356 -2335 -2304 -2331
rect -2164 -2335 -2112 -2330
rect -1587 -2335 -1535 -1053
rect -2360 -2340 -1535 -2335
rect -2360 -2341 -2164 -2340
rect -2360 -2387 -2356 -2341
rect -2304 -2387 -2164 -2341
rect -2356 -2403 -2304 -2393
rect -2112 -2387 -1535 -2340
rect -2164 -2402 -2112 -2392
rect -2357 -2906 -2305 -2896
rect -2165 -2906 -2113 -2897
rect -1926 -2906 -1874 -2896
rect -2305 -2907 -1926 -2906
rect -2305 -2958 -2165 -2907
rect -2357 -2968 -2305 -2958
rect -2113 -2958 -1926 -2907
rect -2165 -2969 -2113 -2959
rect -1926 -2968 -1874 -2958
rect -2356 -3713 -2304 -3705
rect -2164 -3713 -2112 -3707
rect -1587 -3713 -1535 -2387
rect -1416 -194 -1364 -184
rect -1416 -593 -1364 -246
rect -1416 -1528 -1364 -645
rect -1416 -2906 -1364 -1580
rect -2356 -3715 -1532 -3713
rect -2304 -3717 -1532 -3715
rect -2304 -3765 -2164 -3717
rect -2356 -3777 -2304 -3767
rect -2112 -3765 -1532 -3717
rect -2164 -3779 -2112 -3769
rect -2357 -4284 -2305 -4274
rect -2164 -4284 -2112 -4274
rect -1943 -4284 -1891 -4274
rect -2361 -4336 -2357 -4284
rect -2305 -4336 -2164 -4284
rect -2112 -4336 -1943 -4284
rect -2357 -4346 -2305 -4336
rect -2164 -4346 -2112 -4336
rect -1943 -4346 -1891 -4336
rect -2358 -5091 -2306 -5087
rect -2163 -5091 -2111 -5087
rect -1587 -5091 -1535 -3765
rect -1416 -4284 -1364 -2958
rect -1241 -2491 -1187 148
rect -1101 -2388 -1049 148
rect -914 -69 -862 -60
rect -914 -690 -862 -121
rect 425 -186 477 -176
rect -461 -238 425 -193
rect 517 -193 583 -181
rect 1387 -188 1439 -178
rect 477 -238 1387 -193
rect -461 -240 1387 -238
rect 1948 -188 2000 -178
rect 1439 -240 1948 -193
rect 2908 -188 2960 -178
rect 2000 -240 2908 -193
rect -461 -245 2960 -240
rect -461 -584 -409 -245
rect 425 -248 477 -245
rect 517 -247 583 -245
rect 1387 -250 1439 -245
rect 1948 -250 2000 -245
rect 2908 -250 2960 -245
rect -461 -646 -409 -636
rect 1650 -423 1702 -413
rect -914 -752 -862 -742
rect -549 -694 -497 -684
rect -497 -746 -426 -694
rect -549 -756 -426 -746
rect -478 -1000 -426 -756
rect 426 -999 478 -989
rect -478 -1051 426 -1000
rect 1385 -1000 1437 -990
rect 1650 -1000 1702 -475
rect 1946 -1000 1998 -990
rect 2906 -1000 2958 -990
rect 478 -1051 1385 -1000
rect -478 -1052 1385 -1051
rect 1437 -1052 1946 -1000
rect 1998 -1052 2906 -1000
rect 2958 -1052 2972 -1000
rect -478 -1669 -426 -1052
rect 426 -1061 478 -1052
rect 1385 -1062 1437 -1052
rect 1946 -1062 1998 -1052
rect 2906 -1062 2958 -1052
rect 98 -1188 150 -1178
rect -478 -1731 -426 -1721
rect -287 -1303 -235 -1293
rect -592 -1776 -540 -1766
rect -1101 -2450 -1049 -2440
rect -872 -1919 -820 -1909
rect -1241 -2543 -1240 -2491
rect -1188 -2543 -1187 -2491
rect -1241 -2864 -1187 -2543
rect -1098 -2864 -1046 -2855
rect -872 -2864 -820 -1971
rect -592 -2225 -540 -1828
rect -416 -1779 -364 -1769
rect -416 -1919 -364 -1831
rect -416 -1981 -364 -1971
rect -1241 -2865 -1045 -2864
rect -1241 -2917 -1098 -2865
rect -1046 -2917 -1045 -2865
rect -1241 -2918 -1045 -2917
rect -1241 -3485 -1187 -2918
rect -1098 -2927 -1046 -2918
rect -872 -2926 -820 -2916
rect -762 -2388 -710 -2378
rect -762 -2775 -710 -2440
rect -592 -2390 -540 -2277
rect -287 -2261 -235 -1355
rect 98 -1527 150 -1240
rect 425 -1520 477 -1510
rect 98 -1572 425 -1527
rect 517 -1527 583 -1515
rect 1387 -1522 1439 -1512
rect 477 -1572 1387 -1527
rect 98 -1574 1387 -1572
rect 1948 -1522 2000 -1512
rect 1439 -1574 1948 -1527
rect 2908 -1522 2960 -1512
rect 2000 -1574 2908 -1527
rect 98 -1579 2960 -1574
rect 425 -1582 477 -1579
rect 517 -1581 583 -1579
rect 1387 -1584 1439 -1579
rect 1948 -1584 2000 -1579
rect 2908 -1584 2960 -1579
rect 1650 -1757 1702 -1747
rect -235 -2313 148 -2261
rect -287 -2323 -235 -2313
rect 96 -2336 148 -2313
rect 426 -2333 478 -2323
rect 224 -2336 426 -2334
rect -592 -2450 -540 -2442
rect -412 -2385 -360 -2375
rect 96 -2385 426 -2336
rect 1385 -2334 1437 -2324
rect 1650 -2334 1702 -1809
rect 1946 -2334 1998 -2324
rect 2906 -2334 2958 -2324
rect 478 -2385 1385 -2334
rect 96 -2386 1385 -2385
rect 1437 -2386 1946 -2334
rect 1998 -2386 2906 -2334
rect 2958 -2386 2972 -2334
rect 96 -2388 270 -2386
rect 426 -2395 478 -2386
rect 1385 -2396 1437 -2386
rect 1946 -2396 1998 -2386
rect 2906 -2396 2958 -2386
rect -412 -2491 -360 -2437
rect -412 -2553 -360 -2543
rect -762 -3393 -710 -2827
rect -412 -2775 -360 -2765
rect -412 -2866 -360 -2827
rect 425 -2898 477 -2888
rect -412 -2928 -360 -2918
rect -81 -2950 425 -2905
rect 517 -2905 583 -2893
rect 1387 -2900 1439 -2890
rect 477 -2950 1387 -2905
rect -81 -2952 1387 -2950
rect 1948 -2900 2000 -2890
rect 1439 -2952 1948 -2905
rect 2908 -2900 2960 -2890
rect 2000 -2952 2908 -2905
rect -81 -2957 2960 -2952
rect -236 -3026 -184 -3016
rect -762 -3475 -710 -3445
rect -414 -3393 -362 -3383
rect -414 -3474 -362 -3445
rect -414 -3536 -362 -3526
rect -1241 -3549 -1187 -3539
rect -1416 -4346 -1364 -4336
rect -500 -3580 -448 -3570
rect -500 -4555 -448 -3632
rect -236 -3702 -184 -3078
rect -236 -3712 -183 -3702
rect -236 -3764 -235 -3712
rect -236 -3774 -183 -3764
rect -236 -3951 -184 -3774
rect -236 -4013 -184 -4003
rect -81 -4111 -29 -2957
rect 425 -2960 477 -2957
rect 517 -2959 583 -2957
rect 1387 -2962 1439 -2957
rect 1948 -2962 2000 -2957
rect 2908 -2962 2960 -2957
rect 1650 -3135 1702 -3125
rect 140 -3712 192 -3702
rect 426 -3711 478 -3701
rect 192 -3763 426 -3712
rect 1385 -3712 1437 -3702
rect 1650 -3712 1702 -3187
rect 1946 -3712 1998 -3702
rect 2906 -3712 2958 -3702
rect 478 -3763 1385 -3712
rect 192 -3764 1385 -3763
rect 1437 -3764 1946 -3712
rect 1998 -3764 2906 -3712
rect 2958 -3764 2972 -3712
rect 140 -3774 192 -3764
rect 426 -3773 478 -3764
rect 1385 -3774 1437 -3764
rect 1946 -3774 1998 -3764
rect 2906 -3774 2958 -3764
rect -81 -4173 -29 -4163
rect 425 -4276 477 -4266
rect 91 -4328 425 -4283
rect 517 -4283 583 -4271
rect 1387 -4278 1439 -4268
rect 477 -4328 1387 -4283
rect 91 -4330 1387 -4328
rect 1948 -4278 2000 -4268
rect 1439 -4330 1948 -4283
rect 2908 -4278 2960 -4268
rect 2000 -4330 2908 -4283
rect 91 -4335 2960 -4330
rect 91 -4389 144 -4335
rect 425 -4338 477 -4335
rect 517 -4337 583 -4335
rect 1387 -4340 1439 -4335
rect 1948 -4340 2000 -4335
rect 2908 -4340 2960 -4335
rect 92 -4409 144 -4389
rect 92 -4471 144 -4461
rect -548 -4565 -448 -4555
rect -496 -4617 -448 -4565
rect -548 -4627 -448 -4617
rect -2360 -5097 -1535 -5091
rect -2360 -5143 -2358 -5097
rect -2306 -5143 -2163 -5097
rect -2358 -5159 -2306 -5149
rect -2111 -5143 -1535 -5097
rect -500 -5089 -448 -4627
rect 1650 -4513 1702 -4503
rect 426 -5089 478 -5079
rect -500 -5090 245 -5089
rect -500 -5141 426 -5090
rect 1385 -5090 1437 -5080
rect 1650 -5090 1702 -4565
rect 1946 -5090 1998 -5080
rect 2906 -5090 2958 -5080
rect 478 -5141 1385 -5090
rect 224 -5142 1385 -5141
rect 1437 -5142 1946 -5090
rect 1998 -5142 2906 -5090
rect 2958 -5142 2972 -5090
rect -1587 -5148 -1535 -5143
rect -2163 -5159 -2111 -5149
rect 426 -5151 478 -5142
rect 1385 -5152 1437 -5142
rect 1946 -5152 1998 -5142
rect 2906 -5152 2958 -5142
<< labels >>
flabel metal1 3438 -2641 3438 -2641 1 FreeSans 400 0 0 0 out
port 8 n
flabel metal2 -1562 128 -1562 128 1 FreeSans 400 0 0 0 en
port 1 n
flabel metal2 -1216 128 -1216 128 1 FreeSans 400 0 0 0 s1
port 2 n
flabel metal2 -1073 128 -1073 128 1 FreeSans 400 0 0 0 s0
port 3 n
flabel metal1 -3454 -717 -3454 -717 1 FreeSans 400 0 0 0 in0
port 4 n
flabel metal1 -3454 -2051 -3454 -2051 1 FreeSans 400 0 0 0 in1
port 5 n
flabel metal1 -3455 -3430 -3455 -3430 1 FreeSans 400 0 0 0 in2
port 6 n
flabel metal1 -3453 -4807 -3453 -4807 1 FreeSans 400 0 0 0 in3
port 7 n
flabel locali -3783 -5630 -3783 -5630 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel locali -3801 286 -3801 286 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
<< end >>
