magic
tech sky130A
timestamp 1654656593
<< nwell >>
rect -323 -178 324 147
<< pmos >>
rect -223 -68 -208 68
rect -175 -68 -160 68
rect -127 -68 -112 68
rect -79 -68 -64 68
rect -31 -68 -16 68
rect 17 -68 32 68
rect 65 -68 80 68
rect 113 -68 128 68
rect 161 -68 176 68
rect 209 -68 224 68
<< pdiff >>
rect -254 62 -223 68
rect -254 -62 -248 62
rect -231 -62 -223 62
rect -254 -68 -223 -62
rect -208 62 -175 68
rect -208 -62 -200 62
rect -183 -62 -175 62
rect -208 -68 -175 -62
rect -160 62 -127 68
rect -160 -62 -152 62
rect -135 -62 -127 62
rect -160 -68 -127 -62
rect -112 62 -79 68
rect -112 -62 -104 62
rect -87 -62 -79 62
rect -112 -68 -79 -62
rect -64 62 -31 68
rect -64 -62 -56 62
rect -39 -62 -31 62
rect -64 -68 -31 -62
rect -16 62 17 68
rect -16 -62 -8 62
rect 9 -62 17 62
rect -16 -68 17 -62
rect 32 62 65 68
rect 32 -62 40 62
rect 57 -62 65 62
rect 32 -68 65 -62
rect 80 62 113 68
rect 80 -62 88 62
rect 105 -62 113 62
rect 80 -68 113 -62
rect 128 62 161 68
rect 128 -62 136 62
rect 153 -62 161 62
rect 128 -68 161 -62
rect 176 62 209 68
rect 176 -62 184 62
rect 201 -62 209 62
rect 176 -68 209 -62
rect 224 62 255 68
rect 224 -62 232 62
rect 249 -62 255 62
rect 224 -68 255 -62
<< pdiffc >>
rect -248 -62 -231 62
rect -200 -62 -183 62
rect -152 -62 -135 62
rect -104 -62 -87 62
rect -56 -62 -39 62
rect -8 -62 9 62
rect 40 -62 57 62
rect 88 -62 105 62
rect 136 -62 153 62
rect 184 -62 201 62
rect 232 -62 249 62
<< nsubdiff >>
rect -305 112 -257 129
rect 258 112 306 129
rect -305 81 -288 112
rect 289 81 306 112
rect -305 -143 -288 -112
rect 289 -143 306 -112
rect -305 -160 -257 -143
rect 258 -160 306 -143
<< nsubdiffcont >>
rect -257 112 258 129
rect -305 -112 -288 81
rect 289 -112 306 81
rect -257 -160 258 -143
<< poly >>
rect -223 68 -208 81
rect -175 68 -160 81
rect -127 68 -112 81
rect -79 68 -64 81
rect -31 68 -16 81
rect 17 68 32 81
rect 65 68 80 81
rect 113 68 128 81
rect 161 68 176 81
rect 209 68 224 81
rect -223 -84 -208 -68
rect -175 -84 -160 -68
rect -127 -84 -112 -68
rect -79 -84 -64 -68
rect -31 -84 -16 -68
rect 17 -84 32 -68
rect 65 -84 80 -68
rect 113 -84 128 -68
rect 161 -84 176 -68
rect 209 -84 224 -68
rect -256 -92 257 -84
rect -256 -109 -248 -92
rect -231 -109 -152 -92
rect -135 -109 -56 -92
rect -39 -109 40 -92
rect 57 -109 136 -92
rect 153 -109 232 -92
rect 249 -109 257 -92
rect -256 -117 257 -109
<< polycont >>
rect -248 -109 -231 -92
rect -152 -109 -135 -92
rect -56 -109 -39 -92
rect 40 -109 57 -92
rect 136 -109 153 -92
rect 232 -109 249 -92
<< locali >>
rect -305 112 -257 129
rect 258 112 306 129
rect -305 81 -288 112
rect 289 81 306 112
rect -248 62 -231 70
rect -248 -70 -231 -62
rect -200 62 -183 70
rect -200 -70 -183 -62
rect -152 62 -135 70
rect -152 -70 -135 -62
rect -104 62 -87 70
rect -104 -70 -87 -62
rect -56 62 -39 70
rect -56 -70 -39 -62
rect -8 62 9 70
rect -8 -70 9 -62
rect 40 62 57 70
rect 40 -70 57 -62
rect 88 62 105 70
rect 88 -70 105 -62
rect 136 62 153 70
rect 136 -70 153 -62
rect 184 62 201 70
rect 184 -70 201 -62
rect 232 62 249 70
rect 232 -70 249 -62
rect -305 -143 -288 -112
rect -256 -92 257 -88
rect -256 -109 -248 -92
rect -231 -109 -152 -92
rect -135 -109 -56 -92
rect -39 -109 40 -92
rect 57 -109 136 -92
rect 153 -109 232 -92
rect 249 -109 257 -92
rect -256 -113 257 -109
rect 289 -143 306 -112
rect -305 -160 -257 -143
rect 258 -160 306 -143
<< viali >>
rect -248 -62 -231 62
rect -200 -62 -183 62
rect -152 -62 -135 62
rect -104 -62 -87 62
rect -56 -62 -39 62
rect -8 -62 9 62
rect 40 -62 57 62
rect 88 -62 105 62
rect 136 -62 153 62
rect 184 -62 201 62
rect 232 -62 249 62
<< metal1 >>
rect -251 62 -228 68
rect -251 -62 -248 62
rect -231 -62 -228 62
rect -251 -68 -228 -62
rect -203 62 -180 68
rect -203 -62 -200 62
rect -183 -62 -180 62
rect -203 -68 -180 -62
rect -155 62 -132 68
rect -155 -62 -152 62
rect -135 -62 -132 62
rect -155 -68 -132 -62
rect -107 62 -84 68
rect -107 -62 -104 62
rect -87 -62 -84 62
rect -107 -68 -84 -62
rect -59 62 -36 68
rect -59 -62 -56 62
rect -39 -62 -36 62
rect -59 -68 -36 -62
rect -11 62 12 68
rect -11 -62 -8 62
rect 9 -62 12 62
rect -11 -68 12 -62
rect 37 62 60 68
rect 37 -62 40 62
rect 57 -62 60 62
rect 37 -68 60 -62
rect 85 62 108 68
rect 85 -62 88 62
rect 105 -62 108 62
rect 85 -68 108 -62
rect 133 62 156 68
rect 133 -62 136 62
rect 153 -62 156 62
rect 133 -68 156 -62
rect 181 62 204 68
rect 181 -62 184 62
rect 201 -62 204 62
rect 181 -68 204 -62
rect 229 62 252 68
rect 229 -62 232 62
rect 249 -62 252 62
rect 229 -68 252 -62
<< properties >>
string FIXED_BBOX -297 -151 297 151
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.37 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
