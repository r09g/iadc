magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< pwell >>
rect -1020 -166 1020 166
<< nmos >>
rect -936 -140 -816 140
rect -644 -140 -524 140
rect -352 -140 -232 140
rect -60 -140 60 140
rect 232 -140 352 140
rect 524 -140 644 140
rect 816 -140 936 140
<< ndiff >>
rect -994 119 -936 140
rect -994 85 -982 119
rect -948 85 -936 119
rect -994 51 -936 85
rect -994 17 -982 51
rect -948 17 -936 51
rect -994 -17 -936 17
rect -994 -51 -982 -17
rect -948 -51 -936 -17
rect -994 -85 -936 -51
rect -994 -119 -982 -85
rect -948 -119 -936 -85
rect -994 -140 -936 -119
rect -816 119 -758 140
rect -816 85 -804 119
rect -770 85 -758 119
rect -816 51 -758 85
rect -816 17 -804 51
rect -770 17 -758 51
rect -816 -17 -758 17
rect -816 -51 -804 -17
rect -770 -51 -758 -17
rect -816 -85 -758 -51
rect -816 -119 -804 -85
rect -770 -119 -758 -85
rect -816 -140 -758 -119
rect -702 119 -644 140
rect -702 85 -690 119
rect -656 85 -644 119
rect -702 51 -644 85
rect -702 17 -690 51
rect -656 17 -644 51
rect -702 -17 -644 17
rect -702 -51 -690 -17
rect -656 -51 -644 -17
rect -702 -85 -644 -51
rect -702 -119 -690 -85
rect -656 -119 -644 -85
rect -702 -140 -644 -119
rect -524 119 -466 140
rect -524 85 -512 119
rect -478 85 -466 119
rect -524 51 -466 85
rect -524 17 -512 51
rect -478 17 -466 51
rect -524 -17 -466 17
rect -524 -51 -512 -17
rect -478 -51 -466 -17
rect -524 -85 -466 -51
rect -524 -119 -512 -85
rect -478 -119 -466 -85
rect -524 -140 -466 -119
rect -410 119 -352 140
rect -410 85 -398 119
rect -364 85 -352 119
rect -410 51 -352 85
rect -410 17 -398 51
rect -364 17 -352 51
rect -410 -17 -352 17
rect -410 -51 -398 -17
rect -364 -51 -352 -17
rect -410 -85 -352 -51
rect -410 -119 -398 -85
rect -364 -119 -352 -85
rect -410 -140 -352 -119
rect -232 119 -174 140
rect -232 85 -220 119
rect -186 85 -174 119
rect -232 51 -174 85
rect -232 17 -220 51
rect -186 17 -174 51
rect -232 -17 -174 17
rect -232 -51 -220 -17
rect -186 -51 -174 -17
rect -232 -85 -174 -51
rect -232 -119 -220 -85
rect -186 -119 -174 -85
rect -232 -140 -174 -119
rect -118 119 -60 140
rect -118 85 -106 119
rect -72 85 -60 119
rect -118 51 -60 85
rect -118 17 -106 51
rect -72 17 -60 51
rect -118 -17 -60 17
rect -118 -51 -106 -17
rect -72 -51 -60 -17
rect -118 -85 -60 -51
rect -118 -119 -106 -85
rect -72 -119 -60 -85
rect -118 -140 -60 -119
rect 60 119 118 140
rect 60 85 72 119
rect 106 85 118 119
rect 60 51 118 85
rect 60 17 72 51
rect 106 17 118 51
rect 60 -17 118 17
rect 60 -51 72 -17
rect 106 -51 118 -17
rect 60 -85 118 -51
rect 60 -119 72 -85
rect 106 -119 118 -85
rect 60 -140 118 -119
rect 174 119 232 140
rect 174 85 186 119
rect 220 85 232 119
rect 174 51 232 85
rect 174 17 186 51
rect 220 17 232 51
rect 174 -17 232 17
rect 174 -51 186 -17
rect 220 -51 232 -17
rect 174 -85 232 -51
rect 174 -119 186 -85
rect 220 -119 232 -85
rect 174 -140 232 -119
rect 352 119 410 140
rect 352 85 364 119
rect 398 85 410 119
rect 352 51 410 85
rect 352 17 364 51
rect 398 17 410 51
rect 352 -17 410 17
rect 352 -51 364 -17
rect 398 -51 410 -17
rect 352 -85 410 -51
rect 352 -119 364 -85
rect 398 -119 410 -85
rect 352 -140 410 -119
rect 466 119 524 140
rect 466 85 478 119
rect 512 85 524 119
rect 466 51 524 85
rect 466 17 478 51
rect 512 17 524 51
rect 466 -17 524 17
rect 466 -51 478 -17
rect 512 -51 524 -17
rect 466 -85 524 -51
rect 466 -119 478 -85
rect 512 -119 524 -85
rect 466 -140 524 -119
rect 644 119 702 140
rect 644 85 656 119
rect 690 85 702 119
rect 644 51 702 85
rect 644 17 656 51
rect 690 17 702 51
rect 644 -17 702 17
rect 644 -51 656 -17
rect 690 -51 702 -17
rect 644 -85 702 -51
rect 644 -119 656 -85
rect 690 -119 702 -85
rect 644 -140 702 -119
rect 758 119 816 140
rect 758 85 770 119
rect 804 85 816 119
rect 758 51 816 85
rect 758 17 770 51
rect 804 17 816 51
rect 758 -17 816 17
rect 758 -51 770 -17
rect 804 -51 816 -17
rect 758 -85 816 -51
rect 758 -119 770 -85
rect 804 -119 816 -85
rect 758 -140 816 -119
rect 936 119 994 140
rect 936 85 948 119
rect 982 85 994 119
rect 936 51 994 85
rect 936 17 948 51
rect 982 17 994 51
rect 936 -17 994 17
rect 936 -51 948 -17
rect 982 -51 994 -17
rect 936 -85 994 -51
rect 936 -119 948 -85
rect 982 -119 994 -85
rect 936 -140 994 -119
<< ndiffc >>
rect -982 85 -948 119
rect -982 17 -948 51
rect -982 -51 -948 -17
rect -982 -119 -948 -85
rect -804 85 -770 119
rect -804 17 -770 51
rect -804 -51 -770 -17
rect -804 -119 -770 -85
rect -690 85 -656 119
rect -690 17 -656 51
rect -690 -51 -656 -17
rect -690 -119 -656 -85
rect -512 85 -478 119
rect -512 17 -478 51
rect -512 -51 -478 -17
rect -512 -119 -478 -85
rect -398 85 -364 119
rect -398 17 -364 51
rect -398 -51 -364 -17
rect -398 -119 -364 -85
rect -220 85 -186 119
rect -220 17 -186 51
rect -220 -51 -186 -17
rect -220 -119 -186 -85
rect -106 85 -72 119
rect -106 17 -72 51
rect -106 -51 -72 -17
rect -106 -119 -72 -85
rect 72 85 106 119
rect 72 17 106 51
rect 72 -51 106 -17
rect 72 -119 106 -85
rect 186 85 220 119
rect 186 17 220 51
rect 186 -51 220 -17
rect 186 -119 220 -85
rect 364 85 398 119
rect 364 17 398 51
rect 364 -51 398 -17
rect 364 -119 398 -85
rect 478 85 512 119
rect 478 17 512 51
rect 478 -51 512 -17
rect 478 -119 512 -85
rect 656 85 690 119
rect 656 17 690 51
rect 656 -51 690 -17
rect 656 -119 690 -85
rect 770 85 804 119
rect 770 17 804 51
rect 770 -51 804 -17
rect 770 -119 804 -85
rect 948 85 982 119
rect 948 17 982 51
rect 948 -51 982 -17
rect 948 -119 982 -85
<< poly >>
rect -914 212 -838 228
rect -914 194 -893 212
rect -936 178 -893 194
rect -859 194 -838 212
rect -622 212 -546 228
rect -622 194 -601 212
rect -859 178 -816 194
rect -936 140 -816 178
rect -644 178 -601 194
rect -567 194 -546 212
rect -330 212 -254 228
rect -330 194 -309 212
rect -567 178 -524 194
rect -644 140 -524 178
rect -352 178 -309 194
rect -275 194 -254 212
rect -38 212 38 228
rect -38 194 -17 212
rect -275 178 -232 194
rect -352 140 -232 178
rect -60 178 -17 194
rect 17 194 38 212
rect 254 212 330 228
rect 254 194 275 212
rect 17 178 60 194
rect -60 140 60 178
rect 232 178 275 194
rect 309 194 330 212
rect 546 212 622 228
rect 546 194 567 212
rect 309 178 352 194
rect 232 140 352 178
rect 524 178 567 194
rect 601 194 622 212
rect 838 212 914 228
rect 838 194 859 212
rect 601 178 644 194
rect 524 140 644 178
rect 816 178 859 194
rect 893 194 914 212
rect 893 178 936 194
rect 816 140 936 178
rect -936 -178 -816 -140
rect -936 -194 -893 -178
rect -914 -212 -893 -194
rect -859 -194 -816 -178
rect -644 -178 -524 -140
rect -644 -194 -601 -178
rect -859 -212 -838 -194
rect -914 -228 -838 -212
rect -622 -212 -601 -194
rect -567 -194 -524 -178
rect -352 -178 -232 -140
rect -352 -194 -309 -178
rect -567 -212 -546 -194
rect -622 -228 -546 -212
rect -330 -212 -309 -194
rect -275 -194 -232 -178
rect -60 -178 60 -140
rect -60 -194 -17 -178
rect -275 -212 -254 -194
rect -330 -228 -254 -212
rect -38 -212 -17 -194
rect 17 -194 60 -178
rect 232 -178 352 -140
rect 232 -194 275 -178
rect 17 -212 38 -194
rect -38 -228 38 -212
rect 254 -212 275 -194
rect 309 -194 352 -178
rect 524 -178 644 -140
rect 524 -194 567 -178
rect 309 -212 330 -194
rect 254 -228 330 -212
rect 546 -212 567 -194
rect 601 -194 644 -178
rect 816 -178 936 -140
rect 816 -194 859 -178
rect 601 -212 622 -194
rect 546 -228 622 -212
rect 838 -212 859 -194
rect 893 -194 936 -178
rect 893 -212 914 -194
rect 838 -228 914 -212
<< polycont >>
rect -893 178 -859 212
rect -601 178 -567 212
rect -309 178 -275 212
rect -17 178 17 212
rect 275 178 309 212
rect 567 178 601 212
rect 859 178 893 212
rect -893 -212 -859 -178
rect -601 -212 -567 -178
rect -309 -212 -275 -178
rect -17 -212 17 -178
rect 275 -212 309 -178
rect 567 -212 601 -178
rect 859 -212 893 -178
<< locali >>
rect -914 178 -893 212
rect -859 178 -838 212
rect -622 178 -601 212
rect -567 178 -546 212
rect -330 178 -309 212
rect -275 178 -254 212
rect -38 178 -17 212
rect 17 178 38 212
rect 254 178 275 212
rect 309 178 330 212
rect 546 178 567 212
rect 601 178 622 212
rect 838 178 859 212
rect 893 178 914 212
rect -982 125 -948 144
rect -982 53 -948 85
rect -982 -17 -948 17
rect -982 -85 -948 -53
rect -982 -144 -948 -125
rect -804 125 -770 144
rect -804 53 -770 85
rect -804 -17 -770 17
rect -804 -85 -770 -53
rect -804 -144 -770 -125
rect -690 125 -656 144
rect -690 53 -656 85
rect -690 -17 -656 17
rect -690 -85 -656 -53
rect -690 -144 -656 -125
rect -512 125 -478 144
rect -512 53 -478 85
rect -512 -17 -478 17
rect -512 -85 -478 -53
rect -512 -144 -478 -125
rect -398 125 -364 144
rect -398 53 -364 85
rect -398 -17 -364 17
rect -398 -85 -364 -53
rect -398 -144 -364 -125
rect -220 125 -186 144
rect -220 53 -186 85
rect -220 -17 -186 17
rect -220 -85 -186 -53
rect -220 -144 -186 -125
rect -106 125 -72 144
rect -106 53 -72 85
rect -106 -17 -72 17
rect -106 -85 -72 -53
rect -106 -144 -72 -125
rect 72 125 106 144
rect 72 53 106 85
rect 72 -17 106 17
rect 72 -85 106 -53
rect 72 -144 106 -125
rect 186 125 220 144
rect 186 53 220 85
rect 186 -17 220 17
rect 186 -85 220 -53
rect 186 -144 220 -125
rect 364 125 398 144
rect 364 53 398 85
rect 364 -17 398 17
rect 364 -85 398 -53
rect 364 -144 398 -125
rect 478 125 512 144
rect 478 53 512 85
rect 478 -17 512 17
rect 478 -85 512 -53
rect 478 -144 512 -125
rect 656 125 690 144
rect 656 53 690 85
rect 656 -17 690 17
rect 656 -85 690 -53
rect 656 -144 690 -125
rect 770 125 804 144
rect 770 53 804 85
rect 770 -17 804 17
rect 770 -85 804 -53
rect 770 -144 804 -125
rect 948 125 982 144
rect 948 53 982 85
rect 948 -17 982 17
rect 948 -85 982 -53
rect 948 -144 982 -125
rect -914 -212 -893 -178
rect -859 -212 -838 -178
rect -622 -212 -601 -178
rect -567 -212 -546 -178
rect -330 -212 -309 -178
rect -275 -212 -254 -178
rect -38 -212 -17 -178
rect 17 -212 38 -178
rect 254 -212 275 -178
rect 309 -212 330 -178
rect 546 -212 567 -178
rect 601 -212 622 -178
rect 838 -212 859 -178
rect 893 -212 914 -178
<< viali >>
rect -893 178 -859 212
rect -601 178 -567 212
rect -309 178 -275 212
rect -17 178 17 212
rect 275 178 309 212
rect 567 178 601 212
rect 859 178 893 212
rect -982 119 -948 125
rect -982 91 -948 119
rect -982 51 -948 53
rect -982 19 -948 51
rect -982 -51 -948 -19
rect -982 -53 -948 -51
rect -982 -119 -948 -91
rect -982 -125 -948 -119
rect -804 119 -770 125
rect -804 91 -770 119
rect -804 51 -770 53
rect -804 19 -770 51
rect -804 -51 -770 -19
rect -804 -53 -770 -51
rect -804 -119 -770 -91
rect -804 -125 -770 -119
rect -690 119 -656 125
rect -690 91 -656 119
rect -690 51 -656 53
rect -690 19 -656 51
rect -690 -51 -656 -19
rect -690 -53 -656 -51
rect -690 -119 -656 -91
rect -690 -125 -656 -119
rect -512 119 -478 125
rect -512 91 -478 119
rect -512 51 -478 53
rect -512 19 -478 51
rect -512 -51 -478 -19
rect -512 -53 -478 -51
rect -512 -119 -478 -91
rect -512 -125 -478 -119
rect -398 119 -364 125
rect -398 91 -364 119
rect -398 51 -364 53
rect -398 19 -364 51
rect -398 -51 -364 -19
rect -398 -53 -364 -51
rect -398 -119 -364 -91
rect -398 -125 -364 -119
rect -220 119 -186 125
rect -220 91 -186 119
rect -220 51 -186 53
rect -220 19 -186 51
rect -220 -51 -186 -19
rect -220 -53 -186 -51
rect -220 -119 -186 -91
rect -220 -125 -186 -119
rect -106 119 -72 125
rect -106 91 -72 119
rect -106 51 -72 53
rect -106 19 -72 51
rect -106 -51 -72 -19
rect -106 -53 -72 -51
rect -106 -119 -72 -91
rect -106 -125 -72 -119
rect 72 119 106 125
rect 72 91 106 119
rect 72 51 106 53
rect 72 19 106 51
rect 72 -51 106 -19
rect 72 -53 106 -51
rect 72 -119 106 -91
rect 72 -125 106 -119
rect 186 119 220 125
rect 186 91 220 119
rect 186 51 220 53
rect 186 19 220 51
rect 186 -51 220 -19
rect 186 -53 220 -51
rect 186 -119 220 -91
rect 186 -125 220 -119
rect 364 119 398 125
rect 364 91 398 119
rect 364 51 398 53
rect 364 19 398 51
rect 364 -51 398 -19
rect 364 -53 398 -51
rect 364 -119 398 -91
rect 364 -125 398 -119
rect 478 119 512 125
rect 478 91 512 119
rect 478 51 512 53
rect 478 19 512 51
rect 478 -51 512 -19
rect 478 -53 512 -51
rect 478 -119 512 -91
rect 478 -125 512 -119
rect 656 119 690 125
rect 656 91 690 119
rect 656 51 690 53
rect 656 19 690 51
rect 656 -51 690 -19
rect 656 -53 690 -51
rect 656 -119 690 -91
rect 656 -125 690 -119
rect 770 119 804 125
rect 770 91 804 119
rect 770 51 804 53
rect 770 19 804 51
rect 770 -51 804 -19
rect 770 -53 804 -51
rect 770 -119 804 -91
rect 770 -125 804 -119
rect 948 119 982 125
rect 948 91 982 119
rect 948 51 982 53
rect 948 19 982 51
rect 948 -51 982 -19
rect 948 -53 982 -51
rect 948 -119 982 -91
rect 948 -125 982 -119
rect -893 -212 -859 -178
rect -601 -212 -567 -178
rect -309 -212 -275 -178
rect -17 -212 17 -178
rect 275 -212 309 -178
rect 567 -212 601 -178
rect 859 -212 893 -178
<< metal1 >>
rect -914 212 -838 228
rect -914 178 -893 212
rect -859 178 -838 212
rect -914 172 -838 178
rect -622 212 -546 228
rect -622 178 -601 212
rect -567 178 -546 212
rect -622 172 -546 178
rect -330 212 -254 228
rect -330 178 -309 212
rect -275 178 -254 212
rect -330 172 -254 178
rect -38 212 38 228
rect -38 178 -17 212
rect 17 178 38 212
rect -38 172 38 178
rect 254 212 330 228
rect 254 178 275 212
rect 309 178 330 212
rect 254 172 330 178
rect 546 212 622 228
rect 546 178 567 212
rect 601 178 622 212
rect 546 172 622 178
rect 838 212 914 228
rect 838 178 859 212
rect 893 178 914 212
rect 838 172 914 178
rect -988 125 -942 140
rect -988 91 -982 125
rect -948 91 -942 125
rect -988 53 -942 91
rect -988 19 -982 53
rect -948 19 -942 53
rect -988 -19 -942 19
rect -988 -53 -982 -19
rect -948 -53 -942 -19
rect -988 -91 -942 -53
rect -988 -125 -982 -91
rect -948 -125 -942 -91
rect -988 -140 -942 -125
rect -810 125 -764 140
rect -810 91 -804 125
rect -770 91 -764 125
rect -810 53 -764 91
rect -810 19 -804 53
rect -770 19 -764 53
rect -810 -19 -764 19
rect -810 -53 -804 -19
rect -770 -53 -764 -19
rect -810 -91 -764 -53
rect -810 -125 -804 -91
rect -770 -125 -764 -91
rect -810 -140 -764 -125
rect -696 125 -650 140
rect -696 91 -690 125
rect -656 91 -650 125
rect -696 53 -650 91
rect -696 19 -690 53
rect -656 19 -650 53
rect -696 -19 -650 19
rect -696 -53 -690 -19
rect -656 -53 -650 -19
rect -696 -91 -650 -53
rect -696 -125 -690 -91
rect -656 -125 -650 -91
rect -696 -140 -650 -125
rect -518 125 -472 140
rect -518 91 -512 125
rect -478 91 -472 125
rect -518 53 -472 91
rect -518 19 -512 53
rect -478 19 -472 53
rect -518 -19 -472 19
rect -518 -53 -512 -19
rect -478 -53 -472 -19
rect -518 -91 -472 -53
rect -518 -125 -512 -91
rect -478 -125 -472 -91
rect -518 -140 -472 -125
rect -404 125 -358 140
rect -404 91 -398 125
rect -364 91 -358 125
rect -404 53 -358 91
rect -404 19 -398 53
rect -364 19 -358 53
rect -404 -19 -358 19
rect -404 -53 -398 -19
rect -364 -53 -358 -19
rect -404 -91 -358 -53
rect -404 -125 -398 -91
rect -364 -125 -358 -91
rect -404 -140 -358 -125
rect -226 125 -180 140
rect -226 91 -220 125
rect -186 91 -180 125
rect -226 53 -180 91
rect -226 19 -220 53
rect -186 19 -180 53
rect -226 -19 -180 19
rect -226 -53 -220 -19
rect -186 -53 -180 -19
rect -226 -91 -180 -53
rect -226 -125 -220 -91
rect -186 -125 -180 -91
rect -226 -140 -180 -125
rect -112 125 -66 140
rect -112 91 -106 125
rect -72 91 -66 125
rect -112 53 -66 91
rect -112 19 -106 53
rect -72 19 -66 53
rect -112 -19 -66 19
rect -112 -53 -106 -19
rect -72 -53 -66 -19
rect -112 -91 -66 -53
rect -112 -125 -106 -91
rect -72 -125 -66 -91
rect -112 -140 -66 -125
rect 66 125 112 140
rect 66 91 72 125
rect 106 91 112 125
rect 66 53 112 91
rect 66 19 72 53
rect 106 19 112 53
rect 66 -19 112 19
rect 66 -53 72 -19
rect 106 -53 112 -19
rect 66 -91 112 -53
rect 66 -125 72 -91
rect 106 -125 112 -91
rect 66 -140 112 -125
rect 180 125 226 140
rect 180 91 186 125
rect 220 91 226 125
rect 180 53 226 91
rect 180 19 186 53
rect 220 19 226 53
rect 180 -19 226 19
rect 180 -53 186 -19
rect 220 -53 226 -19
rect 180 -91 226 -53
rect 180 -125 186 -91
rect 220 -125 226 -91
rect 180 -140 226 -125
rect 358 125 404 140
rect 358 91 364 125
rect 398 91 404 125
rect 358 53 404 91
rect 358 19 364 53
rect 398 19 404 53
rect 358 -19 404 19
rect 358 -53 364 -19
rect 398 -53 404 -19
rect 358 -91 404 -53
rect 358 -125 364 -91
rect 398 -125 404 -91
rect 358 -140 404 -125
rect 472 125 518 140
rect 472 91 478 125
rect 512 91 518 125
rect 472 53 518 91
rect 472 19 478 53
rect 512 19 518 53
rect 472 -19 518 19
rect 472 -53 478 -19
rect 512 -53 518 -19
rect 472 -91 518 -53
rect 472 -125 478 -91
rect 512 -125 518 -91
rect 472 -140 518 -125
rect 650 125 696 140
rect 650 91 656 125
rect 690 91 696 125
rect 650 53 696 91
rect 650 19 656 53
rect 690 19 696 53
rect 650 -19 696 19
rect 650 -53 656 -19
rect 690 -53 696 -19
rect 650 -91 696 -53
rect 650 -125 656 -91
rect 690 -125 696 -91
rect 650 -140 696 -125
rect 764 125 810 140
rect 764 91 770 125
rect 804 91 810 125
rect 764 53 810 91
rect 764 19 770 53
rect 804 19 810 53
rect 764 -19 810 19
rect 764 -53 770 -19
rect 804 -53 810 -19
rect 764 -91 810 -53
rect 764 -125 770 -91
rect 804 -125 810 -91
rect 764 -140 810 -125
rect 942 125 988 140
rect 942 91 948 125
rect 982 91 988 125
rect 942 53 988 91
rect 942 19 948 53
rect 982 19 988 53
rect 942 -19 988 19
rect 942 -53 948 -19
rect 982 -53 988 -19
rect 942 -91 988 -53
rect 942 -125 948 -91
rect 982 -125 988 -91
rect 942 -140 988 -125
rect -914 -178 -838 -172
rect -914 -212 -893 -178
rect -859 -212 -838 -178
rect -914 -228 -838 -212
rect -622 -178 -546 -172
rect -622 -212 -601 -178
rect -567 -212 -546 -178
rect -622 -228 -546 -212
rect -330 -178 -254 -172
rect -330 -212 -309 -178
rect -275 -212 -254 -178
rect -330 -228 -254 -212
rect -38 -178 38 -172
rect -38 -212 -17 -178
rect 17 -212 38 -178
rect -38 -228 38 -212
rect 254 -178 330 -172
rect 254 -212 275 -178
rect 309 -212 330 -178
rect 254 -228 330 -212
rect 546 -178 622 -172
rect 546 -212 567 -178
rect 601 -212 622 -178
rect 546 -228 622 -212
rect 838 -178 914 -172
rect 838 -212 859 -178
rect 893 -212 914 -178
rect 838 -228 914 -212
<< end >>
