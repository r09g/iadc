magic
tech sky130A
timestamp 1654865385
<< nwell >>
rect 81 234 1488 559
<< pwell >>
rect 81 3 1488 234
rect 715 2 843 3
<< nmos >>
rect 181 108 196 160
rect 229 108 244 160
rect 277 108 292 160
rect 325 108 340 160
rect 373 108 388 160
rect 421 108 436 160
rect 469 108 484 160
rect 517 108 532 160
rect 565 108 580 160
rect 613 108 628 160
rect 769 111 784 161
rect 941 108 956 160
rect 989 108 1004 160
rect 1037 108 1052 160
rect 1085 108 1100 160
rect 1133 108 1148 160
rect 1181 108 1196 160
rect 1229 108 1244 160
rect 1277 108 1292 160
rect 1325 108 1340 160
rect 1373 108 1388 160
<< pmos >>
rect 181 313 196 449
rect 229 313 244 449
rect 277 313 292 449
rect 325 313 340 449
rect 373 313 388 449
rect 421 313 436 449
rect 469 313 484 449
rect 517 313 532 449
rect 565 313 580 449
rect 613 313 628 449
rect 941 313 956 449
rect 989 313 1004 449
rect 1037 313 1052 449
rect 1085 313 1100 449
rect 1133 313 1148 449
rect 1181 313 1196 449
rect 1229 313 1244 449
rect 1277 313 1292 449
rect 1325 313 1340 449
rect 1373 313 1388 449
<< ndiff >>
rect 150 154 181 160
rect 150 114 156 154
rect 173 114 181 154
rect 150 108 181 114
rect 196 154 229 160
rect 196 114 204 154
rect 221 114 229 154
rect 196 108 229 114
rect 244 154 277 160
rect 244 114 252 154
rect 269 114 277 154
rect 244 108 277 114
rect 292 154 325 160
rect 292 114 300 154
rect 317 114 325 154
rect 292 108 325 114
rect 340 154 373 160
rect 340 114 348 154
rect 365 114 373 154
rect 340 108 373 114
rect 388 154 421 160
rect 388 114 396 154
rect 413 114 421 154
rect 388 108 421 114
rect 436 154 469 160
rect 436 114 444 154
rect 461 114 469 154
rect 436 108 469 114
rect 484 154 517 160
rect 484 114 492 154
rect 509 114 517 154
rect 484 108 517 114
rect 532 154 565 160
rect 532 114 540 154
rect 557 114 565 154
rect 532 108 565 114
rect 580 154 613 160
rect 580 114 588 154
rect 605 114 613 154
rect 580 108 613 114
rect 628 154 659 160
rect 628 114 636 154
rect 653 114 659 154
rect 628 108 659 114
rect 740 155 769 161
rect 740 117 746 155
rect 763 117 769 155
rect 740 111 769 117
rect 784 155 813 161
rect 784 117 790 155
rect 807 117 813 155
rect 784 111 813 117
rect 910 154 941 160
rect 910 114 916 154
rect 933 114 941 154
rect 910 108 941 114
rect 956 154 989 160
rect 956 114 964 154
rect 981 114 989 154
rect 956 108 989 114
rect 1004 154 1037 160
rect 1004 114 1012 154
rect 1029 114 1037 154
rect 1004 108 1037 114
rect 1052 154 1085 160
rect 1052 114 1060 154
rect 1077 114 1085 154
rect 1052 108 1085 114
rect 1100 154 1133 160
rect 1100 114 1108 154
rect 1125 114 1133 154
rect 1100 108 1133 114
rect 1148 154 1181 160
rect 1148 114 1156 154
rect 1173 114 1181 154
rect 1148 108 1181 114
rect 1196 154 1229 160
rect 1196 114 1204 154
rect 1221 114 1229 154
rect 1196 108 1229 114
rect 1244 154 1277 160
rect 1244 114 1252 154
rect 1269 114 1277 154
rect 1244 108 1277 114
rect 1292 154 1325 160
rect 1292 114 1300 154
rect 1317 114 1325 154
rect 1292 108 1325 114
rect 1340 154 1373 160
rect 1340 114 1348 154
rect 1365 114 1373 154
rect 1340 108 1373 114
rect 1388 154 1419 160
rect 1388 114 1396 154
rect 1413 114 1419 154
rect 1388 108 1419 114
<< pdiff >>
rect 150 443 181 449
rect 150 319 156 443
rect 173 319 181 443
rect 150 313 181 319
rect 196 443 229 449
rect 196 319 204 443
rect 221 319 229 443
rect 196 313 229 319
rect 244 443 277 449
rect 244 319 252 443
rect 269 319 277 443
rect 244 313 277 319
rect 292 443 325 449
rect 292 319 300 443
rect 317 319 325 443
rect 292 313 325 319
rect 340 443 373 449
rect 340 319 348 443
rect 365 319 373 443
rect 340 313 373 319
rect 388 443 421 449
rect 388 319 396 443
rect 413 319 421 443
rect 388 313 421 319
rect 436 443 469 449
rect 436 319 444 443
rect 461 319 469 443
rect 436 313 469 319
rect 484 443 517 449
rect 484 319 492 443
rect 509 319 517 443
rect 484 313 517 319
rect 532 443 565 449
rect 532 319 540 443
rect 557 319 565 443
rect 532 313 565 319
rect 580 443 613 449
rect 580 319 588 443
rect 605 319 613 443
rect 580 313 613 319
rect 628 443 659 449
rect 628 319 636 443
rect 653 319 659 443
rect 628 313 659 319
rect 910 443 941 449
rect 910 319 916 443
rect 933 319 941 443
rect 910 313 941 319
rect 956 443 989 449
rect 956 319 964 443
rect 981 319 989 443
rect 956 313 989 319
rect 1004 443 1037 449
rect 1004 319 1012 443
rect 1029 319 1037 443
rect 1004 313 1037 319
rect 1052 443 1085 449
rect 1052 319 1060 443
rect 1077 319 1085 443
rect 1052 313 1085 319
rect 1100 443 1133 449
rect 1100 319 1108 443
rect 1125 319 1133 443
rect 1100 313 1133 319
rect 1148 443 1181 449
rect 1148 319 1156 443
rect 1173 319 1181 443
rect 1148 313 1181 319
rect 1196 443 1229 449
rect 1196 319 1204 443
rect 1221 319 1229 443
rect 1196 313 1229 319
rect 1244 443 1277 449
rect 1244 319 1252 443
rect 1269 319 1277 443
rect 1244 313 1277 319
rect 1292 443 1325 449
rect 1292 319 1300 443
rect 1317 319 1325 443
rect 1292 313 1325 319
rect 1340 443 1373 449
rect 1340 319 1348 443
rect 1365 319 1373 443
rect 1340 313 1373 319
rect 1388 443 1419 449
rect 1388 319 1396 443
rect 1413 319 1419 443
rect 1388 313 1419 319
<< ndiffc >>
rect 156 114 173 154
rect 204 114 221 154
rect 252 114 269 154
rect 300 114 317 154
rect 348 114 365 154
rect 396 114 413 154
rect 444 114 461 154
rect 492 114 509 154
rect 540 114 557 154
rect 588 114 605 154
rect 636 114 653 154
rect 746 117 763 155
rect 790 117 807 155
rect 916 114 933 154
rect 964 114 981 154
rect 1012 114 1029 154
rect 1060 114 1077 154
rect 1108 114 1125 154
rect 1156 114 1173 154
rect 1204 114 1221 154
rect 1252 114 1269 154
rect 1300 114 1317 154
rect 1348 114 1365 154
rect 1396 114 1413 154
<< pdiffc >>
rect 156 319 173 443
rect 204 319 221 443
rect 252 319 269 443
rect 300 319 317 443
rect 348 319 365 443
rect 396 319 413 443
rect 444 319 461 443
rect 492 319 509 443
rect 540 319 557 443
rect 588 319 605 443
rect 636 319 653 443
rect 916 319 933 443
rect 964 319 981 443
rect 1012 319 1029 443
rect 1060 319 1077 443
rect 1108 319 1125 443
rect 1156 319 1173 443
rect 1204 319 1221 443
rect 1252 319 1269 443
rect 1300 319 1317 443
rect 1348 319 1365 443
rect 1396 319 1413 443
<< psubdiff >>
rect 99 199 147 216
rect 662 199 710 216
rect 99 168 116 199
rect 693 168 710 199
rect 859 199 907 216
rect 1422 199 1470 216
rect 99 38 116 69
rect 859 168 876 199
rect 693 38 710 69
rect 99 21 147 38
rect 662 21 710 38
rect 1453 168 1470 199
rect 859 38 876 69
rect 1453 38 1470 69
rect 859 21 907 38
rect 1422 21 1470 38
<< nsubdiff >>
rect 99 524 147 541
rect 662 524 710 541
rect 99 493 116 524
rect 693 493 710 524
rect 99 269 116 300
rect 693 269 710 300
rect 99 252 147 269
rect 662 252 710 269
rect 859 524 907 541
rect 1422 524 1470 541
rect 859 493 876 524
rect 1453 493 1470 524
rect 859 269 876 300
rect 1453 269 1470 300
rect 859 252 907 269
rect 1422 252 1470 269
<< psubdiffcont >>
rect 147 199 662 216
rect 99 69 116 168
rect 907 199 1422 216
rect 693 69 710 168
rect 147 21 662 38
rect 859 69 876 168
rect 1453 69 1470 168
rect 907 21 1422 38
<< nsubdiffcont >>
rect 147 524 662 541
rect 99 300 116 493
rect 693 300 710 493
rect 147 252 662 269
rect 907 524 1422 541
rect 859 300 876 493
rect 1453 300 1470 493
rect 907 252 1422 269
<< poly >>
rect 148 490 661 498
rect 148 473 156 490
rect 173 473 252 490
rect 269 473 348 490
rect 365 473 444 490
rect 461 473 540 490
rect 557 473 636 490
rect 653 473 661 490
rect 148 465 661 473
rect 181 449 196 465
rect 229 449 244 465
rect 277 449 292 465
rect 325 449 340 465
rect 373 449 388 465
rect 421 449 436 465
rect 469 449 484 465
rect 517 449 532 465
rect 565 449 580 465
rect 613 449 628 465
rect 181 300 196 313
rect 229 300 244 313
rect 277 300 292 313
rect 325 300 340 313
rect 373 300 388 313
rect 421 300 436 313
rect 469 300 484 313
rect 517 300 532 313
rect 565 300 580 313
rect 613 300 628 313
rect 908 490 1421 498
rect 908 473 916 490
rect 933 473 1012 490
rect 1029 473 1108 490
rect 1125 473 1204 490
rect 1221 473 1300 490
rect 1317 473 1396 490
rect 1413 473 1421 490
rect 908 465 1421 473
rect 941 449 956 465
rect 989 449 1004 465
rect 1037 449 1052 465
rect 1085 449 1100 465
rect 1133 449 1148 465
rect 1181 449 1196 465
rect 1229 449 1244 465
rect 1277 449 1292 465
rect 1325 449 1340 465
rect 1373 449 1388 465
rect 941 300 956 313
rect 989 300 1004 313
rect 1037 300 1052 313
rect 1085 300 1100 313
rect 1133 300 1148 313
rect 1181 300 1196 313
rect 1229 300 1244 313
rect 1277 300 1292 313
rect 1325 300 1340 313
rect 1373 300 1388 313
rect 181 160 196 173
rect 229 160 244 173
rect 277 160 292 173
rect 325 160 340 173
rect 373 160 388 173
rect 421 160 436 173
rect 469 160 484 173
rect 517 160 532 173
rect 565 160 580 173
rect 613 160 628 173
rect 760 197 793 205
rect 760 180 768 197
rect 785 180 793 197
rect 760 172 793 180
rect 181 92 196 108
rect 229 92 244 108
rect 277 92 292 108
rect 325 92 340 108
rect 373 92 388 108
rect 421 92 436 108
rect 469 92 484 108
rect 517 92 532 108
rect 565 92 580 108
rect 613 92 628 108
rect 148 84 661 92
rect 148 67 156 84
rect 173 67 252 84
rect 269 67 348 84
rect 365 67 444 84
rect 461 67 540 84
rect 557 67 636 84
rect 653 67 661 84
rect 148 59 661 67
rect 769 161 784 172
rect 769 98 784 111
rect 941 160 956 173
rect 989 160 1004 173
rect 1037 160 1052 173
rect 1085 160 1100 173
rect 1133 160 1148 173
rect 1181 160 1196 173
rect 1229 160 1244 173
rect 1277 160 1292 173
rect 1325 160 1340 173
rect 1373 160 1388 173
rect 941 92 956 108
rect 989 92 1004 108
rect 1037 92 1052 108
rect 1085 92 1100 108
rect 1133 92 1148 108
rect 1181 92 1196 108
rect 1229 92 1244 108
rect 1277 92 1292 108
rect 1325 92 1340 108
rect 1373 92 1388 108
rect 908 84 1421 92
rect 908 67 916 84
rect 933 67 1012 84
rect 1029 67 1108 84
rect 1125 67 1204 84
rect 1221 67 1300 84
rect 1317 67 1396 84
rect 1413 67 1421 84
rect 908 59 1421 67
<< polycont >>
rect 156 473 173 490
rect 252 473 269 490
rect 348 473 365 490
rect 444 473 461 490
rect 540 473 557 490
rect 636 473 653 490
rect 916 473 933 490
rect 1012 473 1029 490
rect 1108 473 1125 490
rect 1204 473 1221 490
rect 1300 473 1317 490
rect 1396 473 1413 490
rect 768 180 785 197
rect 156 67 173 84
rect 252 67 269 84
rect 348 67 365 84
rect 444 67 461 84
rect 540 67 557 84
rect 636 67 653 84
rect 916 67 933 84
rect 1012 67 1029 84
rect 1108 67 1125 84
rect 1204 67 1221 84
rect 1300 67 1317 84
rect 1396 67 1413 84
<< locali >>
rect 99 524 147 541
rect 662 524 907 541
rect 1422 524 1470 541
rect 99 493 116 524
rect 693 507 879 524
rect 148 490 661 494
rect 148 473 156 490
rect 173 473 252 490
rect 269 473 348 490
rect 365 473 444 490
rect 461 473 540 490
rect 557 473 636 490
rect 653 473 661 490
rect 148 469 661 473
rect 693 493 710 507
rect 156 443 173 451
rect 156 311 173 319
rect 204 443 221 451
rect 204 311 221 319
rect 252 443 269 451
rect 252 311 269 319
rect 300 443 317 451
rect 300 311 317 319
rect 348 443 365 451
rect 348 311 365 319
rect 396 443 413 451
rect 396 311 413 319
rect 444 443 461 451
rect 444 311 461 319
rect 492 443 509 451
rect 492 311 509 319
rect 540 443 557 451
rect 540 311 557 319
rect 588 443 605 451
rect 588 311 605 319
rect 636 443 653 451
rect 636 311 653 319
rect 99 269 116 300
rect 693 269 710 300
rect 99 252 147 269
rect 662 252 710 269
rect 859 493 876 507
rect 908 490 1421 494
rect 908 473 916 490
rect 933 473 1012 490
rect 1029 473 1108 490
rect 1125 473 1204 490
rect 1221 473 1300 490
rect 1317 473 1396 490
rect 1413 473 1421 490
rect 908 469 1421 473
rect 1453 493 1470 524
rect 916 443 933 451
rect 916 311 933 319
rect 964 443 981 451
rect 964 311 981 319
rect 1012 443 1029 451
rect 1012 311 1029 319
rect 1060 443 1077 451
rect 1060 311 1077 319
rect 1108 443 1125 451
rect 1108 311 1125 319
rect 1156 443 1173 451
rect 1156 311 1173 319
rect 1204 443 1221 451
rect 1204 311 1221 319
rect 1252 443 1269 451
rect 1252 311 1269 319
rect 1300 443 1317 451
rect 1300 311 1317 319
rect 1348 443 1365 451
rect 1348 311 1365 319
rect 1396 443 1413 451
rect 1396 311 1413 319
rect 859 269 876 300
rect 1453 269 1470 300
rect 859 252 907 269
rect 1422 252 1470 269
rect 99 199 147 216
rect 662 199 710 216
rect 99 168 116 199
rect 693 168 710 199
rect 859 199 907 216
rect 1422 199 1470 216
rect 760 180 768 197
rect 785 180 793 197
rect 156 154 173 162
rect 156 106 173 114
rect 204 154 221 162
rect 204 106 221 114
rect 252 154 269 162
rect 252 106 269 114
rect 300 154 317 162
rect 300 106 317 114
rect 348 154 365 162
rect 348 106 365 114
rect 396 154 413 162
rect 396 106 413 114
rect 444 154 461 162
rect 444 106 461 114
rect 492 154 509 162
rect 492 106 509 114
rect 540 154 557 162
rect 540 106 557 114
rect 588 154 605 162
rect 588 106 605 114
rect 636 154 653 162
rect 636 106 653 114
rect 859 168 876 199
rect 99 38 116 69
rect 148 84 661 88
rect 148 67 156 84
rect 173 67 252 84
rect 269 67 348 84
rect 365 67 444 84
rect 461 67 540 84
rect 557 67 636 84
rect 653 67 661 84
rect 148 63 661 67
rect 746 155 763 163
rect 746 109 763 117
rect 790 155 807 163
rect 790 109 807 117
rect 693 54 710 69
rect 1453 168 1470 199
rect 916 154 933 162
rect 916 106 933 114
rect 964 154 981 162
rect 964 106 981 114
rect 1012 154 1029 162
rect 1012 106 1029 114
rect 1060 154 1077 162
rect 1060 106 1077 114
rect 1108 154 1125 162
rect 1108 106 1125 114
rect 1156 154 1173 162
rect 1156 106 1173 114
rect 1204 154 1221 162
rect 1204 106 1221 114
rect 1252 154 1269 162
rect 1252 106 1269 114
rect 1300 154 1317 162
rect 1300 106 1317 114
rect 1348 154 1365 162
rect 1348 106 1365 114
rect 1396 154 1413 162
rect 1396 106 1413 114
rect 859 54 876 69
rect 908 84 1421 88
rect 908 67 916 84
rect 933 67 1012 84
rect 1029 67 1108 84
rect 1125 67 1204 84
rect 1221 67 1300 84
rect 1317 67 1396 84
rect 1413 67 1421 84
rect 908 63 1421 67
rect 693 38 876 54
rect 1453 38 1470 69
rect 99 21 147 38
rect 662 21 907 38
rect 1422 21 1470 38
rect 684 20 883 21
<< viali >>
rect 156 473 173 490
rect 636 473 653 490
rect 156 319 173 443
rect 204 319 221 443
rect 252 319 269 443
rect 300 319 317 443
rect 348 319 365 443
rect 396 319 413 443
rect 444 319 461 443
rect 492 319 509 443
rect 540 319 557 443
rect 588 319 605 443
rect 636 319 653 443
rect 916 473 933 490
rect 1396 473 1413 490
rect 916 319 933 443
rect 964 319 981 443
rect 1012 319 1029 443
rect 1060 319 1077 443
rect 1108 319 1125 443
rect 1156 319 1173 443
rect 1204 319 1221 443
rect 1252 319 1269 443
rect 1300 319 1317 443
rect 1348 319 1365 443
rect 1396 319 1413 443
rect 768 180 785 197
rect 156 114 173 154
rect 204 114 221 154
rect 252 114 269 154
rect 300 114 317 154
rect 348 114 365 154
rect 396 114 413 154
rect 444 114 461 154
rect 492 114 509 154
rect 540 114 557 154
rect 588 114 605 154
rect 636 114 653 154
rect 693 111 710 161
rect 156 67 173 84
rect 636 67 653 84
rect 746 117 763 155
rect 790 117 807 155
rect 916 114 933 154
rect 964 114 981 154
rect 1012 114 1029 154
rect 1060 114 1077 154
rect 1108 114 1125 154
rect 1156 114 1173 154
rect 1204 114 1221 154
rect 1252 114 1269 154
rect 1300 114 1317 154
rect 1348 114 1365 154
rect 1396 114 1413 154
rect 916 67 933 84
rect 1396 67 1413 84
<< metal1 >>
rect 81 524 605 541
rect 81 246 98 524
rect 146 468 151 494
rect 177 468 182 494
rect 204 449 221 524
rect 300 449 317 524
rect 396 449 413 524
rect 492 449 509 524
rect 588 449 605 524
rect 841 524 1365 541
rect 626 469 631 495
rect 657 469 662 495
rect 153 443 176 449
rect 153 319 156 443
rect 173 319 176 443
rect 153 313 176 319
rect 201 443 224 449
rect 201 319 204 443
rect 221 319 224 443
rect 201 313 224 319
rect 249 443 272 449
rect 249 319 252 443
rect 269 319 272 443
rect 249 313 272 319
rect 297 443 320 449
rect 297 319 300 443
rect 317 319 320 443
rect 297 313 320 319
rect 345 443 368 449
rect 345 319 348 443
rect 365 319 368 443
rect 345 313 368 319
rect 393 443 416 449
rect 393 319 396 443
rect 413 319 416 443
rect 393 313 416 319
rect 441 443 464 449
rect 441 319 444 443
rect 461 319 464 443
rect 441 313 464 319
rect 489 443 512 449
rect 489 319 492 443
rect 509 319 512 443
rect 489 313 512 319
rect 537 443 560 449
rect 537 319 540 443
rect 557 319 560 443
rect 537 313 560 319
rect 585 443 608 449
rect 585 319 588 443
rect 605 319 608 443
rect 585 313 608 319
rect 633 443 656 449
rect 633 319 636 443
rect 653 319 656 443
rect 633 313 656 319
rect 46 220 98 246
rect 81 37 98 220
rect 156 242 173 313
rect 252 242 269 313
rect 348 242 365 313
rect 444 242 461 313
rect 540 242 557 313
rect 636 242 653 313
rect 841 242 858 524
rect 906 469 911 495
rect 937 469 942 495
rect 964 449 981 524
rect 1060 449 1077 524
rect 1156 449 1173 524
rect 1252 449 1269 524
rect 1348 449 1365 524
rect 1386 469 1391 495
rect 1417 469 1422 495
rect 913 443 936 449
rect 913 319 916 443
rect 933 319 936 443
rect 913 313 936 319
rect 961 443 984 449
rect 961 319 964 443
rect 981 319 984 443
rect 961 313 984 319
rect 1009 443 1032 449
rect 1009 319 1012 443
rect 1029 319 1032 443
rect 1009 313 1032 319
rect 1057 443 1080 449
rect 1057 319 1060 443
rect 1077 319 1080 443
rect 1057 313 1080 319
rect 1105 443 1128 449
rect 1105 319 1108 443
rect 1125 319 1128 443
rect 1105 313 1128 319
rect 1153 443 1176 449
rect 1153 319 1156 443
rect 1173 319 1176 443
rect 1153 313 1176 319
rect 1201 443 1224 449
rect 1201 319 1204 443
rect 1221 319 1224 443
rect 1201 313 1224 319
rect 1249 443 1272 449
rect 1249 319 1252 443
rect 1269 319 1272 443
rect 1249 313 1272 319
rect 1297 443 1320 449
rect 1297 319 1300 443
rect 1317 319 1320 443
rect 1297 313 1320 319
rect 1345 443 1368 449
rect 1345 319 1348 443
rect 1365 319 1368 443
rect 1345 313 1368 319
rect 1393 443 1416 449
rect 1393 319 1396 443
rect 1413 319 1416 443
rect 1393 313 1416 319
rect 156 225 858 242
rect 156 160 173 225
rect 252 160 269 225
rect 348 160 365 225
rect 444 160 461 225
rect 540 160 557 225
rect 636 160 653 225
rect 758 180 763 206
rect 789 180 794 206
rect 762 177 791 180
rect 690 161 713 167
rect 841 161 858 225
rect 153 154 176 160
rect 153 114 156 154
rect 173 114 176 154
rect 153 108 176 114
rect 201 154 224 160
rect 201 114 204 154
rect 221 114 224 154
rect 201 108 224 114
rect 249 154 272 160
rect 249 114 252 154
rect 269 114 272 154
rect 249 108 272 114
rect 297 154 320 160
rect 297 114 300 154
rect 317 114 320 154
rect 297 108 320 114
rect 345 154 368 160
rect 345 114 348 154
rect 365 114 368 154
rect 345 108 368 114
rect 393 154 416 160
rect 393 114 396 154
rect 413 114 416 154
rect 393 108 416 114
rect 441 154 464 160
rect 441 114 444 154
rect 461 114 464 154
rect 441 108 464 114
rect 489 154 512 160
rect 489 114 492 154
rect 509 114 512 154
rect 489 108 512 114
rect 537 154 560 160
rect 537 114 540 154
rect 557 114 560 154
rect 537 108 560 114
rect 585 154 608 160
rect 585 114 588 154
rect 605 114 608 154
rect 585 108 608 114
rect 633 154 656 160
rect 633 114 636 154
rect 653 114 656 154
rect 633 108 656 114
rect 690 111 693 161
rect 710 155 766 161
rect 710 117 746 155
rect 763 117 766 155
rect 710 111 766 117
rect 787 155 858 161
rect 916 242 933 313
rect 1012 242 1029 313
rect 1108 242 1125 313
rect 1204 242 1221 313
rect 1300 242 1317 313
rect 1396 242 1413 313
rect 916 225 1471 242
rect 916 160 933 225
rect 1012 160 1029 225
rect 1108 160 1125 225
rect 1204 160 1221 225
rect 1300 160 1317 225
rect 1396 160 1413 225
rect 787 117 790 155
rect 807 117 858 155
rect 787 111 858 117
rect 146 62 151 88
rect 177 62 182 88
rect 204 37 221 108
rect 300 37 317 108
rect 396 37 413 108
rect 492 37 509 108
rect 588 37 605 108
rect 690 105 713 111
rect 627 63 632 89
rect 658 63 663 89
rect 81 20 605 37
rect 841 37 858 111
rect 913 154 936 160
rect 913 114 916 154
rect 933 114 936 154
rect 913 108 936 114
rect 961 154 984 160
rect 961 114 964 154
rect 981 114 984 154
rect 961 108 984 114
rect 1009 154 1032 160
rect 1009 114 1012 154
rect 1029 114 1032 154
rect 1009 108 1032 114
rect 1057 154 1080 160
rect 1057 114 1060 154
rect 1077 114 1080 154
rect 1057 108 1080 114
rect 1105 154 1128 160
rect 1105 114 1108 154
rect 1125 114 1128 154
rect 1105 108 1128 114
rect 1153 154 1176 160
rect 1153 114 1156 154
rect 1173 114 1176 154
rect 1153 108 1176 114
rect 1201 154 1224 160
rect 1201 114 1204 154
rect 1221 114 1224 154
rect 1201 108 1224 114
rect 1249 154 1272 160
rect 1249 114 1252 154
rect 1269 114 1272 154
rect 1249 108 1272 114
rect 1297 154 1320 160
rect 1297 114 1300 154
rect 1317 114 1320 154
rect 1297 108 1320 114
rect 1345 154 1368 160
rect 1345 114 1348 154
rect 1365 114 1368 154
rect 1345 108 1368 114
rect 1393 154 1416 160
rect 1393 114 1396 154
rect 1413 114 1416 154
rect 1393 108 1416 114
rect 907 63 912 89
rect 938 63 943 89
rect 964 37 981 108
rect 1060 37 1077 108
rect 1156 37 1173 108
rect 1252 37 1269 108
rect 1348 37 1365 108
rect 1387 63 1392 89
rect 1418 63 1423 89
rect 841 20 1365 37
<< via1 >>
rect 151 490 177 494
rect 151 473 156 490
rect 156 473 173 490
rect 173 473 177 490
rect 151 468 177 473
rect 631 490 657 495
rect 631 473 636 490
rect 636 473 653 490
rect 653 473 657 490
rect 631 469 657 473
rect 911 490 937 495
rect 911 473 916 490
rect 916 473 933 490
rect 933 473 937 490
rect 911 469 937 473
rect 1391 490 1417 495
rect 1391 473 1396 490
rect 1396 473 1413 490
rect 1413 473 1417 490
rect 1391 469 1417 473
rect 763 197 789 206
rect 763 180 768 197
rect 768 180 785 197
rect 785 180 789 197
rect 151 84 177 88
rect 151 67 156 84
rect 156 67 173 84
rect 173 67 177 84
rect 151 62 177 67
rect 632 84 658 89
rect 632 67 636 84
rect 636 67 653 84
rect 653 67 658 84
rect 632 63 658 67
rect 912 84 938 89
rect 912 67 916 84
rect 916 67 933 84
rect 933 67 938 84
rect 912 63 938 67
rect 1392 84 1418 89
rect 1392 67 1396 84
rect 1396 67 1413 84
rect 1413 67 1418 84
rect 1392 63 1418 67
<< metal2 >>
rect 151 495 177 499
rect 631 495 657 500
rect 911 495 937 500
rect 1391 495 1417 500
rect 50 494 631 495
rect 50 469 151 494
rect 177 469 631 494
rect 657 469 911 495
rect 937 469 1391 495
rect 1417 469 1424 495
rect 151 463 177 468
rect 631 464 657 469
rect 763 206 789 469
rect 911 464 937 469
rect 1391 464 1417 469
rect 763 175 789 180
rect 151 91 177 93
rect 197 91 230 92
rect 632 91 658 94
rect 912 91 938 94
rect 1392 91 1418 94
rect 46 89 1418 91
rect 46 88 632 89
rect 46 65 151 88
rect 177 65 632 88
rect 151 57 177 62
rect 197 59 230 65
rect 658 65 912 89
rect 632 58 658 63
rect 938 65 1392 89
rect 912 58 938 63
rect 1392 58 1418 63
<< labels >>
flabel locali 776 528 776 528 1 FreeSans 200 0 0 0 VDD
port 5 n power bidirectional
flabel locali 776 33 776 33 1 FreeSans 200 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 57 234 57 234 1 FreeSans 200 0 0 0 in
port 1 n
flabel metal2 60 482 60 482 1 FreeSans 200 0 0 0 en_b
port 4 n
flabel metal2 57 79 57 79 1 FreeSans 200 0 0 0 en
port 3 n
flabel metal1 1463 232 1463 232 1 FreeSans 200 0 0 0 out
port 2 n
<< end >>
