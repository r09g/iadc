magic
tech sky130A
magscale 1 2
timestamp 1653696673
<< nwell >>
rect -53 413 1241 1063
<< pwell >>
rect -53 -51 1241 411
<< nmos >>
rect 147 159 177 263
rect 243 159 273 263
rect 339 159 369 263
rect 435 159 465 263
rect 531 159 561 263
rect 627 159 657 263
rect 723 159 753 263
rect 819 159 849 263
rect 915 159 945 263
rect 1011 159 1041 263
<< pmos >>
rect 147 571 177 843
rect 243 571 273 843
rect 339 571 369 843
rect 435 571 465 843
rect 531 571 561 843
rect 627 571 657 843
rect 723 571 753 843
rect 819 571 849 843
rect 915 571 945 843
rect 1011 571 1041 843
<< ndiff >>
rect 85 251 147 263
rect 85 171 97 251
rect 131 171 147 251
rect 85 159 147 171
rect 177 251 243 263
rect 177 171 193 251
rect 227 171 243 251
rect 177 159 243 171
rect 273 251 339 263
rect 273 171 289 251
rect 323 171 339 251
rect 273 159 339 171
rect 369 251 435 263
rect 369 171 385 251
rect 419 171 435 251
rect 369 159 435 171
rect 465 251 531 263
rect 465 171 481 251
rect 515 171 531 251
rect 465 159 531 171
rect 561 251 627 263
rect 561 171 577 251
rect 611 171 627 251
rect 561 159 627 171
rect 657 251 723 263
rect 657 171 673 251
rect 707 171 723 251
rect 657 159 723 171
rect 753 251 819 263
rect 753 171 769 251
rect 803 171 819 251
rect 753 159 819 171
rect 849 251 915 263
rect 849 171 865 251
rect 899 171 915 251
rect 849 159 915 171
rect 945 251 1011 263
rect 945 171 961 251
rect 995 171 1011 251
rect 945 159 1011 171
rect 1041 251 1103 263
rect 1041 171 1057 251
rect 1091 171 1103 251
rect 1041 159 1103 171
<< pdiff >>
rect 85 831 147 843
rect 85 583 97 831
rect 131 583 147 831
rect 85 571 147 583
rect 177 831 243 843
rect 177 583 193 831
rect 227 583 243 831
rect 177 571 243 583
rect 273 831 339 843
rect 273 583 289 831
rect 323 583 339 831
rect 273 571 339 583
rect 369 831 435 843
rect 369 583 385 831
rect 419 583 435 831
rect 369 571 435 583
rect 465 831 531 843
rect 465 583 481 831
rect 515 583 531 831
rect 465 571 531 583
rect 561 831 627 843
rect 561 583 577 831
rect 611 583 627 831
rect 561 571 627 583
rect 657 831 723 843
rect 657 583 673 831
rect 707 583 723 831
rect 657 571 723 583
rect 753 831 819 843
rect 753 583 769 831
rect 803 583 819 831
rect 753 571 819 583
rect 849 831 915 843
rect 849 583 865 831
rect 899 583 915 831
rect 849 571 915 583
rect 945 831 1011 843
rect 945 583 961 831
rect 995 583 1011 831
rect 945 571 1011 583
rect 1041 831 1103 843
rect 1041 583 1057 831
rect 1091 583 1103 831
rect 1041 571 1103 583
<< ndiffc >>
rect 97 171 131 251
rect 193 171 227 251
rect 289 171 323 251
rect 385 171 419 251
rect 481 171 515 251
rect 577 171 611 251
rect 673 171 707 251
rect 769 171 803 251
rect 865 171 899 251
rect 961 171 995 251
rect 1057 171 1091 251
<< pdiffc >>
rect 97 583 131 831
rect 193 583 227 831
rect 289 583 323 831
rect 385 583 419 831
rect 481 583 515 831
rect 577 583 611 831
rect 673 583 707 831
rect 769 583 803 831
rect 865 583 899 831
rect 961 583 995 831
rect 1057 583 1091 831
<< psubdiff >>
rect -17 341 79 375
rect 1109 341 1205 375
rect -17 279 17 341
rect 1171 279 1205 341
rect -17 19 17 81
rect 1171 19 1205 81
rect -17 -15 79 19
rect 1109 -15 1205 19
<< nsubdiff >>
rect -17 993 79 1027
rect 1109 993 1205 1027
rect -17 931 17 993
rect 1171 931 1205 993
rect -17 483 17 545
rect 1171 483 1205 545
rect -17 449 79 483
rect 1109 449 1205 483
<< psubdiffcont >>
rect 79 341 1109 375
rect -17 81 17 279
rect 1171 81 1205 279
rect 79 -15 1109 19
<< nsubdiffcont >>
rect 79 993 1109 1027
rect -17 545 17 931
rect 1171 545 1205 931
rect 79 449 1109 483
<< poly >>
rect 81 925 1107 941
rect 81 891 97 925
rect 131 891 289 925
rect 323 891 481 925
rect 515 891 673 925
rect 707 891 865 925
rect 899 891 1057 925
rect 1091 891 1107 925
rect 81 875 1107 891
rect 147 843 177 875
rect 243 843 273 875
rect 339 843 369 875
rect 435 843 465 875
rect 531 843 561 875
rect 627 843 657 875
rect 723 843 753 875
rect 819 843 849 875
rect 915 843 945 875
rect 1011 843 1041 875
rect 147 545 177 571
rect 243 545 273 571
rect 339 545 369 571
rect 435 545 465 571
rect 531 545 561 571
rect 627 545 657 571
rect 723 545 753 571
rect 819 545 849 571
rect 915 545 945 571
rect 1011 545 1041 571
rect 147 263 177 289
rect 243 263 273 289
rect 339 263 369 289
rect 435 263 465 289
rect 531 263 561 289
rect 627 263 657 289
rect 723 263 753 289
rect 819 263 849 289
rect 915 263 945 289
rect 1011 263 1041 289
rect 147 137 177 159
rect 243 137 273 159
rect 339 137 369 159
rect 435 137 465 159
rect 531 137 561 159
rect 627 137 657 159
rect 723 137 753 159
rect 819 137 849 159
rect 915 137 945 159
rect 1011 137 1041 159
rect 81 117 1107 137
rect 81 83 97 117
rect 131 83 289 117
rect 323 83 481 117
rect 515 83 673 117
rect 707 83 865 117
rect 899 83 1057 117
rect 1091 83 1107 117
rect 81 71 1107 83
<< polycont >>
rect 97 891 131 925
rect 289 891 323 925
rect 481 891 515 925
rect 673 891 707 925
rect 865 891 899 925
rect 1057 891 1091 925
rect 97 83 131 117
rect 289 83 323 117
rect 481 83 515 117
rect 673 83 707 117
rect 865 83 899 117
rect 1057 83 1091 117
<< locali >>
rect -17 993 79 1027
rect 1109 993 1205 1027
rect -17 931 17 993
rect 1171 931 1205 993
rect 81 891 97 925
rect 131 891 147 925
rect 273 891 289 925
rect 323 891 339 925
rect 465 891 481 925
rect 515 891 531 925
rect 657 891 673 925
rect 707 891 723 925
rect 849 891 865 925
rect 899 891 915 925
rect 1041 891 1057 925
rect 1091 891 1107 925
rect 97 831 131 847
rect 97 567 131 583
rect 193 831 227 847
rect 193 567 227 583
rect 289 831 323 847
rect 289 567 323 583
rect 385 831 419 847
rect 385 567 419 583
rect 481 831 515 847
rect 481 567 515 583
rect 577 831 611 847
rect 577 567 611 583
rect 673 831 707 847
rect 673 567 707 583
rect 769 831 803 847
rect 769 567 803 583
rect 865 831 899 847
rect 865 567 899 583
rect 961 831 995 847
rect 961 567 995 583
rect 1057 831 1091 847
rect 1057 567 1091 583
rect -17 483 17 545
rect 1171 483 1205 545
rect -17 449 79 483
rect 1109 449 1205 483
rect -17 341 79 375
rect 1109 341 1205 375
rect -17 279 17 341
rect 1171 281 1205 341
rect 97 251 131 267
rect 97 155 131 171
rect 193 251 227 267
rect 193 155 227 171
rect 289 251 323 267
rect 289 155 323 171
rect 385 251 419 267
rect 385 155 419 171
rect 481 251 515 267
rect 481 155 515 171
rect 577 251 611 267
rect 577 155 611 171
rect 673 251 707 267
rect 673 155 707 171
rect 769 251 803 267
rect 769 155 803 171
rect 865 251 899 267
rect 865 155 899 171
rect 961 251 995 267
rect 961 155 995 171
rect 1057 251 1091 267
rect 1057 155 1091 171
rect 81 83 97 117
rect 131 83 147 117
rect 273 83 289 117
rect 323 83 339 117
rect 465 83 481 117
rect 515 83 531 117
rect 657 83 673 117
rect 707 83 723 117
rect 849 83 865 117
rect 899 83 915 117
rect 1041 83 1057 117
rect 1091 83 1107 117
rect -17 19 17 81
rect 1171 19 1205 81
rect -17 -15 79 19
rect 1109 -15 1205 19
<< viali >>
rect 97 891 131 925
rect 289 891 323 925
rect 481 891 515 925
rect 673 891 707 925
rect 865 891 899 925
rect 1057 891 1091 925
rect 97 583 131 831
rect 193 583 227 831
rect 289 583 323 831
rect 385 583 419 831
rect 481 583 515 831
rect 577 583 611 831
rect 673 583 707 831
rect 769 583 803 831
rect 865 583 899 831
rect 961 583 995 831
rect 1057 583 1091 831
rect 1171 545 1205 931
rect 1171 279 1205 281
rect 97 171 131 251
rect 193 171 227 251
rect 289 171 323 251
rect 385 171 419 251
rect 481 171 515 251
rect 577 171 611 251
rect 673 171 707 251
rect 769 171 803 251
rect 865 171 899 251
rect 961 171 995 251
rect 1057 171 1091 251
rect 97 83 131 117
rect 289 83 323 117
rect 481 83 515 117
rect 673 83 707 117
rect 865 83 899 117
rect 1057 83 1091 117
rect 1171 81 1205 279
<< metal1 >>
rect -87 993 995 1027
rect -216 883 -189 935
rect -137 883 -127 935
rect -87 430 -53 993
rect 78 883 88 935
rect 140 883 150 935
rect 193 843 227 993
rect 271 883 281 935
rect 333 883 343 935
rect 385 843 419 993
rect 462 883 472 935
rect 524 883 534 935
rect 577 843 611 993
rect 654 883 664 935
rect 716 883 726 935
rect 769 843 803 993
rect 846 883 856 935
rect 908 883 918 935
rect 961 843 995 993
rect 1038 883 1048 935
rect 1100 883 1110 935
rect 1165 931 1211 1063
rect 91 831 137 843
rect 91 583 97 831
rect 131 583 137 831
rect 91 571 137 583
rect 187 831 233 843
rect 187 583 193 831
rect 227 583 233 831
rect 187 571 233 583
rect 283 831 329 843
rect 283 583 289 831
rect 323 583 329 831
rect 283 571 329 583
rect 379 831 425 843
rect 379 583 385 831
rect 419 583 425 831
rect 379 571 425 583
rect 475 831 521 843
rect 475 583 481 831
rect 515 583 521 831
rect 475 571 521 583
rect 571 831 617 843
rect 571 583 577 831
rect 611 583 617 831
rect 571 571 617 583
rect 667 831 713 843
rect 667 583 673 831
rect 707 583 713 831
rect 667 571 713 583
rect 763 831 809 843
rect 763 583 769 831
rect 803 583 809 831
rect 763 571 809 583
rect 859 831 905 843
rect 859 583 865 831
rect 899 583 905 831
rect 859 571 905 583
rect 955 831 1001 843
rect 955 583 961 831
rect 995 583 1001 831
rect 955 571 1001 583
rect 1051 831 1097 843
rect 1051 583 1057 831
rect 1091 583 1097 831
rect 1051 571 1097 583
rect -216 396 -53 430
rect -216 76 -189 128
rect -137 76 -127 128
rect -87 19 -53 396
rect 97 430 131 571
rect 289 430 323 571
rect 481 430 515 571
rect 673 430 707 571
rect 865 430 899 571
rect 1057 430 1091 571
rect 1165 545 1171 931
rect 1205 545 1211 931
rect 1165 533 1211 545
rect 97 396 1283 430
rect 97 263 131 396
rect 289 263 323 396
rect 481 263 515 396
rect 673 263 707 396
rect 865 263 899 396
rect 1057 263 1091 396
rect 1165 281 1211 293
rect 91 251 137 263
rect 91 171 97 251
rect 131 171 137 251
rect 91 159 137 171
rect 187 251 233 263
rect 187 171 193 251
rect 227 171 233 251
rect 187 159 233 171
rect 283 251 329 263
rect 283 171 289 251
rect 323 171 329 251
rect 283 159 329 171
rect 379 251 425 263
rect 379 171 385 251
rect 419 171 425 251
rect 379 159 425 171
rect 475 251 521 263
rect 475 171 481 251
rect 515 171 521 251
rect 475 159 521 171
rect 571 251 617 263
rect 571 171 577 251
rect 611 171 617 251
rect 571 159 617 171
rect 667 251 713 263
rect 667 171 673 251
rect 707 171 713 251
rect 667 159 713 171
rect 763 251 809 263
rect 763 171 769 251
rect 803 171 809 251
rect 763 159 809 171
rect 859 251 905 263
rect 859 171 865 251
rect 899 171 905 251
rect 859 159 905 171
rect 955 251 1001 263
rect 955 171 961 251
rect 995 171 1001 251
rect 955 159 1001 171
rect 1051 251 1097 263
rect 1051 171 1057 251
rect 1091 171 1097 251
rect 1051 159 1097 171
rect 81 128 147 131
rect 78 76 88 128
rect 140 76 150 128
rect 81 71 147 76
rect 193 19 227 159
rect 273 128 339 131
rect 269 76 279 128
rect 331 76 341 128
rect 273 71 339 76
rect 385 19 419 159
rect 465 128 531 131
rect 461 76 471 128
rect 523 76 533 128
rect 465 71 531 76
rect 577 19 611 159
rect 657 128 723 131
rect 653 76 663 128
rect 715 76 725 128
rect 657 71 723 76
rect 769 19 803 159
rect 849 127 915 131
rect 846 75 856 127
rect 908 75 918 127
rect 849 71 915 75
rect 961 19 995 159
rect 1041 127 1107 131
rect 1038 75 1048 127
rect 1100 75 1110 127
rect 1165 81 1171 281
rect 1205 81 1211 281
rect 1041 71 1107 75
rect -87 -15 995 19
rect 1165 -51 1211 81
<< via1 >>
rect -189 883 -137 935
rect 88 925 140 935
rect 88 891 97 925
rect 97 891 131 925
rect 131 891 140 925
rect 88 883 140 891
rect 281 925 333 935
rect 281 891 289 925
rect 289 891 323 925
rect 323 891 333 925
rect 281 883 333 891
rect 472 925 524 935
rect 472 891 481 925
rect 481 891 515 925
rect 515 891 524 925
rect 472 883 524 891
rect 664 925 716 935
rect 664 891 673 925
rect 673 891 707 925
rect 707 891 716 925
rect 664 883 716 891
rect 856 925 908 935
rect 856 891 865 925
rect 865 891 899 925
rect 899 891 908 925
rect 856 883 908 891
rect 1048 925 1100 935
rect 1048 891 1057 925
rect 1057 891 1091 925
rect 1091 891 1100 925
rect 1048 883 1100 891
rect -189 76 -137 128
rect 88 117 140 128
rect 88 83 97 117
rect 97 83 131 117
rect 131 83 140 117
rect 88 76 140 83
rect 279 117 331 128
rect 279 83 289 117
rect 289 83 323 117
rect 323 83 331 117
rect 279 76 331 83
rect 471 117 523 128
rect 471 83 481 117
rect 481 83 515 117
rect 515 83 523 117
rect 471 76 523 83
rect 663 117 715 128
rect 663 83 673 117
rect 673 83 707 117
rect 707 83 715 117
rect 663 76 715 83
rect 856 117 908 127
rect 856 83 865 117
rect 865 83 899 117
rect 899 83 908 117
rect 856 75 908 83
rect 1048 117 1100 127
rect 1048 83 1057 117
rect 1057 83 1091 117
rect 1091 83 1100 117
rect 1048 75 1100 83
<< metal2 >>
rect -189 935 -137 945
rect 88 935 140 945
rect 281 935 333 945
rect 472 935 524 945
rect 664 935 716 945
rect 856 935 908 945
rect 1048 935 1100 945
rect -137 883 88 935
rect 140 883 281 935
rect 333 883 472 935
rect 524 883 664 935
rect 716 883 856 935
rect 908 883 1048 935
rect 1100 883 1107 935
rect -189 873 -137 883
rect 88 873 140 883
rect 281 873 333 883
rect 472 873 524 883
rect 664 873 716 883
rect 856 873 908 883
rect 1048 873 1100 883
rect -189 128 -137 138
rect 88 128 140 138
rect 279 128 331 138
rect 471 128 523 138
rect 663 128 715 138
rect 856 128 908 137
rect 1048 128 1100 137
rect -137 76 88 128
rect 140 76 279 128
rect 331 76 471 128
rect 523 76 663 128
rect 715 127 1107 128
rect 715 76 856 127
rect -189 66 -137 76
rect 88 66 140 76
rect 279 66 331 76
rect 471 66 523 76
rect 663 66 715 76
rect 908 76 1048 127
rect 856 65 908 75
rect 1100 76 1107 127
rect 1048 65 1100 75
<< labels >>
flabel metal1 -211 909 -211 909 3 FreeSans 400 0 0 0 en_b
port 4 e
flabel metal1 -212 413 -212 413 3 FreeSans 400 0 0 0 in
port 1 e
flabel metal1 -212 102 -212 102 3 FreeSans 400 0 0 0 en
port 3 e
flabel metal1 1279 412 1279 412 7 FreeSans 400 0 0 0 out
port 2 w
flabel metal1 1188 1058 1188 1058 5 FreeSans 400 0 0 0 VDD
port 5 s power bidirectional
flabel metal1 1188 -48 1188 -48 1 FreeSans 400 0 0 0 VSS
port 6 n ground bidirectional
<< end >>
