magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< pwell >>
rect -104 -146 104 146
<< nmoslvt >>
rect -20 -120 20 120
<< ndiff >>
rect -78 85 -20 120
rect -78 51 -66 85
rect -32 51 -20 85
rect -78 17 -20 51
rect -78 -17 -66 17
rect -32 -17 -20 17
rect -78 -51 -20 -17
rect -78 -85 -66 -51
rect -32 -85 -20 -51
rect -78 -120 -20 -85
rect 20 85 78 120
rect 20 51 32 85
rect 66 51 78 85
rect 20 17 78 51
rect 20 -17 32 17
rect 66 -17 78 17
rect 20 -51 78 -17
rect 20 -85 32 -51
rect 66 -85 78 -51
rect 20 -120 78 -85
<< ndiffc >>
rect -66 51 -32 85
rect -66 -17 -32 17
rect -66 -85 -32 -51
rect 32 51 66 85
rect 32 -17 66 17
rect 32 -85 66 -51
<< poly >>
rect -33 192 33 208
rect -33 158 -17 192
rect 17 158 33 192
rect -33 142 33 158
rect -20 120 20 142
rect -20 -142 20 -120
rect -33 -158 33 -142
rect -33 -192 -17 -158
rect 17 -192 33 -158
rect -33 -208 33 -192
<< polycont >>
rect -17 158 17 192
rect -17 -192 17 -158
<< locali >>
rect -33 158 -17 192
rect 17 158 33 192
rect -66 89 -32 124
rect -66 17 -32 51
rect -66 -51 -32 -17
rect -66 -124 -32 -89
rect 32 89 66 124
rect 32 17 66 51
rect 32 -51 66 -17
rect 32 -124 66 -89
rect -33 -192 -17 -158
rect 17 -192 33 -158
<< viali >>
rect -17 158 17 192
rect -66 85 -32 89
rect -66 55 -32 85
rect -66 -17 -32 17
rect -66 -85 -32 -55
rect -66 -89 -32 -85
rect 32 85 66 89
rect 32 55 66 85
rect 32 -17 66 17
rect 32 -85 66 -55
rect 32 -89 66 -85
rect -17 -192 17 -158
<< metal1 >>
rect -33 192 33 208
rect -33 158 -17 192
rect 17 158 33 192
rect -33 152 33 158
rect -72 89 -26 120
rect -72 55 -66 89
rect -32 55 -26 89
rect -72 17 -26 55
rect -72 -17 -66 17
rect -32 -17 -26 17
rect -72 -55 -26 -17
rect -72 -89 -66 -55
rect -32 -89 -26 -55
rect -72 -120 -26 -89
rect 26 89 72 120
rect 26 55 32 89
rect 66 55 72 89
rect 26 17 72 55
rect 26 -17 32 17
rect 66 -17 72 17
rect 26 -55 72 -17
rect 26 -89 32 -55
rect 66 -89 72 -55
rect 26 -120 72 -89
rect -33 -158 33 -152
rect -33 -192 -17 -158
rect 17 -192 33 -158
rect -33 -208 33 -192
<< end >>
