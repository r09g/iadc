* NGSPICE file created from sc_cmfb.ext - technology: sky130A

.subckt pmos_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136#
M0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36 l=0.15
M1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36 l=0.15
M2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36 l=0.15
M3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# pmos ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36 l=0.15
M4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36 l=0.15
M5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# pmos ad=0p pd=0u as=0p ps=0u w=1.36 l=0.15
M6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36 l=0.15
M7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# pmos ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36 l=0.15
M8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36 l=0.15
M9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# pmos ad=0p pd=0u as=0p ps=0u w=1.36 l=0.15
.ends

.subckt nmos_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
M0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=0.52 l=0.15
M1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=0.52 l=0.15
M2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=0.52 l=0.15
M3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
M4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
M5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=0.52 l=0.15
M6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=0.52 l=0.15
M7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
M8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# nmos ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=0.52 l=0.15
M9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
.ends

.subckt transmission_gate out en_b en VSS VDD in
Xpmos_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ pmos_UNG2NQ
Xnmos_6J4AMR_0 out in in out in in VSS out en in out out out nmos_6J4AMR
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580#
C0 c1_n530_n480# m3_n630_n580# cm3m4 l=4.8 w=4.8
.ends

.subckt sc_cmfb on cm bias_a op cmc p2_b p2 p1_b p1 VDD VSS
Xtransmission_gate_10 on p1_b p1 VSS VDD transmission_gate_3_out transmission_gate
Xtransmission_gate_11 op p1_b p1 VSS VDD transmission_gate_4_out transmission_gate
Xtransmission_gate_0 transmission_gate_7_in p1_b p1 VSS VDD cm transmission_gate
Xtransmission_gate_1 transmission_gate_6_in p1_b p1 VSS VDD cm transmission_gate
Xtransmission_gate_2 transmission_gate_8_in p1_b p1 VSS VDD bias_a transmission_gate
Xtransmission_gate_3 transmission_gate_3_out p2_b p2 VSS VDD cm transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4_out transmission_gate_9_in unit_cap_mim_m3m4
Xtransmission_gate_4 transmission_gate_4_out p2_b p2 VSS VDD cm transmission_gate
Xunit_cap_mim_m3m4_1 on cmc unit_cap_mim_m3m4
Xtransmission_gate_5 transmission_gate_9_in p2_b p2 VSS VDD bias_a transmission_gate
Xunit_cap_mim_m3m4_2 op cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30_c1_n530_n480# unit_cap_mim_m3m4_30_m3_n630_n580#
+ unit_cap_mim_m3m4
Xtransmission_gate_6 op p2_b p2 VSS VDD transmission_gate_6_in transmission_gate
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20_c1_n530_n480# unit_cap_mim_m3m4_20_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_3 transmission_gate_7_in transmission_gate_8_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31_c1_n530_n480# unit_cap_mim_m3m4_31_m3_n630_n580#
+ unit_cap_mim_m3m4
Xtransmission_gate_7 on p2_b p2 VSS VDD transmission_gate_7_in transmission_gate
Xunit_cap_mim_m3m4_10 transmission_gate_6_in transmission_gate_8_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21_c1_n530_n480# unit_cap_mim_m3m4_21_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_4 on cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32_c1_n530_n480# unit_cap_mim_m3m4_32_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4_out transmission_gate_9_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc unit_cap_mim_m3m4
Xtransmission_gate_8 cmc p2_b p2 VSS VDD transmission_gate_8_in transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6_in transmission_gate_8_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22_c1_n530_n480# unit_cap_mim_m3m4_22_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23_c1_n530_n480# unit_cap_mim_m3m4_23_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34_c1_n530_n480# unit_cap_mim_m3m4_34_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33_c1_n530_n480# unit_cap_mim_m3m4_33_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24_c1_n530_n480# unit_cap_mim_m3m4_24_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_6 transmission_gate_3_out transmission_gate_9_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc unit_cap_mim_m3m4
Xtransmission_gate_9 cmc p1_b p1 VSS VDD transmission_gate_9_in transmission_gate
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35_c1_n530_n480# unit_cap_mim_m3m4_35_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25_c1_n530_n480# unit_cap_mim_m3m4_25_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26_c1_n530_n480# unit_cap_mim_m3m4_26_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7_in transmission_gate_8_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3_out transmission_gate_9_in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27_c1_n530_n480# unit_cap_mim_m3m4_27_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16_c1_n530_n480# unit_cap_mim_m3m4_16_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28_c1_n530_n480# unit_cap_mim_m3m4_28_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17_c1_n530_n480# unit_cap_mim_m3m4_17_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29_c1_n530_n480# unit_cap_mim_m3m4_29_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18_c1_n530_n480# unit_cap_mim_m3m4_18_m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19_c1_n530_n480# unit_cap_mim_m3m4_19_m3_n630_n580#
+ unit_cap_mim_m3m4
.ends

