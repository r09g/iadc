magic
tech sky130A
timestamp 1654711401
<< error_p >>
rect -38 69 -9 72
rect 9 69 38 72
rect -38 52 -32 69
rect 9 52 15 69
rect -38 49 -9 52
rect 9 49 38 52
rect -38 -51 -9 -48
rect 9 -51 38 -48
rect -38 -68 -32 -51
rect 9 -68 15 -51
rect -38 -71 -9 -68
rect 9 -71 38 -68
<< pwell >>
rect -155 -137 155 138
<< nmos >>
rect -55 -32 -40 33
rect -7 -32 7 33
rect 40 -32 55 33
<< ndiff >>
rect -86 27 -55 33
rect -86 -26 -80 27
rect -63 -26 -55 27
rect -86 -32 -55 -26
rect -40 27 -7 33
rect -40 -26 -32 27
rect -15 -26 -7 27
rect -40 -32 -7 -26
rect 7 27 40 33
rect 7 -26 15 27
rect 32 -26 40 27
rect 7 -32 40 -26
rect 55 27 86 33
rect 55 -26 63 27
rect 80 -26 86 27
rect 55 -32 86 -26
<< ndiffc >>
rect -80 -26 -63 27
rect -32 -26 -15 27
rect 15 -26 32 27
rect 63 -26 80 27
<< psubdiff >>
rect -137 103 -89 120
rect 89 103 137 120
rect -137 72 -120 103
rect 120 72 137 103
rect -137 -102 -120 -71
rect 120 -102 137 -71
rect -137 -119 -89 -102
rect 89 -119 137 -102
<< psubdiffcont >>
rect -89 103 89 120
rect -137 -71 -120 72
rect 120 -71 137 72
rect -89 -119 89 -102
<< poly >>
rect -64 69 64 77
rect -64 52 -32 69
rect -15 52 15 69
rect 32 52 64 69
rect -64 44 64 52
rect -55 33 -40 44
rect -7 33 7 44
rect 40 33 55 44
rect -55 -43 -40 -32
rect -7 -43 7 -32
rect 40 -43 55 -32
rect -64 -51 64 -43
rect -64 -68 -32 -51
rect -15 -68 15 -51
rect 32 -68 64 -51
rect -64 -76 64 -68
<< polycont >>
rect -32 52 -15 69
rect 15 52 32 69
rect -32 -68 -15 -51
rect 15 -68 32 -51
<< locali >>
rect -137 103 -89 120
rect 89 103 137 120
rect -137 72 -120 103
rect 120 72 137 103
rect -40 52 -32 69
rect -15 52 15 69
rect 32 52 40 69
rect -80 27 -63 35
rect -80 -34 -63 -26
rect -32 27 -15 35
rect -32 -34 -15 -26
rect 15 27 32 35
rect 15 -34 32 -26
rect 63 27 80 35
rect 63 -34 80 -26
rect -40 -68 -32 -51
rect -15 -68 15 -51
rect 32 -68 40 -51
rect -137 -102 -120 -71
rect 120 -102 137 -71
rect -137 -119 -89 -102
rect 89 -119 137 -102
<< viali >>
rect -32 52 -15 69
rect 15 52 32 69
rect -80 -26 -63 27
rect -32 -26 -15 27
rect 15 -26 32 27
rect 63 -26 80 27
rect -32 -68 -15 -51
rect 15 -68 32 -51
<< metal1 >>
rect -38 69 -9 72
rect -38 52 -32 69
rect -15 52 -9 69
rect -38 49 -9 52
rect 9 69 38 72
rect 9 52 15 69
rect 32 52 38 69
rect 9 49 38 52
rect -83 27 -60 33
rect -83 9 -80 27
rect -138 -9 -80 9
rect -83 -26 -80 -9
rect -63 9 -60 27
rect -35 27 -12 33
rect -35 9 -32 27
rect -63 -9 -32 9
rect -63 -26 -60 -9
rect -83 -32 -60 -26
rect -35 -26 -32 -9
rect -15 9 -12 27
rect 12 27 35 33
rect 12 9 15 27
rect -15 -9 15 9
rect -15 -26 -12 -9
rect -35 -32 -12 -26
rect 12 -26 15 -9
rect 32 9 35 27
rect 60 27 83 33
rect 60 9 63 27
rect 32 -9 63 9
rect 32 -26 35 -9
rect 12 -32 35 -26
rect 60 -26 63 -9
rect 80 9 83 27
rect 80 -9 138 9
rect 80 -26 83 -9
rect 60 -32 83 -26
rect -38 -51 -9 -48
rect -38 -68 -32 -51
rect -15 -68 -9 -51
rect -38 -71 -9 -68
rect 9 -51 38 -48
rect 9 -68 15 -51
rect 32 -68 38 -51
rect 9 -71 38 -68
<< properties >>
string FIXED_BBOX -129 -111 129 111
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.65 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
