* NGSPICE file created from clock_flat.ext - technology: sky130A

.subckt clock_flat clk p2d_b p2d p2_b p2 p1d_b p1d p1_b p1 Ad_b Ad A_b A Bd_b Bd B_b
+ B VDD VSS
X0 VSS a_6941_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS sky130_fd_pr__nfet_01v8 ad=2.2138e+14p pd=2.39592e+09u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1 VDD a_5653_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD sky130_fd_pr__pfet_01v8_hvt ad=3.8151e+14p pd=3.51993e+09u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2 a_9876_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X5 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6 VSS a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X7 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X8 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X9 a_n1738_n6671# a_n2602_n7037# a_n1995_n6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X10 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X11 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X12 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X13 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X14 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X15 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_4661_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X16 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X17 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X18 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X19 a_9876_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X21 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X23 a_3077_n1909# a_3176_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X24 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u
X25 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X26 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_7237_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_9517_n4709# a_9616_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X28 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X29 VDD a_2148_n3799# a_1888_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X30 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X31 VDD a_7130_n10301# a_7237_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X32 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X33 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6874_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X34 VDD sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X35 VDD a_8418_n6493# a_8525_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X36 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X37 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X38 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X39 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X40 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X41 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X42 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X43 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X44 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X45 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 a_6012_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X47 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X48 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X49 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X50 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X51 VSS a_3436_n9783# a_3176_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X52 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X53 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X54 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X55 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X56 a_9706_n8125# a_9450_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X57 a_8418_n1597# a_8162_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X58 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X59 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X60 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X61 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X62 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_3373_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X63 a_3077_n3621# a_3176_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X64 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X65 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X67 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X68 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X69 VSS sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X70 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X71 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X72 VSS sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X73 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X74 VDD a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X75 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X76 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X77 VSS a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X78 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X79 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X80 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X81 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X82 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X84 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X85 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X86 VSS sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X87 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X88 VDD sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X89 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X90 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X91 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X92 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X95 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X96 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X97 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X99 VSS sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X100 VDD clk sky130_fd_sc_hd__clkinv_1_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X101 a_7130_n509# a_6874_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X102 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X103 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X104 VDD a_3436_n13591# a_3176_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X105 a_5842_n11933# a_5586_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X106 VDD sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X107 a_3077_n8437# a_3176_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X108 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X109 VDD a_9706_n5405# a_9813_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X110 a_3266_n10301# a_3010_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X111 VDD a_6012_n8695# a_5752_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X112 VSS a_7130_n8125# a_7237_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X113 a_10805_n5797# a_10904_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X114 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X115 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X116 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X117 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 VDD a_8588_n8695# a_8328_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X119 VDD a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X120 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X121 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X122 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X123 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X124 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_3373_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X125 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X126 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X127 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4298_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X128 VSS a_n1995_n6925# a_n2037_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X129 VSS a_5842_n13021# a_5949_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X130 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X131 a_5653_n12325# a_5752_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X132 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X133 sky130_fd_sc_hd__nand2_4_2/B a_9813_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X134 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X135 a_501_n3621# a_600_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X136 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_8525_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X137 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X138 VDD a_5653_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X139 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_10738_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X140 a_4365_n11237# a_4464_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X141 VDD a_4554_n10301# a_4661_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X142 VSS a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X143 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X144 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X145 VDD a_9706_n2685# a_9813_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X146 a_8418_n5405# a_8162_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X147 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X148 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X149 a_7130_n4317# a_6874_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X150 VDD a_3436_n12503# a_3176_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X151 VDD a_690_n10301# a_797_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X152 a_8229_n821# a_8328_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X153 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_6874_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X154 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_3373_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X155 VDD sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 VSS a_6012_n13591# a_5752_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X157 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_2085_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X158 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X159 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_9813_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X160 VDD a_4554_n5405# a_4661_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X161 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u
X162 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X163 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X164 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X165 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X166 a_860_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X167 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_797_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X168 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X169 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_8525_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X171 VSS sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X173 VDD a_3436_n8695# a_3176_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X174 VDD sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X175 a_1978_n10301# a_1722_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X176 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_9813_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X177 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8525_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X178 VDD a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X179 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X180 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X181 a_8418_n14109# a_8162_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X182 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X183 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X184 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X185 a_2622_n509# a_2366_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X186 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X187 VSS sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X188 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X189 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_1722_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X190 VDD a_4554_n2685# a_4661_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X191 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X192 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X193 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_9813_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X194 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X195 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X196 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X197 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X198 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X199 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X200 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X201 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X202 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_5949_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X203 VDD a_690_n4317# a_797_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X204 a_690_n9213# a_434_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X205 VDD sky130_fd_sc_hd__clkinv_1_0/Y a_2366_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X206 a_4554_n4317# a_4298_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X207 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X208 VSS a_5842_n4317# a_5949_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X209 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 VSS a_501_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X211 VDD a_3077_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X212 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_6006_n7607# a_6101_n7254# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X214 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X216 a_5842_n2685# a_5586_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X217 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_n2436_n7037# a_n2602_n7037# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X219 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X220 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X221 VSS a_8418_n4317# a_8525_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X222 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X223 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X224 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X225 VSS sky130_fd_sc_hd__nand2_4_0/B a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X226 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X227 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X228 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X229 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X230 VDD a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X231 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X232 a_10994_n5405# a_10738_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X233 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_8525_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X234 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X235 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X236 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X237 a_n2436_n7037# a_n2602_n7037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X238 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X239 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_7237_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X240 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X241 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 VDD a_10994_n9213# a_11101_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X243 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9450_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X244 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X245 VDD a_5842_n11933# a_5949_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X246 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X247 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X248 VSS a_n428_n4887# a_n688_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X249 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_434_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X250 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X251 VDD a_7300_n3799# a_7040_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X252 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_797_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X253 VSS a_501_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_59/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X254 a_n787_n12325# a_n688_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X255 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X256 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X258 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X259 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X260 a_1789_n11237# a_1888_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X261 VDD a_9876_n3799# a_9616_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X262 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X263 VDD sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X264 a_5653_n2997# a_5752_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X265 VDD a_8588_n13591# a_8328_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X266 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X267 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X268 a_1978_n4317# a_1722_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X269 a_10994_n2685# a_10738_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X270 VSS a_3266_n4317# a_3373_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X271 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_9706_n9213# a_9450_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X273 VDD a_7300_n11415# a_7040_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X274 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X275 a_1789_n10613# a_1888_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X276 VSS a_3077_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X277 sky130_fd_sc_hd__dfxbp_1_1/D a_n1139_n6715# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X278 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_9450_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X279 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X280 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X281 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X282 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X283 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X284 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X285 VSS a_7130_n14109# a_7237_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X286 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X287 VDD a_6006_n7607# sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X288 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X289 VSS a_n428_n9783# a_n688_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X290 VDD a_501_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_59/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X291 a_11164_n5975# sky130_fd_sc_hd__clkinv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X292 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X293 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11101_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X294 VSS a_7300_n10871# a_7040_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X295 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X296 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X297 VDD a_10994_n10301# a_11101_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X298 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X299 VDD a_9706_n10301# a_9813_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X300 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X301 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3373_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X302 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X304 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X305 VDD sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X306 sky130_fd_sc_hd__nand2_4_2/B a_9813_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X307 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6874_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X309 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X310 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_8525_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X311 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X312 a_5653_n1909# a_5752_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X313 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X314 VDD a_8588_n12503# a_8328_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X315 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X317 VDD a_4724_n3799# a_4464_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X318 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X319 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X320 VSS sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X321 VDD a_6012_n5975# a_5752_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X322 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7237_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X323 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X324 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X325 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X326 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X327 VSS sky130_fd_sc_hd__nand2_4_3/B a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X328 VSS sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X329 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X330 VDD sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X331 a_8588_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X332 VDD sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X333 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_5949_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X334 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X335 VDD a_7130_n9213# a_7237_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X336 VDD a_4623_n7349# sky130_fd_sc_hd__mux2_1_0/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X337 VSS sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 VDD a_8588_n5975# a_8328_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X339 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X340 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X341 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X342 a_11164_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X343 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_10738_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X344 VDD sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X345 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X346 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X347 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X348 VSS sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X349 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3373_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X350 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 VSS a_5842_n9213# a_5949_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X352 a_5653_n3621# a_5752_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X353 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X354 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X355 a_6794_n7203# a_6658_n7363# a_6373_n7349# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X356 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X357 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X358 VSS a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X359 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X360 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_3373_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X361 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X362 VSS a_8418_n9213# a_8525_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X363 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X364 a_7130_n1597# a_6874_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X365 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X366 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X367 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X368 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X369 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 VDD sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X371 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X372 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X373 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X374 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X375 VDD sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 a_n860_n6173# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X377 a_1978_n13021# a_1722_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X378 a_6941_n10613# a_7040_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X379 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3010_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X380 a_11164_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X381 a_7300_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X382 VDD a_3436_n5975# a_3176_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X383 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X386 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X387 a_10805_n13413# a_10904_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X388 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X389 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X390 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X391 VDD a_2622_n8125# a_2729_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X392 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X393 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_5653_n8437# a_5752_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X395 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X396 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X397 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X398 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X399 a_8418_n5405# a_8162_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X400 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X401 VSS a_n1738_n6671# a_n1570_n6769# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X402 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X403 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X404 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11101_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X405 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X406 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5586_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X407 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X408 VSS a_1978_n2685# a_2085_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X409 a_n428_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X410 VSS a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X411 VSS a_3266_n9213# a_3373_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X412 VSS a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X413 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X414 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X415 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X416 VSS a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X417 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 VSS a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X419 VDD a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X420 VDD a_690_n1597# a_797_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X421 VDD a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X422 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X423 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X424 a_n2037_n7037# a_n2436_n7037# a_n2163_n6671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X425 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X426 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X427 a_4554_n1597# a_4298_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X428 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X429 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X430 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X431 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X432 a_8418_n10301# a_8162_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X433 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X434 VDD a_2148_n10871# a_1888_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X435 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X436 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X437 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9450_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X438 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X439 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X440 a_8418_n2685# a_8162_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X441 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X442 VSS a_n787_n12325# sky130_fd_sc_hd__nand2_1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X443 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X444 a_3077_n4709# a_3176_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X445 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X446 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X447 VDD sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X448 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X449 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11101_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X450 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X452 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X453 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_n428_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X455 VDD a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X456 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X457 VDD a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X458 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X460 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X461 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X462 a_n787_n1909# a_n688_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X463 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 VSS a_11164_n5975# a_10904_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X465 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X466 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 VDD a_2148_n3255# a_1888_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X468 VDD a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X469 a_6941_n2997# a_7040_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X470 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_434_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X471 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X472 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X473 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X474 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X475 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X476 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X477 VDD a_4365_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X478 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4298_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X479 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X480 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X481 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X482 VDD a_n787_n12325# sky130_fd_sc_hd__nand2_1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X483 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X484 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X485 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X486 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_5949_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X487 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X488 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_4661_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X489 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X490 a_2622_n6493# a_2366_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X491 VDD sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X492 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X493 a_9517_n5797# a_9616_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X494 a_6941_n821# a_7040_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X495 a_1978_n1597# a_1722_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X496 a_4724_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X497 a_501_n10613# a_600_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X498 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X499 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X500 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7237_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X501 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6874_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X502 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_8525_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X503 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X504 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X505 VSS sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 a_2622_n14109# a_2366_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X507 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9813_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X508 VSS a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X509 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X510 VSS a_11164_n4887# a_10904_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X511 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8162_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X512 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_1_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X513 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X515 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X516 VDD a_2148_n2167# a_1888_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X517 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X518 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X519 a_6941_n1909# a_7040_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X520 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X521 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=0p ps=0u w=840000u l=150000u
X522 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X523 a_5653_n13413# a_5752_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X524 a_6941_n9525# a_7040_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X525 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X526 VSS a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X527 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X528 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X529 VDD a_9706_n8125# a_9813_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X530 VSS sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X531 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X532 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X533 VSS a_860_n3255# a_600_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X534 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X535 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__mux2_1_0/X a_3832_n7261# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X536 a_7130_n509# a_6874_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X537 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X539 a_8229_n11237# a_8328_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X540 a_4365_n2997# a_4464_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X541 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X542 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X543 a_4724_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X544 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7237_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X545 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X546 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X547 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X548 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_797_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X549 a_9517_n4709# a_9616_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X550 VDD sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X551 VSS a_2148_n3799# a_1888_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X552 VSS a_7130_n10301# a_7237_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X553 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X554 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X555 VDD a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X556 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X557 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X558 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_8525_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X559 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9450_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X560 a_8229_n10613# a_8328_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X561 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X562 a_7130_n11933# a_6874_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X563 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X564 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X565 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_2085_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X566 VSS a_11164_n9783# a_10904_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X567 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X568 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X569 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X570 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X571 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X572 a_5653_n12325# a_5752_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X573 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_4661_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X574 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X575 a_501_n2997# a_600_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X576 a_8229_n3621# a_8328_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X577 VSS a_9706_n14109# a_9813_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X578 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X579 a_6941_n12325# a_7040_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X580 VDD a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X581 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X582 VSS a_860_n2167# a_600_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X583 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X584 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_7237_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X585 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X586 a_4365_n1909# a_4464_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X587 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X588 VDD a_860_n9783# a_600_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X589 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X590 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X591 VDD a_5842_n10301# a_5949_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X592 a_4365_n9525# a_4464_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X593 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X595 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X596 a_9517_n9525# a_9616_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X597 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X598 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 VSS a_2148_n8695# a_1888_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X600 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X601 VSS a_3266_n13021# a_3373_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X602 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_2085_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X603 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X604 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X605 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X607 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X608 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X609 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X610 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6874_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X611 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X612 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X613 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X614 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X615 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8162_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X616 a_1789_n2997# a_1888_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X617 a_8418_n14109# a_8162_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X618 a_1789_n11237# a_1888_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X619 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X620 VSS a_n1570_n6769# a_n1612_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X621 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_11101_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X622 VSS a_1978_n11933# a_2085_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X623 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X625 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X626 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X627 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X628 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_4661_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X629 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X630 a_n2248_n7037# sky130_fd_sc_hd__dfxbp_1_1/D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X631 VSS sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X633 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X634 a_501_n1909# a_600_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X635 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_9450_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X636 VSS a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X637 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6874_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X638 VSS a_2622_n6493# a_2729_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X639 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X640 VSS a_3436_n13591# a_3176_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X641 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X642 VSS a_7300_n11415# a_7040_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X643 a_2622_n509# a_2366_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X644 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X645 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X646 a_3266_n10301# a_3010_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X647 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X648 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X649 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X650 VDD sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X651 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X652 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_5586_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X653 a_9706_n6493# a_9450_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X654 VSS a_2148_n12503# a_1888_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X655 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X656 VSS sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X657 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X658 a_n860_n509# sky130_fd_sc_hd__nand2_1_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X659 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X660 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X661 VSS a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X662 VDD a_5842_n4317# a_5949_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X663 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X664 VDD a_10805_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X665 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X666 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X667 VSS a_3077_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X668 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X669 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X670 a_1789_n1909# a_1888_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X671 a_501_n3621# a_600_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X672 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X673 a_8418_n13021# a_8162_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X674 VDD a_8418_n4317# a_8525_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X675 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X676 VSS a_4554_n10301# a_4661_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X677 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X678 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X679 a_1789_n9525# a_1888_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X680 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X681 VSS a_9706_n2685# a_9813_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X682 VDD a_9517_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X683 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X684 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_3373_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X685 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X686 VDD a_8229_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X687 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X688 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X689 a_9517_n10613# a_9616_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X690 VSS a_690_n10301# a_797_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X691 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X692 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X693 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_2729_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X694 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X695 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X696 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X697 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X698 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3010_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X699 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X700 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X702 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X703 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_5949_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X704 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X705 VDD a_11164_n8695# a_10904_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X706 VSS a_1789_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X707 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X708 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4298_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X709 VSS sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X710 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_5586_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X711 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6874_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X712 VDD a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X713 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X714 VDD a_7130_n6493# a_7237_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X715 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X716 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X717 VSS sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X718 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X719 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X720 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X721 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X722 VDD sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X723 a_501_n12325# a_600_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X724 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 a_501_n8437# a_600_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X726 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X727 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_434_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X728 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X729 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X730 sky130_fd_sc_hd__clkinv_1_6/Y clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X731 VDD a_7300_n3255# a_7040_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X732 a_7130_n1597# a_6874_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X733 VDD a_3266_n4317# a_3373_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X734 a_3266_n9213# a_3010_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X735 VDD a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X736 VDD a_6101_n7254# sky130_fd_sc_hd__dfxbp_1_0/Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X737 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X738 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X739 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_2085_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X740 VDD a_9876_n3255# a_9616_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X741 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X742 a_6865_n7304# a_6665_n7459# a_7014_n7215# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.392e+11p ps=1.53e+06u w=360000u l=150000u
X743 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X744 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X745 VSS a_4554_n2685# a_4661_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X746 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X747 a_9517_n8437# a_9616_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X748 VSS a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X749 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 VDD a_7130_n14109# a_7237_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X751 VDD a_3266_n11933# a_3373_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X752 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X753 VDD a_1789_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X754 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4298_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X755 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X756 a_3077_n11237# a_3176_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X757 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X758 VDD a_6941_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X759 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X760 VDD a_5653_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X761 a_10994_n13021# a_10738_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X762 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X763 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_797_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X764 VSS a_9517_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X765 a_3077_n10613# a_3176_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X766 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X768 VDD a_7300_n2167# a_7040_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X769 a_10805_n2997# a_10904_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X770 a_5653_n4709# a_5752_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X771 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X772 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1722_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X774 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X775 a_690_n4317# a_434_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X776 VSS a_9706_n6493# a_9813_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X777 VSS sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X778 VSS a_9517_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X779 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X780 VDD a_4724_n11415# a_4464_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X781 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X782 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X783 VDD a_9876_n2167# a_9616_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X784 VDD a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X785 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_6874_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X786 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X787 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X789 VDD a_7130_n13021# a_7237_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X790 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X791 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X792 VSS a_690_n1597# a_797_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X793 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X794 VDD a_4724_n3255# a_4464_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X795 VDD a_860_n11415# a_600_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X796 a_4554_n1597# a_4298_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X797 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X798 VSS a_8418_n13021# a_8525_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X799 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X800 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_797_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X801 VSS a_4724_n10871# a_4464_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X802 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_9813_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X803 VDD a_6941_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X804 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_8525_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X805 VSS a_7300_n3799# a_7040_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X806 VDD sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X807 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X808 VDD a_9517_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X809 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4298_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X810 VSS a_8229_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X811 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X812 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X813 VSS a_860_n10871# a_600_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X814 VDD sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X815 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1722_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X816 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X817 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8525_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X818 VSS a_10994_n4317# a_11101_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X819 a_10805_n1909# a_10904_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X820 VSS a_9876_n3799# a_9616_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X821 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3010_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X822 a_7130_n5405# a_6874_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X823 VSS a_8588_n13591# a_8328_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X824 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X825 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_5949_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X826 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_4661_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X827 a_10805_n9525# a_10904_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X828 a_10994_n2685# a_10738_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X829 VDD sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X830 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X831 a_6941_n821# a_7040_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X832 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X833 VSS a_6941_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X834 a_6373_n7349# a_6665_n7459# a_6616_n7581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X835 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X836 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9450_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X837 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X838 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X839 VDD a_4724_n2167# a_4464_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X840 sky130_fd_sc_hd__nand2_4_1/B a_9813_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X841 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 a_9876_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X843 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X844 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X845 a_9706_n4317# a_9450_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X846 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X847 VSS a_7300_n8695# a_7040_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X848 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X849 VSS a_10805_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X850 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X851 VSS a_10994_n10301# a_11101_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X852 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X853 VSS a_9706_n10301# a_9813_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X854 a_8418_n8125# a_8162_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X855 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X856 a_9706_n11933# a_9450_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X857 VSS sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X858 a_1978_n1597# a_1722_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X859 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_5/A a_n860_n6173# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X860 VSS a_9876_n8695# a_9616_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X861 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X862 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_1_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=0p ps=0u w=840000u l=150000u
X863 a_3266_n13021# a_3010_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X864 a_n860_n8125# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X865 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X866 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X867 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X868 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X869 VSS a_4724_n3799# a_4464_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X870 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X871 VDD a_6941_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X872 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_797_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X873 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9450_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X875 VSS a_9517_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X876 VDD a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X877 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X878 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X879 a_4365_n10613# a_4464_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X880 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X881 a_10994_n11933# a_10738_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X882 VSS a_690_n5405# a_797_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X883 a_9517_n12325# a_9616_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X884 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X885 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_5949_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X886 VDD a_5842_n1597# a_5949_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X887 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X888 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3010_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X889 a_4554_n5405# a_4298_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X890 VSS sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X891 VSS clk a_n2602_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X892 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X893 VDD a_860_n1079# a_600_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X894 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X895 VSS a_n1570_n6769# a_n1139_n6715# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X896 a_4365_n821# a_4464_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X897 VDD sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X898 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X899 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X900 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X901 VDD a_4554_n13021# a_4661_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X902 a_8229_n11237# a_8328_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X903 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X904 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X905 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X906 VDD a_8418_n1597# a_8525_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X907 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6874_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X908 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X909 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X910 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X911 VSS a_7130_n4317# a_7237_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X912 VDD a_690_n13021# a_797_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X913 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X914 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_7237_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X915 VDD clk a_n2602_n7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X916 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X917 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X918 VSS a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X919 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X920 a_n787_n4709# a_n688_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X921 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X922 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X923 a_690_n9213# a_434_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X924 VSS a_4724_n8695# a_4464_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X925 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X926 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X927 VDD a_8418_n11933# a_8525_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X928 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X929 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X931 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X932 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X933 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X934 VDD a_11164_n5975# a_10904_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X935 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X936 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X937 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X938 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X939 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X940 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X941 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_797_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X942 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X943 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6874_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X944 VSS a_6941_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X945 a_3436_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X946 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X947 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X948 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X949 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X950 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X951 a_3077_n5797# a_3176_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X952 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X953 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_2085_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X954 a_1978_n5405# a_1722_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X955 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X956 VSS a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X957 VDD a_3266_n1597# a_3373_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X958 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X959 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X960 VDD a_11164_n11415# a_10904_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X961 VDD a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X962 VSS a_10994_n9213# a_11101_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X963 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X964 a_2622_n14109# a_2366_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X965 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X966 VDD a_9876_n11415# a_9616_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X967 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X968 a_1789_n821# a_1888_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X969 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X970 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X971 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X972 a_9517_n5797# a_9616_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X973 VDD a_2148_n4887# a_1888_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X974 a_n2163_n6671# a_n2436_n7037# a_n2248_n7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X975 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X976 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X977 VDD sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X978 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X979 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X980 VSS a_11164_n10871# a_10904_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X981 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X982 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_5949_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X983 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X984 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X985 VSS a_9876_n10871# a_9616_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X986 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_10738_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X987 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X988 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X989 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X990 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X991 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X992 a_8418_n2685# a_8162_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X993 VDD sky130_fd_sc_hd__clkinv_1_5/A a_7212_n7203# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X994 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X995 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_3373_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X996 a_9706_n9213# a_9450_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X997 VSS a_6012_n3255# a_5752_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X998 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5586_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X999 a_3077_n4709# a_3176_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1000 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1001 a_6941_n13413# a_7040_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1002 VSS sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1003 VSS sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1004 VSS a_4724_n1079# a_4464_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1005 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1006 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3010_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1007 VSS a_8588_n3255# a_8328_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1008 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8525_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1009 VDD a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1010 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1011 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_434_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1012 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1013 a_3832_n7261# sky130_fd_sc_hd__nand2_1_4/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1014 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1015 VSS a_501_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1016 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1017 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1018 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1019 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1020 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1021 VSS a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1022 VSS a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1023 VDD a_9706_n14109# a_9813_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1024 a_5842_n9213# a_5586_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1025 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1026 a_9876_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1027 sky130_fd_sc_hd__nand2_4_0/B a_9813_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1028 VSS a_3436_n1079# a_3176_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1029 VSS a_6012_n2167# a_5752_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1030 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1031 a_5842_n13021# a_5586_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1032 VDD sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1034 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1035 a_3077_n9525# a_3176_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1036 a_8229_n2997# a_8328_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1037 a_6941_n12325# a_7040_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1038 VDD a_6012_n9783# a_5752_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1039 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1040 VSS a_7130_n9213# a_7237_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1041 a_n1995_n6925# a_n2163_n6671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X1042 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1043 VSS a_8588_n2167# a_8328_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1044 VDD a_2148_n13591# a_1888_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1045 a_4554_n11933# a_4298_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1046 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1047 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1048 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1049 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1050 VDD a_501_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1051 VDD a_8588_n9783# a_8328_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1052 VSS a_3436_n3255# a_3176_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1053 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1055 VDD a_501_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1056 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1057 VSS a_2148_n1079# a_1888_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1058 a_690_n11933# a_434_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1059 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1060 a_860_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1061 VDD sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1062 a_5653_n13413# a_5752_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1063 a_7041_n7581# a_6794_n7203# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1064 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3010_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1065 VDD a_10994_n13021# a_11101_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1066 a_501_n4709# a_600_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1067 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1068 VDD a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1069 VDD a_9706_n13021# a_9813_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1070 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1071 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1072 a_4365_n12325# a_4464_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1073 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_5949_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1074 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_7237_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1075 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1076 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_7237_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1077 a_8418_n6493# a_8162_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1078 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1079 a_7130_n5405# a_6874_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1080 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1081 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1082 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1083 a_3077_n11237# a_3176_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1084 VDD a_3266_n10301# a_3373_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1085 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1086 a_8229_n1909# a_8328_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1087 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1088 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1089 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1090 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1091 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9813_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1092 VDD a_2148_n12503# a_1888_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1093 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1094 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1095 VSS sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1096 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_434_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1097 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 a_10805_n821# a_10904_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1099 VSS a_3436_n2167# a_3176_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1100 a_6865_n7304# a_6658_n7363# a_7041_n7581# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1101 VSS a_2622_n8125# a_2729_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1102 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_797_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1103 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1104 VSS a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1105 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1106 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1107 a_860_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1108 VSS sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1109 VDD a_3436_n9783# a_3176_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1110 VDD a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1111 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1112 a_501_n13413# a_600_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1113 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1114 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1115 VSS a_4724_n11415# a_4464_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1116 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_5949_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1117 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1118 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_8525_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1119 a_8229_n3621# a_8328_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1120 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1121 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1122 a_7130_n2685# a_6874_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1123 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1124 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1125 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7237_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1126 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1127 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1128 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1129 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 VSS a_860_n11415# a_600_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1131 a_n2163_n6671# a_n2602_n7037# a_n2248_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X1132 VDD a_n1570_n6769# a_n1139_n6715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1133 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1134 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_797_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1135 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1136 VSS sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1137 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1138 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1139 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1140 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1141 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9813_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1142 VSS a_5842_n10301# a_5949_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1143 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1144 VDD sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkinv_1_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1145 a_11164_n5975# sky130_fd_sc_hd__clkinv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1146 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1147 VSS sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1148 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1149 VDD a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1150 VDD a_690_n5405# a_797_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1151 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1152 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1153 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1154 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1155 a_4554_n5405# a_4298_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1156 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1157 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1158 VDD a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1159 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1160 a_501_n12325# a_600_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1161 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1162 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1163 a_5842_n11933# a_5586_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1164 VDD a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1165 a_3077_n8437# a_3176_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1166 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1167 a_8229_n8437# a_8328_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1168 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1169 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_797_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1170 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1171 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1173 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1174 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1175 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1176 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1177 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1178 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5586_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1179 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_8525_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1180 VDD sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 VDD a_690_n2685# a_797_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1182 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1183 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1184 a_4554_n2685# a_4298_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1185 VSS a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1186 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9450_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1187 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A a_11101_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1188 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1189 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8162_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1190 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u
X1191 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1192 VSS a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1193 VSS a_4365_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1194 a_n1995_n6925# a_n2163_n6671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1195 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1196 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1197 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_434_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1198 VDD a_7300_n4887# a_7040_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1199 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1200 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1201 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1202 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1203 a_690_n4317# a_434_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1204 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1205 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1206 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1207 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1208 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1209 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1210 VDD a_9876_n4887# a_9616_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1211 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1212 VSS a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1213 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1214 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1215 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X1216 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1217 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1218 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1219 a_1978_n5405# a_1722_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1220 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1221 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1222 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1223 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1225 VSS a_5842_n1597# a_5949_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1226 a_10994_n10301# a_10738_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1227 VDD a_1978_n9213# a_2085_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1228 a_8588_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1229 VDD a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1230 a_7300_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1231 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1232 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1233 VDD a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1234 VDD a_6012_n11415# a_5752_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1235 VSS a_8418_n1597# a_8525_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1236 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1237 VSS a_9706_n8125# a_9813_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1238 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1239 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8162_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1240 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1241 VDD a_10994_n4317# a_11101_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1242 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1243 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1244 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_2729_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1245 VDD sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1246 VSS sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1247 a_5653_n5797# a_5752_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1248 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_3373_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1249 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X1250 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1251 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1254 VSS sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1255 VSS a_6012_n10871# a_5752_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1256 a_6941_n3621# a_7040_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1257 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5586_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1258 a_1978_n2685# a_1722_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1259 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6874_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1260 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1261 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1262 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3010_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1263 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1264 VDD a_8418_n10301# a_8525_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1265 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1266 VDD a_4724_n4887# a_4464_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1267 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1268 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1269 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_7237_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1270 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1272 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1273 a_3266_n4317# a_3010_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1274 a_9706_n4317# a_9450_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1275 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1276 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1722_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1277 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_5949_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1278 a_9517_n13413# a_9616_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1279 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1280 VDD a_8229_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1281 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1282 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1283 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X1284 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1285 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10738_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1286 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1287 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1288 VSS a_3266_n1597# a_3373_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1289 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_3373_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1290 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X1291 VSS a_11164_n11415# a_10904_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1292 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1293 VSS a_9876_n11415# a_9616_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1294 a_3436_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1295 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1296 a_5653_n4709# a_5752_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1297 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1298 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1299 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1300 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1301 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3010_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1302 VSS a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1303 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5586_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1304 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1305 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1306 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1307 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1308 VSS a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1309 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1310 a_8588_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1311 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1312 VDD sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1313 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_434_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1314 VSS a_5842_n5405# a_5949_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1315 VDD a_860_n3799# a_600_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1316 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 VSS sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1318 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1319 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1320 a_4365_n3621# a_4464_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1321 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1322 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1323 VDD a_6012_n1079# a_5752_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1324 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1326 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_4/Y a_n860_n8125# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1327 a_9517_n12325# a_9616_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1328 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1329 VSS a_8418_n5405# a_8525_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1330 VDD a_7130_n4317# a_7237_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1331 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1332 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1333 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1334 VDD a_8588_n1079# a_8328_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1335 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1336 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1337 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1338 a_5653_n9525# a_5752_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1339 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1340 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1341 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9450_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1342 VDD a_5653_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1343 a_8588_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1344 a_n2248_n7037# sky130_fd_sc_hd__dfxbp_1_1/D VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1345 VDD a_5842_n13021# a_5949_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1346 a_1789_n10613# a_1888_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1347 VSS a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1348 VSS a_n428_n2167# a_n688_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1349 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X1350 VSS a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1351 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1352 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1353 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_89/A a_2366_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1354 VSS sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1355 VDD a_n428_n9783# a_n688_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1356 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_5586_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1357 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1358 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1359 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1360 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1361 VDD a_7300_n10871# a_7040_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1362 VSS sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1363 VSS a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1364 VSS a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1365 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1366 VDD a_501_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1367 a_6101_n7254# a_6373_n7349# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1368 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1369 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1370 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_8525_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1371 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_434_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1373 VSS a_3266_n5405# a_3373_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1374 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1375 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_4661_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1376 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1377 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1378 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1379 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1380 VDD a_3436_n1079# a_3176_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1381 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1382 a_1789_n3621# a_1888_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1383 VSS sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1384 a_3077_n5797# a_3176_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1385 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1386 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1387 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1388 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1389 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1390 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_8525_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1391 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1392 VDD a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1393 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1394 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1395 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1396 VSS a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1397 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_11101_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1398 VSS a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1399 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1400 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1401 VDD a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1402 VDD a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1403 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1404 a_7212_n7203# a_6658_n7363# a_6865_n7304# VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=360000u l=150000u
X1405 VDD sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1406 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1407 a_3266_n9213# a_3010_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1408 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1409 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1410 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1411 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_8525_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1412 a_8588_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1413 VSS a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1414 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1415 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_7237_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1416 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1417 VSS a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1418 VSS a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1419 a_690_n1597# a_434_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1420 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3010_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1421 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1422 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1423 VDD sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1424 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_5949_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1425 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1426 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1427 a_n787_n4709# a_n688_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1428 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1429 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6874_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1430 VSS a_2148_n5975# a_1888_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1431 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1432 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1433 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1434 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1435 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1436 VSS a_4365_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1437 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1438 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1439 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8162_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1440 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1441 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1442 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1443 a_11164_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1444 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1445 a_5653_n8437# a_5752_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1446 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1447 VDD a_10994_n1597# a_11101_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1448 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1449 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1450 a_4365_n13413# a_4464_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1451 VDD a_9706_n9213# a_9813_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1452 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1453 VSS sky130_fd_sc_hd__nand2_4_2/B a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1454 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1455 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1456 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1457 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1458 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1459 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1460 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1461 VDD a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1462 VSS a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1463 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 a_10805_n11237# a_10904_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1465 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1466 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1467 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1468 a_n787_n9525# a_n688_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1469 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1470 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_797_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1471 VSS a_2148_n4887# a_1888_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1472 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1473 VSS a_5653_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1474 VDD a_4365_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1475 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1476 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1477 VSS a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1478 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1479 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1480 a_7130_n13021# a_6874_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1481 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1482 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1483 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1484 a_10805_n10613# a_10904_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1485 a_9706_n1597# a_9450_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1486 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1487 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1488 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1489 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1490 a_5842_n10301# a_5586_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1491 VSS sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1492 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1493 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1494 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_2729_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1495 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1496 a_7130_n8125# a_6874_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1497 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1498 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1499 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1500 a_8229_n4709# a_8328_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1501 a_4365_n12325# a_4464_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1502 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1503 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1504 a_6941_n13413# a_7040_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1505 a_1978_n11933# a_1722_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1506 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X1507 sky130_fd_sc_hd__nand2_4_3/A clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1508 VDD a_4554_n9213# a_4661_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1509 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1510 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1511 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1512 VSS a_8418_n14109# a_8525_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1513 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1514 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1515 a_10805_n3621# a_10904_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1516 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1517 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1518 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9450_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1519 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1520 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkinv_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1521 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1522 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1523 VSS a_2148_n9783# a_1888_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1524 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1525 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1526 a_8418_n8125# a_8162_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1527 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1528 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1529 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1530 VSS a_9706_n509# a_9813_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1531 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1532 a_501_n5797# a_600_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1533 VSS a_1978_n13021# a_2085_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1534 a_1789_n12325# a_1888_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1535 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1536 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1537 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1538 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1539 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1540 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1541 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_2085_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1542 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1543 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1544 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1545 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1546 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1547 VDD a_7130_n1597# a_7237_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1548 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5586_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1549 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1550 VSS sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1551 VSS a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1552 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1553 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1554 VSS a_7300_n12503# a_7040_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1555 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1556 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1557 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1558 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1559 VSS sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1560 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1561 VSS a_11164_n3255# a_10904_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1562 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1563 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_42/X a_434_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1564 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1565 VSS a_2148_n13591# a_1888_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1566 VSS a_6012_n11415# a_5752_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1567 a_5842_n4317# a_5586_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1568 VSS a_8418_n509# a_8525_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1569 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10738_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1570 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1571 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1572 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1573 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1574 VDD a_5842_n5405# a_5949_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1575 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4298_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1576 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1577 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1578 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1579 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1580 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1581 a_501_n4709# a_600_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1582 VDD a_8418_n5405# a_8525_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1583 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1585 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1586 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_4661_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1587 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5586_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1588 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1589 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1590 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1591 VDD sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1592 VDD a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1593 a_9517_n2997# a_9616_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1594 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1595 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1596 VSS a_3266_n10301# a_3373_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1597 a_10994_n9213# a_10738_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1598 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1599 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/X a_434_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1600 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1601 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3010_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1602 VSS a_10805_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1603 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1604 VSS a_11164_n2167# a_10904_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1605 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1606 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1607 VDD a_5842_n2685# a_5949_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1608 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1610 a_7130_n11933# a_6874_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1611 a_8229_n10613# a_8328_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1612 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1613 VDD a_4365_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1614 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1615 VDD a_11164_n9783# a_10904_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1616 VSS sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1617 VSS sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1618 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1619 VDD a_8418_n2685# a_8525_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1620 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1621 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1622 a_7014_n7215# a_6794_n7203# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1623 VSS a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1624 VDD a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1625 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1626 a_501_n13413# a_600_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1627 a_501_n9525# a_600_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1628 sky130_fd_sc_hd__nand2_4_3/B a_9813_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1629 a_7130_n2685# a_6874_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1630 VDD a_3266_n5405# a_3373_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1631 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1632 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1633 VDD a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1634 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1635 a_9517_n1909# a_9616_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1636 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1637 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1638 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1639 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1640 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1641 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1642 a_9517_n9525# a_9616_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1643 VSS a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1644 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_7237_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1645 VDD sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1646 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1647 VDD a_2148_n8695# a_1888_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1648 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_797_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1649 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9450_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1650 VDD sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1651 VSS a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1652 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1653 a_6012_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1654 VDD a_1978_n11933# a_2085_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1655 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1656 VSS a_7300_n5975# a_7040_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1657 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1658 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1659 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1660 VSS a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1661 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1662 a_1789_n821# a_1888_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1663 VDD a_3266_n2685# a_3373_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1664 VDD a_2622_n6493# a_2729_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1665 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1666 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1667 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1668 a_5653_n5797# a_5752_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1669 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1670 VSS a_9876_n5975# a_9616_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1671 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1672 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8162_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1673 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1674 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1675 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1676 a_6941_n2997# a_7040_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1677 VDD a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1678 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1679 a_3266_n4317# a_3010_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1680 VSS a_6941_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1681 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1682 VDD a_3436_n11415# a_3176_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1683 VSS a_690_n2685# a_797_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1684 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1685 a_4554_n2685# a_4298_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1686 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1687 a_5842_n9213# a_5586_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1688 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1689 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1690 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_1_6/Y a_n860_n13789# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1691 VSS a_501_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1692 VSS a_7300_n4887# a_7040_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1693 VDD a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1694 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1695 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1696 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1697 VSS a_3436_n10871# a_3176_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1698 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_7237_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1699 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1700 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1701 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1702 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1703 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1704 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1705 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1706 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_8525_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1707 VSS a_6658_n7363# a_6665_n7459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1708 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3010_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1709 VSS a_9876_n4887# a_9616_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1710 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_7237_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1711 a_11164_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1712 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1713 a_7130_n6493# a_6874_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1714 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9813_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1715 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_8525_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1716 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1717 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8162_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1718 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1719 VSS a_4724_n5975# a_4464_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1720 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_1_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1721 a_6941_n1909# a_7040_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1722 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1723 sky130_fd_sc_hd__clkinv_1_5/A a_n1570_n6769# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1724 a_10994_n10301# a_10738_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1725 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1726 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1727 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1728 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1729 VDD a_6012_n3799# a_5752_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1730 VSS a_6941_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1731 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1732 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1733 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1734 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1735 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1736 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1737 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1738 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1739 VSS a_n428_n12503# a_n688_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1740 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1741 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1742 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1743 VDD a_860_n3255# a_600_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1744 VDD a_8588_n3799# a_8328_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1745 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1746 a_501_n8437# a_600_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1747 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1748 a_690_n1597# a_434_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1749 a_4365_n2997# a_4464_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1750 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10738_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1751 VSS a_7300_n9783# a_7040_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1752 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1753 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1754 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1755 VSS a_1978_n4317# a_2085_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1756 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1757 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1758 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1759 a_8418_n9213# a_8162_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1760 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1761 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1762 a_6941_n3621# a_7040_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1763 a_9706_n13021# a_9450_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1764 a_1978_n2685# a_1722_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1765 VSS a_9876_n9783# a_9616_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1766 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1767 VSS a_8418_n10301# a_8525_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1768 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1769 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1770 VSS a_4724_n4887# a_4464_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1771 a_8418_n11933# a_8162_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1772 VDD a_6941_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1773 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1774 VSS a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1775 a_9876_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1776 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1777 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1778 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1779 VDD a_1789_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1780 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1781 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1782 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1783 VDD a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1784 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1785 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1786 a_9517_n13413# a_9616_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1787 VSS a_10994_n1597# a_11101_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1788 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1789 VDD a_860_n2167# a_600_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1790 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1791 a_3077_n10613# a_3176_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1792 a_11164_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1793 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1794 a_4365_n1909# a_4464_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1795 a_8229_n12325# a_8328_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1796 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1797 VDD a_3436_n3799# a_3176_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1798 VSS sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1799 a_10805_n11237# a_10904_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1800 VSS sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1801 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6874_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1802 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1803 VDD a_9706_n6493# a_9813_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1804 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6874_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1805 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1806 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1807 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1808 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1809 VDD a_3266_n13021# a_3373_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1810 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1811 a_6941_n8437# a_7040_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1812 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1813 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1814 a_7300_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1815 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1816 VDD a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1817 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1818 VDD a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1819 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1820 VSS a_6941_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1821 a_1789_n2997# a_1888_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1822 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1823 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1824 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1825 VSS a_4724_n9783# a_4464_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1826 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1827 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1828 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_5949_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1829 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1830 a_9706_n1597# a_9450_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1831 VDD a_4724_n10871# a_4464_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1832 VSS a_860_n3799# a_600_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1833 VSS a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1834 a_4365_n3621# a_4464_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1835 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1836 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1837 VSS sky130_fd_sc_hd__nand2_4_1/B a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1838 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1839 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1840 sky130_fd_sc_hd__nand2_4_0/B a_9813_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1841 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1842 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1843 VSS a_3077_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1844 VDD a_860_n10871# a_600_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1845 VSS a_2622_n14109# a_2729_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1846 VDD a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1847 a_690_n5405# a_434_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1848 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1849 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6874_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1850 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1851 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1852 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1853 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=0p ps=0u w=840000u l=150000u
X1854 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1855 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1856 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1857 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1858 VDD a_6941_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1859 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1860 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1861 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1862 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_797_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1863 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1864 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1865 a_1789_n1909# a_1888_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1866 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1867 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1868 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1869 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1870 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1871 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1872 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10738_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1873 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1874 VDD sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1875 VDD a_8588_n11415# a_8328_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1876 VDD a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1877 VDD a_2148_n5975# a_1888_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1878 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1879 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1880 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1881 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1882 VSS a_860_n8695# a_600_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1883 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1884 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1885 a_4365_n8437# a_4464_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1886 VDD a_7300_n8695# a_7040_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1887 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1888 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1889 VSS a_7130_n1597# a_7237_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1890 VSS a_10994_n5405# a_11101_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1891 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1892 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1893 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1894 VSS a_8588_n10871# a_8328_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1895 VDD a_11164_n1079# a_10904_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1896 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1897 a_9706_n11933# a_9450_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1898 VSS a_7130_n11933# a_7237_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1899 VDD sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_4_1/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1900 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1901 VDD a_9876_n8695# a_9616_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1902 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_11101_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1903 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1904 VSS a_1978_n9213# a_2085_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1905 a_1789_n3621# a_1888_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1906 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5586_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1907 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1908 VDD a_n1570_n6769# a_n1654_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X1909 VDD sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1910 VDD a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1911 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1912 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1913 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1914 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1915 VDD a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1916 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1917 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1918 a_3266_n1597# a_3010_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1919 a_6012_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1920 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_434_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1921 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1922 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8162_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1923 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_3373_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1924 a_9706_n5405# a_9450_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1925 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1926 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1927 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1928 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1929 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1930 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1931 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1932 a_9517_n821# a_9616_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1933 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1934 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1935 a_n1612_n7037# a_n2602_n7037# a_n1738_n6671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X1936 a_1789_n13413# a_1888_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1937 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1938 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10738_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1939 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1940 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1941 VSS a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1942 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1943 VDD a_8418_n14109# a_8525_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1944 VSS clk sky130_fd_sc_hd__clkinv_1_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1945 VSS a_9876_n1079# a_9616_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1946 a_1789_n8437# a_1888_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1947 VDD a_7300_n13591# a_7040_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1948 VDD a_4724_n8695# a_4464_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1949 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1950 a_10994_n13021# a_10738_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1951 a_7130_n10301# a_6874_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1952 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1953 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1954 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1955 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1956 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1957 a_4554_n13021# a_4298_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1958 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1959 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1960 a_6012_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1961 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1962 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1963 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1964 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1965 a_10805_n2997# a_10904_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1966 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1967 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1968 VDD sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1969 a_3266_n11933# a_3010_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1970 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1971 a_690_n13021# a_434_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1972 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1973 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1974 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1975 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1976 VDD sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1977 VSS a_8588_n1079# a_8328_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1978 VSS a_7130_n5405# a_7237_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1979 VDD a_9706_n509# a_9813_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1980 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1981 a_501_n5797# a_600_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1982 a_1789_n12325# a_1888_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1983 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1984 a_8229_n5797# a_8328_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1985 a_4365_n13413# a_4464_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1986 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1987 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_5949_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1988 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_7237_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1989 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1990 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1991 VDD a_8418_n13021# a_8525_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1992 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1993 a_5842_n4317# a_5586_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1994 VDD a_7300_n12503# a_7040_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1995 a_3077_n12325# a_3176_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1996 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1997 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6874_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1998 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/A a_n860_n509# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1999 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A a_11101_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2000 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2001 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2002 VSS a_4554_n11933# a_4661_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2003 VDD a_11164_n10871# a_10904_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2004 VDD a_1978_n10301# a_2085_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2005 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2006 VSS a_860_n1079# a_600_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2007 VSS a_9706_n4317# a_9813_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2008 VDD a_9876_n10871# a_9616_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2009 VDD a_8418_n509# a_8525_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2010 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2011 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2012 a_10805_n1909# a_10904_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2013 VDD a_8418_n8125# a_8525_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2014 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2015 VSS a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2016 VSS a_690_n11933# a_797_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2017 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2018 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2019 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2020 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2021 a_5842_n10301# a_5586_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2022 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2023 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2024 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2025 a_3077_n2997# a_3176_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2026 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2027 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2028 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2029 VSS a_4724_n12503# a_4464_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2030 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_5949_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2031 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_8525_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2032 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2033 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2034 a_8229_n4709# a_8328_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2035 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_434_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2036 VDD sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2037 VSS a_7300_n1079# a_7040_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2038 VDD a_6658_n7363# a_6665_n7459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2039 VSS sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2040 VSS a_3436_n11415# a_3176_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2041 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8162_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2042 VSS a_860_n12503# a_600_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2043 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2044 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_797_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2045 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_2085_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2046 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2047 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2048 a_10805_n3621# a_10904_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2049 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2050 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1722_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2051 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_5949_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2052 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2053 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2054 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2055 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2056 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_1_4/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2057 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_2729_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2058 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2059 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2060 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2061 VSS a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2062 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2063 VDD a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2064 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_4661_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2065 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2067 VSS a_6012_n1079# a_5752_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2068 VSS a_4554_n4317# a_4661_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2069 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2070 VDD a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2071 VDD sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 a_3077_n1909# a_3176_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2073 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2074 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2075 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2076 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2077 a_3077_n9525# a_3176_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2078 a_4765_n7542# sky130_fd_sc_hd__dfxbp_1_0/Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2079 a_8229_n9525# a_8328_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2080 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_797_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2081 a_4554_n11933# a_4298_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2082 VDD a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2083 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2084 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2085 a_4765_n7215# sky130_fd_sc_hd__dfxbp_1_0/Q VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2086 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 a_6012_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2088 a_10805_n8437# a_10904_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2089 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2090 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2091 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2092 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2093 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2094 a_690_n11933# a_434_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2095 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2096 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2097 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2098 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2099 VSS a_3077_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2100 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8162_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2101 VSS a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2102 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2103 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2104 VDD a_7300_n5975# a_7040_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2105 a_6593_n7215# a_6101_n7254# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X2106 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2107 a_4623_n7349# Ad_b a_4765_n7542# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X2108 a_690_n5405# a_434_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2109 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2110 a_8418_n6493# a_8162_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2111 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2112 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2113 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2114 a_5653_n11237# a_5752_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2115 VDD a_9876_n5975# a_9616_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2116 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2117 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2118 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2119 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2120 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2121 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2122 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2123 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2124 VSS a_5842_n2685# a_5949_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2125 VSS a_1789_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2126 a_5653_n10613# a_5752_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2127 VDD sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2128 VDD sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__nand2_4_2/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2129 VDD a_3077_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2130 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2131 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2132 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2133 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2134 VDD a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2135 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2136 VSS a_8418_n2685# a_8525_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2137 VDD a_8229_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2138 a_10994_n4317# a_10738_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2139 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2140 VSS a_9706_n9213# a_9813_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2141 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2142 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2143 a_690_n2685# a_434_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2144 VDD a_10994_n5405# a_11101_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2145 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2146 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2147 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2148 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2149 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2150 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2151 VDD sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2152 a_5082_n7542# Bd_b a_4623_n7349# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2153 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2154 VSS sky130_fd_sc_hd__clkinv_1_3/Y a_2366_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2155 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2156 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2157 a_6941_n4709# a_7040_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2158 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2159 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2160 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2161 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2162 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4298_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2163 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2164 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3010_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2165 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2166 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2167 VSS a_5052_n7283# a_4986_n7215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2168 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2169 a_8588_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2170 VDD a_4724_n5975# a_4464_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2171 VSS a_10994_n11933# a_11101_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2172 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2173 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2174 VSS a_9706_n11933# a_9813_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2175 VSS sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2176 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2177 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2178 VDD a_6012_n3255# a_5752_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2179 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11101_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2180 a_9706_n5405# a_9450_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2181 VDD a_n428_n12503# a_n688_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2182 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5586_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2183 VDD a_1978_n4317# a_2085_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2184 a_7130_n8125# a_6874_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2185 VDD a_10994_n2685# a_11101_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2186 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_4661_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2187 VDD a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2188 a_4986_n7215# Ad_b a_4623_n7349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X2189 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2190 VDD a_8588_n3255# a_8328_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2191 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2192 VSS a_11164_n12503# a_10904_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2193 VSS a_4554_n9213# a_4661_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2194 VSS a_3266_n2685# a_3373_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2195 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2196 a_8229_n13413# a_8328_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2197 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2198 a_8229_n8437# a_8328_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2199 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2200 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2201 VSS a_9876_n12503# a_9616_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2202 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2203 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2204 VSS a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2205 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2206 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3010_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2207 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2208 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2209 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2210 VSS a_8588_n11415# a_8328_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2211 VDD a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2212 a_10805_n821# a_10904_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2213 VDD a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2214 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2215 a_5842_n1597# a_5586_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2216 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2217 a_7130_n14109# a_6874_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2218 sky130_fd_sc_hd__nand2_4_1/B a_9813_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2219 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2220 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2221 VDD sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2222 a_9706_n2685# a_9450_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2223 VSS a_8229_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2224 VDD a_860_n4887# a_600_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2225 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2226 VDD a_6012_n2167# a_5752_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2227 VDD sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2228 a_4365_n4709# a_4464_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2229 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 a_5842_n13021# a_5586_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2231 a_9706_n10301# a_9450_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2232 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1722_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2233 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2234 VSS a_8418_n6493# a_8525_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2235 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2236 VDD a_7130_n5405# a_7237_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2237 VDD a_8588_n2167# a_8328_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2238 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2239 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2240 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2241 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2242 a_8229_n12325# a_8328_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2243 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2244 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2245 VDD a_3436_n3255# a_3176_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2246 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2247 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 a_3266_n1597# a_3010_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2249 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2250 a_6616_n7581# a_6101_n7254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2251 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2252 VDD a_5653_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2253 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2254 a_6101_n7254# a_6373_n7349# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2255 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2256 VSS a_6012_n3799# a_5752_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2257 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8162_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2258 VDD a_8229_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2259 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2260 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2261 VSS a_9517_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2262 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2263 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2264 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2265 VDD a_3077_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2266 VDD a_2622_n14109# a_2729_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2267 VDD a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2268 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2269 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7237_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2270 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2271 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2272 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2273 VSS a_8588_n3799# a_8328_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2274 VDD a_7130_n2685# a_7237_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2275 VSS a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2276 a_11164_n13591# sky130_fd_sc_hd__clkinv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2277 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2278 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8525_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2279 VSS sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2280 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2281 a_10994_n9213# a_10738_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2282 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2283 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2284 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2285 VDD a_5052_n7283# a_5082_n7542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 VDD a_6012_n10871# a_5752_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2287 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2288 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2289 VSS a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2290 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2291 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8162_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2292 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2293 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2294 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2295 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9450_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2296 sky130_fd_sc_hd__nand2_4_3/B a_9813_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2297 a_1789_n4709# a_1888_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2298 VDD a_3436_n2167# a_3176_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2299 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2300 VSS sky130_fd_sc_hd__nand2_4_3/B a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2301 a_n1738_n6671# a_n2436_n7037# a_n1995_n6925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2302 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2303 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2304 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2305 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2306 VDD a_9517_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2307 VSS a_6012_n8695# a_5752_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2308 a_8418_n4317# a_8162_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2309 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2310 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2311 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2312 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2313 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2314 a_5653_n2997# a_5752_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2315 VDD a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2316 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2317 VDD sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2318 VDD a_11164_n3799# a_10904_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2319 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2320 a_11164_n13591# sky130_fd_sc_hd__clkinv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2321 VSS a_8588_n8695# a_8328_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2322 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2323 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2324 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2325 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8525_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2327 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2328 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_2085_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2329 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2330 VSS a_3436_n3799# a_3176_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2331 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2332 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2333 VDD a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2334 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8162_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2335 VSS a_8229_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2336 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2337 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2338 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2340 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2341 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2342 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2343 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_4661_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2344 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2345 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9813_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2346 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2347 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_8525_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2348 a_3266_n5405# a_3010_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2349 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2350 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2351 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2352 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2353 a_3077_n821# a_3176_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2354 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2355 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2356 a_9517_n3621# a_9616_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2357 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2358 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2359 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2360 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2361 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6874_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2362 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2363 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2364 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2365 a_5653_n1909# a_5752_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2366 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2367 a_6658_n7363# p2 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2368 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2369 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2370 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2371 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2372 a_5653_n9525# a_5752_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2373 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11101_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2374 VSS a_3436_n8695# a_3176_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2375 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2376 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2377 VDD a_n1738_n6671# a_n1570_n6769# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2378 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2379 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2380 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2381 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2382 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2383 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 a_3077_n13413# a_3176_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2385 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2386 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2387 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2388 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2389 VSS sky130_fd_sc_hd__nand2_4_0/B a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2390 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2391 VSS sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2392 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2393 VSS a_11164_n1079# a_10904_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2394 VSS a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2395 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2396 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2397 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2398 VSS a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2399 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2400 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2401 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2402 VDD a_1978_n1597# a_2085_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2403 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2404 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2405 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2406 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2407 VSS sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2408 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2409 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2410 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2411 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2412 VDD a_4724_n13591# a_4464_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2413 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2414 a_7130_n9213# a_6874_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2415 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2416 a_8229_n5797# a_8328_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2417 VDD a_10805_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2418 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2419 a_4554_n10301# a_4298_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2420 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2421 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2422 a_4623_n7349# Bd_b a_4765_n7215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2423 VSS a_6101_n7254# sky130_fd_sc_hd__dfxbp_1_0/Q VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2424 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2425 a_1978_n13021# a_1722_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2426 VDD a_860_n13591# a_600_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2427 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2428 VDD a_9706_n4317# a_9813_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2429 a_3077_n12325# a_3176_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2430 VSS a_7130_n509# a_7237_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2431 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2432 a_690_n10301# a_434_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2433 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2434 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2435 a_10805_n4709# a_10904_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2436 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2437 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2438 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2439 VDD a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2440 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2441 a_9706_n509# a_9450_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2442 VDD a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2443 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2444 a_8418_n9213# a_8162_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2445 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2446 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2447 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8162_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2448 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2449 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2450 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2451 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2452 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2453 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4298_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2454 a_1789_n13413# a_1888_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2455 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2456 VSS a_5842_n11933# a_5949_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2457 a_5653_n11237# a_5752_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2458 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2459 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2460 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2461 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2462 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2463 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7237_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2464 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2465 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5586_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2466 VDD a_4724_n12503# a_4464_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2467 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 VSS a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2469 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2470 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2471 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2472 VSS a_7300_n13591# a_7040_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2473 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_797_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2474 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9450_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2475 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2476 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2477 a_7130_n10301# a_6874_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2478 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2479 a_8418_n509# a_8162_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2480 VDD a_860_n12503# a_600_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2481 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2482 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2483 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2484 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2485 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_434_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2486 a_2622_n8125# a_2366_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2487 VSS a_6012_n12503# a_5752_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2488 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_2085_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2489 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10738_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2490 VDD a_690_n9213# a_797_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2491 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2492 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2493 VDD a_4554_n4317# a_4661_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2494 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2495 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2496 a_4554_n9213# a_4298_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2497 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A a_11101_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2498 VDD a_6865_n7304# a_6794_n7203# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2499 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2500 VDD sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2501 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2502 VDD sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2503 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3010_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2504 a_9706_n14109# a_9450_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2505 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8162_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2506 VDD sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2507 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2508 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2509 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2510 VSS a_6006_n7607# sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2511 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2512 a_11164_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2513 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5586_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2514 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2515 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2516 VDD a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2517 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2518 a_n787_n1909# a_n688_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2519 VDD a_501_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2520 VDD a_6941_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2521 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2522 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2523 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2524 VSS a_2148_n3255# a_1888_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2525 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_2085_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2526 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2527 VSS a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2528 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2529 a_n787_n9525# a_n688_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2530 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2531 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_434_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2532 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1722_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2533 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2534 VSS a_2622_n509# a_2729_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2535 VSS a_10805_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2536 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2537 VSS a_1978_n10301# a_2085_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2538 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_4661_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2539 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2540 VDD a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2541 a_10805_n10613# a_10904_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2542 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_3373_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2543 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2544 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2545 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2546 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2547 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2548 a_9876_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2549 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2551 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2552 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2553 VSS a_4623_n7349# sky130_fd_sc_hd__mux2_1_0/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2554 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2555 VDD a_n428_n2167# a_n688_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2556 a_5842_n1597# a_5586_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2557 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2558 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9813_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2559 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_11101_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2560 a_1978_n11933# a_1722_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2561 VDD a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2562 a_1978_n9213# a_1722_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2563 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2565 VDD a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2566 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2567 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2568 VSS a_2148_n2167# a_1888_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2569 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2570 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2571 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2572 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2574 VDD a_2148_n9783# a_1888_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2575 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2576 a_10994_n4317# a_10738_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2577 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2578 VSS sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2579 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2580 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2581 a_6941_n11237# a_7040_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2582 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_7237_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2583 a_n428_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2584 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2585 a_6794_n7203# a_6665_n7459# a_6373_n7349# VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X2586 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2587 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2588 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2589 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2590 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2591 VSS a_501_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2592 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2366_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2593 VDD a_11164_n13591# a_10904_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2594 a_6941_n10613# a_7040_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2595 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2596 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2597 VDD a_9876_n13591# a_9616_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2598 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2599 a_11164_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2600 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2601 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2602 a_9876_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2603 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X2604 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_2729_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2605 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2606 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2607 a_3266_n5405# a_3010_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2608 a_n1654_n6671# a_n2436_n7037# a_n1738_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2609 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2610 a_9706_n8125# a_9450_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2611 VSS sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2612 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2613 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2614 a_501_n2997# a_600_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2615 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2616 a_n428_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2617 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2618 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2619 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2620 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2621 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2622 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2623 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_2729_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2624 VDD a_2148_n11415# a_1888_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2625 a_5052_n7283# sky130_fd_sc_hd__dfxbp_1_0/Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2626 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2627 VDD a_501_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2628 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_2085_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2629 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2630 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2631 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2632 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2633 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2634 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2635 VDD a_11164_n12503# a_10904_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2636 VSS sky130_fd_sc_hd__clkinv_1_0/Y a_2366_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2637 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2638 a_6941_n5797# a_7040_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2639 a_5052_n7283# sky130_fd_sc_hd__dfxbp_1_0/Q VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2640 VDD a_9876_n12503# a_9616_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2641 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_434_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2642 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4298_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2643 a_5842_n5405# a_5586_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2644 a_7130_n14109# a_6874_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2645 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_7237_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2646 VSS sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2647 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2648 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_4661_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2649 VSS a_2148_n10871# a_1888_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2650 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_9813_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2651 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_5949_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2652 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2653 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8525_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2654 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2655 a_3266_n2685# a_3010_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2656 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8162_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2657 a_5653_n821# a_5752_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2658 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2659 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2660 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2661 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2662 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2663 VDD a_9706_n1597# a_9813_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2664 VSS sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2665 VDD a_6012_n4887# a_5752_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2666 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2667 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_7237_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2668 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2669 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2670 a_501_n1909# a_600_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2671 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2672 VDD a_7130_n8125# a_7237_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2673 VDD a_8588_n4887# a_8328_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2674 a_6658_n7363# p2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2675 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2676 a_501_n9525# a_600_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2677 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2678 a_690_n2685# a_434_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2679 VSS sky130_fd_sc_hd__nand2_4_2/B a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2680 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2681 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2682 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2683 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2684 a_n860_n13789# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2685 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2686 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2687 a_5653_n821# a_5752_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2688 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2689 a_6941_n4709# a_7040_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2690 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2691 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2692 a_7300_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2693 a_7130_n13021# a_6874_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2694 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2695 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2696 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2697 a_501_n11237# a_600_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2698 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_2085_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2699 a_8418_n13021# a_8162_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2700 VSS a_8418_n8125# a_8525_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2701 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2702 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2703 VSS a_501_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2704 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2705 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2706 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_2729_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2707 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2708 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2709 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2710 VSS a_860_n5975# a_600_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2711 a_2622_n6493# a_2366_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2712 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2713 a_4365_n5797# a_4464_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2714 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2715 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1722_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2716 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_3373_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2717 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_4661_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2718 VDD a_4554_n1597# a_4661_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2719 a_501_n10613# a_600_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2720 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2721 VSS a_10994_n2685# a_11101_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2722 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2723 a_4365_n821# a_4464_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2724 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2725 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2726 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2727 a_8229_n13413# a_8328_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2728 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2729 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2730 VDD a_3436_n4887# a_3176_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2731 a_10805_n12325# a_10904_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2732 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2733 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2734 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2735 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2736 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2737 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2738 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2739 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2740 a_6941_n9525# a_7040_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2741 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2742 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2743 a_8418_n4317# a_8162_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2744 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2745 VDD a_10805_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2746 VSS a_6941_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2747 VSS sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2748 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2749 VSS a_n787_n4709# sky130_fd_sc_hd__nand2_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2750 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/A a_2366_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2751 VDD a_1978_n13021# a_2085_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2752 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2753 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2754 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2755 a_3077_n821# a_3176_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2756 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11101_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2757 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2758 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2759 a_9706_n2685# a_9450_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2760 VSS a_7300_n3255# a_7040_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2761 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2762 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2763 VSS a_1978_n1597# a_2085_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2764 VSS a_860_n4887# a_600_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2765 VSS a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2766 a_4365_n4709# a_4464_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2767 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2768 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2769 a_860_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2770 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2771 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2772 a_9706_n10301# a_9450_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2773 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2774 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4298_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2775 VDD a_3436_n10871# a_3176_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2776 VSS a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2777 VDD a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2778 VSS a_9876_n3255# a_9616_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2779 VDD a_11164_n3255# a_10904_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2780 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2781 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2782 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2783 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2784 a_7130_n6493# a_6874_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2785 a_1789_n5797# a_1888_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2786 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2787 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2366_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2788 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2789 a_3077_n3621# a_3176_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2790 VDD a_6941_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2791 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2792 VDD a_n787_n4709# sky130_fd_sc_hd__nand2_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2793 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11101_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2794 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2795 a_11164_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2796 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2797 VDD a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2798 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2799 VSS a_7300_n2167# a_7040_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2800 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2801 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2802 a_860_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2803 VSS a_860_n9783# a_600_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2804 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2805 a_10994_n1597# a_10738_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2806 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_2729_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2807 a_4365_n9525# a_4464_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2808 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2809 a_9517_n2997# a_9616_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2810 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5586_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2811 VDD a_7300_n9783# a_7040_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2812 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2813 VSS a_7130_n2685# a_7237_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2814 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2815 VDD a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2816 VSS a_9876_n2167# a_9616_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2817 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2818 VDD a_4365_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2819 VDD a_11164_n2167# a_10904_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2820 VSS a_7130_n13021# a_7237_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2821 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2822 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2823 VSS a_4724_n3255# a_4464_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2824 VDD a_9876_n9783# a_9616_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2825 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2826 VDD sky130_fd_sc_hd__clkinv_1_3/Y a_2366_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2827 VDD sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2828 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2829 a_1789_n4709# a_1888_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2830 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2831 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2832 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_10738_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2833 a_8418_n11933# a_8162_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2834 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4298_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2835 VSS sky130_fd_sc_hd__clkinv_1_5/A a_7212_n7203# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2836 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2837 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2838 VSS a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2839 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_1722_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2840 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2841 VDD a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2842 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2843 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2844 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2845 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2846 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7237_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2847 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_8525_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2848 a_9706_n6493# a_9450_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2849 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_3373_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2850 VSS sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_9813_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2852 VSS a_1978_n5405# a_2085_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2853 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2854 VSS a_11164_n3799# a_10904_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2855 a_9517_n1909# a_9616_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2856 VDD a_2148_n1079# a_1888_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2857 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2858 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2859 VSS sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2860 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2861 a_9517_n821# a_9616_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2862 a_6941_n8437# a_7040_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2863 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2864 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2865 a_9517_n11237# a_9616_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2866 VSS a_4724_n2167# a_4464_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2867 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2868 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2869 a_1789_n9525# a_1888_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2870 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2871 VDD a_4724_n9783# a_4464_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2872 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2873 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2874 VSS a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2875 VDD a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2876 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2877 VDD a_7130_n509# a_7237_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2878 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2879 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2880 VDD a_6012_n13591# a_5752_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2881 a_9517_n10613# a_9616_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2882 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7237_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2883 a_7300_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2884 a_9517_n3621# a_9616_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2885 VDD sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2886 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2887 sky130_fd_sc_hd__dfxbp_1_1/D a_n1139_n6715# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2888 VSS a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2889 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2890 a_n2068_n6671# a_n2602_n7037# a_n2163_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2891 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2892 a_8229_n821# a_8328_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2893 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2894 VSS a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2895 a_3266_n13021# a_3010_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2896 a_9706_n509# a_9450_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2897 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_2085_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2898 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2899 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2900 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2901 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2902 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1722_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2903 VSS a_11164_n8695# a_10904_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2904 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2905 VSS a_7130_n6493# a_7237_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2906 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2907 a_1978_n10301# a_1722_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2908 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2909 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2910 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_4661_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2911 a_5842_n5405# a_5586_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2912 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2913 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2914 a_3077_n13413# a_3176_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2915 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2916 a_6941_n11237# a_7040_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2917 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2918 a_10805_n5797# a_10904_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2919 VDD a_5842_n9213# a_5949_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2920 a_501_n821# a_600_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2921 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2922 a_9876_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2923 a_8418_n509# a_8162_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2924 a_8588_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2925 VSS a_4554_n13021# a_4661_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2926 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2927 VDD a_860_n8695# a_600_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2928 a_6006_n7607# a_6101_n7254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2929 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2930 VDD a_6012_n12503# a_5752_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2931 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2932 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2933 a_4365_n8437# a_4464_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2934 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_9450_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2935 a_9517_n8437# a_9616_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2936 a_9706_n14109# a_9450_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2937 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2938 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2939 VSS a_3266_n11933# a_3373_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2940 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_2085_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2941 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2942 VSS a_690_n13021# a_797_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2943 VSS a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2944 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2945 VDD a_8418_n9213# a_8525_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2946 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2947 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2948 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2949 VDD a_8588_n10871# a_8328_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2950 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2951 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2952 VDD a_1789_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2953 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2954 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2955 VDD a_7130_n11933# a_7237_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2956 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2957 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11101_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2958 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2959 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2960 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2961 VSS a_4724_n13591# a_4464_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2962 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2963 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_4661_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2964 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2965 VSS a_6865_n7304# a_6794_n7203# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2966 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_434_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2967 a_4554_n10301# a_4298_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2968 a_7300_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2969 a_5842_n2685# a_5586_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2970 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2971 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2972 VSS sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2973 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2974 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9450_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2975 a_501_n821# a_600_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2976 VSS a_4365_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2977 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2978 VSS a_5653_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2979 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2980 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2981 VDD sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2982 VSS a_3436_n12503# a_3176_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2983 VSS a_860_n13591# a_600_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2984 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2985 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2986 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2987 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2988 a_690_n10301# a_434_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2989 a_8418_n1597# a_8162_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2990 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2991 a_10805_n4709# a_10904_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2992 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2993 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2994 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2995 VDD a_2622_n509# a_2729_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2996 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2997 VSS a_2148_n11415# a_1888_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2998 VSS a_6941_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2999 a_7130_n4317# a_6874_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3000 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3001 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3002 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3003 VDD a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3004 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3005 a_9706_n13021# a_9450_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3006 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3007 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3008 a_6012_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3009 VDD a_n428_n4887# a_n688_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3010 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3011 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3012 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X3013 VDD a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3014 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3015 VDD a_3266_n9213# a_3373_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3016 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3017 VDD sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3018 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3019 a_8588_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3020 a_1789_n8437# a_1888_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3021 VSS sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_1_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3022 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3023 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3024 VSS a_9706_n1597# a_9813_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3025 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3026 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3027 VSS a_5653_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3028 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_3373_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3029 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3030 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3031 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3032 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3033 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3034 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3035 a_10805_n9525# a_10904_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3036 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3037 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3038 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3039 a_3266_n11933# a_3010_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3040 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3041 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3042 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3043 VSS a_1789_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3044 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4298_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3045 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3046 sky130_fd_sc_hd__clkinv_1_5/A a_n1570_n6769# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3047 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6874_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3048 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3049 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3050 VDD a_10805_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3051 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3052 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3053 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3054 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3056 VSS a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3057 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X3058 a_6373_n7349# a_6658_n7363# a_6593_n7215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3059 VSS a_4365_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3060 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3061 VSS a_690_n4317# a_797_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3062 VDD sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3063 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3064 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_9813_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3065 a_501_n11237# a_600_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3066 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3067 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3068 a_4554_n4317# a_4298_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3069 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3070 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3071 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3072 VDD a_9517_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3073 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3074 VDD a_4554_n11933# a_4661_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3075 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3076 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3077 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3078 a_4365_n11237# a_4464_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3079 VSS a_4554_n1597# a_4661_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3080 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3081 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3082 VDD a_690_n11933# a_797_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3083 VDD a_1789_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3084 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3085 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4298_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3086 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3087 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3088 a_860_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3089 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3090 VSS sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3091 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3092 VDD a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3093 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3094 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3095 a_4365_n10613# a_4464_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3096 a_8229_n2997# a_8328_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3097 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3098 a_10994_n11933# a_10738_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3099 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3100 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3101 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3102 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3103 a_n787_n12325# a_n688_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3104 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3105 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3106 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3107 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3108 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3109 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3110 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3111 VDD a_7300_n1079# a_7040_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3112 a_5653_n3621# a_5752_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3113 a_3436_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3114 a_6941_n5797# a_7040_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3115 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3116 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1722_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3117 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3118 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3119 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3120 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3121 VSS a_9706_n5405# a_9813_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3122 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3123 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3124 VSS a_10805_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3125 VSS a_10994_n13021# a_11101_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3126 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3127 VSS sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3128 VDD a_9876_n1079# a_9616_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3129 VSS a_9706_n13021# a_9813_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3130 VSS a_8229_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3131 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_2085_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3132 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3133 a_1978_n4317# a_1722_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3134 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3135 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3136 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3137 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3138 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A a_11101_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3139 VSS a_8418_n11933# a_8525_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3140 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_5586_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3141 a_7130_n9213# a_6874_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3142 VSS sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3143 VDD a_1978_n5405# a_2085_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3144 VDD a_6941_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3145 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3146 a_8229_n1909# a_8328_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3147 VSS a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3148 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3149 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3150 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4298_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3151 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3152 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3153 VSS a_11164_n13591# a_10904_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3154 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3155 a_8229_n9525# a_8328_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3156 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3157 VSS a_9876_n13591# a_9616_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3158 VSS sky130_fd_sc_hd__nand2_4_1/B a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3159 a_10805_n13413# a_10904_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3160 a_3436_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3161 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1722_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3162 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3163 VSS a_1789_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3164 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3165 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3166 VSS a_8588_n12503# a_8328_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3167 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3168 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3169 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X3170 VSS sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3171 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_4661_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3172 VDD a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3173 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3174 a_10805_n8437# a_10904_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3175 a_10994_n1597# a_10738_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3176 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3177 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3178 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3179 VSS a_6012_n5975# a_5752_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3180 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3181 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3182 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3183 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3184 VSS a_4554_n5405# a_4661_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3185 VSS a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3186 VDD a_1978_n2685# a_2085_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3187 VDD a_860_n5975# a_600_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3188 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3189 VDD a_4724_n1079# a_4464_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3190 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9813_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3191 VDD sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3192 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3193 a_4365_n5797# a_4464_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3194 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3195 VSS a_8588_n5975# a_8328_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3196 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3197 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3198 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3199 VSS a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3200 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3201 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3202 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3203 a_4554_n13021# a_4298_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3204 a_8418_n10301# a_8162_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3205 VSS a_5653_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3206 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3207 a_2622_n8125# a_2366_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3208 a_10805_n12325# a_10904_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3209 VSS a_690_n9213# a_797_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3210 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3211 a_3266_n2685# a_3010_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3212 a_690_n13021# a_434_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3213 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3214 a_4554_n9213# a_4298_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3215 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3216 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3217 VSS a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3218 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3219 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3220 a_5653_n10613# a_5752_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3221 VSS a_6012_n4887# a_5752_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3222 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3223 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3224 VSS a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3225 VDD a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3226 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_3373_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3227 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3228 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3229 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3230 VDD a_3077_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3231 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3232 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3233 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_7237_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3234 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3235 VSS a_8588_n4887# a_8328_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3236 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3237 a_9517_n11237# a_9616_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3238 a_9876_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3239 VSS a_8229_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3240 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3241 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3242 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3243 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3244 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3245 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3246 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3247 VSS a_3436_n5975# a_3176_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3248 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3249 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3250 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_9813_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3251 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_8525_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3252 VSS a_5653_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3253 a_9876_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3254 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3255 VDD a_n1995_n6925# a_n2068_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3256 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_9450_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3257 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9813_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3258 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 a_1789_n5797# a_1888_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3260 a_7212_n7203# a_6665_n7459# a_6865_n7304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3261 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3262 VDD a_10994_n11933# a_11101_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3263 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3264 VSS sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3265 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3266 VDD a_9706_n11933# a_9813_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3267 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3268 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3269 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3270 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3271 a_3077_n2997# a_3176_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3272 a_10994_n5405# a_10738_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3273 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3274 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3275 VSS a_6012_n9783# a_5752_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3276 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3277 VSS a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3278 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3279 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3280 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3281 VDD a_8229_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3282 VDD a_11164_n4887# a_10904_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3283 a_1978_n9213# a_1722_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3284 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3285 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3286 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3287 VSS a_8588_n9783# a_8328_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3288 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3289 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3290 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3291 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3292 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3293 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3294 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_2085_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3295 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3296 VSS a_3436_n4887# a_3176_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3297 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3298 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3299 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3300 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_4365_n1909# a_4298_n2685# 0.01fF
C1 a_2085_n10301# a_2148_n8695# 0.00fF
C2 B Bd 0.20fF
C3 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C4 a_10738_n509# a_10904_n1079# 0.03fF
C5 a_10805_n5797# a_11164_n5975# 0.05fF
C6 a_4365_n3621# a_4464_n4887# 0.00fF
C7 a_10994_n11933# a_10994_n13021# 0.01fF
C8 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkinv_1_4/Y 0.02fF
C9 a_4464_n3799# a_4365_n4709# 0.00fF
C10 a_501_n1909# a_501_n3621# 0.00fF
C11 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.03fF
C12 a_9616_n2167# a_10805_n1909# 0.01fF
C13 a_9517_n1909# a_10904_n2167# 0.01fF
C14 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.01fF
C15 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C16 a_600_n12503# a_600_n10871# 0.00fF
C17 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_9517_n11237# 0.18fF
C18 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_4661_n4317# 0.01fF
C19 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X a_9616_n3799# 0.05fF
C20 a_2366_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.01fF
C21 a_10994_n2685# a_11101_n2685# 0.55fF
C22 sky130_fd_sc_hd__clkinv_1_5/A a_6373_n7349# 0.01fF
C23 sky130_fd_sc_hd__nand2_4_0/A a_n787_n1909# 0.00fF
C24 sky130_fd_sc_hd__nand2_4_0/Y a_10738_n2685# 0.00fF
C25 a_9706_n509# a_10738_n509# 0.01fF
C26 a_9616_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.03fF
C27 a_10904_n11415# VDD 0.38fF
C28 a_10994_n2685# a_10994_n4317# 0.01fF
C29 a_3077_n11237# a_4464_n11415# 0.01fF
C30 a_3176_n11415# a_4365_n11237# 0.01fF
C31 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_7300_n1079# 0.03fF
C32 a_11101_n11933# a_11101_n10301# 0.01fF
C33 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.68fF
C34 a_4724_n5975# a_4554_n4317# 0.00fF
C35 a_4464_n5975# a_4661_n4317# 0.00fF
C36 a_7237_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C37 a_10738_n4317# a_10994_n4317# 0.19fF
C38 a_1722_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C39 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1789_n2997# 0.00fF
C40 a_1888_n4887# a_3436_n4887# 0.01fF
C41 a_8418_n6493# a_9706_n6493# 0.01fF
C42 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_860_n9783# 0.02fF
C43 a_13765_n11933# p1 0.02fF
C44 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_8162_n5405# 0.03fF
C45 a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C46 sky130_fd_sc_hd__clkinv_1_5/A VDD 12.89fF
C47 p1d_b a_13765_n13565# 0.02fF
C48 a_6941_n8437# a_6012_n8695# 0.02fF
C49 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.02fF
C50 sky130_fd_sc_hd__nand2_1_0/A a_n787_n4709# 0.24fF
C51 a_2085_n5405# a_1722_n5405# 0.05fF
C52 a_5949_n13021# a_6012_n12503# 0.01fF
C53 a_4464_n12503# a_4661_n13021# 0.02fF
C54 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/B 0.11fF
C55 sky130_fd_sc_hd__nand2_4_0/A a_n860_n509# 0.02fF
C56 a_8162_n10301# a_9813_n10301# 0.00fF
C57 a_6941_n10613# a_7130_n10301# 0.02fF
C58 a_7040_n10871# a_6874_n10301# 0.04fF
C59 a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.02fF
C60 a_3176_n12503# a_3436_n12503# 0.28fF
C61 a_9706_n13021# a_10738_n13021# 0.02fF
C62 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_4365_n12325# 0.01fF
C63 a_9450_n13021# a_10994_n13021# 0.01fF
C64 a_2366_n8125# a_2148_n8695# 0.03fF
C65 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C66 a_5586_n2685# a_5949_n2685# 0.05fF
C67 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_4724_n8695# 0.01fF
C68 a_9876_n8695# a_9813_n10301# 0.00fF
C69 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C70 a_600_n1079# a_690_n2685# 0.00fF
C71 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5653_n821# 0.00fF
C72 a_3436_n3255# a_3266_n1597# 0.00fF
C73 a_1789_n1909# a_1722_n1597# 0.01fF
C74 a_3373_n5405# a_4554_n5405# 0.01fF
C75 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4298_n5405# 0.35fF
C76 a_3266_n5405# a_4661_n5405# 0.01fF
C77 B_b a_13765_n1053# 0.12fF
C78 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6658_n7363# 0.01fF
C79 a_6658_n7363# a_7212_n7203# 0.17fF
C80 a_6373_n7349# a_6616_n7581# 0.03fF
C81 a_3077_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C82 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A a_600_n3255# 0.04fF
C83 a_10904_n9783# a_11164_n9783# 0.23fF
C84 a_2148_n9783# a_3436_n9783# 0.01fF
C85 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X a_3176_n9783# 0.05fF
C86 a_4365_n9525# a_3077_n9525# 0.01fF
C87 a_1888_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C88 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_3/A 0.46fF
C89 a_5752_n11415# a_5842_n11933# 0.02fF
C90 a_10738_n11933# a_10805_n12325# 0.01fF
C91 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n5405# 0.01fF
C92 a_7130_n4317# a_7040_n4887# 0.01fF
C93 a_7130_n2685# a_7040_n2167# 0.01fF
C94 a_3010_n5405# a_3010_n4317# 0.02fF
C95 a_6874_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C96 a_9517_n821# a_10805_n821# 0.01fF
C97 a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.18fF
C98 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.08fF
C99 a_6616_n7581# VDD 0.00fF
C100 a_10805_n1909# a_11164_n2167# 0.05fF
C101 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C102 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_7237_n9213# 0.00fF
C103 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_4661_n2685# 0.00fF
C104 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C105 a_860_n11415# a_1789_n11237# 0.02fF
C106 a_501_n11237# a_2148_n11415# 0.00fF
C107 a_600_n12503# sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C108 a_10904_n8695# VDD 0.41fF
C109 a_600_n11415# a_1888_n11415# 0.01fF
C110 a_434_n5405# a_797_n5405# 0.05fF
C111 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C112 a_1888_n10871# VDD 0.46fF
C113 a_n1995_n6925# VDD 0.35fF
C114 a_600_n11415# a_501_n10613# 0.01fF
C115 a_13765_n2685# Bd_b 3.19fF
C116 sky130_fd_sc_hd__nand2_4_0/Y Bd_b 0.00fF
C117 a_4365_n11237# a_4724_n11415# 0.05fF
C118 a_4298_n10301# VDD 0.76fF
C119 a_1888_n10871# a_1978_n10301# 0.02fF
C120 a_5949_n13021# a_4554_n13021# 0.01fF
C121 a_5842_n13021# a_4661_n13021# 0.01fF
C122 Ad_b a_6101_n7254# 0.01fF
C123 a_7300_n4887# a_7130_n4317# 0.04fF
C124 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_4464_n4887# 0.01fF
C125 a_3176_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.03fF
C126 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_7040_n5975# 0.00fF
C127 a_10805_n9525# a_10738_n10301# 0.01fF
C128 a_4298_n1597# a_4298_n2685# 0.02fF
C129 a_8588_n4887# a_8525_n5405# 0.01fF
C130 a_7130_n13021# VDD 0.46fF
C131 a_10994_n5405# a_10904_n3799# 0.00fF
C132 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10805_n9525# 0.01fF
C133 a_10738_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.03fF
C134 a_3373_n5405# a_1978_n5405# 0.01fF
C135 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_1_4/B 0.28fF
C136 a_4298_n4317# a_4298_n2685# 0.01fF
C137 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_4464_n12503# 0.05fF
C138 a_5842_n2685# a_5752_n3255# 0.02fF
C139 a_6941_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C140 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_6874_n11933# 0.00fF
C141 a_13765_n4317# VDD 2.48fF
C142 a_4724_n10871# a_4724_n11415# 0.09fF
C143 a_10738_n8125# a_10738_n9213# 0.01fF
C144 a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.00fF
C145 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_2085_n13021# 0.01fF
C146 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.03fF
C147 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_1722_n2685# 0.00fF
C148 a_5949_n2685# a_6012_n1079# 0.00fF
C149 a_4554_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.05fF
C150 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_5842_n5405# 0.00fF
C151 a_9876_n3799# a_8328_n3799# 0.01fF
C152 a_1722_n4317# a_1722_n5405# 0.02fF
C153 a_3077_n4709# VDD 0.36fF
C154 a_2622_n6493# a_2729_n8125# 0.00fF
C155 a_2729_n6493# a_2622_n8125# 0.00fF
C156 a_4464_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C157 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.29fF
C158 sky130_fd_sc_hd__nand2_1_4/Y Ad_b 0.01fF
C159 a_3436_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.29fF
C160 a_3373_n1597# a_3176_n1079# 0.02fF
C161 a_8162_n14109# a_8525_n14109# 0.05fF
C162 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VDD 0.84fF
C163 a_4464_n5975# sky130_fd_sc_hd__dfxbp_1_0/Q 0.00fF
C164 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n14109# 0.01fF
C165 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.01fF
C166 a_9706_n6493# a_9616_n5975# 0.02fF
C167 a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C168 sky130_fd_sc_hd__dfxbp_1_0/Q a_4554_n9213# 0.00fF
C169 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_6874_n11933# 0.03fF
C170 a_4724_n5975# a_4623_n7349# 0.00fF
C171 a_4623_n7349# a_4661_n9213# 0.00fF
C172 a_10805_n821# a_10904_n1079# 0.48fF
C173 a_7300_n8695# a_6658_n7363# 0.00fF
C174 sky130_fd_sc_hd__nand2_4_2/A a_8525_n14109# 0.02fF
C175 a_7237_n6493# a_7237_n5405# 0.02fF
C176 a_7040_n8695# a_6665_n7459# 0.00fF
C177 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C178 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.00fF
C179 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_10738_n1597# 0.00fF
C180 a_1888_n3255# a_2085_n2685# 0.02fF
C181 a_2148_n12503# a_2148_n10871# 0.01fF
C182 a_690_n1597# a_690_n2685# 0.01fF
C183 a_797_n5405# a_1978_n5405# 0.01fF
C184 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_1722_n5405# 0.35fF
C185 a_3436_n10871# VDD 0.78fF
C186 a_5842_n10301# VDD 0.44fF
C187 a_4661_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.01fF
C188 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C189 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X a_7300_n3799# 0.00fF
C190 a_10738_n6173# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C191 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_10738_n2685# 0.01fF
C192 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD 0.83fF
C193 a_7130_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C194 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_3010_n10301# 0.03fF
C195 a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C196 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2148_n13591# 0.01fF
C197 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.02fF
C198 a_8525_n13021# VDD 0.35fF
C199 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_8588_n5975# 0.29fF
C200 a_3373_n10301# a_4298_n10301# 0.02fF
C201 a_3010_n10301# a_4661_n10301# 0.00fF
C202 a_3266_n10301# a_4554_n10301# 0.01fF
C203 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.08fF
C204 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C205 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C206 a_9876_n8695# a_9813_n8125# 0.01fF
C207 a_11101_n9213# a_11164_n9783# 0.01fF
C208 a_2366_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C209 a_3373_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.02fF
C210 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_2085_n1597# 0.01fF
C211 a_1888_n1079# a_1722_n2685# 0.00fF
C212 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6941_n2997# 0.01fF
C213 a_7130_n1597# a_7040_n1079# 0.01fF
C214 a_7300_n13591# a_7237_n11933# 0.00fF
C215 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6665_n7459# 0.01fF
C216 a_5653_n2997# a_6941_n2997# 0.01fF
C217 a_10738_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C218 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_3436_n8695# 0.03fF
C219 a_11101_n11933# a_10904_n13591# 0.00fF
C220 a_10994_n11933# a_11164_n13591# 0.00fF
C221 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C222 a_6012_n3799# a_6012_n4887# 0.02fF
C223 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_9616_n3799# 0.03fF
C224 a_3176_n2167# a_3266_n1597# 0.02fF
C225 a_10904_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C226 a_7040_n9783# a_8229_n9525# 0.01fF
C227 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_8525_n1597# 0.01fF
C228 a_4298_n1597# a_4365_n1909# 0.01fF
C229 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.03fF
C230 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.04fF
C231 a_8162_n6493# a_8229_n4709# 0.00fF
C232 a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X 0.02fF
C233 a_1888_n2167# a_2148_n2167# 0.28fF
C234 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C235 a_1888_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.03fF
C236 a_8525_n14109# a_9706_n14109# 0.01fF
C237 a_8418_n14109# a_9813_n14109# 0.01fF
C238 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9450_n14109# 0.34fF
C239 a_7237_n13021# a_7237_n14109# 0.02fF
C240 a_7300_n11415# a_7237_n11933# 0.01fF
C241 a_9813_n9213# a_11101_n9213# 0.01fF
C242 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10994_n9213# 0.03fF
C243 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__nand2_4_2/B 0.75fF
C244 a_4554_n5405# a_4554_n4317# 0.01fF
C245 a_1722_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.01fF
C246 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1722_n2685# 0.01fF
C247 a_9813_n1597# a_11101_n1597# 0.01fF
C248 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10994_n1597# 0.03fF
C249 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_4464_n2167# 0.01fF
C250 a_434_n4317# a_600_n3255# 0.00fF
C251 a_501_n4709# a_690_n5405# 0.02fF
C252 a_600_n4887# a_434_n5405# 0.04fF
C253 a_5752_n12503# a_5586_n11933# 0.04fF
C254 a_690_n4317# a_501_n2997# 0.00fF
C255 a_9450_n13021# a_9517_n13413# 0.01fF
C256 a_10994_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.04fF
C257 a_11101_n5405# a_11164_n4887# 0.01fF
C258 a_9616_n4887# a_10805_n4709# 0.01fF
C259 a_8229_n3621# VDD 0.35fF
C260 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.02fF
C261 a_9517_n4709# a_10904_n4887# 0.01fF
C262 a_7237_n10301# VDD 0.35fF
C263 a_11164_n3799# a_11101_n2685# 0.00fF
C264 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.04fF
C265 a_8588_n2167# a_7040_n2167# 0.01fF
C266 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.03fF
C267 a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C268 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_8525_n4317# 0.01fF
C269 a_8328_n2167# a_7300_n2167# 0.02fF
C270 a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.18fF
C271 a_3436_n10871# a_3373_n10301# 0.01fF
C272 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.02fF
C273 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_10738_n4317# 0.02fF
C274 a_11164_n3799# a_10994_n4317# 0.04fF
C275 a_10904_n3799# a_11101_n4317# 0.02fF
C276 sky130_fd_sc_hd__clkinv_1_0/A a_3077_n821# 0.06fF
C277 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_5586_n10301# 0.00fF
C278 a_5842_n1597# a_5842_n2685# 0.01fF
C279 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.29fF
C280 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X a_6941_n2997# 0.18fF
C281 a_6012_n3255# a_7040_n3255# 0.02fF
C282 a_5752_n3255# a_7300_n3255# 0.01fF
C283 a_9706_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C284 a_5752_n11415# a_4365_n11237# 0.01fF
C285 a_5653_n11237# a_4464_n11415# 0.01fF
C286 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5653_n821# 0.01fF
C287 a_10805_n10613# a_10805_n11237# 0.05fF
C288 a_5752_n13591# a_7040_n13591# 0.01fF
C289 sky130_fd_sc_hd__clkinv_1_0/A a_10738_n1597# 0.00fF
C290 a_5653_n13413# a_7300_n13591# 0.00fF
C291 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8229_n821# 0.01fF
C292 a_8162_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.03fF
C293 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.00fF
C294 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__nand2_4_3/Y 0.69fF
C295 a_9450_n13021# a_9517_n11237# 0.00fF
C296 a_1789_n9525# VDD 0.36fF
C297 a_3077_n3621# a_3077_n4709# 0.02fF
C298 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.29fF
C299 a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.00fF
C300 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.04fF
C301 a_10738_n2685# VDD 0.70fF
C302 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.00fF
C303 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_2148_n3799# 0.00fF
C304 a_8229_n12325# a_8418_n11933# 0.02fF
C305 a_8328_n12503# a_8162_n11933# 0.04fF
C306 a_1978_n10301# a_1789_n9525# 0.02fF
C307 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3373_n9213# 0.02fF
C308 a_2085_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C309 a_8418_n8125# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C310 a_1722_n10301# a_1888_n9783# 0.04fF
C311 a_8525_n8125# a_9813_n8125# 0.01fF
C312 a_2148_n2167# a_3436_n2167# 0.01fF
C313 a_1888_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.00fF
C314 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.69fF
C315 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_3176_n2167# 0.05fF
C316 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_3436_n5975# 0.03fF
C317 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.00fF
C318 a_4661_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.01fF
C319 a_501_n11237# a_501_n12325# 0.02fF
C320 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_4724_n1079# 0.03fF
C321 a_9706_n14109# sky130_fd_sc_hd__nand2_4_2/B 0.05fF
C322 a_11101_n9213# sky130_fd_sc_hd__clkinv_4_10/Y 0.01fF
C323 a_1888_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.05fF
C324 a_2148_n13591# a_860_n13591# 0.01fF
C325 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_600_n13591# 0.00fF
C326 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.04fF
C327 a_5586_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C328 a_3436_n3255# VDD 0.78fF
C329 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__clkdlybuf4s50_1_50/X 0.06fF
C330 a_7040_n2167# a_6941_n821# 0.00fF
C331 a_6941_n1909# a_7040_n1079# 0.00fF
C332 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.00fF
C333 a_2085_n1597# a_2085_n2685# 0.02fF
C334 a_10805_n9525# VDD 0.32fF
C335 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_4724_n2167# 0.03fF
C336 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C337 a_8162_n5405# a_8229_n3621# 0.00fF
C338 a_434_n9213# a_2085_n9213# 0.00fF
C339 a_5949_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.12fF
C340 a_3077_n10613# a_3010_n9213# 0.00fF
C341 a_9616_n3799# VDD 0.42fF
C342 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C343 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_9876_n10871# 0.03fF
C344 a_434_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.45fF
C345 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkinv_1_4/Y 0.04fF
C346 sky130_fd_sc_hd__clkinv_4_8/Y a_11101_n13021# 0.01fF
C347 a_797_n4317# a_1722_n4317# 0.02fF
C348 a_434_n4317# a_2085_n4317# 0.00fF
C349 a_5842_n1597# a_5752_n3255# 0.00fF
C350 a_6941_n9525# a_7130_n9213# 0.02fF
C351 a_690_n4317# a_1978_n4317# 0.01fF
C352 a_8418_n1597# a_8328_n3255# 0.00fF
C353 a_7040_n9783# a_6874_n9213# 0.04fF
C354 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_6658_n7363# 0.01fF
C355 a_7130_n8125# a_6865_n7304# 0.02fF
C356 a_7237_n8125# a_6665_n7459# 0.00fF
C357 a_6874_n8125# a_6794_n7203# 0.02fF
C358 sky130_fd_sc_hd__clkinv_1_0/A a_4464_n1079# 0.07fF
C359 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C360 a_6874_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C361 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C362 sky130_fd_sc_hd__nand2_4_0/Y a_10738_n509# 0.49fF
C363 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X a_8328_n3255# 0.01fF
C364 a_7040_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C365 a_6874_n6493# a_8418_n6493# 0.01fF
C366 a_7130_n6493# a_8162_n6493# 0.02fF
C367 a_600_n3799# a_690_n5405# 0.00fF
C368 Bd_b a_6373_n7349# 0.01fF
C369 a_10994_n4317# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C370 a_5949_n1597# a_6012_n1079# 0.01fF
C371 a_1789_n10613# a_1722_n11933# 0.00fF
C372 a_8525_n1597# a_8588_n1079# 0.01fF
C373 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C374 a_9876_n12503# a_9813_n13021# 0.01fF
C375 a_3176_n9783# VDD 0.47fF
C376 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VDD 0.90fF
C377 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_8525_n5405# 0.01fF
C378 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.02fF
C379 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkinv_4_4/A 0.02fF
C380 a_9450_n2685# a_9517_n821# 0.00fF
C381 Bd_b VDD 9.36fF
C382 a_9616_n12503# a_9813_n14109# 0.00fF
C383 a_9876_n12503# a_9706_n14109# 0.00fF
C384 a_5752_n9783# a_5653_n8437# 0.00fF
C385 a_600_n5975# a_860_n5975# 0.28fF
C386 a_5653_n9525# a_5752_n8695# 0.00fF
C387 a_9450_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C388 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkinv_4_7/A 0.11fF
C389 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C390 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.29fF
C391 a_6012_n11415# a_6012_n10871# 0.09fF
C392 a_8229_n9525# a_8229_n8437# 0.02fF
C393 a_1789_n2997# a_1789_n3621# 0.05fF
C394 a_1789_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.02fF
C395 a_1888_n4887# a_2148_n4887# 0.28fF
C396 sky130_fd_sc_hd__clkinv_1_0/A a_6941_n821# 0.06fF
C397 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.08fF
C398 a_4365_n12325# a_4554_n11933# 0.02fF
C399 a_4464_n12503# a_4298_n11933# 0.04fF
C400 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6794_n7203# 0.00fF
C401 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11164_n4887# 0.00fF
C402 a_11101_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C403 sky130_fd_sc_hd__clkinv_4_3/A a_11164_n4887# 0.10fF
C404 a_9706_n1597# a_9876_n3255# 0.00fF
C405 a_6658_n7363# sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C406 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD 0.83fF
C407 a_5586_n5405# a_5653_n4709# 0.01fF
C408 a_9813_n1597# a_9616_n3255# 0.00fF
C409 a_1789_n1909# VDD 0.36fF
C410 a_n428_n4887# a_600_n4887# 0.02fF
C411 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VDD 0.72fF
C412 a_1722_n4317# a_1789_n3621# 0.01fF
C413 a_1722_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C414 a_1978_n9213# a_2085_n9213# 0.55fF
C415 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_3010_n9213# 0.00fF
C416 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.02fF
C417 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8525_n14109# 0.02fF
C418 a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C419 a_4298_n1597# a_5842_n1597# 0.01fF
C420 a_4554_n1597# a_5586_n1597# 0.02fF
C421 a_6874_n1597# a_8418_n1597# 0.01fF
C422 a_1978_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C423 a_3436_n8695# a_3266_n9213# 0.04fF
C424 a_3176_n8695# a_3373_n9213# 0.02fF
C425 a_9616_n11415# a_9450_n11933# 0.04fF
C426 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6874_n8125# 0.33fF
C427 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6941_n2997# 0.00fF
C428 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_3010_n4317# 0.00fF
C429 a_6874_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C430 a_9450_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C431 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9517_n2997# 0.00fF
C432 a_4464_n2167# VDD 0.47fF
C433 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_10904_n3799# 0.05fF
C434 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6874_n509# 0.33fF
C435 a_9876_n3799# a_11164_n3799# 0.01fF
C436 a_8525_n14109# a_8328_n13591# 0.02fF
C437 a_8418_n14109# a_8588_n13591# 0.04fF
C438 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X a_8588_n3255# 0.03fF
C439 a_7300_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C440 a_9706_n8125# a_9616_n9783# 0.00fF
C441 a_9616_n4887# a_9517_n5797# 0.00fF
C442 a_9517_n4709# a_9616_n5975# 0.00fF
C443 a_8162_n6493# a_8525_n6493# 0.05fF
C444 a_1789_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C445 a_9517_n12325# a_9876_n12503# 0.05fF
C446 a_5752_n5975# a_5653_n4709# 0.00fF
C447 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.05fF
C448 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X a_1722_n5405# 0.00fF
C449 a_6874_n13021# a_6874_n11933# 0.02fF
C450 a_5653_n5797# a_5752_n4887# 0.00fF
C451 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.02fF
C452 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_9813_n13021# 0.01fF
C453 a_6941_n10613# a_7040_n12503# 0.00fF
C454 a_7040_n10871# a_6941_n12325# 0.00fF
C455 a_10994_n9213# VDD 0.42fF
C456 a_1888_n5975# a_2085_n5405# 0.02fF
C457 a_9876_n11415# a_9876_n9783# 0.01fF
C458 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_1_5/A 0.37fF
C459 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_501_n4709# 0.18fF
C460 a_10904_n12503# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C461 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.04fF
C462 a_3373_n10301# a_3176_n9783# 0.02fF
C463 a_3266_n10301# a_3436_n9783# 0.04fF
C464 a_5949_n9213# a_4661_n9213# 0.01fF
C465 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_4554_n9213# 0.01fF
C466 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.03fF
C467 a_4661_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.12fF
C468 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_501_n10613# 0.00fF
C469 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C470 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_3373_n2685# 0.00fF
C471 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_3176_n4887# 0.05fF
C472 a_3176_n3799# a_3176_n3255# 0.07fF
C473 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.07fF
C474 a_2148_n3799# VDD 0.77fF
C475 sky130_fd_sc_hd__clkinv_1_0/A a_8328_n1079# 0.07fF
C476 a_501_n5797# VDD 0.37fF
C477 a_2366_n8125# sky130_fd_sc_hd__clkinv_1_3/A 0.01fF
C478 a_8418_n4317# a_8229_n3621# 0.02fF
C479 a_3176_n2167# VDD 0.47fF
C480 a_8162_n4317# a_8328_n3799# 0.04fF
C481 a_8588_n10871# a_8525_n9213# 0.00fF
C482 a_1722_n13021# a_3010_n13021# 0.01fF
C483 a_860_n10871# a_860_n9783# 0.02fF
C484 a_5752_n3799# a_6941_n3621# 0.01fF
C485 a_5653_n3621# a_7040_n3799# 0.01fF
C486 a_1888_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C487 a_1978_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C488 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C489 a_9706_n5405# a_9616_n3799# 0.00fF
C490 a_1888_n13591# a_2085_n11933# 0.00fF
C491 a_9616_n11415# a_9450_n10301# 0.00fF
C492 a_2148_n13591# a_1978_n11933# 0.00fF
C493 a_5586_n1597# a_5949_n1597# 0.05fF
C494 a_7300_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C495 a_10904_n10871# a_11101_n11933# 0.00fF
C496 a_11164_n10871# a_10994_n11933# 0.00fF
C497 sky130_fd_sc_hd__dfxbp_1_0/Q a_6012_n5975# 0.00fF
C498 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_434_n4317# 0.03fF
C499 a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.01fF
C500 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_8418_n8125# 0.00fF
C501 a_6012_n2167# VDD 0.78fF
C502 a_7130_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.05fF
C503 a_4724_n12503# a_6012_n12503# 0.01fF
C504 a_6941_n2997# a_6941_n4709# 0.00fF
C505 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_8418_n509# 0.00fF
C506 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_5752_n12503# 0.05fF
C507 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.37fF
C508 a_3436_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.29fF
C509 a_11164_n1079# a_10994_n2685# 0.00fF
C510 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_10738_n2685# 0.00fF
C511 sky130_fd_sc_hd__nand2_4_0/Y a_10805_n821# 0.02fF
C512 a_860_n8695# a_1888_n8695# 0.02fF
C513 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_1789_n8437# 0.18fF
C514 a_600_n8695# a_2148_n8695# 0.01fF
C515 a_10904_n1079# a_11101_n2685# 0.00fF
C516 a_501_n4709# a_600_n3799# 0.00fF
C517 a_9616_n12503# a_11164_n12503# 0.01fF
C518 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n6493# 0.35fF
C519 a_600_n4887# a_501_n3621# 0.00fF
C520 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_10805_n12325# 0.17fF
C521 a_9876_n12503# a_10904_n12503# 0.02fF
C522 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C523 a_434_n9213# a_1978_n9213# 0.01fF
C524 a_690_n9213# a_1722_n9213# 0.02fF
C525 a_6874_n2685# a_6941_n3621# 0.00fF
C526 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C527 a_3176_n10871# a_3266_n11933# 0.01fF
C528 sky130_fd_sc_hd__clkinv_1_0/Y a_2148_n1079# 0.01fF
C529 a_1722_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.00fF
C530 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.00fF
C531 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C532 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.01fF
C533 sky130_fd_sc_hd__nand2_4_0/A a_11164_n1079# 0.04fF
C534 a_797_n4317# a_860_n4887# 0.01fF
C535 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_1722_n11933# 0.03fF
C536 a_5653_n11237# a_7040_n11415# 0.01fF
C537 a_5752_n11415# a_6941_n11237# 0.01fF
C538 a_6006_n7607# a_6101_n7254# 0.20fF
C539 a_5052_n7283# a_6373_n7349# 0.01fF
C540 a_6012_n3799# a_6941_n3621# 0.02fF
C541 a_3077_n8437# a_4464_n8695# 0.01fF
C542 a_3176_n8695# a_4365_n8437# 0.01fF
C543 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.14fF
C544 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.02fF
C545 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.09fF
C546 a_10904_n3799# VDD 0.38fF
C547 a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C548 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.02fF
C549 a_6941_n13413# a_7300_n13591# 0.05fF
C550 a_1888_n5975# a_1722_n4317# 0.00fF
C551 a_1789_n5797# a_1978_n4317# 0.00fF
C552 sky130_fd_sc_hd__clkinv_4_8/Y a_9616_n13591# 0.00fF
C553 a_6874_n9213# a_7237_n9213# 0.05fF
C554 sky130_fd_sc_hd__nand2_4_0/A a_9813_n509# 0.06fF
C555 a_9706_n8125# a_9813_n9213# 0.00fF
C556 a_9616_n2167# a_9450_n1597# 0.04fF
C557 a_9517_n1909# a_9706_n1597# 0.02fF
C558 a_5052_n7283# VDD 0.55fF
C559 a_3010_n13021# a_3266_n13021# 0.19fF
C560 a_9813_n11933# a_8418_n11933# 0.01fF
C561 a_1888_n12503# a_1722_n13021# 0.04fF
C562 a_1789_n12325# a_1978_n13021# 0.02fF
C563 a_10738_n5405# a_10994_n5405# 0.19fF
C564 a_6012_n9783# a_6012_n10871# 0.02fF
C565 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.08fF
C566 a_8229_n9525# a_8418_n8125# 0.00fF
C567 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkinv_1_0/A 0.00fF
C568 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_0/A 0.33fF
C569 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.00fF
C570 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_6012_n9783# 0.03fF
C571 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.06fF
C572 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C573 a_4724_n12503# a_4554_n13021# 0.04fF
C574 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6874_n1597# 0.35fF
C575 a_6794_n7203# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C576 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C577 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X a_4661_n9213# 0.01fF
C578 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.03fF
C579 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VDD 0.90fF
C580 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A VDD 0.89fF
C581 a_5752_n12503# VDD 0.44fF
C582 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.29fF
C583 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8525_n509# 0.02fF
C584 p2_b p2 0.47fF
C585 a_7237_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C586 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.02fF
C587 a_8229_n8437# a_8418_n9213# 0.02fF
C588 a_8328_n8695# a_8162_n9213# 0.04fF
C589 a_9813_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C590 sky130_fd_sc_hd__nand2_4_2/B a_9876_n13591# 0.03fF
C591 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A Bd_b 0.11fF
C592 a_8418_n13021# a_8418_n11933# 0.01fF
C593 a_10904_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.02fF
C594 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.06fF
C595 a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.00fF
C596 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A sky130_fd_sc_hd__clkinv_4_3/Y 0.03fF
C597 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_4298_n11933# 0.01fF
C598 sky130_fd_sc_hd__dfxbp_1_1/D VDD 1.06fF
C599 a_434_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C600 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_3373_n5405# 0.01fF
C601 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_7300_n13591# 0.03fF
C602 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.03fF
C603 a_1722_n2685# a_1789_n3621# 0.00fF
C604 a_10738_n8125# a_11164_n8695# 0.05fF
C605 a_5842_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C606 a_2148_n11415# a_2085_n11933# 0.01fF
C607 sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1597# 0.04fF
C608 a_6874_n8125# a_6874_n9213# 0.02fF
C609 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.03fF
C610 a_6941_n11237# a_7300_n11415# 0.05fF
C611 a_3077_n13413# a_4464_n13591# 0.01fF
C612 a_3176_n13591# a_4365_n13413# 0.01fF
C613 a_7040_n3799# a_7300_n3799# 0.28fF
C614 a_6941_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C615 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_8229_n3621# 0.01fF
C616 a_9876_n2167# a_9876_n3255# 0.02fF
C617 a_7300_n4887# a_7300_n5975# 0.02fF
C618 a_4365_n8437# a_4724_n8695# 0.05fF
C619 a_4724_n4887# VDD 0.78fF
C620 a_501_n3621# a_860_n3799# 0.05fF
C621 a_2729_n509# a_2366_n509# 0.05fF
C622 a_7300_n13591# a_8328_n13591# 0.02fF
C623 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_8229_n13413# 0.18fF
C624 a_7040_n13591# a_8588_n13591# 0.01fF
C625 a_2148_n3799# a_3077_n3621# 0.02fF
C626 a_7237_n9213# a_8418_n9213# 0.01fF
C627 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8162_n9213# 0.35fF
C628 a_7130_n9213# a_8525_n9213# 0.01fF
C629 a_4724_n3799# a_4724_n3255# 0.09fF
C630 a_3077_n1909# a_3176_n3799# 0.00fF
C631 a_10738_n509# VDD 0.11fF
C632 a_3176_n2167# a_3077_n3621# 0.00fF
C633 a_10904_n11415# a_10738_n13021# 0.00fF
C634 a_10805_n11237# a_10994_n13021# 0.00fF
C635 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/Y 0.05fF
C636 a_3266_n13021# a_4554_n13021# 0.01fF
C637 a_3373_n13021# a_4298_n13021# 0.02fF
C638 a_3010_n13021# a_4661_n13021# 0.00fF
C639 a_797_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C640 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9706_n11933# 0.05fF
C641 a_4464_n10871# a_3077_n10613# 0.01fF
C642 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_860_n3799# 0.03fF
C643 a_10994_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C644 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.04fF
C645 a_5653_n9525# a_5653_n11237# 0.00fF
C646 a_4298_n13021# VDD 0.76fF
C647 a_11164_n11415# a_10994_n10301# 0.00fF
C648 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.00fF
C649 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_3373_n11933# 0.00fF
C650 sky130_fd_sc_hd__nand2_4_2/B a_10738_n13789# 0.36fF
C651 a_10904_n11415# a_11101_n10301# 0.00fF
C652 a_600_n12503# a_1888_n12503# 0.01fF
C653 a_860_n12503# a_1789_n12325# 0.02fF
C654 a_9876_n12503# a_9876_n13591# 0.02fF
C655 a_4464_n9783# a_4298_n10301# 0.04fF
C656 a_1789_n12325# VDD 0.36fF
C657 a_4365_n9525# a_4554_n10301# 0.02fF
C658 a_4464_n3799# a_4464_n2167# 0.00fF
C659 a_3266_n2685# a_4298_n2685# 0.02fF
C660 a_3010_n2685# a_4554_n2685# 0.01fF
C661 a_3436_n12503# a_4724_n12503# 0.01fF
C662 a_3176_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C663 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.06fF
C664 a_8162_n10301# a_8162_n9213# 0.02fF
C665 a_7300_n12503# VDD 0.77fF
C666 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C667 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6874_n9213# 0.03fF
C668 a_8162_n2685# a_9450_n2685# 0.01fF
C669 a_1888_n3255# a_3436_n3255# 0.01fF
C670 sky130_fd_sc_hd__mux2_1_0/X a_4554_n9213# 0.00fF
C671 a_2366_n14109# a_2622_n14109# 0.18fF
C672 a_4464_n5975# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C673 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n11933# 0.01fF
C674 a_9450_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C675 a_9813_n5405# a_9616_n3799# 0.00fF
C676 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A VDD 0.63fF
C677 a_8418_n2685# a_8328_n3799# 0.01fF
C678 a_8328_n9783# a_9616_n9783# 0.01fF
C679 a_8588_n9783# a_9517_n9525# 0.02fF
C680 a_501_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.02fF
C681 a_1722_n10301# a_3010_n10301# 0.01fF
C682 a_600_n9783# a_860_n9783# 0.28fF
C683 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.23fF
C684 a_n428_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.02fF
C685 sky130_fd_sc_hd__clkinv_4_3/A Ad_b 0.00fF
C686 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_4661_n4317# 0.01fF
C687 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.05fF
C688 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.02fF
C689 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.04fF
C690 a_9517_n5797# a_9876_n5975# 0.05fF
C691 a_600_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.04fF
C692 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.03fF
C693 a_600_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.04fF
C694 a_7300_n11415# a_8328_n11415# 0.02fF
C695 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_8229_n11237# 0.18fF
C696 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_3373_n4317# 0.01fF
C697 a_4365_n11237# a_4365_n10613# 0.05fF
C698 a_7040_n11415# a_8588_n11415# 0.01fF
C699 a_7040_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C700 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X a_8328_n3799# 0.05fF
C701 a_4365_n13413# a_4724_n13591# 0.05fF
C702 a_7300_n3799# a_8588_n3799# 0.01fF
C703 a_4464_n8695# a_6012_n8695# 0.01fF
C704 a_4724_n8695# a_5752_n8695# 0.02fF
C705 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X a_5653_n8437# 0.18fF
C706 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VDD 0.86fF
C707 a_2148_n12503# a_2366_n14109# 0.00fF
C708 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_9616_n13591# 0.01fF
C709 a_8328_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C710 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X a_1789_n3621# 0.18fF
C711 a_860_n3799# a_1888_n3799# 0.02fF
C712 a_6874_n14109# VDD 0.73fF
C713 a_1789_n11237# a_3176_n11415# 0.01fF
C714 a_1888_n11415# a_3077_n11237# 0.01fF
C715 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_4365_n3621# 0.01fF
C716 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.84fF
C717 a_3436_n5975# a_3266_n4317# 0.00fF
C718 a_3176_n5975# a_3373_n4317# 0.00fF
C719 a_9813_n11933# a_9813_n10301# 0.01fF
C720 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_9706_n9213# 0.00fF
C721 a_10805_n10613# a_10738_n9213# 0.00fF
C722 a_8418_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.05fF
C723 a_9450_n4317# a_9706_n4317# 0.19fF
C724 a_1888_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.05fF
C725 a_10994_n5405# a_10994_n4317# 0.01fF
C726 a_4554_n13021# a_4661_n13021# 0.55fF
C727 a_4298_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C728 a_8588_n9783# a_8418_n10301# 0.04fF
C729 a_4724_n10871# a_4365_n10613# 0.05fF
C730 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_10738_n10301# 0.00fF
C731 a_11164_n8695# a_10994_n10301# 0.00fF
C732 a_10904_n8695# a_11101_n10301# 0.00fF
C733 a_3176_n12503# a_3373_n13021# 0.02fF
C734 a_6941_n8437# a_8328_n8695# 0.01fF
C735 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C736 a_3436_n12503# a_3266_n13021# 0.04fF
C737 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_3077_n12325# 0.01fF
C738 a_6874_n10301# a_8525_n10301# 0.00fF
C739 a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.02fF
C740 a_1888_n12503# a_2148_n12503# 0.28fF
C741 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.04fF
C742 a_5752_n10871# a_5586_n10301# 0.04fF
C743 a_5653_n10613# a_5842_n10301# 0.02fF
C744 a_8588_n8695# a_8525_n10301# 0.00fF
C745 a_3176_n12503# VDD 0.44fF
C746 a_4298_n2685# a_4661_n2685# 0.05fF
C747 sky130_fd_sc_hd__dfxbp_1_0/Q a_6794_n7203# 0.02fF
C748 a_9876_n4887# a_9876_n3255# 0.01fF
C749 a_9706_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.10fF
C750 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VDD 0.85fF
C751 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VDD 0.85fF
C752 a_9706_n6493# a_9876_n4887# 0.00fF
C753 a_9450_n2685# a_9706_n2685# 0.19fF
C754 a_9450_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.03fF
C755 a_2085_n5405# a_3266_n5405# 0.01fF
C756 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3010_n5405# 0.35fF
C757 a_1789_n1909# a_1888_n3255# 0.00fF
C758 a_9876_n8695# a_9706_n9213# 0.04fF
C759 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_10805_n9525# 0.01fF
C760 a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.02fF
C761 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9517_n3621# 0.00fF
C762 a_9450_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C763 a_9616_n9783# a_9876_n9783# 0.28fF
C764 a_3010_n10301# a_3266_n10301# 0.19fF
C765 a_860_n9783# a_2148_n9783# 0.01fF
C766 a_600_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C767 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X a_1888_n9783# 0.05fF
C768 a_10738_n1597# a_10738_n2685# 0.02fF
C769 a_5842_n4317# a_5752_n4887# 0.01fF
C770 a_5586_n13021# a_5752_n13591# 0.04fF
C771 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_10805_n5797# 0.17fF
C772 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_797_n9213# 0.01fF
C773 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.03fF
C774 a_9876_n5975# a_10904_n5975# 0.02fF
C775 a_9616_n5975# a_11164_n5975# 0.01fF
C776 a_8418_n8125# a_8418_n9213# 0.01fF
C777 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n13021# 0.01fF
C778 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_5949_n9213# 0.00fF
C779 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.00fF
C780 a_8328_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.03fF
C781 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C782 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.08fF
C783 a_9517_n1909# a_9876_n2167# 0.05fF
C784 a_4724_n13591# a_5752_n13591# 0.02fF
C785 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_5653_n13413# 0.18fF
C786 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_3373_n2685# 0.00fF
C787 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C788 a_8588_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.29fF
C789 a_8328_n2167# a_8328_n3799# 0.00fF
C790 a_5752_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.03fF
C791 a_7237_n5405# a_7040_n4887# 0.02fF
C792 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C793 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X a_9876_n13591# 0.03fF
C794 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.29fF
C795 a_3077_n11237# a_3436_n11415# 0.05fF
C796 a_10738_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C797 a_9876_n11415# VDD 0.74fF
C798 a_9813_n4317# a_10738_n4317# 0.02fF
C799 a_9706_n4317# a_10994_n4317# 0.01fF
C800 a_7237_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C801 a_9450_n4317# a_11101_n4317# 0.00fF
C802 a_600_n10871# a_690_n10301# 0.02fF
C803 B a_13765_n1053# 2.54fF
C804 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_10738_n13789# 0.01fF
C805 a_10805_n821# VDD 0.32fF
C806 sky130_fd_sc_hd__clkinv_4_4/A Bd_b 0.46fF
C807 a_797_n1597# a_860_n3255# 0.00fF
C808 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkinv_1_5/A 0.39fF
C809 a_9517_n9525# a_9450_n10301# 0.01fF
C810 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.07fF
C811 a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C812 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X a_501_n9525# 0.01fF
C813 a_7300_n4887# a_7237_n5405# 0.01fF
C814 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A p2d_b 0.04fF
C815 a_2085_n5405# a_690_n5405# 0.01fF
C816 a_7040_n9783# a_7040_n11415# 0.00fF
C817 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.04fF
C818 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n2685# 0.35fF
C819 a_9813_n2685# a_10994_n2685# 0.01fF
C820 a_9706_n2685# a_11101_n2685# 0.01fF
C821 a_3010_n4317# a_3010_n2685# 0.01fF
C822 a_9450_n13021# a_9813_n13021# 0.05fF
C823 a_8162_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.03fF
C824 a_1888_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.00fF
C825 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_3176_n12503# 0.05fF
C826 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X sky130_fd_sc_hd__clkdlybuf4s50_1_50/X 0.05fF
C827 a_2148_n12503# a_3436_n12503# 0.01fF
C828 a_6874_n509# a_6941_n1909# 0.00fF
C829 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_9450_n10301# 0.00fF
C830 a_9616_n8695# a_9450_n8125# 0.04fF
C831 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C832 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5586_n2685# 0.35fF
C833 a_4554_n2685# a_5949_n2685# 0.01fF
C834 a_4661_n2685# a_5842_n2685# 0.01fF
C835 A_b VDD 4.25fF
C836 a_1722_n1597# a_3010_n1597# 0.01fF
C837 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.08fF
C838 a_n787_n1909# a_n688_n2167# 0.49fF
C839 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_4554_n5405# 0.00fF
C840 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.08fF
C841 a_3266_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.05fF
C842 a_6941_n8437# a_7130_n8125# 0.02fF
C843 a_7130_n14109# a_7237_n14109# 0.53fF
C844 a_9706_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C845 a_8418_n10301# a_9450_n10301# 0.02fF
C846 a_1888_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C847 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X a_10904_n9783# 0.05fF
C848 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.29fF
C849 a_9876_n9783# a_11164_n9783# 0.01fF
C850 a_8525_n509# a_8418_n1597# 0.00fF
C851 a_8418_n509# a_8525_n1597# 0.00fF
C852 a_10738_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.01fF
C853 a_10738_n8125# a_10904_n9783# 0.00fF
C854 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6941_n4709# 0.01fF
C855 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.03fF
C856 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C857 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_9876_n12503# 0.00fF
C858 a_9517_n821# a_9616_n1079# 0.49fF
C859 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.03fF
C860 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9450_n9213# 0.01fF
C861 a_9450_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C862 a_9616_n2167# a_11164_n2167# 0.01fF
C863 a_600_n2167# a_600_n3799# 0.00fF
C864 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_10805_n1909# 0.17fF
C865 a_9876_n2167# a_10904_n2167# 0.02fF
C866 a_860_n12503# a_860_n10871# 0.01fF
C867 sky130_fd_sc_hd__clkinv_4_8/A a_10994_n13021# 0.09fF
C868 a_11101_n11933# a_11101_n13021# 0.02fF
C869 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.05fF
C870 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_434_n5405# 0.42fF
C871 a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.02fF
C872 a_860_n10871# VDD 0.78fF
C873 sky130_fd_sc_hd__clkinv_1_5/A a_6665_n7459# 0.40fF
C874 a_10994_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.04fF
C875 sky130_fd_sc_hd__nand2_4_0/Y a_11101_n2685# 0.01fF
C876 a_3176_n11415# a_4724_n11415# 0.01fF
C877 a_4464_n5975# a_4365_n4709# 0.00fF
C878 a_4365_n5797# a_4464_n4887# 0.00fF
C879 a_3436_n11415# a_4464_n11415# 0.02fF
C880 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_4365_n11237# 0.18fF
C881 a_11101_n2685# a_11101_n4317# 0.01fF
C882 sky130_fd_sc_hd__nand2_4_0/B a_10738_n509# 0.38fF
C883 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VDD 0.62fF
C884 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C885 a_10738_n4317# sky130_fd_sc_hd__clkinv_4_3/A 0.00fF
C886 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C887 a_10994_n4317# a_11101_n4317# 0.55fF
C888 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_6012_n3799# 0.00fF
C889 a_11101_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C890 a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C891 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X VDD 0.81fF
C892 a_5842_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C893 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_1722_n10301# 0.03fF
C894 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_3436_n4887# 0.03fF
C895 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.00fF
C896 clk sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.00fF
C897 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9706_n6493# 0.03fF
C898 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.02fF
C899 a_5949_n13021# VDD 0.34fF
C900 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10805_n3621# 0.00fF
C901 a_10738_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C902 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_1978_n5405# 0.05fF
C903 a_3266_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C904 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C905 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_1_4/Y 0.01fF
C906 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.08fF
C907 a_9517_n11237# a_10805_n11237# 0.01fF
C908 a_9813_n9213# a_9876_n9783# 0.01fF
C909 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C910 a_10805_n13413# VDD 0.31fF
C911 a_9450_n13021# a_9517_n12325# 0.01fF
C912 a_7040_n10871# a_7237_n10301# 0.02fF
C913 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.29fF
C914 a_7300_n10871# a_7130_n10301# 0.04fF
C915 a_9706_n13021# a_11101_n13021# 0.01fF
C916 a_6012_n13591# a_5949_n11933# 0.00fF
C917 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C918 a_860_n1079# a_797_n2685# 0.00fF
C919 a_5842_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.05fF
C920 a_5653_n2997# a_5842_n2685# 0.02fF
C921 a_3010_n1597# a_3266_n1597# 0.19fF
C922 a_10994_n5405# sky130_fd_sc_hd__clkinv_4_4/Y 0.01fF
C923 a_1888_n2167# a_1978_n1597# 0.02fF
C924 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4661_n5405# 0.02fF
C925 a_3373_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.01fF
C926 a_1888_n4887# VDD 0.44fF
C927 a_5752_n9783# a_6941_n9525# 0.01fF
C928 a_5653_n9525# a_7040_n9783# 0.01fF
C929 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6865_n7304# 0.00fF
C930 a_6865_n7304# a_7212_n7203# 0.09fF
C931 a_3436_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C932 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C933 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C934 a_8418_n8125# a_9450_n8125# 0.02fF
C935 a_4724_n9783# a_3077_n9525# 0.00fF
C936 a_4365_n9525# a_3436_n9783# 0.02fF
C937 a_4464_n9783# a_3176_n9783# 0.01fF
C938 a_6012_n11415# a_5949_n11933# 0.01fF
C939 a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C940 a_7237_n2685# a_7300_n2167# 0.01fF
C941 a_9876_n1079# a_10805_n821# 0.02fF
C942 a_9616_n1079# a_10904_n1079# 0.01fF
C943 a_3266_n5405# a_3266_n4317# 0.01fF
C944 a_10994_n11933# a_10904_n12503# 0.01fF
C945 a_9517_n821# a_11164_n1079# 0.00fF
C946 sky130_fd_sc_hd__nand2_4_3/A VDD 13.16fF
C947 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD 3.54fF
C948 a_600_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C949 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C950 a_690_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.05fF
C951 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD 0.83fF
C952 a_860_n11415# a_2148_n11415# 0.01fF
C953 a_n1570_n6769# VDD 0.80fF
C954 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_1978_n5405# 0.00fF
C955 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.01fF
C956 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_8588_n10871# 0.01fF
C957 sky130_fd_sc_hd__nand2_4_1/A p2 0.17fF
C958 a_8162_n13021# a_8229_n13413# 0.01fF
C959 a_8229_n4709# a_9616_n4887# 0.01fF
C960 a_8328_n4887# a_9517_n4709# 0.01fF
C961 a_3176_n2167# a_3077_n821# 0.00fF
C962 a_3077_n1909# a_3176_n1079# 0.00fF
C963 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.02fF
C964 a_4464_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C965 a_4661_n10301# VDD 0.35fF
C966 a_9706_n509# a_9616_n1079# 0.02fF
C967 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.03fF
C968 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_7237_n4317# 0.01fF
C969 a_2148_n10871# a_2085_n10301# 0.01fF
C970 a_9876_n3799# a_9706_n4317# 0.04fF
C971 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_4661_n13021# 0.01fF
C972 a_5949_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.02fF
C973 Ad_b a_6658_n7363# 0.06fF
C974 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C975 a_10904_n9783# a_10994_n10301# 0.01fF
C976 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X VDD 0.87fF
C977 a_9450_n6493# a_10738_n6173# 0.01fF
C978 a_4554_n1597# a_4554_n2685# 0.01fF
C979 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_4298_n10301# 0.00fF
C980 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.08fF
C981 a_5752_n8695# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C982 a_11101_n5405# a_11164_n3799# 0.00fF
C983 a_4554_n4317# a_4554_n2685# 0.01fF
C984 a_4464_n1079# a_4464_n2167# 0.01fF
C985 a_4365_n13413# a_6012_n13591# 0.00fF
C986 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.88fF
C987 a_5949_n2685# a_6012_n3255# 0.01fF
C988 a_9706_n2685# a_9876_n3799# 0.00fF
C989 a_10738_n8125# a_11101_n9213# 0.01fF
C990 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.09fF
C991 a_5653_n2997# a_5752_n3255# 0.49fF
C992 a_8162_n13021# a_8229_n11237# 0.00fF
C993 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.00fF
C994 a_690_n10301# a_501_n9525# 0.02fF
C995 a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.01fF
C996 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_3010_n1597# 0.03fF
C997 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.03fF
C998 a_1978_n4317# a_1978_n5405# 0.01fF
C999 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_8588_n3799# 0.00fF
C1000 a_434_n10301# a_600_n9783# 0.04fF
C1001 a_6941_n12325# a_7130_n11933# 0.02fF
C1002 a_7040_n12503# a_6874_n11933# 0.04fF
C1003 a_6941_n9525# a_7300_n9783# 0.05fF
C1004 a_5586_n13021# a_5653_n11237# 0.00fF
C1005 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C1006 a_8328_n10871# a_8418_n10301# 0.02fF
C1007 a_10738_n5405# VDD 0.69fF
C1008 a_3373_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.01fF
C1009 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3436_n1079# 0.03fF
C1010 a_434_n13021# a_1722_n13021# 0.01fF
C1011 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C1012 a_10738_n2685# a_10805_n2997# 0.01fF
C1013 a_8418_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.05fF
C1014 a_7040_n8695# a_6794_n7203# 0.00fF
C1015 a_9813_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.12fF
C1016 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_6665_n7459# 0.00fF
C1017 a_10904_n1079# a_11164_n1079# 0.23fF
C1018 a_10805_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.01fF
C1019 sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# 0.53fF
C1020 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4298_n4317# 0.01fF
C1021 a_4298_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C1022 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.04fF
C1023 a_797_n1597# a_797_n2685# 0.02fF
C1024 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C1025 a_5752_n2167# a_5653_n821# 0.00fF
C1026 a_5653_n1909# a_5752_n1079# 0.00fF
C1027 a_9813_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C1028 a_6874_n5405# a_6941_n3621# 0.00fF
C1029 a_9517_n4709# a_9876_n4887# 0.05fF
C1030 a_7040_n3799# VDD 0.44fF
C1031 sky130_fd_sc_hd__nand2_4_0/B a_10805_n821# 0.03fF
C1032 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A VDD 0.89fF
C1033 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_9706_n4317# 0.01fF
C1034 a_8328_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C1035 a_7130_n1597# a_7040_n3255# 0.00fF
C1036 sky130_fd_sc_hd__clkinv_1_0/A a_1888_n1079# 0.07fF
C1037 a_3373_n10301# a_4661_n10301# 0.01fF
C1038 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4554_n10301# 0.03fF
C1039 a_3266_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C1040 a_5586_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C1041 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5586_n2685# 0.01fF
C1042 a_1789_n8437# a_3077_n8437# 0.01fF
C1043 a_5752_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.03fF
C1044 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.03fF
C1045 a_9706_n509# a_9813_n509# 0.55fF
C1046 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5586_n2685# 0.00fF
C1047 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/B 0.08fF
C1048 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_6941_n13413# 0.01fF
C1049 a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.02fF
C1050 a_5752_n13591# a_6012_n13591# 0.28fF
C1051 a_4623_n7349# a_4464_n8695# 0.00fF
C1052 a_1888_n1079# a_2085_n2685# 0.00fF
C1053 a_7237_n1597# a_7300_n1079# 0.01fF
C1054 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6794_n7203# 0.00fF
C1055 a_2148_n1079# a_1978_n2685# 0.00fF
C1056 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C1057 a_600_n9783# VDD 0.47fF
C1058 a_5653_n2997# a_7300_n3255# 0.00fF
C1059 sky130_fd_sc_hd__clkinv_4_8/A a_11164_n13591# 0.12fF
C1060 a_11101_n5405# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C1061 a_690_n11933# a_600_n10871# 0.01fF
C1062 a_434_n1597# a_501_n821# 0.01fF
C1063 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C1064 a_9616_n3799# a_9517_n2997# 0.01fF
C1065 a_9450_n4317# VDD 0.76fF
C1066 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.04fF
C1067 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_8229_n9525# 0.18fF
C1068 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.13fF
C1069 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X 0.29fF
C1070 a_6874_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C1071 a_8418_n6493# a_8328_n4887# 0.00fF
C1072 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A p2 0.03fF
C1073 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X sky130_fd_sc_hd__clkinv_1_5/A 0.76fF
C1074 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C1075 a_n787_n12325# a_n428_n12503# 0.05fF
C1076 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.05fF
C1077 a_501_n2997# a_501_n3621# 0.05fF
C1078 a_11101_n9213# a_10994_n10301# 0.00fF
C1079 a_10994_n9213# a_11101_n10301# 0.00fF
C1080 a_501_n1909# a_860_n2167# 0.05fF
C1081 a_8525_n14109# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C1082 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.08fF
C1083 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9813_n14109# 0.02fF
C1084 a_9450_n2685# VDD 0.75fF
C1085 a_10738_n6173# a_10805_n5797# 0.03fF
C1086 a_3077_n12325# a_3266_n11933# 0.02fF
C1087 a_3176_n12503# a_3010_n11933# 0.04fF
C1088 a_4298_n5405# a_4365_n4709# 0.01fF
C1089 a_600_n12503# a_434_n13021# 0.04fF
C1090 a_4661_n5405# a_4661_n4317# 0.02fF
C1091 a_9616_n9783# VDD 0.45fF
C1092 a_860_n4887# a_690_n5405# 0.04fF
C1093 a_600_n4887# a_797_n5405# 0.02fF
C1094 a_797_n4317# a_600_n3255# 0.00fF
C1095 a_690_n4317# a_860_n3255# 0.00fF
C1096 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C1097 a_9706_n13021# a_9616_n13591# 0.01fF
C1098 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C1099 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_10805_n4709# 0.17fF
C1100 a_9876_n4887# a_10904_n4887# 0.02fF
C1101 a_8588_n3799# VDD 0.77fF
C1102 a_8418_n1597# a_9450_n1597# 0.02fF
C1103 a_8162_n1597# a_9706_n1597# 0.01fF
C1104 a_5586_n1597# a_7130_n1597# 0.01fF
C1105 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.02fF
C1106 a_10738_n509# a_10738_n1597# 0.01fF
C1107 a_1888_n8695# a_1722_n9213# 0.04fF
C1108 a_1789_n8437# a_1978_n9213# 0.02fF
C1109 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_1722_n4317# 0.00fF
C1110 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C1111 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_7300_n2167# 0.00fF
C1112 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.08fF
C1113 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11101_n4317# 0.12fF
C1114 a_3266_n4317# a_4298_n4317# 0.02fF
C1115 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8229_n2997# 0.00fF
C1116 a_8162_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C1117 a_3010_n4317# a_4554_n4317# 0.01fF
C1118 sky130_fd_sc_hd__clkinv_1_0/A a_3436_n1079# 0.12fF
C1119 a_5949_n1597# a_5949_n2685# 0.02fF
C1120 a_4365_n3621# a_5653_n3621# 0.01fF
C1121 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C1122 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X a_7300_n3255# 0.03fF
C1123 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C1124 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.05fF
C1125 a_8328_n11415# a_8162_n10301# 0.00fF
C1126 a_n787_n1909# VDD 0.35fF
C1127 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.02fF
C1128 sky130_fd_sc_hd__clkinv_1_0/A a_11101_n1597# 0.01fF
C1129 a_501_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.00fF
C1130 a_6874_n6493# a_7237_n6493# 0.05fF
C1131 sky130_fd_sc_hd__nand2_4_3/Y a_10904_n8695# 0.16fF
C1132 a_6012_n11415# a_4464_n11415# 0.01fF
C1133 a_5752_n11415# a_4724_n11415# 0.02fF
C1134 a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.18fF
C1135 a_5752_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C1136 a_5653_n2997# a_5842_n1597# 0.00fF
C1137 a_10904_n10871# a_10904_n11415# 0.07fF
C1138 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A p2 0.00fF
C1139 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.03fF
C1140 a_4661_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C1141 a_2148_n9783# VDD 0.78fF
C1142 a_5653_n10613# a_5752_n12503# 0.00fF
C1143 a_5752_n10871# a_5653_n12325# 0.00fF
C1144 a_3176_n3799# a_3176_n4887# 0.01fF
C1145 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1789_n10613# 0.00fF
C1146 a_11101_n2685# VDD 0.32fF
C1147 a_8328_n12503# a_8525_n11933# 0.02fF
C1148 a_1978_n10301# a_2148_n9783# 0.04fF
C1149 a_2085_n10301# a_1888_n9783# 0.02fF
C1150 a_8588_n12503# a_8418_n11933# 0.04fF
C1151 a_10994_n4317# VDD 0.44fF
C1152 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C1153 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.02fF
C1154 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C1155 a_8418_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C1156 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9517_n4709# 0.00fF
C1157 a_9450_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.00fF
C1158 a_3077_n5797# a_3077_n4709# 0.02fF
C1159 a_10994_n5405# a_9450_n5405# 0.01fF
C1160 a_10738_n5405# a_9706_n5405# 0.02fF
C1161 a_6941_n1909# a_7040_n3255# 0.00fF
C1162 a_7040_n2167# a_6941_n2997# 0.00fF
C1163 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.06fF
C1164 sky130_fd_sc_hd__clkinv_1_0/A a_5752_n1079# 0.07fF
C1165 a_3010_n1597# VDD 0.76fF
C1166 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkinv_4_4/A 0.89fF
C1167 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.02fF
C1168 a_7130_n4317# a_6941_n3621# 0.02fF
C1169 a_6874_n4317# a_7040_n3799# 0.04fF
C1170 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.04fF
C1171 a_11164_n9783# VDD 0.67fF
C1172 a_690_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C1173 a_797_n9213# a_2085_n9213# 0.01fF
C1174 a_8418_n5405# a_8328_n3799# 0.00fF
C1175 a_4298_n1597# a_4661_n1597# 0.05fF
C1176 a_3176_n10871# a_3266_n9213# 0.00fF
C1177 a_600_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.04fF
C1178 B_b a_13765_n2685# 0.06fF
C1179 a_9450_n1597# a_9813_n1597# 0.05fF
C1180 a_9616_n10871# a_9813_n11933# 0.00fF
C1181 a_13765_n1597# Bd_b 0.06fF
C1182 a_6874_n1597# a_7237_n1597# 0.05fF
C1183 a_797_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C1184 a_690_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C1185 a_797_n4317# a_2085_n4317# 0.01fF
C1186 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1978_n4317# 0.03fF
C1187 a_5949_n1597# a_6012_n3255# 0.00fF
C1188 a_4298_n4317# a_4661_n4317# 0.05fF
C1189 a_7040_n9783# a_7237_n9213# 0.02fF
C1190 a_8525_n1597# a_8588_n3255# 0.00fF
C1191 a_7300_n9783# a_7130_n9213# 0.04fF
C1192 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.84fF
C1193 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.29fF
C1194 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X p2 0.02fF
C1195 a_5653_n3621# a_5752_n3799# 0.49fF
C1196 Bd_b a_6665_n7459# 0.06fF
C1197 a_860_n3799# a_797_n5405# 0.00fF
C1198 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y 1.55fF
C1199 a_7040_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C1200 a_7130_n6493# a_8525_n6493# 0.01fF
C1201 a_7237_n6493# a_8418_n6493# 0.01fF
C1202 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n6493# 0.35fF
C1203 a_501_n5797# a_434_n4317# 0.00fF
C1204 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.06fF
C1205 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.08fF
C1206 a_1888_n10871# a_1978_n11933# 0.01fF
C1207 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VDD 0.90fF
C1208 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkinv_1_3/A 0.84fF
C1209 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C1210 a_8229_n12325# a_8162_n14109# 0.00fF
C1211 a_9813_n9213# VDD 0.33fF
C1212 a_9706_n2685# a_9616_n1079# 0.00fF
C1213 a_9876_n12503# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C1214 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_9813_n14109# 0.00fF
C1215 a_2148_n3255# a_501_n2997# 0.00fF
C1216 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.09fF
C1217 a_8162_n2685# a_8162_n4317# 0.01fF
C1218 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.29fF
C1219 sky130_fd_sc_hd__clkinv_1_0/A a_7300_n1079# 0.12fF
C1220 a_5842_n5405# a_5752_n4887# 0.02fF
C1221 a_4464_n12503# a_4661_n11933# 0.02fF
C1222 a_2148_n2167# VDD 0.78fF
C1223 a_1722_n13021# a_1978_n13021# 0.19fF
C1224 a_9813_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1225 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_9876_n3255# 0.00fF
C1226 a_1978_n4317# a_1888_n3799# 0.02fF
C1227 a_501_n4709# a_860_n4887# 0.05fF
C1228 a_n428_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C1229 a_10904_n3799# a_10805_n2997# 0.01fF
C1230 a_10805_n3621# a_10904_n3255# 0.01fF
C1231 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.02fF
C1232 a_5653_n3621# a_6012_n3799# 0.05fF
C1233 a_1888_n3255# a_1888_n4887# 0.00fF
C1234 a_6941_n9525# a_7130_n8125# 0.00fF
C1235 a_7040_n9783# a_6874_n8125# 0.00fF
C1236 a_9450_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C1237 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9517_n3621# 0.00fF
C1238 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5586_n1597# 0.35fF
C1239 a_4661_n1597# a_5842_n1597# 0.01fF
C1240 a_4554_n1597# a_5949_n1597# 0.01fF
C1241 a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.00fF
C1242 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_4298_n9213# 0.00fF
C1243 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C1244 a_10738_n1597# a_10805_n821# 0.01fF
C1245 sky130_fd_sc_hd__clkinv_4_8/Y a_11164_n12503# 0.01fF
C1246 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.01fF
C1247 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_3373_n9213# 0.01fF
C1248 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.03fF
C1249 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD 0.91fF
C1250 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_7237_n509# 0.01fF
C1251 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_7237_n8125# 0.01fF
C1252 a_434_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C1253 a_9876_n11415# a_9706_n11933# 0.04fF
C1254 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.29fF
C1255 a_7040_n8695# a_6874_n9213# 0.04fF
C1256 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.01fF
C1257 A p2 0.02fF
C1258 a_8525_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C1259 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_8588_n13591# 0.03fF
C1260 a_7130_n13021# a_7130_n11933# 0.01fF
C1261 a_9616_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C1262 a_8418_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.05fF
C1263 a_434_n9213# a_797_n9213# 0.05fF
C1264 a_4365_n12325# a_4464_n10871# 0.00fF
C1265 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_3010_n11933# 0.01fF
C1266 a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C1267 a_9706_n8125# a_10738_n8125# 0.01fF
C1268 a_434_n2685# a_501_n3621# 0.00fF
C1269 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.03fF
C1270 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_2085_n5405# 0.01fF
C1271 a_8162_n4317# a_9706_n4317# 0.01fF
C1272 sky130_fd_sc_hd__clkinv_4_10/Y VDD 2.17fF
C1273 a_8418_n4317# a_9450_n4317# 0.02fF
C1274 a_690_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.02fF
C1275 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_860_n4887# 0.02fF
C1276 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10805_n821# 0.00fF
C1277 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.05fF
C1278 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C1279 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_3436_n9783# 0.03fF
C1280 a_6874_n1597# a_7040_n2167# 0.04fF
C1281 a_5653_n11237# a_6012_n11415# 0.05fF
C1282 a_3373_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C1283 a_501_n1909# a_501_n2997# 0.02fF
C1284 a_1789_n13413# a_3176_n13591# 0.01fF
C1285 a_1888_n13591# a_3077_n13413# 0.01fF
C1286 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_1789_n2997# 0.02fF
C1287 a_690_n2685# a_797_n4317# 0.00fF
C1288 a_797_n2685# a_690_n4317# 0.00fF
C1289 a_3077_n8437# a_3436_n8695# 0.05fF
C1290 a_9876_n3799# VDD 0.74fF
C1291 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.08fF
C1292 a_6012_n13591# a_7040_n13591# 0.02fF
C1293 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_6941_n13413# 0.18fF
C1294 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.02fF
C1295 a_5949_n9213# a_7130_n9213# 0.01fF
C1296 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6874_n9213# 0.35fF
C1297 a_9706_n6493# a_10738_n6173# 0.01fF
C1298 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_3010_n5405# 0.00fF
C1299 a_2148_n3255# a_1978_n4317# 0.00fF
C1300 a_3436_n3799# a_3436_n3255# 0.09fF
C1301 a_2729_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.02fF
C1302 a_n787_n9525# a_n428_n9783# 0.05fF
C1303 a_860_n5975# VDD 0.80fF
C1304 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VDD 0.90fF
C1305 a_1978_n13021# a_3266_n13021# 0.01fF
C1306 a_8418_n4317# a_8588_n3799# 0.04fF
C1307 a_8525_n4317# a_8328_n3799# 0.02fF
C1308 a_1722_n13021# a_3373_n13021# 0.00fF
C1309 a_2085_n13021# a_3010_n13021# 0.02fF
C1310 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C1311 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.05fF
C1312 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.02fF
C1313 sky130_fd_sc_hd__clkinv_4_4/Y VDD 2.22fF
C1314 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.04fF
C1315 a_5752_n3799# a_7300_n3799# 0.01fF
C1316 a_9813_n5405# a_10738_n5405# 0.02fF
C1317 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C1318 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_2085_n11933# 0.00fF
C1319 a_1722_n13021# VDD 0.75fF
C1320 a_9616_n11415# a_9813_n10301# 0.00fF
C1321 a_5842_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.05fF
C1322 a_9876_n11415# a_9706_n10301# 0.00fF
C1323 a_5949_n10301# a_5842_n9213# 0.00fF
C1324 a_4724_n12503# VDD 0.78fF
C1325 a_6874_n10301# a_6874_n9213# 0.02fF
C1326 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C1327 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_9706_n11933# 0.01fF
C1328 a_6874_n2685# a_8162_n2685# 0.01fF
C1329 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.02fF
C1330 a_7040_n3255# a_7040_n4887# 0.00fF
C1331 a_11164_n5975# sky130_fd_sc_hd__nand2_4_1/A 0.04fF
C1332 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_2148_n8695# 0.03fF
C1333 a_9517_n12325# a_8229_n12325# 0.01fF
C1334 sky130_fd_sc_hd__nand2_4_3/Y a_10805_n9525# 0.08fF
C1335 sky130_fd_sc_hd__nand2_4_0/Y a_11164_n1079# 0.12fF
C1336 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_11101_n2685# 0.01fF
C1337 a_8162_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C1338 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.00fF
C1339 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_11164_n12503# 0.03fF
C1340 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n11933# 0.01fF
C1341 a_797_n9213# a_1978_n9213# 0.01fF
C1342 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1722_n9213# 0.35fF
C1343 a_3436_n10871# a_3373_n11933# 0.00fF
C1344 a_7130_n2685# a_7040_n3799# 0.01fF
C1345 a_434_n10301# a_1722_n10301# 0.01fF
C1346 a_3077_n9525# a_3266_n9213# 0.02fF
C1347 a_3176_n9783# a_3010_n9213# 0.04fF
C1348 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.06fF
C1349 a_4554_n11933# a_4661_n10301# 0.00fF
C1350 a_9813_n509# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C1351 a_4661_n11933# a_4554_n10301# 0.00fF
C1352 a_9517_n821# a_8229_n821# 0.01fF
C1353 a_5052_n7283# a_6665_n7459# 0.01fF
C1354 a_6012_n11415# a_7040_n11415# 0.02fF
C1355 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_6941_n11237# 0.18fF
C1356 a_5752_n11415# a_7300_n11415# 0.01fF
C1357 a_6006_n7607# a_6658_n7363# 0.03fF
C1358 a_6101_n7254# a_6373_n7349# 0.43fF
C1359 a_3077_n11237# a_3077_n10613# 0.05fF
C1360 a_5586_n10301# a_5653_n8437# 0.00fF
C1361 a_3077_n13413# a_3436_n13591# 0.05fF
C1362 a_501_n10613# a_690_n9213# 0.00fF
C1363 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_7040_n3799# 0.05fF
C1364 a_6012_n3799# a_7300_n3799# 0.01fF
C1365 a_7300_n8695# a_5653_n8437# 0.00fF
C1366 a_7040_n8695# a_5752_n8695# 0.01fF
C1367 a_8162_n6493# a_9813_n6493# 0.00fF
C1368 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A VDD 0.62fF
C1369 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VDD 0.86fF
C1370 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_4365_n8437# 0.18fF
C1371 a_3436_n8695# a_4464_n8695# 0.02fF
C1372 a_3176_n8695# a_4724_n8695# 0.01fF
C1373 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C1374 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_8328_n13591# 0.01fF
C1375 a_8229_n8437# a_9616_n8695# 0.01fF
C1376 a_8328_n8695# a_9517_n8437# 0.01fF
C1377 a_7040_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C1378 a_7130_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.05fF
C1379 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_8418_n9213# 0.00fF
C1380 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C1381 a_2148_n5975# a_1978_n4317# 0.00fF
C1382 a_1888_n5975# a_2085_n4317# 0.00fF
C1383 a_9616_n2167# a_9813_n1597# 0.02fF
C1384 a_9876_n2167# a_9706_n1597# 0.04fF
C1385 a_6101_n7254# VDD 0.83fF
C1386 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_4298_n13021# 0.00fF
C1387 a_3010_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.03fF
C1388 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_8525_n11933# 0.01fF
C1389 a_9813_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.02fF
C1390 a_3266_n13021# a_3373_n13021# 0.55fF
C1391 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_1789_n3621# 0.01fF
C1392 Bd_b sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C1393 sky130_fd_sc_hd__clkinv_1_0/Y a_2622_n509# 0.03fF
C1394 a_1888_n12503# a_2085_n13021# 0.02fF
C1395 a_2148_n12503# a_1978_n13021# 0.04fF
C1396 a_10994_n5405# a_11101_n5405# 0.55fF
C1397 a_10738_n5405# sky130_fd_sc_hd__clkinv_4_4/A 0.00fF
C1398 a_3266_n13021# VDD 0.46fF
C1399 a_4464_n10871# a_4298_n10301# 0.04fF
C1400 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.04fF
C1401 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.00fF
C1402 a_600_n12503# a_860_n12503# 0.28fF
C1403 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1404 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C1405 sky130_fd_sc_hd__clkinv_4_8/Y p1d_b 0.04fF
C1406 a_600_n12503# VDD 0.44fF
C1407 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_4661_n13021# 0.01fF
C1408 a_3010_n2685# a_3373_n2685# 0.05fF
C1409 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VDD 0.86fF
C1410 a_8162_n2685# a_8418_n2685# 0.19fF
C1411 a_10805_n10613# a_10904_n9783# 0.00fF
C1412 a_7237_n10301# a_7130_n11933# 0.00fF
C1413 a_6012_n8695# a_5949_n9213# 0.01fF
C1414 a_7130_n10301# a_7237_n11933# 0.00fF
C1415 a_10904_n10871# a_10805_n9525# 0.00fF
C1416 a_8588_n8695# a_8418_n9213# 0.04fF
C1417 a_8328_n8695# a_8525_n9213# 0.02fF
C1418 a_1722_n10301# VDD 0.76fF
C1419 a_8525_n13021# a_8525_n11933# 0.02fF
C1420 a_8328_n9783# a_8588_n9783# 0.28fF
C1421 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8229_n3621# 0.00fF
C1422 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C1423 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A a_600_n9783# 0.01fF
C1424 a_1722_n10301# a_1978_n10301# 0.19fF
C1425 a_1978_n2685# a_1888_n3799# 0.01fF
C1426 sky130_fd_sc_hd__nand2_1_4/Y VDD 1.03fF
C1427 a_501_n11237# a_600_n10871# 0.01fF
C1428 a_n787_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C1429 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_9517_n5797# 0.18fF
C1430 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.08fF
C1431 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.04fF
C1432 a_7130_n8125# a_7130_n9213# 0.01fF
C1433 a_7040_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.03fF
C1434 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_8328_n11415# 0.01fF
C1435 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_3010_n13021# 0.00fF
C1436 B_b VDD 4.27fF
C1437 a_5949_n5405# a_5752_n4887# 0.02fF
C1438 a_9876_n3799# a_9706_n5405# 0.00fF
C1439 a_3436_n13591# a_4464_n13591# 0.02fF
C1440 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_4365_n13413# 0.18fF
C1441 a_4464_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.03fF
C1442 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.04fF
C1443 a_3176_n13591# a_4724_n13591# 0.01fF
C1444 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.29fF
C1445 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_5752_n8695# 0.01fF
C1446 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_2622_n509# 0.04fF
C1447 a_2622_n14109# VDD 0.47fF
C1448 a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.01fF
C1449 a_9450_n6493# sky130_fd_sc_hd__nand2_4_1/B 0.03fF
C1450 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C1451 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_8588_n13591# 0.03fF
C1452 a_600_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C1453 a_9517_n8437# a_9876_n8695# 0.05fF
C1454 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_3176_n3799# 0.05fF
C1455 a_2148_n3799# a_3436_n3799# 0.01fF
C1456 a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.00fF
C1457 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8525_n9213# 0.02fF
C1458 a_7237_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C1459 a_1789_n11237# a_2148_n11415# 0.05fF
C1460 a_1978_n1597# a_1789_n821# 0.02fF
C1461 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.09fF
C1462 a_10904_n11415# a_11101_n13021# 0.00fF
C1463 sky130_fd_sc_hd__nand2_4_3/Y a_10994_n9213# 0.10fF
C1464 a_8525_n6493# a_8418_n8125# 0.00fF
C1465 a_8418_n6493# a_8525_n8125# 0.00fF
C1466 a_11164_n11415# a_10994_n13021# 0.00fF
C1467 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10738_n4317# 0.01fF
C1468 a_10738_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C1469 a_3373_n13021# a_4661_n13021# 0.01fF
C1470 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.06fF
C1471 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4554_n13021# 0.03fF
C1472 a_3266_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C1473 a_8328_n12503# a_8229_n13413# 0.00fF
C1474 a_8229_n12325# a_8328_n13591# 0.00fF
C1475 a_4464_n10871# a_3436_n10871# 0.02fF
C1476 a_5752_n9783# a_5752_n11415# 0.00fF
C1477 a_4724_n10871# a_3176_n10871# 0.01fF
C1478 a_6941_n8437# a_7300_n8695# 0.05fF
C1479 a_4661_n13021# VDD 0.35fF
C1480 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11101_n10301# 0.00fF
C1481 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__clkinv_1_3/Y 0.12fF
C1482 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.04fF
C1483 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_1888_n12503# 0.05fF
C1484 a_860_n12503# a_2148_n12503# 0.01fF
C1485 a_600_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C1486 a_8328_n8695# a_8162_n8125# 0.04fF
C1487 a_8229_n8437# a_8418_n8125# 0.02fF
C1488 a_4724_n3799# a_4724_n2167# 0.01fF
C1489 a_4464_n9783# a_4661_n10301# 0.02fF
C1490 a_2148_n12503# VDD 0.78fF
C1491 a_4724_n9783# a_4554_n10301# 0.04fF
C1492 a_3373_n2685# a_4554_n2685# 0.01fF
C1493 a_3266_n2685# a_4661_n2685# 0.01fF
C1494 a_10805_n13413# a_10738_n13021# 0.01fF
C1495 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4298_n2685# 0.35fF
C1496 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.02fF
C1497 a_434_n1597# a_1722_n1597# 0.01fF
C1498 a_8525_n2685# a_9450_n2685# 0.02fF
C1499 a_8162_n2685# a_9813_n2685# 0.00fF
C1500 a_8418_n2685# a_9706_n2685# 0.01fF
C1501 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.07fF
C1502 a_3266_n10301# VDD 0.44fF
C1503 a_2622_n14109# a_2729_n14109# 0.52fF
C1504 a_2366_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.02fF
C1505 a_2148_n3255# a_1978_n2685# 0.04fF
C1506 a_501_n1909# a_434_n2685# 0.01fF
C1507 a_600_n12503# a_501_n13413# 0.00fF
C1508 a_4298_n11933# a_5586_n11933# 0.01fF
C1509 a_8588_n9783# a_9876_n9783# 0.01fF
C1510 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_9616_n9783# 0.05fF
C1511 a_8328_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C1512 a_8229_n11237# a_8328_n12503# 0.00fF
C1513 a_8328_n11415# a_8229_n12325# 0.00fF
C1514 a_860_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.29fF
C1515 a_8525_n2685# a_8588_n3799# 0.00fF
C1516 a_8229_n1909# a_8418_n2685# 0.02fF
C1517 a_1722_n10301# a_3373_n10301# 0.00fF
C1518 a_8328_n2167# a_8162_n2685# 0.04fF
C1519 a_1978_n10301# a_3266_n10301# 0.01fF
C1520 a_2085_n10301# a_3010_n10301# 0.02fF
C1521 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_8588_n3255# 0.00fF
C1522 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C1523 a_7130_n509# a_7237_n1597# 0.00fF
C1524 a_7237_n509# a_7130_n1597# 0.00fF
C1525 a_8418_n10301# a_8418_n11933# 0.01fF
C1526 a_9616_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.03fF
C1527 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_10904_n5975# 0.01fF
C1528 a_5586_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.03fF
C1529 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C1530 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.05fF
C1531 a_8162_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C1532 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8162_n9213# 0.01fF
C1533 a_9813_n11933# a_9813_n13021# 0.02fF
C1534 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_8588_n11415# 0.03fF
C1535 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C1536 a_4464_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.03fF
C1537 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C1538 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.00fF
C1539 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X a_6012_n8695# 0.03fF
C1540 a_8162_n4317# a_8229_n5797# 0.00fF
C1541 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_5752_n13591# 0.01fF
C1542 a_9450_n509# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C1543 a_7237_n14109# VDD 0.32fF
C1544 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.02fF
C1545 a_10904_n10871# a_10994_n9213# 0.00fF
C1546 a_2148_n11415# a_3176_n11415# 0.02fF
C1547 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_3077_n11237# 0.18fF
C1548 a_1888_n11415# a_3436_n11415# 0.01fF
C1549 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C1550 a_9450_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.03fF
C1551 sky130_fd_sc_hd__mux2_1_0/X a_4365_n8437# 0.00fF
C1552 a_9706_n4317# a_9813_n4317# 0.55fF
C1553 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_3373_n4317# 0.00fF
C1554 a_10805_n12325# a_10904_n11415# 0.00fF
C1555 a_10904_n12503# a_10805_n11237# 0.00fF
C1556 a_9616_n1079# VDD 0.45fF
C1557 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A 0.81fF
C1558 a_4661_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.12fF
C1559 a_6941_n8437# a_7130_n10301# 0.00fF
C1560 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_11101_n10301# 0.01fF
C1561 a_11101_n5405# a_11101_n4317# 0.02fF
C1562 a_10994_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.10fF
C1563 a_5752_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.01fF
C1564 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_10994_n2685# 0.00fF
C1565 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_3373_n13021# 0.01fF
C1566 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.03fF
C1567 a_9706_n2685# a_9813_n4317# 0.00fF
C1568 a_9813_n2685# a_9706_n4317# 0.00fF
C1569 a_501_n8437# a_600_n9783# 0.00fF
C1570 a_8418_n13021# a_9813_n13021# 0.01fF
C1571 a_600_n8695# a_501_n9525# 0.00fF
C1572 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.29fF
C1573 a_6012_n10871# a_5842_n10301# 0.04fF
C1574 a_5752_n10871# a_5949_n10301# 0.02fF
C1575 a_7237_n10301# a_8525_n10301# 0.01fF
C1576 a_7130_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C1577 a_6874_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.03fF
C1578 a_9450_n5405# VDD 0.75fF
C1579 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VDD 0.86fF
C1580 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C1581 a_4554_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.05fF
C1582 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_5842_n2685# 0.00fF
C1583 a_1722_n1597# a_1978_n1597# 0.19fF
C1584 a_4365_n2997# a_4554_n2685# 0.02fF
C1585 a_4464_n3255# a_4298_n2685# 0.04fF
C1586 a_9706_n2685# a_9813_n2685# 0.55fF
C1587 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1588 a_9450_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.03fF
C1589 a_2085_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.01fF
C1590 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3373_n5405# 0.02fF
C1591 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_7130_n14109# 0.02fF
C1592 sky130_fd_sc_hd__nand2_4_1/B a_10805_n5797# 0.03fF
C1593 a_10738_n11933# sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C1594 a_434_n13021# a_690_n13021# 0.19fF
C1595 a_9876_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.29fF
C1596 a_8229_n4709# a_6941_n4709# 0.01fF
C1597 a_7130_n8125# a_8162_n8125# 0.02fF
C1598 a_6874_n8125# a_8418_n8125# 0.01fF
C1599 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.02fF
C1600 a_3266_n10301# a_3373_n10301# 0.55fF
C1601 a_3010_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.03fF
C1602 a_4365_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C1603 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_11164_n5975# 0.03fF
C1604 a_10994_n1597# a_10994_n2685# 0.01fF
C1605 a_5949_n4317# a_6012_n4887# 0.01fF
C1606 a_8525_n8125# a_8525_n9213# 0.02fF
C1607 sky130_fd_sc_hd__clkinv_4_8/A a_9813_n13021# 0.05fF
C1608 a_9616_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C1609 a_600_n12503# a_434_n11933# 0.04fF
C1610 a_3010_n1597# a_3077_n821# 0.01fF
C1611 a_6874_n13021# a_6941_n13413# 0.01fF
C1612 a_8588_n2167# a_8588_n3799# 0.01fF
C1613 a_8229_n1909# a_8328_n2167# 0.49fF
C1614 a_1789_n1909# a_1888_n1079# 0.00fF
C1615 a_5653_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C1616 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C1617 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_4464_n11415# 0.01fF
C1618 a_3176_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.03fF
C1619 sky130_fd_sc_hd__clkinv_4_8/A a_9706_n14109# 0.02fF
C1620 sky130_fd_sc_hd__nand2_4_0/A a_10994_n1597# 0.00fF
C1621 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10994_n4317# 0.03fF
C1622 sky130_fd_sc_hd__nand2_4_3/B a_10904_n8695# 0.02fF
C1623 a_9813_n4317# a_11101_n4317# 0.01fF
C1624 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.01fF
C1625 a_860_n10871# a_797_n10301# 0.01fF
C1626 a_11164_n1079# VDD 0.67fF
C1627 sky130_fd_sc_hd__dfxbp_1_0/Q a_4765_n7542# 0.02fF
C1628 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.02fF
C1629 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.08fF
C1630 a_9616_n9783# a_9706_n10301# 0.01fF
C1631 a_7300_n9783# a_7300_n11415# 0.01fF
C1632 a_9813_n5405# a_9876_n3799# 0.00fF
C1633 a_9706_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.01fF
C1634 a_9517_n11237# a_9616_n11415# 0.49fF
C1635 a_2085_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C1636 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_797_n5405# 0.01fF
C1637 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_11101_n2685# 0.02fF
C1638 a_501_n11237# a_501_n9525# 0.00fF
C1639 a_3266_n4317# a_3266_n2685# 0.01fF
C1640 a_8162_n4317# VDD 0.76fF
C1641 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_10994_n13021# 0.00fF
C1642 a_9706_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.05fF
C1643 a_7130_n509# a_7040_n2167# 0.00fF
C1644 a_4365_n3621# VDD 0.35fF
C1645 a_8162_n5405# a_9450_n5405# 0.01fF
C1646 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.02fF
C1647 a_9813_n509# VDD 0.35fF
C1648 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C1649 a_4661_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C1650 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5949_n2685# 0.02fF
C1651 a_6874_n13021# a_6941_n11237# 0.00fF
C1652 a_2085_n1597# a_3010_n1597# 0.02fF
C1653 a_1978_n1597# a_3266_n1597# 0.01fF
C1654 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C1655 a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C1656 a_n688_n2167# a_n428_n2167# 0.28fF
C1657 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.02fF
C1658 a_8162_n2685# a_8229_n821# 0.00fF
C1659 a_8328_n2167# sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C1660 a_9706_n13021# a_9813_n14109# 0.00fF
C1661 a_10738_n6173# a_10904_n4887# 0.00fF
C1662 a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.01fF
C1663 a_2729_n6493# sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C1664 sky130_fd_sc_hd__nand2_1_0/A VDD 1.58fF
C1665 a_5653_n12325# a_5842_n11933# 0.02fF
C1666 a_5653_n9525# a_6012_n9783# 0.05fF
C1667 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C1668 a_8418_n10301# a_9813_n10301# 0.01fF
C1669 a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C1670 a_8162_n8125# a_8525_n8125# 0.05fF
C1671 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C1672 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10805_n12325# 0.01fF
C1673 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C1674 a_9616_n1079# a_9876_n1079# 0.28fF
C1675 a_9517_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.02fF
C1676 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_10805_n821# 0.01fF
C1677 sky130_fd_sc_hd__clkinv_4_8/A a_9517_n12325# 0.07fF
C1678 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.03fF
C1679 a_3010_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C1680 a_4464_n3255# a_4365_n1909# 0.00fF
C1681 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3010_n4317# 0.01fF
C1682 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_11164_n2167# 0.03fF
C1683 a_860_n2167# a_860_n3799# 0.01fF
C1684 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_7/A 0.72fF
C1685 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_4724_n4887# 0.01fF
C1686 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C1687 a_10738_n9213# a_9706_n9213# 0.02fF
C1688 a_10994_n9213# a_9450_n9213# 0.01fF
C1689 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.00fF
C1690 a_10805_n13413# a_10904_n13591# 0.47fF
C1691 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.29fF
C1692 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_797_n5405# 0.01fF
C1693 sky130_fd_sc_hd__clkinv_1_5/A a_6794_n7203# 0.04fF
C1694 a_1789_n2997# a_1722_n4317# 0.00fF
C1695 a_8229_n4709# a_8588_n4887# 0.05fF
C1696 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.01fF
C1697 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_3/A 0.03fF
C1698 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11101_n4317# 0.00fF
C1699 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C1700 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_4724_n11415# 0.03fF
C1701 a_11101_n4317# sky130_fd_sc_hd__clkinv_4_3/A 0.01fF
C1702 a_8328_n10871# a_8328_n9783# 0.01fF
C1703 a_10805_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C1704 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X a_10738_n10301# 0.03fF
C1705 a_4298_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C1706 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4298_n2685# 0.01fF
C1707 a_6006_n7607# a_5842_n9213# 0.00fF
C1708 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.08fF
C1709 a_9517_n11237# a_11164_n11415# 0.00fF
C1710 a_8162_n4317# a_8162_n5405# 0.02fF
C1711 a_6941_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C1712 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4298_n2685# 0.00fF
C1713 a_4298_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C1714 a_9706_n13021# a_9616_n12503# 0.02fF
C1715 a_5752_n3799# VDD 0.44fF
C1716 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C1717 a_8162_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C1718 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C1719 a_9450_n5405# a_9706_n5405# 0.19fF
C1720 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.03fF
C1721 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_7237_n10301# 0.01fF
C1722 a_10738_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C1723 a_7130_n6493# a_6941_n4709# 0.00fF
C1724 a_6874_n6493# a_7040_n4887# 0.00fF
C1725 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.00fF
C1726 a_4365_n2997# a_6012_n3255# 0.00fF
C1727 a_4464_n3255# a_5752_n3255# 0.01fF
C1728 sky130_fd_sc_hd__clkinv_4_4/A a_860_n5975# 0.10fF
C1729 a_2148_n2167# a_2085_n1597# 0.01fF
C1730 a_1722_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C1731 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y 1.20fF
C1732 a_8328_n3799# a_8229_n2997# 0.01fF
C1733 a_8229_n3621# a_8328_n3255# 0.01fF
C1734 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_3077_n5797# 0.01fF
C1735 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VDD 0.86fF
C1736 a_5752_n9783# a_7300_n9783# 0.01fF
C1737 a_6012_n9783# a_7040_n9783# 0.02fF
C1738 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6941_n9525# 0.18fF
C1739 a_6665_n7459# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C1740 p2 a_7212_n7203# 0.01fF
C1741 a_6865_n7304# a_7041_n7581# 0.02fF
C1742 a_9450_n10301# a_10738_n10301# 0.01fF
C1743 sky130_fd_sc_hd__nand2_1_0/A a_n688_n4887# 0.04fF
C1744 a_4464_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.05fF
C1745 a_2148_n8695# a_2085_n9213# 0.01fF
C1746 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9450_n8125# 0.35fF
C1747 a_4724_n9783# a_3436_n9783# 0.01fF
C1748 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_3176_n9783# 0.00fF
C1749 a_9813_n9213# a_9706_n10301# 0.00fF
C1750 a_5752_n2167# a_5586_n2685# 0.04fF
C1751 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.03fF
C1752 a_8229_n1909# a_8229_n821# 0.02fF
C1753 a_1722_n2685# a_3266_n2685# 0.01fF
C1754 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.08fF
C1755 a_1978_n2685# a_3010_n2685# 0.02fF
C1756 a_5653_n1909# a_5842_n2685# 0.02fF
C1757 a_6874_n2685# VDD 0.76fF
C1758 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X a_10904_n1079# 0.05fF
C1759 a_1789_n12325# a_1978_n11933# 0.02fF
C1760 a_1888_n12503# a_1722_n11933# 0.04fF
C1761 a_9876_n1079# a_11164_n1079# 0.01fF
C1762 a_11101_n11933# a_11164_n12503# 0.01fF
C1763 a_9616_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.00fF
C1764 sky130_fd_sc_hd__clkinv_4_8/A a_10904_n12503# 0.07fF
C1765 a_3373_n5405# a_3373_n4317# 0.02fF
C1766 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.06fF
C1767 a_4724_n12503# a_4554_n11933# 0.04fF
C1768 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_9706_n9213# 0.01fF
C1769 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_9517_n4709# 0.18fF
C1770 a_8328_n4887# a_9876_n4887# 0.01fF
C1771 a_8588_n4887# a_9616_n4887# 0.02fF
C1772 a_8418_n13021# a_8328_n13591# 0.01fF
C1773 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkinv_1_5/A 0.13fF
C1774 a_6012_n3799# VDD 0.77fF
C1775 a_501_n821# a_860_n1079# 0.05fF
C1776 a_9813_n509# a_9876_n1079# 0.01fF
C1777 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkinv_1_3/A 0.88fF
C1778 sky130_fd_sc_hd__clkinv_1_6/Y clk 0.33fF
C1779 a_7130_n1597# a_8162_n1597# 0.02fF
C1780 a_4365_n1909# a_5653_n1909# 0.01fF
C1781 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_9813_n4317# 0.01fF
C1782 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.03fF
C1783 a_9450_n4317# a_9517_n2997# 0.00fF
C1784 a_6874_n4317# a_8162_n4317# 0.01fF
C1785 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.08fF
C1786 a_1722_n4317# a_3266_n4317# 0.01fF
C1787 a_1978_n4317# a_3010_n4317# 0.02fF
C1788 a_11164_n9783# a_11101_n10301# 0.01fF
C1789 a_4661_n1597# a_4661_n2685# 0.02fF
C1790 a_5653_n3621# a_5586_n4317# 0.01fF
C1791 a_6941_n11237# a_7130_n10301# 0.00fF
C1792 a_7040_n11415# a_6874_n10301# 0.00fF
C1793 a_3077_n3621# a_4365_n3621# 0.01fF
C1794 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.02fF
C1795 a_4661_n4317# a_4661_n2685# 0.01fF
C1796 a_9616_n3255# a_9616_n3799# 0.07fF
C1797 a_9616_n10871# a_9616_n11415# 0.07fF
C1798 a_4724_n1079# a_4724_n2167# 0.02fF
C1799 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.05fF
C1800 a_600_n3255# a_501_n4709# 0.00fF
C1801 a_4724_n13591# a_6012_n13591# 0.01fF
C1802 a_4365_n2997# a_4554_n1597# 0.00fF
C1803 a_501_n2997# a_600_n4887# 0.00fF
C1804 a_4464_n3255# a_4298_n1597# 0.00fF
C1805 a_4464_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C1806 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.08fF
C1807 a_9450_n2685# a_9517_n2997# 0.01fF
C1808 a_9813_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C1809 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9876_n3799# 0.01fF
C1810 a_4365_n2997# a_4554_n4317# 0.00fF
C1811 a_4464_n3255# a_4298_n4317# 0.00fF
C1812 a_8418_n13021# a_8328_n11415# 0.00fF
C1813 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_6941_n2997# 0.01fF
C1814 a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.02fF
C1815 a_9813_n11933# a_9876_n13591# 0.00fF
C1816 a_9706_n6493# sky130_fd_sc_hd__nand2_4_1/B 0.05fF
C1817 a_5653_n12325# a_5653_n13413# 0.02fF
C1818 a_7040_n12503# a_7237_n11933# 0.02fF
C1819 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkinv_1_4/Y 0.02fF
C1820 a_797_n10301# a_600_n9783# 0.02fF
C1821 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4365_n1909# 0.01fF
C1822 a_7300_n12503# a_7130_n11933# 0.04fF
C1823 a_690_n10301# a_860_n9783# 0.04fF
C1824 a_2622_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C1825 a_2622_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.08fF
C1826 a_7040_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.03fF
C1827 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8229_n4709# 0.00fF
C1828 a_8162_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C1829 a_1789_n5797# a_1789_n4709# 0.02fF
C1830 a_10738_n10301# a_10994_n10301# 0.19fF
C1831 a_11101_n5405# VDD 0.32fF
C1832 a_5653_n1909# a_5752_n3255# 0.00fF
C1833 a_434_n13021# a_2085_n13021# 0.00fF
C1834 a_690_n13021# a_1978_n13021# 0.01fF
C1835 a_434_n1597# VDD 0.76fF
C1836 a_10994_n2685# a_10904_n3255# 0.02fF
C1837 a_8418_n2685# VDD 0.44fF
C1838 a_11164_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.32fF
C1839 a_10994_n4317# a_10805_n2997# 0.00fF
C1840 a_10738_n4317# a_10904_n3255# 0.00fF
C1841 a_4298_n11933# VDD 0.76fF
C1842 a_8588_n9783# VDD 0.78fF
C1843 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.04fF
C1844 a_2366_n6493# a_2148_n4887# 0.00fF
C1845 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_10904_n4887# 0.01fF
C1846 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9517_n13413# 0.01fF
C1847 a_9616_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.03fF
C1848 a_9450_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C1849 a_7130_n5405# a_7040_n3799# 0.00fF
C1850 a_13765_n13021# VDD 2.23fF
C1851 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C1852 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD 0.84fF
C1853 sky130_fd_sc_hd__nand2_4_3/B a_10805_n9525# 0.01fF
C1854 a_8162_n1597# a_8525_n1597# 0.05fF
C1855 a_8162_n4317# a_8418_n4317# 0.19fF
C1856 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C1857 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkinv_4_3/A 0.02fF
C1858 a_5752_n9783# a_5949_n9213# 0.02fF
C1859 a_3010_n4317# a_3373_n4317# 0.05fF
C1860 a_7237_n1597# a_7300_n3255# 0.00fF
C1861 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.02fF
C1862 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.03fF
C1863 a_2148_n8695# a_3077_n8437# 0.02fF
C1864 a_1789_n8437# a_3436_n8695# 0.00fF
C1865 a_1888_n8695# a_3176_n8695# 0.01fF
C1866 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.84fF
C1867 a_4365_n3621# a_4464_n3799# 0.49fF
C1868 a_9813_n509# sky130_fd_sc_hd__nand2_4_0/B 0.13fF
C1869 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n6493# 0.33fF
C1870 a_4623_n7349# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C1871 a_5752_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C1872 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.00fF
C1873 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_2085_n2685# 0.00fF
C1874 sky130_fd_sc_hd__dfxbp_1_0/Q a_4724_n8695# 0.01fF
C1875 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.06fF
C1876 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VDD 0.91fF
C1877 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9517_n11237# 0.00fF
C1878 a_9450_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C1879 a_1722_n2685# a_1789_n2997# 0.01fF
C1880 a_797_n11933# a_860_n10871# 0.00fF
C1881 VDD a_9450_n11933# 0.76fF
C1882 B a_13765_n2685# 0.02fF
C1883 a_9813_n4317# VDD 0.33fF
C1884 a_7237_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C1885 a_9813_n5405# a_9450_n5405# 0.05fF
C1886 a_6874_n2685# a_6874_n4317# 0.01fF
C1887 a_6941_n10613# a_8229_n10613# 0.01fF
C1888 a_7040_n9783# a_7040_n8695# 0.01fF
C1889 a_8525_n6493# a_8588_n4887# 0.00fF
C1890 a_n688_n12503# a_501_n12325# 0.01fF
C1891 a_1722_n2685# a_1722_n4317# 0.01fF
C1892 sky130_fd_sc_hd__clkinv_1_0/A a_2366_n509# 0.01fF
C1893 Bd_b sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C1894 a_600_n3255# a_600_n3799# 0.07fF
C1895 a_4661_n13021# a_4554_n11933# 0.00fF
C1896 a_4554_n13021# a_4661_n11933# 0.00fF
C1897 a_600_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X 0.03fF
C1898 a_1978_n1597# VDD 0.45fF
C1899 a_10738_n6173# a_11164_n5975# 0.05fF
C1900 a_9813_n2685# VDD 0.34fF
C1901 sky130_fd_sc_hd__clkinv_4_8/A a_13765_n11933# 0.04fF
C1902 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X p2 0.03fF
C1903 a_3436_n12503# a_3266_n11933# 0.04fF
C1904 a_3176_n12503# a_3373_n11933# 0.02fF
C1905 a_4554_n5405# a_4464_n4887# 0.02fF
C1906 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.04fF
C1907 a_860_n12503# a_690_n13021# 0.04fF
C1908 a_690_n13021# VDD 0.47fF
C1909 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD 0.83fF
C1910 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.03fF
C1911 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_797_n5405# 0.01fF
C1912 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_860_n3255# 0.01fF
C1913 a_797_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C1914 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_3010_n9213# 0.00fF
C1915 a_8162_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C1916 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8229_n3621# 0.00fF
C1917 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.06fF
C1918 a_9450_n509# a_9517_n821# 0.01fF
C1919 a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C1920 a_3373_n1597# a_4554_n1597# 0.01fF
C1921 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4298_n1597# 0.35fF
C1922 a_10738_n8125# VDD 0.13fF
C1923 a_10738_n509# a_11101_n1597# 0.01fF
C1924 a_5949_n1597# a_7130_n1597# 0.01fF
C1925 a_5842_n1597# a_7237_n1597# 0.01fF
C1926 a_8525_n1597# a_9706_n1597# 0.01fF
C1927 a_8418_n1597# a_9813_n1597# 0.01fF
C1928 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9450_n1597# 0.35fF
C1929 a_8328_n2167# VDD 0.46fF
C1930 a_2148_n8695# a_1978_n9213# 0.04fF
C1931 a_9517_n11237# a_9517_n9525# 0.00fF
C1932 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4298_n4317# 0.35fF
C1933 a_3373_n4317# a_4554_n4317# 0.01fF
C1934 a_3266_n4317# a_4661_n4317# 0.01fF
C1935 a_9517_n1909# a_9517_n3621# 0.00fF
C1936 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.04fF
C1937 a_4464_n3799# a_5752_n3799# 0.01fF
C1938 a_4724_n3799# a_5653_n3621# 0.02fF
C1939 a_4365_n821# VDD 0.36fF
C1940 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A 0.97fF
C1941 a_7130_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.05fF
C1942 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_8418_n6493# 0.00fF
C1943 a_n428_n2167# VDD 0.83fF
C1944 sky130_fd_sc_hd__clkinv_4_8/A a_10738_n13789# 0.47fF
C1945 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 1.54fF
C1946 a_5842_n13021# a_5842_n11933# 0.01fF
C1947 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C1948 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_4724_n11415# 0.00fF
C1949 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C1950 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.01fF
C1951 a_11164_n10871# a_11164_n11415# 0.09fF
C1952 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_1722_n11933# 0.01fF
C1953 a_9450_n10301# VDD 0.75fF
C1954 a_4365_n9525# VDD 0.36fF
C1955 a_4365_n12325# a_4365_n13413# 0.02fF
C1956 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C1957 a_6941_n5797# a_8229_n5797# 0.01fF
C1958 a_9450_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.00fF
C1959 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9517_n821# 0.00fF
C1960 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X VDD 0.66fF
C1961 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_2148_n9783# 0.03fF
C1962 a_5842_n1597# a_5653_n1909# 0.02fF
C1963 a_2085_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C1964 a_5586_n1597# a_5752_n2167# 0.04fF
C1965 sky130_fd_sc_hd__clkinv_4_3/A VDD 7.49fF
C1966 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X a_8525_n11933# 0.01fF
C1967 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.03fF
C1968 a_7040_n9783# a_6874_n10301# 0.04fF
C1969 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/A 0.46fF
C1970 sky130_fd_sc_hd__nand2_4_3/B a_10994_n9213# 0.00fF
C1971 a_6941_n9525# a_7130_n10301# 0.02fF
C1972 a_8229_n10613# a_8328_n10871# 0.49fF
C1973 a_3176_n5975# a_3176_n4887# 0.01fF
C1974 a_11101_n5405# a_9706_n5405# 0.01fF
C1975 a_n1738_n6671# a_n2248_n7037# 0.02fF
C1976 a_13765_n5949# a_13765_n4861# 0.07fF
C1977 a_10805_n1909# a_10738_n2685# 0.01fF
C1978 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.84fF
C1979 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5653_n4709# 0.01fF
C1980 a_5586_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.03fF
C1981 a_7130_n4317# a_7300_n3799# 0.04fF
C1982 a_7237_n4317# a_7040_n3799# 0.02fF
C1983 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__clkinv_1_4/Y 0.01fF
C1984 a_797_n13021# a_1722_n13021# 0.02fF
C1985 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VDD 1.94fF
C1986 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X a_7300_n1079# 0.01fF
C1987 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C1988 a_1722_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C1989 a_4464_n3799# a_6012_n3799# 0.01fF
C1990 a_8525_n5405# a_8588_n3799# 0.00fF
C1991 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C1992 sky130_fd_sc_hd__nand2_4_1/B p2 0.04fF
C1993 a_3436_n10871# a_3373_n9213# 0.00fF
C1994 a_4554_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.05fF
C1995 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_5842_n1597# 0.00fF
C1996 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_3077_n2997# 0.18fF
C1997 a_2148_n3255# a_3176_n3255# 0.02fF
C1998 a_7130_n9213# a_7212_n7203# 0.00fF
C1999 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C2000 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C2001 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_9813_n11933# 0.00fF
C2002 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_8418_n1597# 0.00fF
C2003 a_9706_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.05fF
C2004 a_4554_n10301# a_4661_n9213# 0.00fF
C2005 a_4661_n10301# a_4554_n9213# 0.00fF
C2006 a_1789_n1909# a_1789_n3621# 0.00fF
C2007 a_4298_n4317# a_4365_n4709# 0.01fF
C2008 a_434_n13021# a_600_n13591# 0.04fF
C2009 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.02fF
C2010 a_2366_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C2011 a_690_n13021# a_501_n13413# 0.02fF
C2012 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.02fF
C2013 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C2014 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.03fF
C2015 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_7237_n9213# 0.01fF
C2016 a_9450_n509# a_9706_n509# 0.19fF
C2017 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A p2 0.04fF
C2018 a_4554_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.05fF
C2019 a_5752_n3255# a_5752_n4887# 0.00fF
C2020 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8525_n6493# 0.02fF
C2021 a_7237_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C2022 a_600_n5975# a_690_n4317# 0.00fF
C2023 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n11933# 0.01fF
C2024 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C2025 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C2026 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_434_n9213# 0.43fF
C2027 a_1888_n10871# a_1722_n9213# 0.00fF
C2028 a_1789_n10613# a_1978_n9213# 0.00fF
C2029 a_6941_n10613# VDD 0.35fF
C2030 a_10994_n10301# VDD 0.42fF
C2031 a_2148_n10871# a_2085_n11933# 0.00fF
C2032 Ad_b a_4661_n9213# 0.00fF
C2033 a_8229_n5797# a_8328_n5975# 0.49fF
C2034 a_8328_n12503# a_8418_n14109# 0.00fF
C2035 a_4724_n5975# Ad_b 0.00fF
C2036 a_9517_n8437# a_10805_n8437# 0.01fF
C2037 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_501_n4709# 0.01fF
C2038 a_9813_n2685# a_9876_n1079# 0.00fF
C2039 a_9706_n5405# a_9813_n4317# 0.00fF
C2040 a_8162_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.08fF
C2041 a_1789_n11237# a_1789_n10613# 0.05fF
C2042 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6012_n8695# 0.01fF
C2043 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.01fF
C2044 a_1789_n13413# a_2148_n13591# 0.05fF
C2045 a_4298_n10301# a_4365_n8437# 0.00fF
C2046 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_600_n3255# 0.00fF
C2047 a_2148_n3255# a_860_n3255# 0.01fF
C2048 a_n428_n4887# a_n787_n4709# 0.05fF
C2049 a_1888_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C2050 a_8418_n2685# a_8418_n4317# 0.01fF
C2051 a_7040_n8695# a_8229_n8437# 0.01fF
C2052 a_9517_n4709# a_9517_n3621# 0.02fF
C2053 a_6941_n5797# VDD 0.35fF
C2054 a_8229_n821# VDD 0.35fF
C2055 p2 sky130_fd_sc_hd__clkinv_1_3/A 0.24fF
C2056 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_3010_n13021# 0.00fF
C2057 a_1722_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.03fF
C2058 a_1978_n13021# a_2085_n13021# 0.55fF
C2059 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_7040_n3799# 0.01fF
C2060 a_600_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.03fF
C2061 a_5752_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.03fF
C2062 a_1888_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C2063 a_600_n12503# a_797_n13021# 0.02fF
C2064 a_7300_n9783# a_7130_n8125# 0.00fF
C2065 a_7040_n9783# a_7237_n8125# 0.00fF
C2066 a_4365_n12325# a_4464_n11415# 0.00fF
C2067 a_4464_n12503# a_4365_n11237# 0.00fF
C2068 a_9813_n6493# a_9616_n4887# 0.00fF
C2069 a_4661_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C2070 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_4464_n3255# 0.01fF
C2071 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5949_n1597# 0.02fF
C2072 a_2148_n3799# a_1789_n3621# 0.05fF
C2073 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C2074 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_1722_n5405# 0.03fF
C2075 a_10738_n11933# a_11101_n11933# 0.05fF
C2076 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.13fF
C2077 a_10994_n1597# a_10904_n1079# 0.01fF
C2078 a_5842_n10301# a_5949_n11933# 0.00fF
C2079 a_5949_n10301# a_5842_n11933# 0.00fF
C2080 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkinv_1_5/A 0.12fF
C2081 a_9517_n10613# a_9616_n9783# 0.00fF
C2082 a_9616_n10871# a_9517_n9525# 0.00fF
C2083 a_6874_n2685# a_7130_n2685# 0.19fF
C2084 a_7040_n8695# a_7237_n9213# 0.02fF
C2085 a_7300_n8695# a_7130_n9213# 0.04fF
C2086 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C2087 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_9876_n5975# 0.01fF
C2088 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C2089 a_860_n1079# a_1789_n821# 0.02fF
C2090 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Bd_b 0.07fF
C2091 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.09fF
C2092 a_5842_n13021# a_5653_n13413# 0.02fF
C2093 sky130_fd_sc_hd__nand2_4_3/Y a_9616_n9783# 0.05fF
C2094 a_7237_n13021# a_7237_n11933# 0.02fF
C2095 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6012_n4887# 0.01fF
C2096 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C2097 a_690_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.05fF
C2098 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_1978_n9213# 0.00fF
C2099 a_8328_n10871# VDD 0.46fF
C2100 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.01fF
C2101 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9450_n4317# 0.35fF
C2102 a_690_n2685# a_600_n3799# 0.01fF
C2103 a_434_n10301# a_690_n10301# 0.19fF
C2104 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C2105 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_7300_n12503# 0.00fF
C2106 a_8418_n4317# a_9813_n4317# 0.01fF
C2107 a_8525_n4317# a_9706_n4317# 0.01fF
C2108 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X a_9450_n14109# 0.00fF
C2109 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C2110 a_9706_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.08fF
C2111 a_5752_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.03fF
C2112 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.10fF
C2113 a_1888_n13591# a_3436_n13591# 0.01fF
C2114 a_3176_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.03fF
C2115 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.29fF
C2116 a_2148_n13591# a_3176_n13591# 0.02fF
C2117 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_3077_n13413# 0.18fF
C2118 a_600_n2167# a_600_n3255# 0.01fF
C2119 a_9450_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C2120 a_434_n1597# a_600_n1079# 0.04fF
C2121 a_8229_n8437# a_8588_n8695# 0.05fF
C2122 a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.17fF
C2123 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_7300_n13591# 0.03fF
C2124 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C2125 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_7237_n9213# 0.02fF
C2126 a_5949_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C2127 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.01fF
C2128 a_8328_n5975# VDD 0.44fF
C2129 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.09fF
C2130 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C2131 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_2085_n4317# 0.00fF
C2132 a_7237_n6493# a_7130_n8125# 0.00fF
C2133 a_9616_n11415# a_9813_n13021# 0.00fF
C2134 a_7130_n6493# a_7237_n8125# 0.00fF
C2135 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.02fF
C2136 a_2085_n13021# a_3373_n13021# 0.01fF
C2137 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3266_n13021# 0.03fF
C2138 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_600_n3799# 0.04fF
C2139 a_1978_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C2140 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8588_n3799# 0.03fF
C2141 a_8525_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C2142 a_7040_n12503# a_6941_n13413# 0.00fF
C2143 a_6941_n12325# a_7040_n13591# 0.00fF
C2144 a_8525_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.01fF
C2145 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10994_n5405# 0.03fF
C2146 a_9813_n5405# a_11101_n5405# 0.01fF
C2147 a_2085_n13021# VDD 0.34fF
C2148 sky130_fd_sc_hd__nand2_4_1/B a_10904_n4887# 0.00fF
C2149 a_7040_n8695# a_6874_n8125# 0.04fF
C2150 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C2151 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_9813_n10301# 0.00fF
C2152 B VDD 4.22fF
C2153 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11164_n3799# 0.00fF
C2154 a_7130_n10301# a_7130_n9213# 0.01fF
C2155 a_7130_n2685# a_8418_n2685# 0.01fF
C2156 a_7237_n2685# a_8162_n2685# 0.02fF
C2157 a_6874_n2685# a_8525_n2685# 0.00fF
C2158 a_9876_n12503# a_8229_n12325# 0.00fF
C2159 a_9517_n12325# a_8588_n12503# 0.02fF
C2160 a_9616_n12503# a_8328_n12503# 0.01fF
C2161 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.03fF
C2162 a_690_n10301# VDD 0.45fF
C2163 a_3010_n11933# a_4298_n11933# 0.01fF
C2164 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_860_n3799# 0.01fF
C2165 sky130_fd_sc_hd__nand2_4_3/Y a_11164_n9783# 0.11fF
C2166 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C2167 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__clkinv_4_3/A 0.02fF
C2168 a_7040_n11415# a_6941_n12325# 0.00fF
C2169 a_6941_n11237# a_7040_n12503# 0.00fF
C2170 a_7237_n2685# a_7300_n3799# 0.00fF
C2171 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.03fF
C2172 a_797_n10301# a_1722_n10301# 0.02fF
C2173 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1789_n3621# 0.00fF
C2174 a_1722_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C2175 a_690_n10301# a_1978_n10301# 0.01fF
C2176 a_434_n10301# a_2085_n10301# 0.00fF
C2177 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_10994_n4317# 0.00fF
C2178 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C2179 a_3266_n5405# a_3077_n4709# 0.02fF
C2180 a_3010_n5405# a_3176_n4887# 0.04fF
C2181 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_7300_n3255# 0.00fF
C2182 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C2183 a_3436_n9783# a_3266_n9213# 0.04fF
C2184 a_3176_n9783# a_3373_n9213# 0.02fF
C2185 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.10fF
C2186 a_9616_n1079# a_8328_n1079# 0.01fF
C2187 a_9517_n821# a_8588_n1079# 0.02fF
C2188 a_3176_n11415# a_3176_n10871# 0.07fF
C2189 a_9876_n1079# a_8229_n821# 0.00fF
C2190 a_6874_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C2191 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.03fF
C2192 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C2193 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_7300_n11415# 0.03fF
C2194 a_5052_n7283# a_6794_n7203# 0.01fF
C2195 a_6373_n7349# a_6658_n7363# 0.11fF
C2196 a_6101_n7254# a_6665_n7459# 0.13fF
C2197 a_6006_n7607# a_6865_n7304# 0.02fF
C2198 a_5842_n10301# a_5752_n8695# 0.00fF
C2199 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C2200 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_4464_n13591# 0.01fF
C2201 a_3176_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.03fF
C2202 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C2203 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_4724_n8695# 0.03fF
C2204 a_11164_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.00fF
C2205 a_6874_n4317# a_6941_n5797# 0.00fF
C2206 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_5752_n8695# 0.00fF
C2207 a_4365_n11237# a_4554_n10301# 0.00fF
C2208 a_4464_n11415# a_4298_n10301# 0.00fF
C2209 a_8525_n6493# a_9813_n6493# 0.01fF
C2210 a_7300_n8695# a_6012_n8695# 0.01fF
C2211 a_8328_n8695# a_8162_n10301# 0.00fF
C2212 a_8418_n6493# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C2213 a_6874_n509# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C2214 a_7040_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.05fF
C2215 a_8328_n8695# a_9876_n8695# 0.01fF
C2216 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_9517_n8437# 0.18fF
C2217 a_8588_n8695# a_9616_n8695# 0.02fF
C2218 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C2219 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_1789_n11237# 0.18fF
C2220 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_2085_n4317# 0.00fF
C2221 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.02fF
C2222 a_8418_n5405# a_8229_n5797# 0.02fF
C2223 a_8162_n5405# a_8328_n5975# 0.04fF
C2224 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.03fF
C2225 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C2226 a_9517_n12325# a_9616_n11415# 0.00fF
C2227 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_9813_n1597# 0.01fF
C2228 a_10904_n2167# a_10805_n3621# 0.00fF
C2229 sky130_fd_sc_hd__nand2_4_3/Y a_9813_n9213# 0.05fF
C2230 a_6658_n7363# VDD 1.30fF
C2231 a_1722_n9213# a_1789_n9525# 0.01fF
C2232 a_10805_n1909# a_10904_n3799# 0.00fF
C2233 a_3373_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.12fF
C2234 a_9813_n5405# a_9813_n4317# 0.02fF
C2235 a_1888_n5975# a_501_n5797# 0.01fF
C2236 a_4464_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C2237 a_1789_n5797# a_600_n5975# 0.01fF
C2238 a_11101_n5405# sky130_fd_sc_hd__clkinv_4_4/A 0.01fF
C2239 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_2085_n13021# 0.01fF
C2240 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.03fF
C2241 a_5586_n11933# a_6874_n11933# 0.01fF
C2242 a_3077_n8437# a_3077_n9525# 0.02fF
C2243 a_4724_n10871# a_4554_n10301# 0.04fF
C2244 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2245 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X VDD 0.87fF
C2246 a_4464_n10871# a_4661_n10301# 0.02fF
C2247 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.29fF
C2248 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VDD 0.86fF
C2249 a_6874_n5405# VDD 0.76fF
C2250 a_3266_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.05fF
C2251 a_13765_n1597# B_b 2.55fF
C2252 a_434_n1597# a_690_n1597# 0.19fF
C2253 clk sky130_fd_sc_hd__clkinv_1_4/Y 0.09fF
C2254 a_1888_n4887# a_1722_n5405# 0.04fF
C2255 a_1888_n3255# a_1978_n1597# 0.00fF
C2256 a_1789_n4709# a_1978_n5405# 0.02fF
C2257 a_3077_n2997# a_3266_n2685# 0.02fF
C2258 a_3176_n3255# a_3010_n2685# 0.04fF
C2259 a_8418_n2685# a_8525_n2685# 0.55fF
C2260 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.06fF
C2261 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.03fF
C2262 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_9450_n2685# 0.00fF
C2263 a_1789_n821# a_3176_n1079# 0.01fF
C2264 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.04fF
C2265 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n9213# 0.01fF
C2266 a_8162_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C2267 a_5653_n3621# a_5586_n5405# 0.00fF
C2268 a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C2269 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.03fF
C2270 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_8525_n9213# 0.01fF
C2271 a_2085_n10301# VDD 0.35fF
C2272 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2622_n14109# 0.03fF
C2273 a_4298_n11933# a_4554_n11933# 0.19fF
C2274 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.04fF
C2275 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.29fF
C2276 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C2277 a_1722_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C2278 a_1978_n10301# a_2085_n10301# 0.55fF
C2279 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_3010_n10301# 0.00fF
C2280 a_n428_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.27fF
C2281 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_9876_n5975# 0.03fF
C2282 a_434_n9213# sky130_fd_sc_hd__clkinv_1_3/A 0.00fF
C2283 a_13765_n13021# p1_b 2.54fF
C2284 a_7237_n8125# a_7237_n9213# 0.02fF
C2285 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C2286 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.02fF
C2287 a_6874_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.00fF
C2288 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_100/A 0.00fF
C2289 a_3010_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C2290 a_8162_n11933# a_9450_n11933# 0.01fF
C2291 a_9706_n8125# a_9813_n8125# 0.55fF
C2292 a_5949_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C2293 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6012_n4887# 0.03fF
C2294 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_4724_n13591# 0.03fF
C2295 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C2296 a_10805_n10613# a_10738_n10301# 0.01fF
C2297 a_8418_n509# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C2298 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VDD 1.92fF
C2299 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_797_n4317# 0.00fF
C2300 a_3077_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C2301 a_9616_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.03fF
C2302 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.02fF
C2303 a_1888_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.03fF
C2304 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_10738_n9213# 0.00fF
C2305 a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C2306 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_3176_n11415# 0.01fF
C2307 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_3436_n3799# 0.00fF
C2308 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C2309 a_2366_n8125# VDD 0.80fF
C2310 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_10/Y 0.19fF
C2311 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11101_n13021# 0.00fF
C2312 a_9813_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.05fF
C2313 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.02fF
C2314 a_n2436_n7037# a_n1738_n6671# 0.38fF
C2315 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.03fF
C2316 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_3436_n10871# 0.00fF
C2317 a_6012_n9783# a_6012_n11415# 0.01fF
C2318 a_5586_n4317# VDD 0.76fF
C2319 a_10805_n1909# a_10738_n509# 0.01fF
C2320 a_8328_n8695# a_8525_n8125# 0.02fF
C2321 a_8588_n8695# a_8418_n8125# 0.04fF
C2322 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.04fF
C2323 a_6874_n5405# a_8162_n5405# 0.01fF
C2324 a_9517_n9525# a_9706_n9213# 0.02fF
C2325 a_9616_n9783# a_9450_n9213# 0.04fF
C2326 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.02fF
C2327 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C2328 a_8418_n5405# VDD 0.47fF
C2329 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C2330 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_4661_n10301# 0.01fF
C2331 a_3373_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C2332 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4661_n2685# 0.02fF
C2333 a_690_n1597# a_1978_n1597# 0.01fF
C2334 a_797_n1597# a_1722_n1597# 0.02fF
C2335 a_434_n1597# a_2085_n1597# 0.00fF
C2336 a_8525_n2685# a_9813_n2685# 0.01fF
C2337 a_8418_n13021# a_8525_n14109# 0.00fF
C2338 a_8525_n13021# a_8418_n14109# 0.00fF
C2339 a_8418_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C2340 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9706_n2685# 0.03fF
C2341 a_6874_n2685# a_6941_n821# 0.00fF
C2342 a_9813_n6493# a_9876_n5975# 0.01fF
C2343 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2344 a_2729_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.12fF
C2345 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A VDD 0.89fF
C2346 a_4661_n11933# a_5586_n11933# 0.02fF
C2347 a_600_n2167# a_690_n2685# 0.01fF
C2348 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_2085_n2685# 0.01fF
C2349 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.03fF
C2350 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.02fF
C2351 a_600_n13591# VDD 0.46fF
C2352 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.03fF
C2353 a_10904_n4887# a_10805_n3621# 0.00fF
C2354 a_9450_n509# sky130_fd_sc_hd__nand2_4_0/Y 0.01fF
C2355 a_10805_n4709# a_10904_n3799# 0.00fF
C2356 a_6874_n8125# a_7237_n8125# 0.05fF
C2357 a_1978_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.01fF
C2358 a_2085_n10301# a_3373_n10301# 0.01fF
C2359 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3266_n10301# 0.03fF
C2360 a_8588_n2167# a_8418_n2685# 0.04fF
C2361 a_8328_n2167# a_8525_n2685# 0.02fF
C2362 a_2366_n6493# VDD 0.79fF
C2363 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_3436_n4887# 0.01fF
C2364 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.04fF
C2365 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C2366 a_10805_n5797# a_10738_n4317# 0.00fF
C2367 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C2368 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C2369 a_9450_n11933# a_9706_n11933# 0.19fF
C2370 a_8418_n4317# a_8328_n5975# 0.00fF
C2371 a_434_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C2372 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X Ad_b 0.02fF
C2373 a_4464_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C2374 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C2375 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_3436_n11415# 0.03fF
C2376 a_11164_n10871# a_11101_n9213# 0.00fF
C2377 a_9517_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C2378 a_9813_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.12fF
C2379 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VDD 0.76fF
C2380 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_9450_n10301# 0.03fF
C2381 a_3077_n2997# a_1789_n2997# 0.01fF
C2382 a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C2383 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.03fF
C2384 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_3/A 0.73fF
C2385 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.07fF
C2386 a_8229_n11237# a_9876_n11415# 0.00fF
C2387 a_8328_n11415# a_9616_n11415# 0.01fF
C2388 a_7130_n4317# VDD 0.47fF
C2389 a_6874_n4317# a_6874_n5405# 0.02fF
C2390 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__nand2_4_0/Y 0.06fF
C2391 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3010_n2685# 0.00fF
C2392 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6941_n1909# 0.00fF
C2393 a_8525_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C2394 a_6874_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C2395 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.03fF
C2396 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_5949_n10301# 0.01fF
C2397 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9813_n13021# 0.02fF
C2398 a_3176_n3799# VDD 0.44fF
C2399 a_3176_n11415# a_3077_n9525# 0.00fF
C2400 a_3077_n11237# a_3176_n9783# 0.00fF
C2401 a_10805_n13413# a_10805_n12325# 0.02fF
C2402 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.02fF
C2403 a_8162_n5405# a_8418_n5405# 0.19fF
C2404 a_3077_n821# a_4365_n821# 0.01fF
C2405 a_9517_n4709# a_11164_n4887# 0.00fF
C2406 a_1978_n1597# a_2085_n1597# 0.55fF
C2407 a_3077_n1909# a_3010_n2685# 0.01fF
C2408 a_1722_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.03fF
C2409 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_3010_n1597# 0.00fF
C2410 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/A 0.12fF
C2411 a_4724_n3255# a_4554_n2685# 0.04fF
C2412 a_4464_n3255# a_4661_n2685# 0.02fF
C2413 a_9813_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.12fF
C2414 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__nand2_1_0/A 0.19fF
C2415 a_6941_n3621# a_7040_n3255# 0.01fF
C2416 a_7040_n3799# a_6941_n2997# 0.01fF
C2417 a_11101_n11933# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C2418 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_1722_n2685# 0.03fF
C2419 a_8418_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.05fF
C2420 a_8328_n4887# a_7040_n4887# 0.01fF
C2421 a_8588_n4887# a_6941_n4709# 0.00fF
C2422 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8162_n8125# 0.35fF
C2423 a_7130_n8125# a_8525_n8125# 0.01fF
C2424 a_7237_n8125# a_8418_n8125# 0.01fF
C2425 a_600_n3255# a_1789_n2997# 0.01fF
C2426 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C2427 a_3373_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.12fF
C2428 a_4464_n2167# a_4298_n2685# 0.04fF
C2429 sky130_fd_sc_hd__nand2_1_4/Y a_3010_n9213# 0.00fF
C2430 a_1789_n8437# a_2148_n8695# 0.05fF
C2431 sky130_fd_sc_hd__nand2_4_0/Y a_10994_n1597# 0.10fF
C2432 a_3077_n5797# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C2433 a_2085_n5405# a_2085_n4317# 0.02fF
C2434 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_9616_n1079# 0.05fF
C2435 a_9813_n11933# a_9876_n12503# 0.01fF
C2436 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.06fF
C2437 a_11101_n1597# a_11101_n2685# 0.02fF
C2438 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.04fF
C2439 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkinv_1_4/Y 0.21fF
C2440 a_9813_n9213# a_9450_n9213# 0.05fF
C2441 a_3266_n1597# a_3176_n1079# 0.01fF
C2442 a_600_n12503# a_797_n11933# 0.02fF
C2443 a_860_n12503# a_690_n11933# 0.04fF
C2444 a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C2445 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.05fF
C2446 a_690_n11933# VDD 0.48fF
C2447 a_501_n13413# a_600_n13591# 0.48fF
C2448 a_7130_n13021# a_7040_n13591# 0.01fF
C2449 a_7300_n4887# a_8328_n4887# 0.02fF
C2450 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_8229_n4709# 0.18fF
C2451 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C2452 a_8328_n2167# a_8588_n2167# 0.28fF
C2453 a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.02fF
C2454 a_6012_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C2455 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/A 0.82fF
C2456 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1789_n4709# 0.01fF
C2457 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/B 0.44fF
C2458 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.08fF
C2459 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkinv_4_3/A 0.06fF
C2460 a_5752_n10871# a_5586_n11933# 0.00fF
C2461 a_5586_n4317# a_6874_n4317# 0.01fF
C2462 a_9876_n9783# a_9813_n10301# 0.01fF
C2463 a_3373_n1597# a_3373_n2685# 0.02fF
C2464 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C2465 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_10805_n11237# 0.01fF
C2466 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.02fF
C2467 a_600_n11415# a_600_n9783# 0.00fF
C2468 a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C2469 a_5752_n11415# a_5586_n10301# 0.00fF
C2470 a_5653_n11237# a_5842_n10301# 0.00fF
C2471 a_8525_n4317# VDD 0.35fF
C2472 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.01fF
C2473 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9517_n12325# 0.01fF
C2474 a_3373_n4317# a_3373_n2685# 0.01fF
C2475 a_10805_n1909# a_10805_n821# 0.02fF
C2476 a_7237_n509# a_7300_n2167# 0.00fF
C2477 a_4724_n3799# VDD 0.77fF
C2478 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C2479 a_8418_n5405# a_9706_n5405# 0.01fF
C2480 sky130_fd_sc_hd__clkinv_4_4/A a_6941_n5797# 0.07fF
C2481 a_8525_n5405# a_9450_n5405# 0.02fF
C2482 a_3176_n3255# a_3010_n4317# 0.00fF
C2483 a_8162_n2685# a_8229_n2997# 0.01fF
C2484 a_3077_n2997# a_3266_n4317# 0.00fF
C2485 a_4365_n821# a_4464_n1079# 0.49fF
C2486 a_7130_n13021# a_7040_n11415# 0.00fF
C2487 a_10904_n4887# a_11164_n4887# 0.23fF
C2488 a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C2489 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3266_n1597# 0.03fF
C2490 VDD a_4298_n9213# 0.76fF
C2491 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.34fF
C2492 a_4365_n5797# VDD 0.36fF
C2493 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__nand2_4_0/Y 0.69fF
C2494 a_8418_n2685# a_8328_n1079# 0.00fF
C2495 a_4464_n3255# a_5653_n2997# 0.01fF
C2496 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_1888_n5975# 0.05fF
C2497 a_6012_n12503# a_5842_n11933# 0.04fF
C2498 a_5752_n12503# a_5949_n11933# 0.02fF
C2499 a_5752_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.03fF
C2500 a_501_n11237# a_434_n13021# 0.00fF
C2501 a_9450_n10301# a_9706_n10301# 0.19fF
C2502 a_10805_n10613# VDD 0.32fF
C2503 a_8418_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C2504 a_4365_n9525# a_4464_n9783# 0.49fF
C2505 a_8588_n10871# a_8588_n12503# 0.01fF
C2506 a_8229_n10613# a_8418_n11933# 0.00fF
C2507 a_8328_n10871# a_8162_n11933# 0.00fF
C2508 a_9450_n4317# a_9616_n3255# 0.00fF
C2509 a_9876_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.29fF
C2510 a_1888_n4887# a_1789_n3621# 0.00fF
C2511 sky130_fd_sc_hd__clkinv_4_8/A a_9876_n12503# 0.10fF
C2512 a_1789_n4709# a_1888_n3799# 0.00fF
C2513 a_1722_n11933# VDD 0.76fF
C2514 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.00fF
C2515 a_11101_n9213# a_9706_n9213# 0.01fF
C2516 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8229_n13413# 0.01fF
C2517 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_9616_n4887# 0.01fF
C2518 a_8328_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.03fF
C2519 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_3010_n5405# 0.00fF
C2520 a_8162_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C2521 a_9450_n2685# a_9616_n3255# 0.04fF
C2522 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C2523 a_10805_n13413# a_9616_n13591# 0.01fF
C2524 a_4365_n1909# a_4464_n2167# 0.49fF
C2525 a_6874_n4317# a_7130_n4317# 0.19fF
C2526 a_1722_n4317# a_2085_n4317# 0.05fF
C2527 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkinv_1_0/A 0.08fF
C2528 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.02fF
C2529 a_3077_n3621# a_3176_n3799# 0.49fF
C2530 a_434_n11933# a_600_n13591# 0.00fF
C2531 a_690_n11933# a_501_n13413# 0.00fF
C2532 a_8418_n4317# a_8418_n5405# 0.01fF
C2533 a_860_n1079# VDD 0.80fF
C2534 sky130_fd_sc_hd__clkinv_4_4/A a_8328_n5975# 0.07fF
C2535 a_8162_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C2536 a_7237_n6493# a_7040_n4887# 0.00fF
C2537 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8229_n11237# 0.00fF
C2538 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_5752_n3255# 0.05fF
C2539 a_4724_n3255# a_6012_n3255# 0.01fF
C2540 a_4464_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C2541 VDD a_5842_n9213# 0.44fF
C2542 a_434_n2685# a_501_n2997# 0.01fF
C2543 VDD a_6874_n11933# 0.76fF
C2544 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.08fF
C2545 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.05fF
C2546 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_7300_n9783# 0.03fF
C2547 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.00fF
C2548 a_8229_n1909# a_8229_n2997# 0.02fF
C2549 a_7237_n6493# a_7300_n4887# 0.00fF
C2550 a_5653_n10613# a_6941_n10613# 0.01fF
C2551 a_9706_n10301# a_10994_n10301# 0.01fF
C2552 a_9813_n10301# a_10738_n10301# 0.02fF
C2553 a_9450_n10301# a_11101_n10301# 0.00fF
C2554 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VDD 0.84fF
C2555 a_501_n5797# a_690_n5405# 0.02fF
C2556 a_3266_n13021# a_3373_n11933# 0.00fF
C2557 a_600_n5975# a_434_n5405# 0.04fF
C2558 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C2559 a_3373_n13021# a_3266_n11933# 0.00fF
C2560 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_1722_n13021# 0.00fF
C2561 a_434_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.03fF
C2562 a_7237_n2685# VDD 0.35fF
C2563 a_6012_n2167# a_5842_n2685# 0.04fF
C2564 a_690_n13021# a_797_n13021# 0.55fF
C2565 a_5752_n2167# a_5949_n2685# 0.02fF
C2566 a_8328_n2167# a_8328_n1079# 0.01fF
C2567 a_10738_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C2568 a_2085_n2685# a_3266_n2685# 0.01fF
C2569 a_1978_n2685# a_3373_n2685# 0.01fF
C2570 a_2148_n12503# a_1978_n11933# 0.04fF
C2571 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3010_n2685# 0.35fF
C2572 a_1888_n12503# a_2085_n11933# 0.02fF
C2573 a_5653_n2997# a_5653_n1909# 0.02fF
C2574 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.01fF
C2575 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.16fF
C2576 a_3176_n2167# a_4365_n1909# 0.01fF
C2577 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.04fF
C2578 a_3266_n11933# VDD 0.47fF
C2579 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.00fF
C2580 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_4661_n11933# 0.01fF
C2581 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.03fF
C2582 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_9876_n4887# 0.03fF
C2583 a_6874_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C2584 a_13765_n2141# Bd 2.55fF
C2585 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C2586 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6941_n3621# 0.00fF
C2587 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_3436_n1079# 0.01fF
C2588 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.01fF
C2589 a_8525_n13021# a_8588_n13591# 0.01fF
C2590 a_9813_n8125# a_9876_n9783# 0.00fF
C2591 a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C2592 a_7237_n1597# a_8418_n1597# 0.01fF
C2593 a_7130_n1597# a_8525_n1597# 0.01fF
C2594 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8162_n1597# 0.35fF
C2595 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.08fF
C2596 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkinv_1_3/Y 0.02fF
C2597 Ad_b p2 1.13fF
C2598 a_7130_n4317# a_8418_n4317# 0.01fF
C2599 a_7237_n4317# a_8162_n4317# 0.02fF
C2600 a_4365_n1909# a_6012_n2167# 0.00fF
C2601 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3010_n4317# 0.35fF
C2602 a_1978_n4317# a_3373_n4317# 0.01fF
C2603 a_2085_n4317# a_3266_n4317# 0.01fF
C2604 a_6874_n4317# a_8525_n4317# 0.00fF
C2605 a_11164_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.03fF
C2606 a_13765_n9757# a_13765_n10301# 0.31fF
C2607 a_5752_n3799# a_5842_n4317# 0.02fF
C2608 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.04fF
C2609 a_7040_n11415# a_7237_n10301# 0.00fF
C2610 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9450_n5405# 0.01fF
C2611 a_3176_n3799# a_4464_n3799# 0.01fF
C2612 a_7300_n11415# a_7130_n10301# 0.00fF
C2613 a_9450_n509# VDD 0.80fF
C2614 a_3436_n3799# a_4365_n3621# 0.02fF
C2615 a_3077_n3621# a_4724_n3799# 0.00fF
C2616 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.04fF
C2617 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.02fF
C2618 a_4464_n3255# a_4661_n1597# 0.00fF
C2619 a_4724_n3255# a_4554_n1597# 0.00fF
C2620 a_2622_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.04fF
C2621 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_1_5/A 0.03fF
C2622 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.02fF
C2623 a_9876_n10871# a_9876_n11415# 0.09fF
C2624 a_4365_n13413# a_4298_n13021# 0.01fF
C2625 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C2626 a_4464_n3255# a_4661_n4317# 0.00fF
C2627 a_4724_n3255# a_4554_n4317# 0.00fF
C2628 a_8525_n13021# a_8588_n11415# 0.00fF
C2629 sky130_fd_sc_hd__clkinv_4_4/A a_6658_n7363# 0.02fF
C2630 a_5653_n5797# a_6941_n5797# 0.01fF
C2631 a_3077_n12325# a_3077_n13413# 0.02fF
C2632 a_434_n11933# a_690_n11933# 0.19fF
C2633 VDD a_8418_n11933# 0.47fF
C2634 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.09fF
C2635 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C2636 a_5752_n12503# a_5752_n13591# 0.01fF
C2637 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_860_n9783# 0.03fF
C2638 a_5752_n9783# a_5586_n10301# 0.04fF
C2639 a_4298_n1597# a_4464_n2167# 0.04fF
C2640 a_5653_n9525# a_5842_n10301# 0.02fF
C2641 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C2642 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_7237_n11933# 0.01fF
C2643 a_797_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C2644 a_7130_n1597# a_6941_n1909# 0.02fF
C2645 a_6941_n821# a_8229_n821# 0.01fF
C2646 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_3/A 2.16fF
C2647 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_1/A 2.16fF
C2648 a_7130_n6493# sky130_fd_sc_hd__clkinv_1_5/A 0.00fF
C2649 a_1888_n5975# a_1888_n4887# 0.01fF
C2650 a_9813_n5405# a_8418_n5405# 0.01fF
C2651 a_6941_n10613# a_7040_n10871# 0.49fF
C2652 a_10994_n10301# a_11101_n10301# 0.55fF
C2653 a_690_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C2654 a_797_n1597# VDD 0.36fF
C2655 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A VDD 0.89fF
C2656 a_11101_n2685# a_11164_n3255# 0.01fF
C2657 a_10738_n6173# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C2658 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_10805_n2997# 0.01fF
C2659 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_4554_n2685# 0.00fF
C2660 a_4298_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.03fF
C2661 a_10994_n4317# a_11164_n3255# 0.00fF
C2662 a_11101_n4317# a_10904_n3255# 0.00fF
C2663 a_4661_n11933# VDD 0.35fF
C2664 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4365_n4709# 0.01fF
C2665 a_5842_n4317# a_6012_n3799# 0.04fF
C2666 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.01fF
C2667 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_6012_n1079# 0.01fF
C2668 a_501_n821# a_2148_n1079# 0.00fF
C2669 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.95fF
C2670 a_2148_n10871# a_2085_n9213# 0.00fF
C2671 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkinv_4_8/A 0.02fF
C2672 a_7237_n5405# a_7300_n3799# 0.00fF
C2673 a_3266_n10301# a_3373_n11933# 0.00fF
C2674 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_7130_n1597# 0.00fF
C2675 a_3373_n10301# a_3266_n11933# 0.00fF
C2676 a_8418_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.05fF
C2677 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_9706_n1597# 0.00fF
C2678 a_8418_n4317# a_8525_n4317# 0.55fF
C2679 a_8162_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.03fF
C2680 a_10805_n5797# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C2681 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_4554_n4317# 0.00fF
C2682 a_3266_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.05fF
C2683 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.03fF
C2684 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C2685 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_5949_n9213# 0.01fF
C2686 a_690_n10301# a_501_n8437# 0.00fF
C2687 a_434_n10301# a_600_n8695# 0.00fF
C2688 a_2148_n8695# a_3436_n8695# 0.01fF
C2689 a_1888_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.00fF
C2690 a_3176_n1079# VDD 0.49fF
C2691 a_4464_n3799# a_4724_n3799# 0.28fF
C2692 a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.02fF
C2693 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_5653_n3621# 0.01fF
C2694 a_7237_n6493# a_7212_n7203# 0.01fF
C2695 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_7237_n6493# 0.01fF
C2696 a_10738_n11933# a_10904_n11415# 0.04fF
C2697 a_10994_n11933# a_10805_n11237# 0.02fF
C2698 a_600_n10871# a_434_n9213# 0.00fF
C2699 a_10994_n1597# VDD 0.42fF
C2700 a_434_n11933# a_1722_n11933# 0.01fF
C2701 a_6941_n5797# a_7040_n5975# 0.49fF
C2702 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.03fF
C2703 a_8328_n11415# a_8418_n10301# 0.01fF
C2704 a_8229_n821# a_8328_n1079# 0.49fF
C2705 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9706_n5405# 0.05fF
C2706 a_7040_n10871# a_8328_n10871# 0.01fF
C2707 a_7300_n9783# a_7300_n8695# 0.02fF
C2708 a_10994_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.00fF
C2709 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.02fF
C2710 a_1978_n2685# a_1978_n4317# 0.01fF
C2711 a_7300_n10871# a_8229_n10613# 0.02fF
C2712 a_7130_n2685# a_7130_n4317# 0.01fF
C2713 a_11164_n5975# a_11164_n4887# 0.02fF
C2714 a_13765_n10301# p2d_b 2.55fF
C2715 a_501_n5797# a_501_n4709# 0.02fF
C2716 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.04fF
C2717 a_860_n3255# a_860_n3799# 0.09fF
C2718 a_8229_n4709# a_8229_n3621# 0.02fF
C2719 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A VDD 0.89fF
C2720 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.03fF
C2721 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_3373_n11933# 0.01fF
C2722 a_5653_n821# VDD 0.35fF
C2723 a_4661_n5405# a_4724_n4887# 0.01fF
C2724 a_4464_n11415# a_4298_n13021# 0.00fF
C2725 a_4365_n11237# a_4554_n13021# 0.00fF
C2726 a_3077_n12325# a_3176_n11415# 0.00fF
C2727 a_3176_n12503# a_3077_n11237# 0.00fF
C2728 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4661_n1597# 0.02fF
C2729 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_7237_n1597# 0.02fF
C2730 a_3373_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C2731 sky130_fd_sc_hd__nand2_4_2/A a_2366_n14109# 0.03fF
C2732 a_600_n8695# VDD 0.49fF
C2733 a_5949_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C2734 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.15fF
C2735 a_8525_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C2736 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VDD 0.89fF
C2737 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9813_n1597# 0.02fF
C2738 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C2739 a_2366_n6493# sky130_fd_sc_hd__clkinv_4_4/A 0.01fF
C2740 a_501_n11237# a_434_n10301# 0.00fF
C2741 a_3373_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C2742 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4661_n4317# 0.02fF
C2743 a_8418_n509# a_9706_n509# 0.01fF
C2744 a_8162_n509# a_9813_n509# 0.00fF
C2745 a_9616_n2167# a_9616_n3799# 0.00fF
C2746 a_4724_n1079# VDD 0.83fF
C2747 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_5752_n3799# 0.05fF
C2748 a_5586_n5405# VDD 0.76fF
C2749 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.01fF
C2750 a_5949_n13021# a_5949_n11933# 0.02fF
C2751 sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# 0.58fF
C2752 a_501_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.00fF
C2753 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X a_4724_n4887# 0.01fF
C2754 a_5653_n2997# a_5752_n4887# 0.00fF
C2755 sky130_fd_sc_hd__clkinv_1_5/A a_7237_n9213# 0.00fF
C2756 a_5752_n10871# VDD 0.46fF
C2757 a_9813_n10301# VDD 0.34fF
C2758 a_4724_n9783# VDD 0.78fF
C2759 a_10805_n4709# a_10738_n5405# 0.01fF
C2760 a_7040_n5975# a_8328_n5975# 0.01fF
C2761 a_7300_n5975# a_8229_n5797# 0.02fF
C2762 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__dfxbp_1_0/Q 0.10fF
C2763 a_6941_n5797# a_8588_n5975# 0.00fF
C2764 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C2765 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_6012_n12503# 0.00fF
C2766 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.06fF
C2767 a_4464_n12503# a_4464_n13591# 0.01fF
C2768 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_8162_n14109# 0.00fF
C2769 a_6012_n5975# a_6101_n7254# 0.00fF
C2770 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6006_n7607# 0.00fF
C2771 a_4298_n9213# a_5586_n9213# 0.01fF
C2772 a_7130_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.23fF
C2773 a_7300_n9783# a_7130_n10301# 0.04fF
C2774 a_5949_n1597# a_5752_n2167# 0.02fF
C2775 a_5842_n1597# a_6012_n2167# 0.04fF
C2776 a_7040_n9783# a_7237_n10301# 0.02fF
C2777 a_n2602_n7037# a_n1738_n6671# 0.10fF
C2778 a_n1738_n6671# a_n1654_n6671# 0.02fF
C2779 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n4317# 0.00fF
C2780 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C2781 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3010_n4317# 0.00fF
C2782 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C2783 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X a_7300_n3255# 0.01fF
C2784 A Ad 0.20fF
C2785 a_5752_n5975# VDD 0.44fF
C2786 a_10904_n2167# a_10994_n2685# 0.01fF
C2787 a_7040_n1079# VDD 0.46fF
C2788 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7300_n3799# 0.03fF
C2789 a_7237_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C2790 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1978_n13021# 0.03fF
C2791 a_797_n13021# a_2085_n13021# 0.01fF
C2792 a_600_n12503# a_600_n11415# 0.01fF
C2793 a_9706_n8125# a_9706_n9213# 0.01fF
C2794 a_501_n11237# VDD 0.36fF
C2795 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C2796 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_6012_n3799# 0.03fF
C2797 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.02fF
C2798 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_3436_n3255# 0.03fF
C2799 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C2800 a_7130_n14109# a_8162_n14109# 0.02fF
C2801 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C2802 a_6874_n14109# a_8418_n14109# 0.01fF
C2803 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.02fF
C2804 sky130_fd_sc_hd__nand2_4_2/A a_7130_n14109# 0.03fF
C2805 a_2148_n3799# a_600_n3799# 0.01fF
C2806 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n11933# 0.35fF
C2807 a_9813_n11933# a_10994_n11933# 0.01fF
C2808 a_10738_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.03fF
C2809 a_1888_n2167# a_1888_n3799# 0.00fF
C2810 a_4554_n4317# a_4464_n4887# 0.01fF
C2811 a_690_n13021# a_860_n13591# 0.04fF
C2812 a_9450_n509# sky130_fd_sc_hd__nand2_4_0/B 0.03fF
C2813 a_690_n2685# a_1722_n2685# 0.02fF
C2814 a_434_n2685# a_1978_n2685# 0.01fF
C2815 a_10994_n13021# VDD 0.43fF
C2816 a_6012_n3255# a_6012_n4887# 0.01fF
C2817 sky130_fd_sc_hd__nand2_4_3/Y a_8588_n9783# 0.11fF
C2818 a_600_n1079# a_860_n1079# 0.28fF
C2819 a_1789_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C2820 a_1722_n11933# a_3010_n11933# 0.01fF
C2821 a_860_n5975# a_797_n4317# 0.00fF
C2822 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_797_n9213# 0.01fF
C2823 a_2148_n10871# a_1978_n9213# 0.00fF
C2824 a_5752_n11415# a_5653_n12325# 0.00fF
C2825 a_5653_n11237# a_5752_n12503# 0.00fF
C2826 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C2827 a_13765_n10301# VDD 2.20fF
C2828 a_7300_n10871# VDD 0.78fF
C2829 a_3176_n10871# a_4365_n10613# 0.01fF
C2830 a_8229_n9525# a_9616_n9783# 0.01fF
C2831 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_9706_n4317# 0.00fF
C2832 a_8328_n5975# a_8588_n5975# 0.28fF
C2833 a_1888_n9783# a_2085_n9213# 0.02fF
C2834 a_8588_n12503# a_8525_n14109# 0.00fF
C2835 a_5586_n9213# a_5842_n9213# 0.19fF
C2836 a_7040_n5975# a_6658_n7363# 0.00fF
C2837 a_9517_n8437# a_11164_n8695# 0.00fF
C2838 a_9616_n8695# a_10904_n8695# 0.01fF
C2839 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.00fF
C2840 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_860_n4887# 0.00fF
C2841 a_9876_n8695# a_10805_n8437# 0.02fF
C2842 a_1888_n11415# a_1888_n10871# 0.07fF
C2843 a_8525_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.05fF
C2844 a_600_n4887# a_n787_n4709# 0.01fF
C2845 a_5586_n4317# a_5653_n5797# 0.00fF
C2846 a_1888_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.03fF
C2847 a_4554_n10301# a_4464_n8695# 0.00fF
C2848 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.02fF
C2849 a_8229_n2997# VDD 0.35fF
C2850 a_501_n10613# a_1888_n10871# 0.01fF
C2851 a_8525_n2685# a_8525_n4317# 0.01fF
C2852 a_7040_n8695# a_6874_n10301# 0.00fF
C2853 a_8588_n10871# a_8418_n10301# 0.04fF
C2854 a_7040_n8695# a_8588_n8695# 0.01fF
C2855 clk a_n1139_n6715# 0.00fF
C2856 a_7300_n8695# a_8328_n8695# 0.02fF
C2857 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_8229_n8437# 0.18fF
C2858 a_6874_n5405# a_7040_n5975# 0.04fF
C2859 a_7130_n5405# a_6941_n5797# 0.02fF
C2860 a_7300_n5975# VDD 0.78fF
C2861 a_2366_n14109# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C2862 a_4365_n5797# sky130_fd_sc_hd__clkinv_4_4/A 0.07fF
C2863 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C2864 a_9616_n4887# a_9616_n3799# 0.01fF
C2865 a_8588_n1079# VDD 0.77fF
C2866 a_9517_n10613# a_9450_n11933# 0.00fF
C2867 a_7130_n8125# a_7212_n7203# 0.01fF
C2868 a_434_n9213# a_501_n9525# 0.01fF
C2869 a_2085_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.12fF
C2870 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11164_n3255# 0.02fF
C2871 a_8162_n13021# a_9706_n13021# 0.01fF
C2872 a_8418_n13021# a_9450_n13021# 0.02fF
C2873 a_9813_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.12fF
C2874 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_1/A 0.82fF
C2875 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.03fF
C2876 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A VDD 0.87fF
C2877 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_797_n13021# 0.01fF
C2878 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_7237_n8125# 0.00fF
C2879 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C2880 sky130_fd_sc_hd__nand2_4_1/B a_9876_n4887# 0.00fF
C2881 a_9813_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C2882 a_10994_n11933# sky130_fd_sc_hd__clkinv_4_8/A 0.01fF
C2883 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_1888_n3799# 0.03fF
C2884 a_n787_n9525# a_501_n9525# 0.01fF
C2885 a_11101_n1597# a_11164_n1079# 0.01fF
C2886 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkinv_1_5/A 0.02fF
C2887 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5653_n4709# 0.01fF
C2888 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C2889 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.02fF
C2890 a_5586_n13021# a_7130_n13021# 0.01fF
C2891 a_4365_n3621# a_4298_n5405# 0.00fF
C2892 a_7130_n2685# a_7237_n2685# 0.55fF
C2893 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C2894 a_1722_n2685# a_2085_n2685# 0.05fF
C2895 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n9213# 0.01fF
C2896 a_6874_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C2897 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_7237_n9213# 0.01fF
C2898 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.03fF
C2899 a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C2900 a_9813_n8125# VDD 0.36fF
C2901 a_5949_n13021# a_5752_n13591# 0.02fF
C2902 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C2903 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.69fF
C2904 a_3010_n11933# a_3266_n11933# 0.19fF
C2905 sky130_fd_sc_hd__nand2_4_0/B a_10994_n1597# 0.00fF
C2906 a_10904_n4887# a_10738_n4317# 0.04fF
C2907 a_10805_n4709# a_10994_n4317# 0.02fF
C2908 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.04fF
C2909 a_10904_n3255# VDD 0.41fF
C2910 sky130_fd_sc_hd__nand2_4_3/Y a_10738_n8125# 0.49fF
C2911 a_434_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.03fF
C2912 a_690_n10301# a_797_n10301# 0.55fF
C2913 a_8525_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C2914 a_797_n2685# a_860_n3799# 0.00fF
C2915 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9813_n4317# 0.02fF
C2916 a_690_n13021# a_797_n11933# 0.00fF
C2917 a_9450_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.07fF
C2918 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.04fF
C2919 a_9517_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C2920 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_8229_n821# 0.02fF
C2921 a_690_n4317# VDD 0.48fF
C2922 a_860_n2167# a_860_n3255# 0.02fF
C2923 B a_13765_n1597# 0.12fF
C2924 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5653_n8437# 0.00fF
C2925 a_6874_n11933# a_8162_n11933# 0.01fF
C2926 a_5653_n3621# a_5586_n2685# 0.00fF
C2927 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.00fF
C2928 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_3436_n13591# 0.03fF
C2929 a_5586_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C2930 a_9517_n10613# a_9450_n10301# 0.01fF
C2931 a_8328_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.03fF
C2932 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_9616_n8695# 0.01fF
C2933 a_690_n1597# a_860_n1079# 0.04fF
C2934 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.02fF
C2935 a_797_n1597# a_600_n1079# 0.02fF
C2936 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C2937 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C2938 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C2939 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_9813_n13021# 0.00fF
C2940 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C2941 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.02fF
C2942 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C2943 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X 0.01fF
C2944 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_2148_n3255# 0.01fF
C2945 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A 0.02fF
C2946 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkinv_4_4/A 0.04fF
C2947 a_5586_n11933# a_5842_n11933# 0.19fF
C2948 a_600_n2167# a_1789_n1909# 0.01fF
C2949 a_501_n1909# a_1888_n2167# 0.01fF
C2950 a_8328_n9783# a_8162_n9213# 0.04fF
C2951 a_7300_n8695# a_7130_n8125# 0.04fF
C2952 a_7040_n8695# a_7237_n8125# 0.02fF
C2953 a_1789_n821# a_2148_n1079# 0.05fF
C2954 a_13765_n12477# VDD 1.90fF
C2955 a_7237_n2685# a_8525_n2685# 0.01fF
C2956 a_7237_n10301# a_7237_n9213# 0.02fF
C2957 a_7130_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C2958 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8418_n2685# 0.03fF
C2959 a_9616_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.05fF
C2960 a_9876_n12503# a_8588_n12503# 0.01fF
C2961 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_8328_n12503# 0.00fF
C2962 a_797_n13021# a_600_n13591# 0.02fF
C2963 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A VDD 0.89fF
C2964 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2965 a_3373_n11933# a_4298_n11933# 0.02fF
C2966 a_3010_n11933# a_4661_n11933# 0.00fF
C2967 a_3266_n11933# a_4554_n11933# 0.01fF
C2968 a_9616_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C2969 a_13765_n5949# a_13765_n4317# 0.01fF
C2970 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C2971 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD 0.83fF
C2972 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1978_n10301# 0.03fF
C2973 a_7130_n14109# a_6941_n13413# 0.02fF
C2974 a_797_n10301# a_2085_n10301# 0.01fF
C2975 a_3373_n5405# a_3176_n4887# 0.02fF
C2976 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkinv_4_3/A 0.06fF
C2977 a_690_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C2978 a_6874_n14109# a_7040_n13591# 0.04fF
C2979 a_4365_n9525# a_4554_n9213# 0.02fF
C2980 a_3436_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.03fF
C2981 a_4464_n9783# a_4298_n9213# 0.04fF
C2982 a_9517_n8437# a_9517_n9525# 0.02fF
C2983 a_501_n11237# a_434_n11933# 0.01fF
C2984 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A a_3373_n9213# 0.01fF
C2985 a_9876_n1079# a_8588_n1079# 0.01fF
C2986 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C2987 a_3436_n11415# a_3436_n10871# 0.09fF
C2988 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X a_8328_n1079# 0.00fF
C2989 a_6006_n7607# p2 0.00fF
C2990 a_6101_n7254# a_6794_n7203# 0.06fF
C2991 a_7130_n4317# a_7040_n5975# 0.00fF
C2992 a_7130_n10301# a_8162_n10301# 0.02fF
C2993 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VDD 0.66fF
C2994 a_6658_n7363# a_6665_n7459# 1.73fF
C2995 a_6373_n7349# a_6865_n7304# 0.04fF
C2996 a_9517_n5797# a_9450_n4317# 0.00fF
C2997 a_8162_n11933# a_8418_n11933# 0.19fF
C2998 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/B 0.02fF
C2999 a_5949_n10301# a_6012_n8695# 0.00fF
C3000 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_100/A 0.02fF
C3001 a_4724_n11415# a_4554_n10301# 0.00fF
C3002 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.02fF
C3003 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.02fF
C3004 a_7237_n509# sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C3005 a_4464_n11415# a_4661_n10301# 0.00fF
C3006 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_2148_n11415# 0.03fF
C3007 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C3008 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_9876_n8695# 0.03fF
C3009 a_10994_n5405# a_10805_n5797# 0.02fF
C3010 a_10738_n5405# a_10904_n5975# 0.04fF
C3011 a_8525_n5405# a_8328_n5975# 0.02fF
C3012 a_9876_n10871# a_9813_n9213# 0.00fF
C3013 a_11164_n13591# VDD 0.66fF
C3014 a_8418_n5405# a_8588_n5975# 0.04fF
C3015 sky130_fd_sc_hd__nand2_4_3/Y a_10994_n10301# 0.01fF
C3016 a_9706_n6493# a_9706_n8125# 0.00fF
C3017 a_6865_n7304# VDD 0.47fF
C3018 a_4365_n5797# a_5653_n5797# 0.01fF
C3019 a_1978_n9213# a_1888_n9783# 0.02fF
C3020 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.04fF
C3021 a_9450_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C3022 a_9517_n13413# VDD 0.34fF
C3023 a_8229_n1909# a_8418_n509# 0.00fF
C3024 a_8328_n2167# a_8162_n509# 0.00fF
C3025 a_2148_n5975# a_600_n5975# 0.01fF
C3026 a_1888_n5975# a_860_n5975# 0.02fF
C3027 a_3176_n8695# a_3176_n9783# 0.01fF
C3028 a_5586_n11933# a_7237_n11933# 0.00fF
C3029 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C3030 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_4661_n10301# 0.01fF
C3031 a_1888_n11415# a_1789_n9525# 0.00fF
C3032 a_1789_n11237# a_1888_n9783# 0.00fF
C3033 a_6874_n5405# a_7130_n5405# 0.19fF
C3034 a_7237_n5405# VDD 0.35fF
C3035 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C3036 a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C3037 a_2148_n4887# a_1978_n5405# 0.04fF
C3038 a_3436_n3255# a_3266_n2685# 0.04fF
C3039 a_434_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.03fF
C3040 a_5653_n4709# a_7040_n4887# 0.01fF
C3041 a_5752_n4887# a_6941_n4709# 0.01fF
C3042 a_3176_n3255# a_3373_n2685# 0.02fF
C3043 a_690_n1597# a_797_n1597# 0.55fF
C3044 a_5752_n3799# a_5842_n5405# 0.00fF
C3045 a_n1139_n6715# sky130_fd_sc_hd__clkinv_1_5/A 0.31fF
C3046 a_8525_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.12fF
C3047 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkinv_1_0/A 0.02fF
C3048 a_7130_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.05fF
C3049 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.01fF
C3050 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_5586_n11933# 0.00fF
C3051 a_4298_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.03fF
C3052 a_4554_n11933# a_4661_n11933# 0.55fF
C3053 a_9517_n11237# VDD 0.34fF
C3054 a_7300_n4887# a_5653_n4709# 0.00fF
C3055 a_n688_n12503# sky130_fd_sc_hd__nand2_1_4/B 0.14fF
C3056 a_5653_n10613# a_5842_n9213# 0.00fF
C3057 a_5752_n10871# a_5586_n9213# 0.00fF
C3058 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.01fF
C3059 a_2085_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.12fF
C3060 a_8418_n4317# a_8229_n2997# 0.00fF
C3061 a_8162_n4317# a_8328_n3255# 0.00fF
C3062 a_8418_n10301# a_8525_n9213# 0.00fF
C3063 a_690_n11933# a_797_n13021# 0.00fF
C3064 sky130_fd_sc_hd__clkinv_4_3/Y p2 0.03fF
C3065 a_n688_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3066 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.04fF
C3067 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8229_n5797# 0.00fF
C3068 a_8162_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C3069 a_1978_n1597# a_1888_n1079# 0.01fF
C3070 a_8418_n11933# a_9706_n11933# 0.01fF
C3071 a_8525_n11933# a_9450_n11933# 0.02fF
C3072 a_9616_n10871# a_8229_n10613# 0.01fF
C3073 a_9517_n10613# a_8328_n10871# 0.01fF
C3074 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/A 0.46fF
C3075 a_3436_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C3076 a_10904_n10871# a_10994_n10301# 0.02fF
C3077 a_8328_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C3078 a_3077_n4709# a_3266_n4317# 0.02fF
C3079 a_3176_n4887# a_3010_n4317# 0.04fF
C3080 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.02fF
C3081 a_4464_n10871# a_4298_n11933# 0.00fF
C3082 a_2729_n8125# VDD 0.36fF
C3083 a_8588_n9783# a_8525_n10301# 0.01fF
C3084 p2d a_13765_n10301# 0.12fF
C3085 a_n2163_n6671# a_n1738_n6671# 0.04fF
C3086 a_n2436_n7037# a_n2248_n7037# 0.22fF
C3087 a_n1995_n6925# a_n1139_n6715# 0.02fF
C3088 a_5842_n5405# a_6012_n3799# 0.00fF
C3089 a_13765_n8669# a_13765_n9213# 0.31fF
C3090 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X a_8588_n13591# 0.01fF
C3091 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C3092 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.00fF
C3093 a_5949_n4317# VDD 0.35fF
C3094 a_5653_n13413# a_5586_n11933# 0.00fF
C3095 a_11164_n2167# a_10738_n509# 0.01fF
C3096 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C3097 a_9517_n1909# a_9517_n821# 0.02fF
C3098 a_9876_n9783# a_9706_n9213# 0.04fF
C3099 a_6874_n5405# a_8525_n5405# 0.00fF
C3100 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C3101 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_8525_n8125# 0.01fF
C3102 a_7130_n5405# a_8418_n5405# 0.01fF
C3103 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A VDD 0.87fF
C3104 a_7237_n5405# a_8162_n5405# 0.02fF
C3105 a_6874_n2685# a_6941_n2997# 0.01fF
C3106 a_3077_n821# a_3176_n1079# 0.49fF
C3107 a_5842_n13021# a_5752_n11415# 0.00fF
C3108 a_501_n4709# a_1888_n4887# 0.01fF
C3109 Bd_b a_4724_n8695# 0.01fF
C3110 a_600_n4887# a_1789_n4709# 0.01fF
C3111 a_797_n1597# a_2085_n1597# 0.01fF
C3112 a_690_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.01fF
C3113 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.04fF
C3114 a_1789_n5797# VDD 0.37fF
C3115 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1978_n1597# 0.03fF
C3116 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.02fF
C3117 Ad_b a_4986_n7215# 0.02fF
C3118 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C3119 a_3176_n3255# a_4365_n2997# 0.01fF
C3120 a_3077_n2997# a_4464_n3255# 0.01fF
C3121 a_7130_n2685# a_7040_n1079# 0.00fF
C3122 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.08fF
C3123 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_860_n13591# 0.01fF
C3124 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C3125 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_690_n13021# 0.02fF
C3126 a_10738_n1597# a_10994_n1597# 0.19fF
C3127 a_860_n2167# a_797_n2685# 0.01fF
C3128 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VDD 0.83fF
C3129 a_7130_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.05fF
C3130 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C3131 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_8588_n12503# 0.01fF
C3132 a_7300_n4887# a_7040_n4887# 0.28fF
C3133 a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C3134 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_6941_n4709# 0.02fF
C3135 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.03fF
C3136 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.02fF
C3137 sky130_fd_sc_hd__nand2_4_1/A a_n787_n4709# 0.00fF
C3138 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_8525_n2685# 0.01fF
C3139 a_501_n2997# a_860_n3255# 0.05fF
C3140 a_7040_n10871# a_6874_n11933# 0.00fF
C3141 a_6941_n10613# a_7130_n11933# 0.00fF
C3142 a_2366_n8125# a_2622_n8125# 0.19fF
C3143 a_9450_n10301# a_9450_n9213# 0.02fF
C3144 a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3145 a_9813_n9213# a_8418_n9213# 0.01fF
C3146 a_600_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.04fF
C3147 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3077_n821# 0.01fF
C3148 a_8525_n4317# a_8588_n5975# 0.00fF
C3149 a_3010_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.03fF
C3150 a_10904_n5975# a_10994_n4317# 0.00fF
C3151 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.03fF
C3152 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6941_n13413# 0.01fF
C3153 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkinv_1_3/A 0.84fF
C3154 a_8162_n509# a_8229_n821# 0.01fF
C3155 a_9876_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C3156 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_501_n3621# 0.00fF
C3157 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_3436_n4887# 0.01fF
C3158 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C3159 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_1888_n4887# 0.01fF
C3160 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.03fF
C3161 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_11164_n11415# 0.01fF
C3162 a_5586_n4317# a_5842_n4317# 0.19fF
C3163 a_9450_n8125# a_9616_n9783# 0.00fF
C3164 a_690_n11933# a_797_n10301# 0.00fF
C3165 a_797_n11933# a_690_n10301# 0.00fF
C3166 a_3436_n3255# a_1789_n2997# 0.00fF
C3167 a_501_n1909# a_501_n821# 0.02fF
C3168 a_8328_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C3169 a_8588_n11415# a_9876_n11415# 0.01fF
C3170 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_9616_n11415# 0.05fF
C3171 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VDD 0.88fF
C3172 a_7130_n4317# a_7130_n5405# 0.01fF
C3173 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_860_n9783# 0.01fF
C3174 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VDD 0.84fF
C3175 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C3176 sky130_fd_sc_hd__clkinv_4_4/A a_5752_n5975# 0.07fF
C3177 a_8162_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.03fF
C3178 a_8418_n5405# a_8525_n5405# 0.55fF
C3179 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_9450_n5405# 0.00fF
C3180 a_3077_n821# a_4724_n1079# 0.00fF
C3181 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkinv_1_3/Y 0.04fF
C3182 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6941_n11237# 0.00fF
C3183 a_3436_n1079# a_4365_n821# 0.02fF
C3184 a_3176_n1079# a_4464_n1079# 0.01fF
C3185 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_3010_n2685# 0.01fF
C3186 sky130_fd_sc_hd__nand2_4_1/A a_11164_n4887# 0.01fF
C3187 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.00fF
C3188 a_9876_n4887# a_11164_n4887# 0.01fF
C3189 a_9616_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.00fF
C3190 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.02fF
C3191 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkinv_1_5/A 0.09fF
C3192 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_4661_n2685# 0.01fF
C3193 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C3194 a_2085_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.12fF
C3195 sky130_fd_sc_hd__nand2_4_0/A a_2622_n509# 0.08fF
C3196 VDD a_3266_n9213# 0.45fF
C3197 a_3176_n2167# a_3266_n2685# 0.01fF
C3198 a_3176_n5975# VDD 0.47fF
C3199 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkinv_1_0/A 0.03fF
C3200 a_9517_n1909# a_9706_n509# 0.00fF
C3201 a_4365_n2997# a_4724_n3255# 0.05fF
C3202 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.00fF
C3203 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8229_n821# 0.00fF
C3204 sky130_fd_sc_hd__nand2_4_3/Y a_6658_n7363# 0.01fF
C3205 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.04fF
C3206 a_8525_n10301# a_9450_n10301# 0.02fF
C3207 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.02fF
C3208 a_7237_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C3209 a_4365_n9525# a_4464_n10871# 0.00fF
C3210 a_9616_n10871# VDD 0.45fF
C3211 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8525_n8125# 0.02fF
C3212 a_2085_n13021# a_1978_n11933# 0.00fF
C3213 a_1978_n13021# a_2085_n11933# 0.00fF
C3214 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_7040_n4887# 0.00fF
C3215 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X a_1789_n2997# 0.18fF
C3216 a_4464_n2167# a_4661_n2685# 0.02fF
C3217 a_4724_n2167# a_4554_n2685# 0.04fF
C3218 a_8229_n10613# a_8162_n9213# 0.00fF
C3219 a_11101_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.00fF
C3220 a_9813_n10301# a_9706_n11933# 0.00fF
C3221 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_1/Y 0.19fF
C3222 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.04fF
C3223 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.02fF
C3224 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.06fF
C3225 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9706_n9213# 0.05fF
C3226 a_10994_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.00fF
C3227 a_13765_n5949# Bd_b 0.10fF
C3228 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.03fF
C3229 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_797_n11933# 0.01fF
C3230 a_2148_n3799# a_2085_n5405# 0.00fF
C3231 a_501_n8437# a_600_n8695# 0.49fF
C3232 a_4464_n1079# a_5653_n821# 0.01fF
C3233 a_4365_n821# a_5752_n1079# 0.01fF
C3234 a_501_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.02fF
C3235 a_600_n13591# a_860_n13591# 0.28fF
C3236 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A VDD 0.88fF
C3237 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X a_1722_n4317# 0.01fF
C3238 a_7237_n13021# a_7300_n13591# 0.01fF
C3239 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_2148_n1079# 0.01fF
C3240 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.01fF
C3241 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.00fF
C3242 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_8588_n4887# 0.03fF
C3243 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.29fF
C3244 a_5949_n4317# a_6874_n4317# 0.02fF
C3245 a_5842_n4317# a_7130_n4317# 0.01fF
C3246 a_5586_n4317# a_7237_n4317# 0.00fF
C3247 a_1789_n1909# a_1789_n2997# 0.02fF
C3248 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.06fF
C3249 sky130_fd_sc_hd__nand2_1_4/B a_4623_n7349# 0.01fF
C3250 a_6874_n2685# a_6874_n1597# 0.02fF
C3251 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.04fF
C3252 a_9450_n2685# a_9450_n1597# 0.02fF
C3253 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8162_n5405# 0.01fF
C3254 a_8162_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C3255 a_860_n11415# a_860_n9783# 0.01fF
C3256 a_6012_n11415# a_5842_n10301# 0.00fF
C3257 a_5752_n11415# a_5949_n10301# 0.00fF
C3258 a_6874_n509# VDD 0.78fF
C3259 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.02fF
C3260 a_5752_n3799# a_5949_n5405# 0.00fF
C3261 a_3176_n3255# a_3373_n1597# 0.00fF
C3262 a_8418_n2685# a_8328_n3255# 0.02fF
C3263 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C3264 a_10904_n2167# a_10904_n1079# 0.01fF
C3265 a_3077_n13413# a_3010_n13021# 0.01fF
C3266 a_3436_n3255# a_3266_n4317# 0.00fF
C3267 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9706_n5405# 0.03fF
C3268 a_3176_n3255# a_3373_n4317# 0.00fF
C3269 a_4464_n1079# a_4724_n1079# 0.28fF
C3270 a_4365_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.02fF
C3271 sky130_fd_sc_hd__clkinv_4_4/A a_7300_n5975# 0.11fF
C3272 a_7237_n13021# a_7300_n11415# 0.00fF
C3273 a_1789_n12325# a_1789_n13413# 0.02fF
C3274 VDD a_4661_n9213# 0.35fF
C3275 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_4298_n2685# 0.03fF
C3276 a_4724_n5975# VDD 0.83fF
C3277 a_2148_n2167# a_2366_n509# 0.00fF
C3278 VDD a_5842_n11933# 0.47fF
C3279 a_13765_n4317# a_13765_n4861# 0.31fF
C3280 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_4_3/A 0.80fF
C3281 a_5653_n821# a_6941_n821# 0.01fF
C3282 a_8525_n2685# a_8588_n1079# 0.00fF
C3283 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_5653_n2997# 0.18fF
C3284 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.03fF
C3285 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_5949_n11933# 0.01fF
C3286 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C3287 a_4623_n7349# Ad_b 0.16fF
C3288 a_3373_n10301# a_3266_n9213# 0.00fF
C3289 a_3266_n10301# a_3373_n9213# 0.00fF
C3290 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_10738_n10301# 0.00fF
C3291 a_5653_n10613# a_5752_n10871# 0.49fF
C3292 a_9706_n10301# a_9813_n10301# 0.55fF
C3293 a_9450_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C3294 a_600_n11415# a_690_n13021# 0.00fF
C3295 a_11164_n10871# VDD 0.67fF
C3296 a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.02fF
C3297 a_4464_n9783# a_4724_n9783# 0.28fF
C3298 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C3299 a_8328_n10871# a_8525_n11933# 0.00fF
C3300 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_3266_n2685# 0.00fF
C3301 a_9450_n6493# VDD 0.77fF
C3302 a_9813_n4317# a_9616_n3255# 0.00fF
C3303 a_9706_n4317# a_9876_n3255# 0.00fF
C3304 a_2085_n11933# VDD 0.35fF
C3305 a_5586_n5405# a_5653_n5797# 0.01fF
C3306 a_5949_n5405# a_6012_n3799# 0.00fF
C3307 a_434_n13021# sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C3308 a_1722_n10301# a_1722_n9213# 0.02fF
C3309 a_1978_n10301# a_2085_n11933# 0.00fF
C3310 a_9813_n2685# a_9616_n3255# 0.02fF
C3311 a_2085_n10301# a_1978_n11933# 0.00fF
C3312 a_9706_n2685# a_9876_n3255# 0.04fF
C3313 a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.17fF
C3314 a_7130_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.05fF
C3315 a_7130_n4317# a_7237_n4317# 0.55fF
C3316 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_8162_n4317# 0.00fF
C3317 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.03fF
C3318 a_4365_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C3319 a_1978_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.05fF
C3320 a_9450_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C3321 a_3010_n10301# a_3077_n8437# 0.00fF
C3322 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_5586_n4317# 0.03fF
C3323 a_8162_n13021# a_8328_n12503# 0.04fF
C3324 a_8418_n13021# a_8229_n12325# 0.02fF
C3325 a_8525_n4317# a_8525_n5405# 0.02fF
C3326 a_4298_n1597# a_3010_n1597# 0.01fF
C3327 a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.02fF
C3328 a_3176_n3799# a_3436_n3799# 0.28fF
C3329 a_690_n11933# a_860_n13591# 0.00fF
C3330 a_8418_n509# VDD 0.47fF
C3331 a_797_n11933# a_600_n13591# 0.00fF
C3332 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.09fF
C3333 a_13765_n2141# a_13765_n1053# 0.07fF
C3334 a_9450_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C3335 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9517_n2997# 0.01fF
C3336 a_5653_n5797# a_5752_n5975# 0.49fF
C3337 a_5586_n13021# a_5752_n12503# 0.04fF
C3338 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.02fF
C3339 a_690_n2685# a_600_n3255# 0.02fF
C3340 VDD a_7237_n11933# 0.35fF
C3341 a_8162_n9213# VDD 0.76fF
C3342 a_8588_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C3343 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X a_8588_n3255# 0.01fF
C3344 a_6941_n821# a_7040_n1079# 0.49fF
C3345 a_8328_n2167# a_8328_n3255# 0.01fF
C3346 a_10738_n1597# a_10904_n3255# 0.00fF
C3347 a_10994_n1597# a_10805_n2997# 0.00fF
C3348 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.02fF
C3349 a_9813_n10301# a_11101_n10301# 0.01fF
C3350 a_8328_n10871# a_8525_n10301# 0.02fF
C3351 a_5653_n10613# a_7300_n10871# 0.00fF
C3352 a_6012_n10871# a_6941_n10613# 0.02fF
C3353 a_5752_n10871# a_7040_n10871# 0.01fF
C3354 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_10994_n10301# 0.03fF
C3355 Bd_b sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C3356 a_860_n5975# a_690_n5405# 0.04fF
C3357 a_600_n5975# a_797_n5405# 0.02fF
C3358 a_2148_n3255# a_2148_n4887# 0.01fF
C3359 a_6012_n8695# a_6006_n7607# 0.01fF
C3360 sky130_fd_sc_hd__clkinv_4_8/A a_8229_n12325# 0.07fF
C3361 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.03fF
C3362 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_5949_n2685# 0.01fF
C3363 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_9616_n3255# 0.00fF
C3364 a_8588_n2167# a_8588_n1079# 0.02fF
C3365 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3373_n2685# 0.02fF
C3366 a_2085_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C3367 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C3368 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_2085_n11933# 0.01fF
C3369 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_4365_n1909# 0.18fF
C3370 a_3373_n5405# a_3436_n4887# 0.01fF
C3371 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A VDD 0.88fF
C3372 a_3176_n11415# a_3010_n13021# 0.00fF
C3373 a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.18fF
C3374 a_3077_n11237# a_3266_n13021# 0.00fF
C3375 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.06fF
C3376 a_5653_n8437# VDD 0.36fF
C3377 a_1789_n12325# a_1888_n11415# 0.00fF
C3378 a_1888_n12503# a_1789_n11237# 0.00fF
C3379 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.02fF
C3380 a_13765_n12477# p1_b 0.15fF
C3381 p1d a_13765_n13021# 0.15fF
C3382 a_7237_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C3383 a_8328_n11415# a_8328_n9783# 0.00fF
C3384 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8525_n1597# 0.02fF
C3385 a_7130_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C3386 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8418_n4317# 0.03fF
C3387 a_7237_n4317# a_8525_n4317# 0.01fF
C3388 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3373_n4317# 0.02fF
C3389 a_2085_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C3390 a_9616_n5975# sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C3391 sky130_fd_sc_hd__nand2_4_3/B a_10738_n8125# 0.38fF
C3392 a_2148_n1079# VDD 0.79fF
C3393 a_5586_n13021# a_4298_n13021# 0.01fF
C3394 a_3436_n3799# a_4724_n3799# 0.01fF
C3395 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C3396 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_7237_n10301# 0.00fF
C3397 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_4464_n3799# 0.05fF
C3398 a_3010_n5405# VDD 0.76fF
C3399 a_3176_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C3400 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_3010_n4317# 0.03fF
C3401 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkinv_4_3/A 0.09fF
C3402 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_4661_n1597# 0.00fF
C3403 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C3404 a_10738_n13021# a_10994_n13021# 0.19fF
C3405 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X a_860_n4887# 0.00fF
C3406 a_4464_n3255# a_4365_n4709# 0.00fF
C3407 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C3408 a_4365_n2997# a_4464_n4887# 0.00fF
C3409 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.09fF
C3410 a_4464_n13591# a_4554_n13021# 0.01fF
C3411 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C3412 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_4661_n4317# 0.00fF
C3413 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.02fF
C3414 a_6012_n5975# a_6941_n5797# 0.02fF
C3415 a_10805_n5797# VDD 0.32fF
C3416 a_5752_n5975# a_7040_n5975# 0.01fF
C3417 a_5653_n5797# a_7300_n5975# 0.00fF
C3418 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C3419 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_4724_n12503# 0.00fF
C3420 a_3176_n12503# a_3176_n13591# 0.01fF
C3421 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1789_n2997# 0.01fF
C3422 a_1722_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C3423 a_5653_n13413# VDD 0.35fF
C3424 a_434_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.03fF
C3425 a_690_n11933# a_797_n11933# 0.55fF
C3426 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.88fF
C3427 a_3010_n9213# a_4298_n9213# 0.01fF
C3428 a_9706_n9213# VDD 0.43fF
C3429 sky130_fd_sc_hd__nand2_4_1/B a_10738_n6173# 0.39fF
C3430 a_6941_n821# a_8588_n1079# 0.00fF
C3431 a_7300_n1079# a_8229_n821# 0.02fF
C3432 a_7040_n1079# a_8328_n1079# 0.01fF
C3433 a_6012_n9783# a_5842_n10301# 0.04fF
C3434 a_5752_n9783# a_5949_n10301# 0.02fF
C3435 a_7130_n1597# a_7300_n2167# 0.04fF
C3436 a_3077_n5797# a_4365_n5797# 0.01fF
C3437 a_7237_n1597# a_7040_n2167# 0.02fF
C3438 a_4554_n1597# a_4724_n2167# 0.04fF
C3439 a_4661_n1597# a_4464_n2167# 0.02fF
C3440 a_13765_n13565# a_13765_n13021# 0.31fF
C3441 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.00fF
C3442 a_10994_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.04fF
C3443 a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C3444 a_7040_n10871# a_7300_n10871# 0.28fF
C3445 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_1/A 0.31fF
C3446 a_9813_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.02fF
C3447 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_8525_n5405# 0.01fF
C3448 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_8229_n10613# 0.01fF
C3449 a_2148_n5975# a_2148_n4887# 0.02fF
C3450 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1722_n4317# 0.00fF
C3451 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C3452 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_6012_n3255# 0.01fF
C3453 a_5586_n2685# VDD 0.76fF
C3454 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkinv_4_3/A 0.00fF
C3455 a_9450_n13021# a_9616_n11415# 0.00fF
C3456 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11164_n3255# 0.35fF
C3457 a_4464_n12503# a_4365_n10613# 0.00fF
C3458 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6012_n3799# 0.03fF
C3459 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.01fF
C3460 a_1789_n1909# a_1722_n2685# 0.01fF
C3461 a_10738_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.02fF
C3462 a_9450_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.03fF
C3463 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C3464 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9517_n821# 0.01fF
C3465 a_434_n5405# VDD 0.76fF
C3466 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C3467 a_9517_n10613# a_10805_n10613# 0.01fF
C3468 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C3469 a_9616_n2167# a_9450_n2685# 0.04fF
C3470 a_9517_n1909# a_9706_n2685# 0.02fF
C3471 a_4365_n11237# VDD 0.35fF
C3472 sky130_fd_sc_hd__nand2_4_1/A Ad_b 0.48fF
C3473 a_8525_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.12fF
C3474 a_5752_n2167# a_6941_n1909# 0.01fF
C3475 a_5653_n1909# a_7040_n2167# 0.01fF
C3476 a_11164_n5975# sky130_fd_sc_hd__clkinv_4_3/Y 0.31fF
C3477 a_3077_n11237# a_3266_n10301# 0.00fF
C3478 a_3176_n11415# a_3010_n10301# 0.00fF
C3479 a_797_n10301# a_600_n8695# 0.00fF
C3480 a_690_n10301# a_860_n8695# 0.00fF
C3481 a_6941_n8437# VDD 0.36fF
C3482 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VDD 0.83fF
C3483 a_8229_n1909# a_9517_n1909# 0.01fF
C3484 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.29fF
C3485 a_4554_n5405# VDD 0.47fF
C3486 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_4298_n1597# 0.03fF
C3487 a_9517_n13413# a_9706_n11933# 0.00fF
C3488 a_9616_n13591# a_9450_n11933# 0.00fF
C3489 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.02fF
C3490 a_10994_n11933# a_11164_n11415# 0.04fF
C3491 a_11101_n11933# a_10904_n11415# 0.02fF
C3492 a_860_n10871# a_690_n9213# 0.00fF
C3493 a_8162_n14109# VDD 0.75fF
C3494 sky130_fd_sc_hd__clkinv_4_1/Y VDD 2.17fF
C3495 a_600_n10871# a_797_n9213# 0.00fF
C3496 a_4724_n10871# VDD 0.78fF
C3497 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A VDD 0.89fF
C3498 a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C3499 a_797_n11933# a_1722_n11933# 0.02fF
C3500 a_690_n11933# a_1978_n11933# 0.01fF
C3501 a_9517_n5797# a_9450_n5405# 0.01fF
C3502 a_1789_n10613# a_3176_n10871# 0.01fF
C3503 a_1888_n10871# a_3077_n10613# 0.01fF
C3504 a_6941_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C3505 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_8229_n5797# 0.01fF
C3506 a_434_n11933# a_2085_n11933# 0.00fF
C3507 a_7040_n5975# a_7300_n5975# 0.28fF
C3508 a_9517_n8437# a_9706_n8125# 0.02fF
C3509 a_6941_n9525# a_8328_n9783# 0.01fF
C3510 sky130_fd_sc_hd__nand2_4_2/A VDD 7.13fF
C3511 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.00fF
C3512 a_4298_n9213# a_4554_n9213# 0.19fF
C3513 a_1789_n8437# a_1888_n9783# 0.00fF
C3514 a_10738_n11933# a_10805_n13413# 0.00fF
C3515 a_8328_n1079# a_8588_n1079# 0.28fF
C3516 a_1888_n8695# a_1789_n9525# 0.00fF
C3517 a_4365_n5797# a_4464_n5975# 0.49fF
C3518 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.04fF
C3519 a_7237_n2685# a_7237_n4317# 0.01fF
C3520 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_8328_n10871# 0.05fF
C3521 a_2085_n2685# a_2085_n4317# 0.01fF
C3522 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.04fF
C3523 Bd_b a_13765_n4861# 0.10fF
C3524 a_600_n5975# a_600_n4887# 0.01fF
C3525 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.09fF
C3526 a_9517_n11237# a_9706_n11933# 0.02fF
C3527 a_9517_n1909# sky130_fd_sc_hd__nand2_4_0/Y 0.08fF
C3528 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_10738_n2685# 0.03fF
C3529 a_8328_n4887# a_8328_n3799# 0.01fF
C3530 a_1789_n5797# sky130_fd_sc_hd__clkinv_4_4/A 0.07fF
C3531 sky130_fd_sc_hd__dfxbp_1_0/Q Bd_b 0.37fF
C3532 a_6012_n1079# VDD 0.78fF
C3533 a_600_n12503# a_n787_n12325# 0.01fF
C3534 a_797_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.12fF
C3535 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.08fF
C3536 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C3537 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_9876_n3255# 0.01fF
C3538 a_7130_n13021# a_8162_n13021# 0.02fF
C3539 a_6874_n13021# a_8418_n13021# 0.01fF
C3540 a_4464_n11415# a_4661_n13021# 0.00fF
C3541 a_4724_n11415# a_4554_n13021# 0.00fF
C3542 a_10805_n10613# a_10904_n10871# 0.48fF
C3543 a_1978_n5405# VDD 0.47fF
C3544 a_5052_n7283# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.02fF
C3545 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VDD 0.84fF
C3546 sky130_fd_sc_hd__nand2_4_2/A a_2729_n14109# 0.02fF
C3547 a_600_n11415# a_690_n10301# 0.01fF
C3548 a_6941_n1909# a_7300_n2167# 0.05fF
C3549 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_600_n13591# 0.04fF
C3550 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4365_n4709# 0.01fF
C3551 a_4298_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.03fF
C3552 a_434_n2685# a_797_n2685# 0.05fF
C3553 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9706_n509# 0.03fF
C3554 a_8229_n2997# a_9517_n2997# 0.01fF
C3555 a_3077_n3621# a_3010_n5405# 0.00fF
C3556 a_9813_n13021# VDD 0.33fF
C3557 a_8418_n509# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C3558 a_8525_n509# a_9813_n509# 0.01fF
C3559 a_5586_n5405# a_7130_n5405# 0.01fF
C3560 a_5842_n5405# a_6874_n5405# 0.02fF
C3561 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C3562 a_1722_n11933# a_1978_n11933# 0.19fF
C3563 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.04fF
C3564 a_9517_n4709# a_9706_n4317# 0.02fF
C3565 a_9616_n4887# a_9450_n4317# 0.04fF
C3566 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.02fF
C3567 a_9706_n14109# VDD 0.45fF
C3568 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VDD 0.83fF
C3569 a_7300_n5975# a_8588_n5975# 0.01fF
C3570 a_3077_n10613# a_3436_n10871# 0.05fF
C3571 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X a_8328_n5975# 0.05fF
C3572 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_3010_n11933# 0.00fF
C3573 a_8229_n9525# a_8588_n9783# 0.05fF
C3574 a_10904_n4887# a_10994_n5405# 0.02fF
C3575 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.04fF
C3576 a_4365_n10613# a_4554_n10301# 0.02fF
C3577 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.04fF
C3578 a_4661_n9213# a_5586_n9213# 0.02fF
C3579 a_4554_n9213# a_5842_n9213# 0.01fF
C3580 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_10805_n8437# 0.01fF
C3581 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkinv_4_3/A 0.44fF
C3582 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6012_n2167# 0.03fF
C3583 a_9517_n11237# a_9706_n10301# 0.00fF
C3584 a_5949_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C3585 a_4298_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.00fF
C3586 a_10805_n2997# a_10904_n3255# 0.48fF
C3587 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.03fF
C3588 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_7237_n10301# 0.01fF
C3589 a_501_n10613# a_860_n10871# 0.05fF
C3590 a_4365_n3621# a_4298_n2685# 0.00fF
C3591 a_n2602_n7037# a_n2248_n7037# 0.17fF
C3592 a_13765_n9757# p2 0.06fF
C3593 a_7040_n3255# VDD 0.46fF
C3594 sky130_fd_sc_hd__dfxbp_1_1/D a_n1139_n6715# 0.21fF
C3595 sky130_fd_sc_hd__nand2_1_4/B a_n428_n9783# 0.15fF
C3596 a_n1738_n6671# a_n1612_n7037# 0.03fF
C3597 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_1722_n4317# 0.00fF
C3598 a_7040_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.03fF
C3599 a_8162_n8125# a_9706_n8125# 0.01fF
C3600 a_10904_n2167# sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C3601 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VDD 0.84fF
C3602 a_11164_n2167# a_11101_n2685# 0.01fF
C3603 a_3176_n5975# sky130_fd_sc_hd__clkinv_4_4/A 0.07fF
C3604 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Ad_b 0.04fF
C3605 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.04fF
C3606 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VDD 0.83fF
C3607 a_10904_n13591# a_10994_n13021# 0.01fF
C3608 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.02fF
C3609 a_10904_n3255# a_9517_n2997# 0.01fF
C3610 a_860_n12503# a_860_n11415# 0.02fF
C3611 a_n428_n4887# VDD 0.83fF
C3612 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_3010_n1597# 0.00fF
C3613 a_8162_n13021# a_8525_n13021# 0.05fF
C3614 a_860_n11415# VDD 0.78fF
C3615 a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C3616 a_7237_n14109# a_8418_n14109# 0.01fF
C3617 a_7130_n14109# a_8525_n14109# 0.01fF
C3618 a_434_n4317# a_690_n4317# 0.19fF
C3619 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.06fF
C3620 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C3621 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_860_n3799# 0.00fF
C3622 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_11101_n11933# 0.02fF
C3623 a_860_n12503# sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C3624 a_5949_n10301# a_5949_n9213# 0.02fF
C3625 a_5586_n13021# a_5949_n13021# 0.05fF
C3626 a_9517_n12325# VDD 0.35fF
C3627 a_4661_n4317# a_4724_n4887# 0.01fF
C3628 a_797_n2685# a_1978_n2685# 0.01fF
C3629 a_690_n2685# a_2085_n2685# 0.01fF
C3630 a_7237_n8125# sky130_fd_sc_hd__clkinv_1_5/A 0.00fF
C3631 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C3632 sky130_fd_sc_hd__clkinv_4_7/A VDD 5.79fF
C3633 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1722_n2685# 0.35fF
C3634 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.29fF
C3635 a_2148_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C3636 a_1978_n11933# a_3266_n11933# 0.01fF
C3637 a_1722_n11933# a_3373_n11933# 0.00fF
C3638 a_2085_n11933# a_3010_n11933# 0.02fF
C3639 a_9876_n3255# VDD 0.74fF
C3640 a_9706_n6493# VDD 0.47fF
C3641 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_4365_n10613# 0.18fF
C3642 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.02fF
C3643 a_501_n1909# a_n688_n2167# 0.01fF
C3644 a_600_n2167# a_n787_n1909# 0.01fF
C3645 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C3646 a_2085_n5405# a_1888_n4887# 0.02fF
C3647 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X a_2085_n9213# 0.01fF
C3648 a_8418_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.07fF
C3649 a_6941_n5797# a_6794_n7203# 0.00fF
C3650 a_13765_n5405# A 0.12fF
C3651 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X a_6658_n7363# 0.00fF
C3652 a_7300_n5975# a_6665_n7459# 0.00fF
C3653 a_7040_n5975# a_6865_n7304# 0.00fF
C3654 A_b a_13765_n5949# 0.12fF
C3655 a_9876_n8695# a_11164_n8695# 0.01fF
C3656 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_10904_n8695# 0.05fF
C3657 a_9616_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.00fF
C3658 a_5586_n1597# VDD 0.76fF
C3659 a_2148_n11415# a_2148_n10871# 0.09fF
C3660 a_8229_n11237# a_8328_n10871# 0.01fF
C3661 a_8328_n11415# a_8229_n10613# 0.01fF
C3662 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.02fF
C3663 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_7040_n1079# 0.00fF
C3664 a_5842_n4317# a_5752_n5975# 0.00fF
C3665 a_4661_n10301# a_4724_n8695# 0.00fF
C3666 a_5842_n10301# a_6874_n10301# 0.02fF
C3667 a_5586_n10301# a_7130_n10301# 0.01fF
C3668 a_7040_n8695# a_7237_n10301# 0.00fF
C3669 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.02fF
C3670 a_6874_n11933# a_7130_n11933# 0.19fF
C3671 a_7300_n8695# a_7130_n10301# 0.00fF
C3672 a_8588_n3255# VDD 0.77fF
C3673 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C3674 a_7237_n5405# a_7040_n5975# 0.02fF
C3675 a_7130_n5405# a_7300_n5975# 0.04fF
C3676 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_8588_n8695# 0.03fF
C3677 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.00fF
C3678 a_4724_n5975# sky130_fd_sc_hd__clkinv_4_4/A 0.11fF
C3679 a_690_n9213# a_600_n9783# 0.02fF
C3680 a_6874_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C3681 a_9616_n10871# a_9706_n11933# 0.01fF
C3682 a_6941_n13413# VDD 0.35fF
C3683 a_8525_n13021# a_9706_n13021# 0.01fF
C3684 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Ad_b 0.02fF
C3685 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n13021# 0.35fF
C3686 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__clkinv_1_5/A 0.05fF
C3687 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/Y 0.73fF
C3688 a_4298_n11933# a_5949_n11933# 0.00fF
C3689 a_3077_n2997# a_3077_n4709# 0.00fF
C3690 a_4554_n11933# a_5842_n11933# 0.01fF
C3691 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X 0.01fF
C3692 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_2148_n3255# 0.01fF
C3693 a_4365_n3621# a_4365_n1909# 0.00fF
C3694 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C3695 a_n688_n4887# a_n428_n4887# 0.28fF
C3696 a_5653_n8437# a_5586_n9213# 0.01fF
C3697 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.14fF
C3698 a_n688_n9783# a_600_n9783# 0.01fF
C3699 sky130_fd_sc_hd__dfxbp_1_0/Q a_5052_n7283# 0.37fF
C3700 a_n428_n9783# a_501_n9525# 0.02fF
C3701 a_4623_n7349# a_6006_n7607# 0.01fF
C3702 a_8162_n509# a_9450_n509# 0.01fF
C3703 a_n787_n9525# a_860_n9783# 0.00fF
C3704 a_4464_n4887# a_5653_n4709# 0.01fF
C3705 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C3706 a_4365_n4709# a_5752_n4887# 0.01fF
C3707 p2d_b p2 0.08fF
C3708 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C3709 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_9876_n9783# 0.01fF
C3710 a_600_n1079# a_2148_n1079# 0.01fF
C3711 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C3712 a_860_n1079# a_1888_n1079# 0.02fF
C3713 a_10904_n12503# VDD 0.39fF
C3714 a_1978_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.05fF
C3715 a_4464_n3799# a_4554_n5405# 0.00fF
C3716 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.12fF
C3717 a_9450_n1597# a_9616_n1079# 0.04fF
C3718 a_6941_n11237# VDD 0.35fF
C3719 a_9706_n1597# a_9517_n821# 0.02fF
C3720 a_3010_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.03fF
C3721 a_3266_n11933# a_3373_n11933# 0.55fF
C3722 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_4298_n11933# 0.00fF
C3723 a_10904_n4887# a_11101_n4317# 0.02fF
C3724 a_501_n3621# VDD 0.36fF
C3725 a_10805_n4709# sky130_fd_sc_hd__clkinv_4_3/A 0.07fF
C3726 a_4365_n5797# a_4298_n5405# 0.01fF
C3727 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Ad_b 0.02fF
C3728 a_4464_n10871# a_4298_n9213# 0.00fF
C3729 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C3730 a_797_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.12fF
C3731 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3732 a_13765_n11933# p2d_b 0.02fF
C3733 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.02fF
C3734 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C3735 a_6874_n4317# a_7040_n3255# 0.00fF
C3736 a_7130_n4317# a_6941_n2997# 0.00fF
C3737 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.00fF
C3738 a_10805_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.05fF
C3739 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C3740 a_1789_n2997# a_1888_n4887# 0.00fF
C3741 a_10994_n13021# sky130_fd_sc_hd__clkinv_4_7/Y 0.01fF
C3742 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A VDD 0.88fF
C3743 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_8588_n1079# 0.29fF
C3744 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.04fF
C3745 a_6874_n10301# a_7237_n10301# 0.05fF
C3746 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6941_n5797# 0.00fF
C3747 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C3748 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VDD 0.87fF
C3749 a_7130_n11933# a_8418_n11933# 0.01fF
C3750 a_7237_n11933# a_8162_n11933# 0.02fF
C3751 a_5752_n3799# a_5842_n2685# 0.01fF
C3752 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__nand2_4_0/A 2.16fF
C3753 a_10738_n6173# a_11164_n4887# 0.01fF
C3754 a_6874_n11933# a_8525_n11933# 0.00fF
C3755 a_9616_n10871# a_9706_n10301# 0.02fF
C3756 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_860_n1079# 0.03fF
C3757 a_797_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.01fF
C3758 a_1888_n4887# a_1722_n4317# 0.04fF
C3759 a_1789_n4709# a_1978_n4317# 0.02fF
C3760 a_1722_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C3761 a_8418_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C3762 a_8328_n13591# VDD 0.43fF
C3763 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1789_n9525# 0.01fF
C3764 a_3176_n10871# a_3077_n9525# 0.00fF
C3765 a_3077_n10613# a_3176_n9783# 0.00fF
C3766 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_7300_n13591# 0.01fF
C3767 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C3768 a_10805_n8437# a_10738_n9213# 0.01fF
C3769 a_4365_n13413# a_4298_n11933# 0.00fF
C3770 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Bd_b 0.05fF
C3771 a_5586_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.03fF
C3772 a_8328_n8695# a_8418_n10301# 0.00fF
C3773 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_6874_n11933# 0.00fF
C3774 a_8328_n9783# a_8525_n9213# 0.02fF
C3775 a_8588_n9783# a_8418_n9213# 0.04fF
C3776 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_1789_n1909# 0.18fF
C3777 a_860_n2167# a_1888_n2167# 0.02fF
C3778 a_600_n2167# a_2148_n2167# 0.01fF
C3779 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_860_n4887# 0.01fF
C3780 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.03fF
C3781 a_5949_n5405# a_6874_n5405# 0.02fF
C3782 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_7237_n8125# 0.01fF
C3783 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A VDD 0.88fF
C3784 a_6874_n2685# a_5842_n2685# 0.02fF
C3785 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkinv_1_4/Y 0.31fF
C3786 a_7130_n2685# a_5586_n2685# 0.01fF
C3787 a_501_n10613# a_600_n9783# 0.00fF
C3788 a_6941_n12325# a_8328_n12503# 0.01fF
C3789 a_7040_n12503# a_8229_n12325# 0.01fF
C3790 a_5653_n4709# a_6012_n4887# 0.05fF
C3791 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.04fF
C3792 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_3176_n1079# 0.01fF
C3793 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.02fF
C3794 a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.00fF
C3795 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_5586_n5405# 0.00fF
C3796 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.02fF
C3797 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_860_n13591# 0.03fF
C3798 a_797_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C3799 a_8328_n11415# VDD 0.44fF
C3800 a_9517_n1909# VDD 0.34fF
C3801 a_3266_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C3802 a_3373_n11933# a_4661_n11933# 0.01fF
C3803 a_5842_n2685# a_6012_n3799# 0.00fF
C3804 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4554_n11933# 0.03fF
C3805 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_7300_n12503# 0.01fF
C3806 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C3807 a_1888_n3799# VDD 0.44fF
C3808 a_9706_n6493# a_9706_n5405# 0.01fF
C3809 A Ad_b 0.26fF
C3810 a_501_n12325# a_600_n10871# 0.00fF
C3811 a_10904_n13591# a_11164_n13591# 0.22fF
C3812 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.02fF
C3813 a_4464_n9783# a_4661_n9213# 0.02fF
C3814 a_4724_n9783# a_4554_n9213# 0.04fF
C3815 a_9706_n1597# a_9706_n509# 0.01fF
C3816 a_7130_n14109# a_7300_n13591# 0.04fF
C3817 a_7237_n14109# a_7040_n13591# 0.02fF
C3818 a_5653_n10613# a_5842_n11933# 0.00fF
C3819 a_9616_n8695# a_9616_n9783# 0.01fF
C3820 a_600_n11415# a_690_n11933# 0.02fF
C3821 a_4365_n3621# a_4298_n4317# 0.01fF
C3822 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C3823 a_10904_n13591# a_9517_n13413# 0.01fF
C3824 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.03fF
C3825 a_6373_n7349# p2 0.01fF
C3826 a_6658_n7363# a_6794_n7203# 0.30fF
C3827 a_6665_n7459# a_6865_n7304# 0.26fF
C3828 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.09fF
C3829 a_5752_n3799# a_5752_n3255# 0.07fF
C3830 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.00fF
C3831 a_7237_n4317# a_7300_n5975# 0.00fF
C3832 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n10301# 0.35fF
C3833 a_9616_n5975# a_9706_n4317# 0.00fF
C3834 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C3835 a_8588_n10871# a_8229_n10613# 0.05fF
C3836 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_9450_n11933# 0.00fF
C3837 a_8162_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.03fF
C3838 a_8418_n11933# a_8525_n11933# 0.55fF
C3839 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_10738_n10301# 0.03fF
C3840 a_6874_n509# a_6941_n821# 0.01fF
C3841 a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C3842 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X a_4661_n10301# 0.00fF
C3843 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C3844 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_8588_n5975# 0.03fF
C3845 a_10994_n5405# a_11164_n5975# 0.04fF
C3846 sky130_fd_sc_hd__clkinv_4_4/A a_10805_n5797# 0.07fF
C3847 a_11101_n5405# a_10904_n5975# 0.02fF
C3848 a_7300_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C3849 sky130_fd_sc_hd__nand2_4_3/Y a_13765_n10301# 0.04fF
C3850 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.02fF
C3851 p1 VDD 4.14fF
C3852 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C3853 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_9876_n11415# 0.01fF
C3854 sky130_fd_sc_hd__clkinv_4_8/Y a_10805_n13413# 0.01fF
C3855 a_4724_n5975# a_5653_n5797# 0.02fF
C3856 a_4464_n5975# a_5752_n5975# 0.01fF
C3857 a_4365_n5797# a_6012_n5975# 0.00fF
C3858 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.00fF
C3859 a_8162_n8125# a_8328_n9783# 0.00fF
C3860 a_9876_n13591# VDD 0.73fF
C3861 p2 VDD 7.12fF
C3862 a_8328_n2167# a_8525_n509# 0.00fF
C3863 a_8588_n2167# a_8418_n509# 0.00fF
C3864 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_860_n5975# 0.00fF
C3865 a_8162_n10301# a_8418_n10301# 0.19fF
C3866 a_8229_n9525# a_8328_n10871# 0.00fF
C3867 a_3436_n8695# a_3436_n9783# 0.02fF
C3868 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_10738_n509# 0.00fF
C3869 a_4365_n9525# a_4365_n8437# 0.02fF
C3870 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_3176_n2167# 0.01fF
C3871 a_1888_n1079# a_3176_n1079# 0.01fF
C3872 a_6874_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.03fF
C3873 a_7130_n5405# a_7237_n5405# 0.55fF
C3874 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_8162_n5405# 0.00fF
C3875 a_2148_n1079# a_3077_n821# 0.02fF
C3876 a_8229_n12325# a_8588_n12503# 0.05fF
C3877 sky130_fd_sc_hd__nand2_1_0/A a_501_n4709# 0.01fF
C3878 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X a_6941_n4709# 0.18fF
C3879 a_6012_n4887# a_7040_n4887# 0.02fF
C3880 a_13765_n11933# VDD 2.48fF
C3881 a_797_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.12fF
C3882 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_3373_n2685# 0.01fF
C3883 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C3884 sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.33fF
C3885 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.00fF
C3886 a_3077_n2997# a_3436_n3255# 0.05fF
C3887 a_2148_n3255# VDD 0.78fF
C3888 a_6373_n7349# a_6593_n7215# 0.01fF
C3889 sky130_fd_sc_hd__clkinv_4_4/A a_434_n5405# 0.00fF
C3890 a_10904_n2167# VDD 0.41fF
C3891 a_4661_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.12fF
C3892 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X sky130_fd_sc_hd__clkinv_1_5/A 0.04fF
C3893 a_501_n12325# sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C3894 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_5752_n4887# 0.00fF
C3895 a_7300_n4887# a_6012_n4887# 0.01fF
C3896 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.06fF
C3897 a_6012_n10871# a_5842_n9213# 0.00fF
C3898 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C3899 a_4365_n11237# a_4554_n11933# 0.02fF
C3900 a_4464_n11415# a_4298_n11933# 0.04fF
C3901 a_8418_n4317# a_8588_n3255# 0.00fF
C3902 a_8525_n4317# a_8328_n3255# 0.00fF
C3903 a_8525_n10301# a_8418_n11933# 0.00fF
C3904 a_6941_n10613# a_6874_n9213# 0.00fF
C3905 a_4365_n821# a_4298_n2685# 0.00fF
C3906 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X Bd_b 0.03fF
C3907 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6658_n7363# 0.02fF
C3908 a_2085_n1597# a_2148_n1079# 0.01fF
C3909 a_10805_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C3910 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_10738_n4317# 0.00fF
C3911 a_10738_n13789# VDD 0.11fF
C3912 a_9876_n10871# a_8328_n10871# 0.01fF
C3913 a_5949_n13021# a_6012_n13591# 0.01fF
C3914 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_9706_n11933# 0.03fF
C3915 a_6941_n9525# VDD 0.35fF
C3916 a_9813_n8125# sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C3917 a_11164_n10871# a_11101_n10301# 0.01fF
C3918 a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.01fF
C3919 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkinv_1_3/A 0.84fF
C3920 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.03fF
C3921 a_3176_n4887# a_3373_n4317# 0.02fF
C3922 a_n2602_n7037# a_n2436_n7037# 1.73fF
C3923 a_9517_n4709# VDD 0.35fF
C3924 a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C3925 a_4724_n10871# a_4554_n11933# 0.00fF
C3926 a_4464_n10871# a_4661_n11933# 0.00fF
C3927 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.06fF
C3928 a_n2163_n6671# a_n2248_n7037# 0.09fF
C3929 a_n1570_n6769# a_n1139_n6715# 0.24fF
C3930 a_8162_n2685# a_8162_n1597# 0.02fF
C3931 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6874_n5405# 0.01fF
C3932 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C3933 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.06fF
C3934 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C3935 a_7237_n5405# a_8525_n5405# 0.01fF
C3936 a_7130_n2685# a_7040_n3255# 0.02fF
C3937 a_9616_n2167# a_9616_n1079# 0.01fF
C3938 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8418_n5405# 0.03fF
C3939 a_7130_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C3940 a_9616_n8695# a_9813_n9213# 0.02fF
C3941 a_1789_n13413# a_1722_n13021# 0.01fF
C3942 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_4365_n821# 0.01fF
C3943 a_3176_n1079# a_3436_n1079# 0.28fF
C3944 a_3077_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.02fF
C3945 a_5949_n13021# a_6012_n11415# 0.00fF
C3946 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_1789_n4709# 0.18fF
C3947 a_600_n4887# a_2148_n4887# 0.01fF
C3948 a_860_n4887# a_1888_n4887# 0.02fF
C3949 VDD a_2085_n9213# 0.36fF
C3950 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Bd_b 0.02fF
C3951 a_8418_n6493# a_8229_n5797# 0.02fF
C3952 a_8162_n6493# a_8328_n5975# 0.04fF
C3953 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_3010_n2685# 0.03fF
C3954 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.02fF
C3955 a_2148_n5975# VDD 0.79fF
C3956 clk sky130_fd_sc_hd__clkinv_1_5/A 0.06fF
C3957 a_7237_n2685# a_7300_n1079# 0.00fF
C3958 a_3176_n3255# a_4724_n3255# 0.01fF
C3959 a_3436_n3255# a_4464_n3255# 0.02fF
C3960 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_4365_n2997# 0.18fF
C3961 a_501_n1909# VDD 0.36fF
C3962 a_3176_n3799# a_1789_n3621# 0.01fF
C3963 a_3077_n3621# a_1888_n3799# 0.01fF
C3964 a_10738_n1597# sky130_fd_sc_hd__clkinv_4_1/Y 0.00fF
C3965 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.06fF
C3966 a_10994_n1597# a_11101_n1597# 0.55fF
C3967 a_1978_n10301# a_2085_n9213# 0.00fF
C3968 a_13765_n5405# Ad 0.15fF
C3969 A_b a_13765_n4861# 0.15fF
C3970 a_8588_n10871# VDD 0.78fF
C3971 a_600_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C3972 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C3973 a_10805_n10613# a_10805_n12325# 0.00fF
C3974 a_9706_n10301# a_9706_n9213# 0.01fF
C3975 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_3010_n9213# 0.03fF
C3976 a_7300_n10871# a_7130_n11933# 0.00fF
C3977 a_7040_n10871# a_7237_n11933# 0.00fF
C3978 a_6874_n6493# VDD 0.76fF
C3979 a_2366_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C3980 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C3981 a_2622_n8125# a_2729_n8125# 0.54fF
C3982 a_9813_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.02fF
C3983 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_8525_n9213# 0.01fF
C3984 a_10904_n5975# sky130_fd_sc_hd__clkinv_4_3/A 0.16fF
C3985 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C3986 a_11164_n5975# a_11101_n4317# 0.00fF
C3987 a_9706_n6493# a_9813_n5405# 0.00fF
C3988 a_434_n10301# a_434_n9213# 0.02fF
C3989 a_6941_n1909# a_6941_n3621# 0.00fF
C3990 a_8418_n509# a_8328_n1079# 0.02fF
C3991 a_3077_n4709# a_4365_n4709# 0.01fF
C3992 a_5586_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.03fF
C3993 a_5842_n4317# a_5949_n4317# 0.55fF
C3994 a_10904_n4887# VDD 0.39fF
C3995 a_6874_n13021# a_7040_n12503# 0.04fF
C3996 a_7130_n13021# a_6941_n12325# 0.02fF
C3997 clk a_n1995_n6925# 0.01fF
C3998 a_7237_n4317# a_7237_n5405# 0.02fF
C3999 a_4365_n821# a_4365_n1909# 0.02fF
C4000 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C4001 a_5949_n9213# a_6006_n7607# 0.00fF
C4002 a_9450_n8125# a_10738_n8125# 0.01fF
C4003 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C4004 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8229_n2997# 0.01fF
C4005 a_8525_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.12fF
C4006 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C4007 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_3436_n9783# 0.00fF
C4008 a_3176_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C4009 a_4464_n9783# a_4365_n11237# 0.00fF
C4010 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_4464_n1079# 0.05fF
C4011 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkinv_1_3/A 0.08fF
C4012 a_4365_n9525# a_4464_n11415# 0.00fF
C4013 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.85fF
C4014 a_3436_n1079# a_4724_n1079# 0.01fF
C4015 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C4016 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.89fF
C4017 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_3176_n4887# 0.01fF
C4018 a_3436_n2167# a_3373_n2685# 0.01fF
C4019 a_4298_n5405# a_5586_n5405# 0.01fF
C4020 a_8229_n1909# a_8162_n1597# 0.01fF
C4021 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VDD 0.85fF
C4022 a_9616_n2167# a_9813_n509# 0.00fF
C4023 a_9876_n2167# a_9706_n509# 0.00fF
C4024 sky130_fd_sc_hd__mux2_1_0/X Bd_b 0.05fF
C4025 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X a_7300_n3255# 0.01fF
C4026 a_4464_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.03fF
C4027 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C4028 a_3077_n1909# a_3176_n3255# 0.00fF
C4029 a_3176_n2167# a_3077_n2997# 0.00fF
C4030 a_5653_n821# a_5752_n1079# 0.49fF
C4031 a_9616_n11415# a_10805_n11237# 0.01fF
C4032 a_9813_n13021# a_9706_n11933# 0.00fF
C4033 a_4724_n10871# a_5653_n10613# 0.02fF
C4034 a_4464_n10871# a_5752_n10871# 0.01fF
C4035 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD 0.84fF
C4036 a_8525_n10301# a_9813_n10301# 0.01fF
C4037 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9706_n10301# 0.03fF
C4038 a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C4039 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_4661_n2685# 0.01fF
C4040 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C4041 a_8328_n10871# a_8418_n9213# 0.00fF
C4042 a_8418_n6493# VDD 0.48fF
C4043 a_434_n9213# VDD 0.77fF
C4044 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Bd_b 0.03fF
C4045 a_4464_n3255# a_4464_n2167# 0.01fF
C4046 a_9517_n11237# a_9517_n10613# 0.05fF
C4047 a_1888_n11415# a_1722_n13021# 0.00fF
C4048 a_1789_n11237# a_1978_n13021# 0.00fF
C4049 a_860_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.29fF
C4050 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.06fF
C4051 a_4464_n1079# a_6012_n1079# 0.01fF
C4052 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_5653_n821# 0.18fF
C4053 a_4724_n1079# a_5752_n1079# 0.02fF
C4054 a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.02fF
C4055 a_600_n8695# a_860_n8695# 0.28fF
C4056 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C4057 a_3077_n8437# VDD 0.36fF
C4058 a_8229_n4709# a_8162_n4317# 0.01fF
C4059 a_8162_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.07fF
C4060 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.73fF
C4061 a_9616_n5975# a_8229_n5797# 0.01fF
C4062 a_n787_n9525# VDD 0.35fF
C4063 a_9517_n5797# a_8328_n5975# 0.01fF
C4064 a_5949_n4317# a_7237_n4317# 0.01fF
C4065 a_5842_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C4066 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_7130_n4317# 0.03fF
C4067 a_9517_n4709# a_9706_n5405# 0.02fF
C4068 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__nand2_4_3/A 0.11fF
C4069 a_9616_n4887# a_9450_n5405# 0.04fF
C4070 a_9706_n2685# a_9706_n1597# 0.01fF
C4071 a_7237_n509# VDD 0.34fF
C4072 a_6874_n9213# a_6658_n7363# 0.00fF
C4073 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_5949_n10301# 0.00fF
C4074 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C4075 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_3373_n1597# 0.00fF
C4076 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C4077 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_3373_n4317# 0.00fF
C4078 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C4079 a_11164_n2167# a_11164_n1079# 0.02fF
C4080 a_8525_n2685# a_8588_n3255# 0.01fF
C4081 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.29fF
C4082 a_3176_n13591# a_3266_n13021# 0.01fF
C4083 a_10738_n9213# sky130_fd_sc_hd__clkinv_1_3/A 0.00fF
C4084 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.02fF
C4085 a_1888_n12503# a_1888_n13591# 0.01fF
C4086 a_3077_n13413# VDD 0.35fF
C4087 a_5586_n5405# a_5842_n5405# 0.19fF
C4088 a_10805_n3621# a_9517_n3621# 0.01fF
C4089 a_4724_n12503# a_4724_n13591# 0.02fF
C4090 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.88fF
C4091 a_10904_n2167# sky130_fd_sc_hd__nand2_4_0/B 0.00fF
C4092 a_7130_n9213# VDD 0.44fF
C4093 a_5653_n821# a_7300_n1079# 0.00fF
C4094 Ad_b Ad 0.60fF
C4095 a_5752_n1079# a_7040_n1079# 0.01fF
C4096 a_1789_n5797# a_3077_n5797# 0.01fF
C4097 a_6012_n1079# a_6941_n821# 0.02fF
C4098 a_9616_n12503# a_9450_n11933# 0.04fF
C4099 a_9517_n12325# a_9706_n11933# 0.02fF
C4100 a_10805_n11237# a_11164_n11415# 0.05fF
C4101 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_6941_n10613# 0.01fF
C4102 p2d p2 0.20fF
C4103 a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.02fF
C4104 a_5752_n10871# a_6012_n10871# 0.28fF
C4105 a_9813_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.12fF
C4106 a_4298_n1597# a_4365_n821# 0.01fF
C4107 a_600_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.04fF
C4108 a_3010_n2685# VDD 0.76fF
C4109 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.01fF
C4110 sky130_fd_sc_hd__clkinv_4_8/A a_7040_n12503# 0.04fF
C4111 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.29fF
C4112 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_9876_n3255# 0.01fF
C4113 a_3176_n12503# a_3077_n10613# 0.00fF
C4114 a_3077_n12325# a_3176_n10871# 0.00fF
C4115 a_1978_n9213# VDD 0.45fF
C4116 a_9813_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C4117 a_5842_n5405# a_5752_n5975# 0.01fF
C4118 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_7040_n1079# 0.01fF
C4119 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.02fF
C4120 a_4464_n8695# VDD 0.51fF
C4121 a_9706_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.08fF
C4122 a_1978_n10301# a_1978_n9213# 0.01fF
C4123 a_1789_n11237# VDD 0.35fF
C4124 a_9517_n8437# VDD 0.34fF
C4125 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9876_n3255# 0.03fF
C4126 a_5752_n11415# a_5586_n11933# 0.04fF
C4127 a_600_n12503# a_501_n10613# 0.00fF
C4128 a_9813_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C4129 a_1888_n3255# a_1888_n3799# 0.07fF
C4130 a_7237_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.12fF
C4131 a_4464_n2167# a_5653_n1909# 0.01fF
C4132 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C4133 a_3266_n10301# a_3176_n8695# 0.00fF
C4134 a_1789_n11237# a_1978_n10301# 0.00fF
C4135 a_1888_n11415# a_1722_n10301# 0.00fF
C4136 a_8418_n13021# a_8588_n12503# 0.04fF
C4137 p2_b a_13765_n9757# 0.15fF
C4138 a_8525_n13021# a_8328_n12503# 0.02fF
C4139 a_4554_n1597# a_3266_n1597# 0.01fF
C4140 a_4661_n1597# a_3010_n1597# 0.00fF
C4141 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.04fF
C4142 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_860_n13591# 0.00fF
C4143 a_797_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.00fF
C4144 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C4145 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.29fF
C4146 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VDD 0.92fF
C4147 a_8229_n13413# a_8418_n11933# 0.00fF
C4148 a_8328_n13591# a_8162_n11933# 0.00fF
C4149 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.02fF
C4150 a_2148_n3799# a_2085_n4317# 0.01fF
C4151 a_9813_n11933# a_9616_n11415# 0.02fF
C4152 a_9813_n13021# a_10738_n13021# 0.02fF
C4153 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_4298_n13021# 0.03fF
C4154 a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C4155 a_600_n10871# a_1789_n10613# 0.01fF
C4156 a_5752_n5975# a_6012_n5975# 0.28fF
C4157 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X a_6941_n5797# 0.01fF
C4158 a_5653_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.02fF
C4159 a_9616_n5975# VDD 0.42fF
C4160 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkinv_1_3/A 0.01fF
C4161 Bd a_13765_n1053# 0.06fF
C4162 a_434_n4317# a_434_n5405# 0.02fF
C4163 a_4464_n13591# VDD 0.48fF
C4164 a_7040_n3799# a_6941_n4709# 0.00fF
C4165 a_6941_n3621# a_7040_n4887# 0.00fF
C4166 a_797_n2685# a_860_n3255# 0.01fF
C4167 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_690_n11933# 0.02fF
C4168 a_8525_n9213# VDD 0.35fF
C4169 a_3010_n9213# a_3266_n9213# 0.19fF
C4170 a_3077_n5797# a_3176_n5975# 0.49fF
C4171 a_7040_n1079# a_7300_n1079# 0.28fF
C4172 a_6941_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.02fF
C4173 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X a_8229_n821# 0.01fF
C4174 a_8588_n2167# a_8588_n3255# 0.02fF
C4175 a_5752_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C4176 a_10994_n1597# a_11164_n3255# 0.00fF
C4177 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_7040_n10871# 0.05fF
C4178 a_6012_n10871# a_7300_n10871# 0.01fF
C4179 a_11101_n1597# a_10904_n3255# 0.00fF
C4180 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.04fF
C4181 a_n1995_n6925# sky130_fd_sc_hd__clkinv_1_5/A 0.11fF
C4182 a_9813_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.01fF
C4183 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.03fF
C4184 a_8229_n11237# a_8418_n11933# 0.02fF
C4185 a_8328_n11415# a_8162_n11933# 0.04fF
C4186 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C4187 a_4554_n2685# VDD 0.44fF
C4188 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6101_n7254# 0.00fF
C4189 a_501_n11237# a_600_n11415# 0.49fF
C4190 sky130_fd_sc_hd__clkinv_4_8/A a_8588_n12503# 0.10fF
C4191 a_10738_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.02fF
C4192 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C4193 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.08fF
C4194 sky130_fd_sc_hd__mux2_1_0/X a_5052_n7283# 0.02fF
C4195 a_5842_n13021# a_6874_n13021# 0.02fF
C4196 a_1888_n3255# a_2148_n3255# 0.28fF
C4197 a_3436_n11415# a_3266_n13021# 0.00fF
C4198 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C4199 a_3176_n11415# a_3373_n13021# 0.00fF
C4200 a_6012_n8695# VDD 0.78fF
C4201 a_9517_n10613# a_9616_n10871# 0.49fF
C4202 a_3176_n11415# VDD 0.44fF
C4203 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X a_4724_n12503# 0.01fF
C4204 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C4205 a_8588_n11415# a_8588_n9783# 0.01fF
C4206 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.02fF
C4207 a_5653_n1909# a_6012_n2167# 0.05fF
C4208 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4365_n8437# 0.00fF
C4209 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C4210 a_6941_n2997# a_8229_n2997# 0.01fF
C4211 a_5586_n13021# a_4661_n13021# 0.02fF
C4212 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.02fF
C4213 a_3436_n2167# a_3373_n1597# 0.01fF
C4214 a_3373_n5405# VDD 0.35fF
C4215 a_10994_n13021# a_11101_n13021# 0.55fF
C4216 a_10738_n13021# sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C4217 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.02fF
C4218 a_10805_n8437# a_11164_n8695# 0.05fF
C4219 a_8162_n8125# VDD 0.78fF
C4220 a_n2436_n7037# a_n2163_n6671# 0.25fF
C4221 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C4222 a_4724_n13591# a_4661_n13021# 0.01fF
C4223 a_1789_n10613# a_2148_n10871# 0.05fF
C4224 a_5752_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C4225 a_6012_n5975# a_7300_n5975# 0.01fF
C4226 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_7040_n5975# 0.05fF
C4227 a_11164_n5975# VDD 0.67fF
C4228 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_1722_n11933# 0.00fF
C4229 sky130_fd_sc_hd__clkinv_4_4/A p2 0.16fF
C4230 a_3436_n12503# a_3436_n13591# 0.02fF
C4231 a_501_n1909# a_600_n1079# 0.00fF
C4232 a_797_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.12fF
C4233 a_3010_n9213# a_4661_n9213# 0.00fF
C4234 a_3266_n9213# a_4554_n9213# 0.01fF
C4235 a_3373_n9213# a_4298_n9213# 0.02fF
C4236 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_4724_n2167# 0.03fF
C4237 a_3176_n5975# a_4464_n5975# 0.01fF
C4238 a_3436_n5975# a_4365_n5797# 0.02fF
C4239 a_3077_n5797# a_4724_n5975# 0.00fF
C4240 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A a_8328_n1079# 0.05fF
C4241 a_7300_n1079# a_8588_n1079# 0.01fF
C4242 a_2148_n9783# sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C4243 a_4661_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C4244 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.03fF
C4245 a_7237_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C4246 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_5949_n10301# 0.01fF
C4247 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7300_n2167# 0.03fF
C4248 p1 p1_b 0.47fF
C4249 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.29fF
C4250 a_3077_n3621# a_3010_n2685# 0.00fF
C4251 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.04fF
C4252 p2_b p2d_b 0.20fF
C4253 a_2622_n509# VDD 0.50fF
C4254 a_5949_n2685# VDD 0.35fF
C4255 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Ad_b 0.12fF
C4256 a_9706_n13021# a_9876_n11415# 0.00fF
C4257 a_860_n11415# a_797_n13021# 0.00fF
C4258 a_11101_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.12fF
C4259 a_1888_n2167# a_1978_n2685# 0.01fF
C4260 sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# 0.58fF
C4261 a_9616_n3255# a_8229_n2997# 0.01fF
C4262 a_6874_n13021# a_7237_n13021# 0.05fF
C4263 a_9876_n2167# a_9706_n2685# 0.04fF
C4264 a_797_n5405# VDD 0.36fF
C4265 a_9616_n10871# a_10904_n10871# 0.01fF
C4266 a_9616_n2167# a_9813_n2685# 0.02fF
C4267 a_9517_n10613# a_11164_n10871# 0.00fF
C4268 a_9876_n10871# a_10805_n10613# 0.02fF
C4269 a_4724_n11415# VDD 0.77fF
C4270 a_13765_n11933# p1_b 0.06fF
C4271 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/A 0.69fF
C4272 p1d_b a_13765_n13021# 0.06fF
C4273 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A a_2366_n8125# 0.00fF
C4274 a_5752_n2167# a_7300_n2167# 0.01fF
C4275 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_6941_n1909# 0.18fF
C4276 a_6012_n2167# a_7040_n2167# 0.02fF
C4277 a_3373_n4317# a_3436_n4887# 0.01fF
C4278 a_8229_n2997# a_8328_n3255# 0.49fF
C4279 a_797_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.00fF
C4280 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_860_n8695# 0.00fF
C4281 a_3436_n11415# a_3266_n10301# 0.00fF
C4282 a_3176_n11415# a_3373_n10301# 0.00fF
C4283 a_5586_n5405# a_5949_n5405# 0.05fF
C4284 a_10805_n12325# a_10994_n13021# 0.02fF
C4285 a_8588_n2167# a_9517_n1909# 0.02fF
C4286 a_8328_n2167# a_9616_n2167# 0.01fF
C4287 a_6874_n1597# a_7040_n1079# 0.04fF
C4288 a_9876_n13591# a_9706_n11933# 0.00fF
C4289 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VDD 0.88fF
C4290 a_8229_n1909# a_9876_n2167# 0.00fF
C4291 a_10904_n12503# a_10738_n13021# 0.04fF
C4292 a_11101_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.12fF
C4293 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4294 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C4295 a_9876_n8695# a_9706_n8125# 0.04fF
C4296 a_1888_n10871# a_3436_n10871# 0.01fF
C4297 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_797_n9213# 0.00fF
C4298 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C4299 a_9616_n5975# a_9706_n5405# 0.01fF
C4300 a_2148_n10871# a_3176_n10871# 0.02fF
C4301 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_3077_n10613# 0.18fF
C4302 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.04fF
C4303 a_8525_n14109# VDD 0.33fF
C4304 a_797_n11933# a_2085_n11933# 0.01fF
C4305 a_690_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C4306 a_10994_n5405# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C4307 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1978_n11933# 0.03fF
C4308 a_7300_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.29fF
C4309 a_7040_n9783# a_8588_n9783# 0.01fF
C4310 a_7300_n9783# a_8328_n9783# 0.02fF
C4311 a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.01fF
C4312 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_10738_n5405# 0.03fF
C4313 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_5586_n9213# 0.00fF
C4314 a_4298_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.03fF
C4315 a_4554_n9213# a_4661_n9213# 0.55fF
C4316 a_8162_n1597# VDD 0.76fF
C4317 a_4464_n5975# a_4724_n5975# 0.28fF
C4318 a_10805_n1909# a_10994_n1597# 0.02fF
C4319 a_10904_n2167# a_10738_n1597# 0.04fF
C4320 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C4321 a_3010_n4317# VDD 0.76fF
C4322 a_7040_n11415# a_6941_n10613# 0.01fF
C4323 a_6941_n11237# a_7040_n10871# 0.01fF
C4324 a_4298_n10301# a_5842_n10301# 0.01fF
C4325 a_4554_n10301# a_5586_n10301# 0.02fF
C4326 a_9616_n3255# a_10904_n3255# 0.01fF
C4327 a_9876_n3255# a_10805_n2997# 0.02fF
C4328 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.02fF
C4329 a_6012_n3255# VDD 0.78fF
C4330 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.02fF
C4331 a_5949_n5405# a_5752_n5975# 0.02fF
C4332 a_860_n5975# a_860_n4887# 0.02fF
C4333 a_2366_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.34fF
C4334 a_9876_n2167# sky130_fd_sc_hd__nand2_4_0/Y 0.11fF
C4335 a_8588_n4887# a_8588_n3799# 0.02fF
C4336 a_860_n12503# a_n688_n12503# 0.01fF
C4337 a_2148_n3799# a_2085_n2685# 0.00fF
C4338 a_2148_n5975# sky130_fd_sc_hd__clkinv_4_4/A 0.11fF
C4339 a_600_n12503# a_n428_n12503# 0.02fF
C4340 a_n688_n12503# VDD 0.48fF
C4341 a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.01fF
C4342 sky130_fd_sc_hd__nand2_4_3/Y a_8162_n9213# 0.07fF
C4343 a_501_n1909# a_690_n1597# 0.02fF
C4344 a_600_n2167# a_434_n1597# 0.04fF
C4345 a_9876_n3255# a_9517_n2997# 0.05fF
C4346 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n13021# 0.35fF
C4347 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C4348 a_2148_n3255# a_2085_n1597# 0.00fF
C4349 a_7130_n13021# a_8525_n13021# 0.01fF
C4350 a_7237_n13021# a_8418_n13021# 0.01fF
C4351 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X a_4661_n13021# 0.00fF
C4352 a_4365_n9525# a_5653_n9525# 0.01fF
C4353 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_8418_n14109# 0.00fF
C4354 a_10904_n10871# a_11164_n10871# 0.23fF
C4355 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C4356 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_3436_n11415# 0.01fF
C4357 a_6101_n7254# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.03fF
C4358 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4359 a_4365_n8437# a_4298_n9213# 0.01fF
C4360 a_860_n11415# a_797_n10301# 0.00fF
C4361 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C4362 a_6874_n509# a_8162_n509# 0.01fF
C4363 a_7040_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C4364 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C4365 a_9450_n14109# a_9517_n13413# 0.01fF
C4366 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.01fF
C4367 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/B 0.02fF
C4368 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8588_n9783# 0.01fF
C4369 a_8588_n3255# a_9517_n2997# 0.02fF
C4370 a_3176_n3799# a_3266_n5405# 0.00fF
C4371 a_690_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.05fF
C4372 a_5842_n5405# a_7237_n5405# 0.01fF
C4373 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_10805_n1909# 0.01fF
C4374 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4375 a_1722_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C4376 a_1978_n11933# a_2085_n11933# 0.55fF
C4377 a_9876_n4887# a_9706_n4317# 0.04fF
C4378 a_9616_n4887# a_9813_n4317# 0.02fF
C4379 a_8229_n4709# sky130_fd_sc_hd__clkinv_4_3/A 0.07fF
C4380 a_n1738_n6671# VDD 0.38fF
C4381 a_3077_n5797# a_3010_n5405# 0.01fF
C4382 a_9813_n8125# sky130_fd_sc_hd__nand2_4_3/B 0.13fF
C4383 a_3176_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.03fF
C4384 sky130_fd_sc_hd__nand2_4_2/B VDD 1.22fF
C4385 p2_b VDD 4.27fF
C4386 a_10904_n11415# a_10805_n9525# 0.00fF
C4387 a_10805_n11237# a_10904_n9783# 0.00fF
C4388 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_9616_n9783# 0.01fF
C4389 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C4390 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6665_n7459# 0.01fF
C4391 a_4554_n1597# VDD 0.45fF
C4392 a_7237_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.05fF
C4393 a_5586_n4317# a_5752_n3255# 0.00fF
C4394 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_5842_n9213# 0.03fF
C4395 a_9706_n1597# VDD 0.43fF
C4396 a_4554_n4317# VDD 0.47fF
C4397 a_10904_n3255# a_11164_n3255# 0.23fF
C4398 a_5586_n10301# a_5949_n10301# 0.05fF
C4399 a_5586_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C4400 a_7130_n9213# a_5586_n9213# 0.01fF
C4401 a_6874_n9213# a_5842_n9213# 0.02fF
C4402 a_4464_n3799# a_4554_n2685# 0.01fF
C4403 a_5949_n11933# a_6874_n11933# 0.02fF
C4404 a_5842_n11933# a_7130_n11933# 0.01fF
C4405 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VDD 0.83fF
C4406 a_13765_n2141# a_13765_n2685# 0.31fF
C4407 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.03fF
C4408 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y 0.53fF
C4409 a_8525_n8125# a_9706_n8125# 0.01fF
C4410 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_501_n2997# 0.01fF
C4411 a_1888_n12503# a_501_n12325# 0.01fF
C4412 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkinv_4_7/A 0.62fF
C4413 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkinv_4_4/A 0.85fF
C4414 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_9450_n11933# 0.01fF
C4415 a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C4416 a_501_n821# a_434_n2685# 0.00fF
C4417 a_434_n4317# a_501_n3621# 0.01fF
C4418 a_434_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C4419 a_9616_n10871# a_9450_n9213# 0.00fF
C4420 a_9517_n10613# a_9706_n9213# 0.00fF
C4421 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_501_n9525# 0.01fF
C4422 a_1789_n10613# a_1888_n9783# 0.00fF
C4423 a_11164_n13591# a_11101_n13021# 0.01fF
C4424 a_1888_n10871# a_1789_n9525# 0.00fF
C4425 a_10904_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.05fF
C4426 sky130_fd_sc_hd__nand2_4_3/Y a_9706_n9213# 0.08fF
C4427 a_3077_n13413# a_3010_n11933# 0.00fF
C4428 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_6012_n13591# 0.01fF
C4429 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C4430 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_9706_n13021# 0.00fF
C4431 a_8418_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.05fF
C4432 a_600_n4887# VDD 0.44fF
C4433 a_7237_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C4434 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X Ad_b 0.02fF
C4435 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C4436 a_434_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.03fF
C4437 a_690_n4317# a_797_n4317# 0.55fF
C4438 a_1789_n5797# a_1722_n5405# 0.01fF
C4439 a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C4440 a_8162_n509# a_8418_n509# 0.19fF
C4441 a_5653_n12325# a_7040_n12503# 0.01fF
C4442 a_5752_n12503# a_6941_n12325# 0.01fF
C4443 a_5842_n5405# a_5949_n4317# 0.00fF
C4444 a_4365_n4709# a_4724_n4887# 0.05fF
C4445 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.04fF
C4446 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.06fF
C4447 a_9876_n12503# VDD 0.74fF
C4448 a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.00fF
C4449 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_4298_n5405# 0.00fF
C4450 a_797_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.01fF
C4451 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_2085_n2685# 0.02fF
C4452 a_5752_n11415# VDD 0.44fF
C4453 Bd_b sky130_fd_sc_hd__clkinv_1_5/A 1.60fF
C4454 a_10904_n8695# a_10805_n9525# 0.00fF
C4455 a_1978_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C4456 a_10805_n8437# a_10904_n9783# 0.00fF
C4457 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3266_n11933# 0.03fF
C4458 a_2085_n11933# a_3373_n11933# 0.01fF
C4459 a_9616_n4887# sky130_fd_sc_hd__clkinv_4_3/A 0.07fF
C4460 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.01fF
C4461 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_6012_n12503# 0.01fF
C4462 a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C4463 a_600_n2167# a_n428_n2167# 0.02fF
C4464 a_860_n2167# a_n688_n2167# 0.01fF
C4465 a_5586_n4317# a_4298_n4317# 0.01fF
C4466 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_2148_n4887# 0.03fF
C4467 a_2085_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C4468 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C4469 a_3077_n3621# a_3010_n4317# 0.01fF
C4470 a_8328_n8695# a_8328_n9783# 0.01fF
C4471 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkinv_4_8/A 0.44fF
C4472 a_5949_n1597# VDD 0.35fF
C4473 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.01fF
C4474 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.02fF
C4475 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.09fF
C4476 a_5949_n4317# a_6012_n5975# 0.00fF
C4477 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C4478 a_5842_n10301# a_7237_n10301# 0.01fF
C4479 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n10301# 0.35fF
C4480 a_5949_n10301# a_7130_n10301# 0.01fF
C4481 a_6874_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C4482 a_7130_n11933# a_7237_n11933# 0.55fF
C4483 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_8162_n11933# 0.00fF
C4484 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_7237_n10301# 0.00fF
C4485 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C4486 a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C4487 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_5586_n2685# 0.01fF
C4488 a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C4489 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_9450_n10301# 0.03fF
C4490 clk sky130_fd_sc_hd__dfxbp_1_1/D 0.08fF
C4491 a_9813_n5405# a_9616_n5975# 0.02fF
C4492 a_7237_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C4493 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_7300_n5975# 0.03fF
C4494 a_10738_n13789# a_10738_n13021# 0.01fF
C4495 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.06fF
C4496 a_10738_n11933# a_9450_n11933# 0.01fF
C4497 a_797_n9213# a_860_n9783# 0.01fF
C4498 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_9876_n3799# 0.00fF
C4499 a_10904_n13591# a_10904_n12503# 0.01fF
C4500 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11164_n3255# 0.01fF
C4501 a_7237_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C4502 a_7300_n13591# VDD 0.76fF
C4503 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C4504 a_9517_n1909# a_9517_n2997# 0.02fF
C4505 a_6941_n9525# a_7040_n10871# 0.00fF
C4506 a_7040_n9783# a_6941_n10613# 0.00fF
C4507 a_3176_n3255# a_3176_n4887# 0.00fF
C4508 a_4661_n11933# a_5949_n11933# 0.01fF
C4509 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5842_n11933# 0.03fF
C4510 a_4554_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C4511 a_n428_n9783# a_860_n9783# 0.01fF
C4512 a_n688_n4887# a_600_n4887# 0.01fF
C4513 a_5752_n8695# a_5842_n9213# 0.01fF
C4514 a_n688_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C4515 sky130_fd_sc_hd__dfxbp_1_0/Q a_6101_n7254# 0.31fF
C4516 a_8525_n509# a_9450_n509# 0.02fF
C4517 sky130_fd_sc_hd__nand2_4_1/B Ad_b 0.06fF
C4518 a_10738_n6173# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C4519 a_4623_n7349# a_6373_n7349# 0.00fF
C4520 a_6941_n12325# a_7300_n12503# 0.05fF
C4521 a_4464_n4887# a_6012_n4887# 0.01fF
C4522 a_4724_n4887# a_5752_n4887# 0.02fF
C4523 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X a_5653_n4709# 0.18fF
C4524 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_2148_n1079# 0.03fF
C4525 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.00fF
C4526 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VDD 0.63fF
C4527 a_4724_n3799# a_4661_n5405# 0.00fF
C4528 a_9706_n1597# a_9876_n1079# 0.04fF
C4529 a_9813_n1597# a_9616_n1079# 0.02fF
C4530 a_13765_n12477# p1d 2.55fF
C4531 a_3373_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.12fF
C4532 a_7300_n11415# VDD 0.77fF
C4533 a_860_n3799# VDD 0.78fF
C4534 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Ad_b 0.03fF
C4535 a_4464_n5975# a_4554_n5405# 0.01fF
C4536 a_4623_n7349# VDD 0.37fF
C4537 Bd_b a_13765_n4317# 0.14fF
C4538 a_4464_n10871# a_4661_n9213# 0.00fF
C4539 a_4724_n10871# a_4554_n9213# 0.00fF
C4540 a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C4541 a_501_n8437# a_434_n9213# 0.01fF
C4542 a_3176_n11415# a_3010_n11933# 0.04fF
C4543 a_3077_n11237# a_3266_n11933# 0.02fF
C4544 sky130_fd_sc_hd__clkinv_4_7/A a_860_n13591# 0.09fF
C4545 a_8162_n10301# a_8328_n9783# 0.04fF
C4546 a_8229_n4709# a_8328_n5975# 0.00fF
C4547 a_7237_n4317# a_7040_n3255# 0.00fF
C4548 a_8328_n4887# a_8229_n5797# 0.00fF
C4549 a_7130_n4317# a_7300_n3255# 0.00fF
C4550 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y 1.20fF
C4551 a_11164_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.11fF
C4552 a_3077_n821# a_3010_n2685# 0.00fF
C4553 a_10904_n2167# a_10805_n2997# 0.00fF
C4554 a_10805_n1909# a_10904_n3255# 0.00fF
C4555 a_7130_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.05fF
C4556 a_8229_n13413# a_9517_n13413# 0.01fF
C4557 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_9450_n4317# 0.00fF
C4558 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_4_3/A 0.07fF
C4559 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C4560 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8418_n11933# 0.03fF
C4561 a_7130_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C4562 a_8588_n10871# a_7040_n10871# 0.01fF
C4563 a_7237_n11933# a_8525_n11933# 0.01fF
C4564 a_8162_n9213# a_9450_n9213# 0.01fF
C4565 a_6874_n14109# a_6941_n12325# 0.00fF
C4566 a_9876_n10871# a_9813_n10301# 0.01fF
C4567 sky130_fd_sc_hd__clkinv_4_4/A a_9616_n5975# 0.07fF
C4568 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__dfxbp_1_0/Q 0.02fF
C4569 a_5752_n3799# a_5653_n2997# 0.01fF
C4570 a_2148_n4887# a_1978_n4317# 0.04fF
C4571 a_1888_n4887# a_2085_n4317# 0.02fF
C4572 a_13765_n13565# a_13765_n12477# 0.07fF
C4573 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/A 0.46fF
C4574 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VDD 0.82fF
C4575 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_5653_n5797# 0.01fF
C4576 a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.02fF
C4577 a_10904_n8695# a_10994_n9213# 0.01fF
C4578 a_4464_n13591# a_4554_n11933# 0.00fF
C4579 a_7130_n10301# a_8418_n10301# 0.01fF
C4580 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkinv_1_0/Y 0.00fF
C4581 Ad_b sky130_fd_sc_hd__clkinv_1_3/A 0.25fF
C4582 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X 0.00fF
C4583 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_2148_n2167# 0.03fF
C4584 a_4365_n12325# a_5752_n12503# 0.01fF
C4585 a_4464_n12503# a_5653_n12325# 0.01fF
C4586 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_8525_n9213# 0.01fF
C4587 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_7130_n5405# 0.03fF
C4588 a_5949_n5405# a_7237_n5405# 0.01fF
C4589 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.03fF
C4590 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C4591 a_1888_n1079# a_2148_n1079# 0.28fF
C4592 a_7130_n2685# a_5949_n2685# 0.01fF
C4593 a_7237_n2685# a_5842_n2685# 0.01fF
C4594 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.35fF
C4595 a_7040_n12503# a_8588_n12503# 0.01fF
C4596 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X a_7040_n4887# 0.01fF
C4597 a_5752_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.03fF
C4598 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Bd_b 0.02fF
C4599 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_8229_n12325# 0.18fF
C4600 a_7300_n12503# a_8328_n12503# 0.02fF
C4601 a_7130_n6493# a_6941_n5797# 0.02fF
C4602 a_6874_n6493# a_7040_n5975# 0.04fF
C4603 a_1789_n8437# VDD 0.36fF
C4604 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.02fF
C4605 a_9876_n2167# VDD 0.74fF
C4606 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VDD 0.83fF
C4607 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6012_n3799# 0.01fF
C4608 a_5949_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C4609 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_9876_n3799# 0.01fF
C4610 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C4611 a_9517_n4709# a_9517_n2997# 0.00fF
C4612 a_9517_n10613# a_9517_n12325# 0.00fF
C4613 a_7237_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C4614 a_1978_n10301# a_1789_n8437# 0.00fF
C4615 a_1722_n10301# a_1888_n8695# 0.00fF
C4616 a_5752_n10871# a_5949_n11933# 0.00fF
C4617 a_6012_n10871# a_5842_n11933# 0.00fF
C4618 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_4661_n9213# 0.01fF
C4619 a_9813_n1597# a_9813_n509# 0.02fF
C4620 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.03fF
C4621 a_860_n11415# a_797_n11933# 0.01fF
C4622 a_10904_n13591# a_9876_n13591# 0.02fF
C4623 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_434_n2685# 0.45fF
C4624 a_9876_n8695# a_9876_n9783# 0.02fF
C4625 a_8229_n11237# a_9517_n11237# 0.01fF
C4626 a_4464_n3799# a_4554_n4317# 0.02fF
C4627 a_11164_n13591# a_9616_n13591# 0.01fF
C4628 a_8229_n3621# a_9616_n3799# 0.01fF
C4629 a_n688_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.04fF
C4630 a_8328_n3799# a_9517_n3621# 0.01fF
C4631 a_6665_n7459# p2 0.08fF
C4632 a_6865_n7304# a_6794_n7203# 0.47fF
C4633 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C4634 a_9876_n5975# a_9813_n4317# 0.00fF
C4635 a_9517_n13413# a_9616_n13591# 0.48fF
C4636 a_4365_n5797# a_4298_n4317# 0.00fF
C4637 a_9450_n9213# a_9706_n9213# 0.19fF
C4638 a_9616_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C4639 a_8525_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.12fF
C4640 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8328_n10871# 0.03fF
C4641 a_9616_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C4642 a_5752_n9783# VDD 0.46fF
C4643 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.00fF
C4644 sky130_fd_sc_hd__clkinv_4_4/A a_11164_n5975# 0.10fF
C4645 a_7130_n509# a_7040_n1079# 0.02fF
C4646 sky130_fd_sc_hd__clkinv_1_0/A a_10805_n821# 0.05fF
C4647 a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C4648 a_4464_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C4649 p2d p2_b 0.53fF
C4650 a_8418_n8125# a_8588_n9783# 0.00fF
C4651 a_8525_n8125# a_8328_n9783# 0.00fF
C4652 a_4724_n5975# a_6012_n5975# 0.01fF
C4653 a_8328_n4887# VDD 0.44fF
C4654 a_4365_n12325# a_4298_n13021# 0.01fF
C4655 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.03fF
C4656 a_5842_n13021# a_5653_n12325# 0.02fF
C4657 a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C4658 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_5586_n11933# 0.00fF
C4659 a_5949_n4317# a_5949_n5405# 0.02fF
C4660 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_8525_n509# 0.00fF
C4661 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.00fF
C4662 a_4464_n9783# a_4464_n8695# 0.01fF
C4663 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.04fF
C4664 a_9517_n8437# a_9706_n10301# 0.00fF
C4665 a_9616_n8695# a_9450_n10301# 0.00fF
C4666 a_7237_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.12fF
C4667 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.03fF
C4668 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_2148_n9783# 0.00fF
C4669 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C4670 a_2148_n1079# a_3436_n1079# 0.01fF
C4671 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_3176_n1079# 0.05fF
C4672 a_1888_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.00fF
C4673 a_8418_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C4674 a_10904_n4887# a_10805_n2997# 0.00fF
C4675 a_3266_n1597# a_3373_n2685# 0.00fF
C4676 a_10805_n4709# a_10904_n3255# 0.00fF
C4677 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__clkinv_1_5/A 0.97fF
C4678 a_8328_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C4679 a_3010_n5405# a_4298_n5405# 0.01fF
C4680 a_3077_n2997# a_3010_n1597# 0.00fF
C4681 a_n2037_n7037# sky130_fd_sc_hd__clkinv_1_5/A 0.01fF
C4682 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C4683 a_3176_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.03fF
C4684 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C4685 a_6006_n7607# a_7212_n7203# 0.01fF
C4686 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_6012_n3255# 0.01fF
C4687 a_13765_n2141# VDD 2.19fF
C4688 a_10904_n13591# a_10738_n13789# 0.03fF
C4689 a_1888_n9783# a_3077_n9525# 0.01fF
C4690 a_1789_n9525# a_3176_n9783# 0.01fF
C4691 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.02fF
C4692 a_4724_n11415# a_4554_n11933# 0.04fF
C4693 a_2622_n6493# VDD 0.50fF
C4694 a_4464_n11415# a_4661_n11933# 0.02fF
C4695 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n9213# 0.01fF
C4696 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8588_n3255# 0.01fF
C4697 a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C4698 a_7040_n10871# a_7130_n9213# 0.00fF
C4699 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_1978_n2685# 0.00fF
C4700 a_8525_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C4701 a_9450_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C4702 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6865_n7304# 0.01fF
C4703 a_4464_n1079# a_4554_n2685# 0.00fF
C4704 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkinv_4_4/A 0.04fF
C4705 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.06fF
C4706 a_7300_n9783# VDD 0.78fF
C4707 a_600_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C4708 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.06fF
C4709 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.35fF
C4710 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.02fF
C4711 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8229_n821# 0.01fF
C4712 a_8162_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.03fF
C4713 a_1978_n1597# a_1789_n2997# 0.00fF
C4714 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C4715 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_4661_n11933# 0.00fF
C4716 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_1789_n9525# 0.01fF
C4717 a_8229_n4709# a_8418_n5405# 0.02fF
C4718 a_8328_n4887# a_8162_n5405# 0.04fF
C4719 sky130_fd_sc_hd__nand2_4_1/A VDD 13.21fF
C4720 a_n2602_n7037# a_n2163_n6671# 0.53fF
C4721 a_9876_n4887# VDD 0.74fF
C4722 a_3010_n5405# a_1722_n5405# 0.01fF
C4723 a_2729_n6493# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C4724 sky130_fd_sc_hd__dfxbp_1_1/D a_n1995_n6925# 0.14fF
C4725 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C4726 a_8418_n2685# a_8418_n1597# 0.01fF
C4727 a_3077_n12325# a_4464_n12503# 0.01fF
C4728 a_3176_n12503# a_4365_n12325# 0.01fF
C4729 a_4464_n10871# a_4365_n11237# 0.01fF
C4730 a_9876_n2167# a_9876_n1079# 0.02fF
C4731 a_7237_n2685# a_7300_n3255# 0.01fF
C4732 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.02fF
C4733 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.29fF
C4734 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_9813_n9213# 0.01fF
C4735 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.03fF
C4736 a_1888_n13591# a_1978_n13021# 0.01fF
C4737 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.02fF
C4738 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.02fF
C4739 a_2366_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.00fF
C4740 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C4741 a_5842_n2685# a_5653_n821# 0.00fF
C4742 a_5586_n2685# a_5752_n1079# 0.00fF
C4743 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_2148_n4887# 0.03fF
C4744 a_4298_n5405# a_4554_n5405# 0.19fF
C4745 a_8525_n6493# a_8328_n5975# 0.02fF
C4746 a_8418_n6493# a_8588_n5975# 0.04fF
C4747 sky130_fd_sc_hd__clkinv_1_0/Y VDD 1.17fF
C4748 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.00fF
C4749 a_860_n2167# VDD 0.78fF
C4750 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_4724_n3255# 0.03fF
C4751 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C4752 a_3436_n3799# a_1888_n3799# 0.01fF
C4753 a_7130_n6493# a_6658_n7363# 0.00fF
C4754 a_6874_n6493# a_6665_n7459# 0.00fF
C4755 a_11101_n1597# sky130_fd_sc_hd__clkinv_4_1/Y 0.01fF
C4756 a_3077_n9525# a_3436_n9783# 0.05fF
C4757 a_4464_n10871# a_4724_n10871# 0.28fF
C4758 a_8525_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.12fF
C4759 a_6874_n509# a_6874_n1597# 0.02fF
C4760 a_9450_n509# a_9450_n1597# 0.02fF
C4761 a_10904_n10871# a_10904_n12503# 0.00fF
C4762 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C4763 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_7237_n11933# 0.00fF
C4764 a_7237_n6493# VDD 0.34fF
C4765 a_1888_n12503# a_1789_n10613# 0.00fF
C4766 a_1789_n12325# a_1888_n10871# 0.00fF
C4767 a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C4768 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_8162_n9213# 0.00fF
C4769 a_5653_n3621# a_5653_n4709# 0.02fF
C4770 a_434_n5405# a_1722_n5405# 0.01fF
C4771 a_2729_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.12fF
C4772 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_5586_n2685# 0.00fF
C4773 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_5752_n1079# 0.01fF
C4774 a_7040_n2167# a_7040_n3799# 0.00fF
C4775 a_690_n10301# a_690_n9213# 0.01fF
C4776 a_7130_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.23fF
C4777 a_8525_n509# a_8588_n1079# 0.01fF
C4778 a_3077_n4709# a_4724_n4887# 0.00fF
C4779 a_3176_n4887# a_4464_n4887# 0.01fF
C4780 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.12fF
C4781 a_10994_n9213# a_10805_n9525# 0.02fF
C4782 a_10738_n9213# a_10904_n9783# 0.04fF
C4783 a_7130_n13021# a_7300_n12503# 0.04fF
C4784 a_2366_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C4785 clk sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C4786 a_7237_n13021# a_7040_n12503# 0.02fF
C4787 a_3373_n1597# a_1722_n1597# 0.00fF
C4788 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.04fF
C4789 clk a_n1570_n6769# 0.01fF
C4790 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C4791 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkinv_1_5/A 0.03fF
C4792 a_8229_n10613# a_8162_n10301# 0.01fF
C4793 a_9450_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C4794 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n1597# 0.01fF
C4795 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VDD 2.08fF
C4796 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.02fF
C4797 a_6941_n13413# a_7130_n11933# 0.00fF
C4798 a_7040_n13591# a_6874_n11933# 0.00fF
C4799 a_1789_n821# a_1978_n2685# 0.00fF
C4800 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_3010_n13021# 0.03fF
C4801 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.02fF
C4802 a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C4803 a_4661_n5405# a_5586_n5405# 0.02fF
C4804 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.06fF
C4805 a_4554_n5405# a_5842_n5405# 0.01fF
C4806 a_1888_n13591# VDD 0.45fF
C4807 a_8328_n2167# a_8418_n1597# 0.02fF
C4808 a_9876_n2167# sky130_fd_sc_hd__nand2_4_0/B 0.00fF
C4809 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_9813_n509# 0.00fF
C4810 sky130_fd_sc_hd__nand2_4_3/Y p2 0.09fF
C4811 a_5949_n9213# VDD 0.35fF
C4812 a_5752_n1079# a_6012_n1079# 0.28fF
C4813 a_5653_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.02fF
C4814 a_1789_n5797# a_1888_n5975# 0.49fF
C4815 a_501_n12325# a_434_n13021# 0.01fF
C4816 a_9616_n11415# a_11164_n11415# 0.01fF
C4817 a_9876_n11415# a_10904_n11415# 0.02fF
C4818 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_10805_n11237# 0.17fF
C4819 a_4724_n10871# a_6012_n10871# 0.01fF
C4820 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_5752_n10871# 0.05fF
C4821 a_4464_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C4822 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C4823 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_4724_n10871# 0.01fF
C4824 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.02fF
C4825 a_10994_n11933# VDD 0.44fF
C4826 a_6941_n11237# a_7130_n11933# 0.02fF
C4827 a_7040_n11415# a_6874_n11933# 0.04fF
C4828 a_8162_n14109# a_9450_n14109# 0.01fF
C4829 sky130_fd_sc_hd__nand2_4_2/A a_9450_n14109# 0.03fF
C4830 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VDD 0.98fF
C4831 a_4724_n3255# a_4724_n2167# 0.02fF
C4832 a_9706_n1597# a_10738_n1597# 0.02fF
C4833 a_797_n9213# VDD 0.36fF
C4834 a_9450_n1597# a_10994_n1597# 0.01fF
C4835 a_1722_n5405# a_1978_n5405# 0.19fF
C4836 a_4365_n10613# VDD 0.35fF
C4837 a_2366_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C4838 a_2148_n11415# a_1978_n13021# 0.00fF
C4839 a_1888_n11415# a_2085_n13021# 0.00fF
C4840 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.29fF
C4841 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5653_n5797# 0.01fF
C4842 a_5586_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.03fF
C4843 a_10738_n6173# a_10994_n5405# 0.01fF
C4844 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C4845 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.00fF
C4846 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_6012_n1079# 0.03fF
C4847 a_3436_n8695# VDD 0.80fF
C4848 a_8525_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C4849 a_1722_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C4850 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n9213# 0.01fF
C4851 a_10805_n3621# a_10994_n2685# 0.00fF
C4852 a_10904_n3799# a_10738_n2685# 0.00fF
C4853 a_8328_n4887# a_8418_n4317# 0.01fF
C4854 a_8328_n8695# VDD 0.47fF
C4855 a_2366_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C4856 a_3077_n10613# a_3266_n10301# 0.02fF
C4857 a_3176_n10871# a_3010_n10301# 0.04fF
C4858 a_10805_n3621# a_10738_n4317# 0.01fF
C4859 a_8229_n1909# a_6941_n1909# 0.01fF
C4860 a_n428_n9783# VDD 0.83fF
C4861 a_9876_n5975# a_8328_n5975# 0.01fF
C4862 a_9616_n5975# a_8588_n5975# 0.02fF
C4863 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.02fF
C4864 a_9876_n4887# a_9706_n5405# 0.04fF
C4865 a_9450_n13021# VDD 0.75fF
C4866 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_10904_n9783# 0.02fF
C4867 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3077_n8437# 0.00fF
C4868 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3010_n1597# 0.03fF
C4869 a_4298_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.00fF
C4870 a_3373_n1597# a_3266_n1597# 0.55fF
C4871 a_9813_n2685# a_9813_n1597# 0.02fF
C4872 a_7130_n9213# a_6665_n7459# 0.00fF
C4873 a_6874_n9213# a_6865_n7304# 0.00fF
C4874 a_7237_n9213# a_6658_n7363# 0.00fF
C4875 a_501_n10613# a_690_n10301# 0.02fF
C4876 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_4365_n8437# 0.01fF
C4877 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.01fF
C4878 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.08fF
C4879 a_3436_n13591# a_3373_n13021# 0.01fF
C4880 a_6941_n9525# sky130_fd_sc_hd__nand2_4_3/Y 0.08fF
C4881 a_11101_n9213# sky130_fd_sc_hd__clkinv_1_3/A 0.01fF
C4882 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X a_5752_n5975# 0.05fF
C4883 a_2148_n12503# a_2148_n13591# 0.02fF
C4884 a_3436_n13591# VDD 0.78fF
C4885 a_10904_n3799# a_9616_n3799# 0.01fF
C4886 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_9450_n1597# 0.03fF
C4887 a_11164_n3799# a_9517_n3621# 0.00fF
C4888 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.04fF
C4889 a_1888_n2167# a_3077_n1909# 0.01fF
C4890 a_1789_n1909# a_3176_n2167# 0.01fF
C4891 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VDD 0.88fF
C4892 a_2085_n9213# a_3010_n9213# 0.02fF
C4893 sky130_fd_sc_hd__nand2_4_0/Y a_6941_n1909# 0.08fF
C4894 a_5752_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.00fF
C4895 a_1789_n5797# a_3436_n5975# 0.00fF
C4896 a_6012_n1079# a_7300_n1079# 0.01fF
C4897 a_1888_n5975# a_3176_n5975# 0.01fF
C4898 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X a_7040_n1079# 0.05fF
C4899 sky130_fd_sc_hd__nand2_4_2/A a_11101_n13021# 0.00fF
C4900 a_2148_n5975# a_3077_n5797# 0.02fF
C4901 a_9876_n12503# a_9706_n11933# 0.04fF
C4902 a_10904_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.02fF
C4903 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.29fF
C4904 a_4554_n1597# a_4464_n1079# 0.01fF
C4905 a_3373_n2685# VDD 0.35fF
C4906 a_9450_n14109# a_9706_n14109# 0.19fF
C4907 a_1888_n13591# a_501_n13413# 0.01fF
C4908 a_1789_n13413# a_600_n13591# 0.01fF
C4909 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.70fF
C4910 a_10738_n9213# a_11101_n9213# 0.05fF
C4911 a_8418_n6493# a_8525_n5405# 0.00fF
C4912 a_8525_n6493# a_8418_n5405# 0.00fF
C4913 a_3176_n2167# a_4464_n2167# 0.01fF
C4914 a_3077_n1909# a_4724_n2167# 0.00fF
C4915 a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.01fF
C4916 a_8162_n10301# VDD 0.76fF
C4917 a_8588_n10871# a_9517_n10613# 0.02fF
C4918 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD 0.85fF
C4919 a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C4920 a_5752_n9783# a_5586_n9213# 0.04fF
C4921 a_5653_n9525# a_5842_n9213# 0.02fF
C4922 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__nand2_4_0/Y 0.44fF
C4923 a_9876_n8695# VDD 0.74fF
C4924 a_2148_n11415# VDD 0.77fF
C4925 a_6874_n8125# a_6658_n7363# 0.01fF
C4926 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_5653_n1909# 0.18fF
C4927 a_4724_n2167# a_5752_n2167# 0.02fF
C4928 a_4464_n2167# a_6012_n2167# 0.01fF
C4929 a_3373_n10301# a_3436_n8695# 0.00fF
C4930 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_3266_n1597# 0.01fF
C4931 Bd_b a_5052_n7283# 0.20fF
C4932 a_6941_n2997# a_7040_n3255# 0.49fF
C4933 a_1888_n11415# a_2085_n10301# 0.00fF
C4934 a_8525_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C4935 a_2148_n11415# a_1978_n10301# 0.00fF
C4936 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8588_n12503# 0.03fF
C4937 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C4938 a_5842_n1597# a_5653_n821# 0.02fF
C4939 a_5586_n1597# a_5752_n1079# 0.04fF
C4940 a_8162_n1597# a_8328_n1079# 0.04fF
C4941 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VDD 0.87fF
C4942 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.08fF
C4943 a_8328_n13591# a_8525_n11933# 0.00fF
C4944 a_8588_n13591# a_8418_n11933# 0.00fF
C4945 a_8418_n1597# a_8229_n821# 0.02fF
C4946 a_9813_n13021# a_11101_n13021# 0.01fF
C4947 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9876_n11415# 0.03fF
C4948 a_9813_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C4949 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_10994_n13021# 0.03fF
C4950 A_b a_13765_n4317# 0.06fF
C4951 a_13765_n5405# Ad_b 0.16fF
C4952 a_7130_n8125# VDD 0.44fF
C4953 a_600_n10871# a_2148_n10871# 0.01fF
C4954 a_860_n10871# a_1888_n10871# 0.02fF
C4955 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_1789_n10613# 0.18fF
C4956 a_501_n2997# VDD 0.36fF
C4957 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD 0.78fF
C4958 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.29fF
C4959 a_9616_n2167# a_9450_n509# 0.00fF
C4960 a_690_n4317# a_690_n5405# 0.01fF
C4961 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.08fF
C4962 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VDD 0.84fF
C4963 a_9517_n12325# a_9450_n14109# 0.00fF
C4964 a_9450_n8125# a_9813_n8125# 0.05fF
C4965 sky130_fd_sc_hd__nand2_4_2/B a_10738_n13021# 0.01fF
C4966 a_3077_n1909# a_3436_n2167# 0.05fF
C4967 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.01fF
C4968 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_4298_n9213# 0.00fF
C4969 a_3266_n9213# a_3373_n9213# 0.55fF
C4970 a_3010_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.03fF
C4971 a_3176_n5975# a_3436_n5975# 0.28fF
C4972 a_7300_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.29fF
C4973 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkinv_1_3/Y 0.02fF
C4974 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_4365_n5797# 0.01fF
C4975 a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.02fF
C4976 a_5752_n11415# a_5653_n10613# 0.01fF
C4977 a_5653_n11237# a_5752_n10871# 0.01fF
C4978 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.04fF
C4979 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_4_3/A 0.30fF
C4980 a_5586_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.03fF
C4981 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C4982 a_n1570_n6769# sky130_fd_sc_hd__clkinv_1_5/A 0.25fF
C4983 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VDD 0.89fF
C4984 a_8328_n11415# a_8525_n11933# 0.02fF
C4985 a_8588_n11415# a_8418_n11933# 0.04fF
C4986 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6658_n7363# 0.01fF
C4987 a_7300_n4887# a_7300_n3799# 0.02fF
C4988 sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# 0.58fF
C4989 a_11101_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.12fF
C4990 a_600_n11415# a_860_n11415# 0.28fF
C4991 a_4365_n2997# VDD 0.35fF
C4992 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_5653_n1909# 0.01fF
C4993 a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.01fF
C4994 a_5842_n13021# a_7237_n13021# 0.01fF
C4995 a_5949_n13021# a_7130_n13021# 0.01fF
C4996 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_3373_n13021# 0.00fF
C4997 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n13021# 0.35fF
C4998 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C4999 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A VDD 0.84fF
C5000 a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.02fF
C5001 a_9616_n10871# a_9876_n10871# 0.28fF
C5002 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C5003 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_2148_n11415# 0.01fF
C5004 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_10805_n10613# 0.01fF
C5005 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.08fF
C5006 a_3077_n8437# a_3010_n9213# 0.01fF
C5007 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VDD 0.84fF
C5008 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C5009 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.00fF
C5010 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_7040_n2167# 0.01fF
C5011 a_5752_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.03fF
C5012 a_8162_n14109# a_8229_n13413# 0.01fF
C5013 a_7040_n3255# a_8328_n3255# 0.01fF
C5014 a_7300_n3255# a_8229_n2997# 0.02fF
C5015 a_6941_n2997# a_8588_n3255# 0.00fF
C5016 a_4554_n5405# a_5949_n5405# 0.01fF
C5017 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.08fF
C5018 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C5019 a_11101_n13021# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C5020 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C5021 a_10904_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.02fF
C5022 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.06fF
C5023 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.00fF
C5024 a_8525_n8125# VDD 0.35fF
C5025 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_4724_n4887# 0.00fF
C5026 a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C5027 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_3176_n10871# 0.01fF
C5028 a_1888_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.03fF
C5029 a_n1995_n6925# a_n1570_n6769# 0.06fF
C5030 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_9450_n5405# 0.03fF
C5031 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C5032 a_9876_n4887# a_9813_n5405# 0.01fF
C5033 a_9616_n11415# a_9517_n9525# 0.00fF
C5034 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_8328_n9783# 0.01fF
C5035 A VDD 4.21fF
C5036 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.04fF
C5037 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__mux2_1_0/X 0.20fF
C5038 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1722_n5405# 0.01fF
C5039 a_3010_n10301# a_3077_n9525# 0.01fF
C5040 a_3266_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C5041 a_3373_n9213# a_4661_n9213# 0.01fF
C5042 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4554_n9213# 0.03fF
C5043 a_7130_n1597# VDD 0.44fF
C5044 a_3436_n5975# a_4724_n5975# 0.01fF
C5045 a_9616_n3255# a_9876_n3255# 0.28fF
C5046 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10805_n13413# 0.00fF
C5047 a_8328_n11415# a_8525_n10301# 0.00fF
C5048 a_1978_n4317# VDD 0.47fF
C5049 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_4464_n5975# 0.05fF
C5050 a_3176_n3799# a_3266_n2685# 0.01fF
C5051 a_4298_n10301# a_4661_n10301# 0.05fF
C5052 a_1789_n4709# a_3176_n4887# 0.01fF
C5053 a_1888_n4887# a_3077_n4709# 0.01fF
C5054 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.00fF
C5055 sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# 0.53fF
C5056 sky130_fd_sc_hd__nand2_1_4/B Ad_b 0.02fF
C5057 a_600_n10871# a_501_n9525# 0.00fF
C5058 a_2148_n2167# a_2085_n2685# 0.01fF
C5059 sky130_fd_sc_hd__nand2_4_3/Y a_7130_n9213# 0.23fF
C5060 a_7130_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.05fF
C5061 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_8418_n13021# 0.00fF
C5062 a_1789_n13413# a_1722_n11933# 0.00fF
C5063 a_9876_n3255# a_8328_n3255# 0.01fF
C5064 a_9616_n3255# a_8588_n3255# 0.02fF
C5065 a_1722_n9213# a_3266_n9213# 0.01fF
C5066 a_1978_n9213# a_3010_n9213# 0.02fF
C5067 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_9450_n14109# 0.00fF
C5068 a_9876_n10871# a_11164_n10871# 0.01fF
C5069 a_10805_n10613# a_10738_n11933# 0.00fF
C5070 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.03fF
C5071 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_10904_n10871# 0.05fF
C5072 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_9813_n2685# 0.01fF
C5073 a_6941_n8437# a_6794_n7203# 0.00fF
C5074 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C5075 sky130_fd_sc_hd__clkinv_4_3/A a_6941_n4709# 0.08fF
C5076 a_6874_n1597# a_7040_n3255# 0.00fF
C5077 a_6874_n509# a_7130_n509# 0.19fF
C5078 a_10805_n3621# a_11164_n3799# 0.05fF
C5079 a_8229_n9525# a_8162_n9213# 0.01fF
C5080 a_2622_n6493# sky130_fd_sc_hd__clkinv_4_4/A 0.01fF
C5081 a_9706_n1597# a_9517_n2997# 0.00fF
C5082 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_7300_n2167# 0.03fF
C5083 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C5084 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.06fF
C5085 a_501_n8437# a_1789_n8437# 0.01fF
C5086 a_10805_n821# a_10738_n2685# 0.00fF
C5087 a_8162_n6493# a_9450_n6493# 0.01fF
C5088 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.01fF
C5089 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_3373_n10301# 0.00fF
C5090 a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C5091 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X a_9517_n2997# 0.01fF
C5092 a_8229_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C5093 a_8328_n3255# a_8588_n3255# 0.28fF
C5094 a_9517_n12325# a_10805_n12325# 0.01fF
C5095 a_8588_n2167# a_9876_n2167# 0.01fF
C5096 a_5842_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.05fF
C5097 a_8328_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C5098 a_1888_n3799# a_1722_n5405# 0.00fF
C5099 a_1789_n3621# a_1978_n5405# 0.00fF
C5100 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_9616_n2167# 0.05fF
C5101 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_7130_n5405# 0.00fF
C5102 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_10738_n13021# 0.02fF
C5103 a_11164_n12503# a_10994_n13021# 0.04fF
C5104 a_10904_n12503# a_11101_n13021# 0.02fF
C5105 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A 2.39fF
C5106 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.02fF
C5107 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.00fF
C5108 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_3436_n10871# 0.03fF
C5109 a_690_n4317# a_501_n4709# 0.02fF
C5110 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_8588_n9783# 0.03fF
C5111 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.00fF
C5112 a_434_n4317# a_600_n4887# 0.04fF
C5113 a_3373_n1597# VDD 0.35fF
C5114 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C5115 a_4661_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.12fF
C5116 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.09fF
C5117 a_8525_n1597# VDD 0.35fF
C5118 a_10904_n2167# a_11101_n1597# 0.02fF
C5119 a_11164_n2167# a_10994_n1597# 0.04fF
C5120 a_9876_n3255# a_11164_n3255# 0.01fF
C5121 a_5949_n9213# a_5586_n9213# 0.05fF
C5122 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X a_10904_n3255# 0.05fF
C5123 a_3373_n4317# VDD 0.35fF
C5124 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C5125 a_5842_n4317# a_5949_n2685# 0.00fF
C5126 a_5949_n4317# a_5842_n2685# 0.00fF
C5127 a_4661_n10301# a_5842_n10301# 0.01fF
C5128 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5586_n10301# 0.35fF
C5129 a_4554_n10301# a_5949_n10301# 0.01fF
C5130 a_5842_n11933# a_5949_n11933# 0.55fF
C5131 a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C5132 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_4298_n2685# 0.01fF
C5133 a_5653_n2997# a_5586_n4317# 0.00fF
C5134 a_690_n11933# a_501_n10613# 0.00fF
C5135 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6012_n5975# 0.03fF
C5136 a_5949_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.01fF
C5137 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_9706_n8125# 0.00fF
C5138 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkinv_1_0/A 0.02fF
C5139 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.04fF
C5140 a_860_n12503# a_501_n12325# 0.05fF
C5141 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.03fF
C5142 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_n428_n12503# 0.00fF
C5143 a_8588_n10871# a_8525_n11933# 0.00fF
C5144 a_501_n12325# VDD 0.36fF
C5145 sky130_fd_sc_hd__nand2_4_3/Y a_8525_n9213# 0.05fF
C5146 a_5752_n9783# a_5653_n10613# 0.00fF
C5147 a_7237_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C5148 a_5653_n9525# a_5752_n10871# 0.00fF
C5149 a_600_n2167# a_797_n1597# 0.02fF
C5150 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8525_n13021# 0.02fF
C5151 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.02fF
C5152 a_860_n2167# a_690_n1597# 0.04fF
C5153 a_10904_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C5154 a_4464_n9783# a_5752_n9783# 0.01fF
C5155 a_4724_n9783# a_5653_n9525# 0.02fF
C5156 a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.01fF
C5157 a_4365_n9525# a_6012_n9783# 0.00fF
C5158 a_5586_n1597# a_6874_n1597# 0.01fF
C5159 a_8229_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C5160 sky130_fd_sc_hd__nand2_4_2/A a_n860_n13789# 0.01fF
C5161 a_9616_n13591# a_9813_n13021# 0.02fF
C5162 a_4464_n8695# a_4554_n9213# 0.01fF
C5163 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_690_n4317# 0.02fF
C5164 a_6658_n7363# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.02fF
C5165 a_10904_n13591# sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C5166 a_6941_n1909# VDD 0.35fF
C5167 a_6874_n509# a_8525_n509# 0.00fF
C5168 a_7130_n509# a_8418_n509# 0.01fF
C5169 a_7237_n509# a_8162_n509# 0.02fF
C5170 a_434_n2685# VDD 0.76fF
C5171 a_5653_n12325# a_6012_n12503# 0.05fF
C5172 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X a_4365_n4709# 0.18fF
C5173 a_3436_n4887# a_4464_n4887# 0.02fF
C5174 a_10805_n4709# a_10805_n5797# 0.02fF
C5175 a_9706_n14109# a_9616_n13591# 0.02fF
C5176 a_3436_n3799# a_3373_n5405# 0.00fF
C5177 a_6941_n5797# a_6941_n4709# 0.02fF
C5178 a_10805_n12325# a_10904_n12503# 0.48fF
C5179 a_2085_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.12fF
C5180 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_9813_n4317# 0.01fF
C5181 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.03fF
C5182 a_8588_n4887# sky130_fd_sc_hd__clkinv_4_3/A 0.10fF
C5183 a_n2248_n7037# VDD 0.23fF
C5184 a_8229_n10613# a_8229_n12325# 0.00fF
C5185 a_3176_n5975# a_3266_n5405# 0.01fF
C5186 a_1888_n11415# a_1722_n11933# 0.04fF
C5187 a_1789_n11237# a_1978_n11933# 0.02fF
C5188 a_5949_n4317# a_5752_n3255# 0.00fF
C5189 a_5842_n4317# a_6012_n3255# 0.00fF
C5190 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VDD 0.89fF
C5191 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6794_n7203# 0.00fF
C5192 a_9517_n1909# a_9616_n3255# 0.00fF
C5193 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VDD 0.84fF
C5194 a_7237_n9213# a_5842_n9213# 0.01fF
C5195 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VDD 0.88fF
C5196 a_4724_n3799# a_4661_n2685# 0.00fF
C5197 a_5842_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.05fF
C5198 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_7130_n11933# 0.03fF
C5199 a_5949_n11933# a_7237_n11933# 0.01fF
C5200 a_5842_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C5201 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_7130_n10301# 0.00fF
C5202 a_6941_n13413# a_8229_n13413# 0.01fF
C5203 a_8588_n10871# a_8525_n10301# 0.01fF
C5204 a_6874_n9213# a_8162_n9213# 0.01fF
C5205 a_4365_n3621# a_4464_n3255# 0.01fF
C5206 a_4464_n3799# a_4365_n2997# 0.01fF
C5207 a_9876_n10871# a_9706_n9213# 0.00fF
C5208 a_11164_n3799# a_11164_n4887# 0.02fF
C5209 a_690_n4317# a_600_n3799# 0.02fF
C5210 a_9450_n6493# a_9517_n5797# 0.01fF
C5211 Bd a_13765_n2685# 0.12fF
C5212 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_501_n5797# 0.02fF
C5213 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VDD 0.82fF
C5214 sky130_fd_sc_hd__nand2_4_0/Y Bd 0.01fF
C5215 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A 0.51fF
C5216 a_3176_n13591# a_3266_n11933# 0.00fF
C5217 a_9616_n12503# a_9517_n13413# 0.00fF
C5218 a_9517_n12325# a_9616_n13591# 0.00fF
C5219 a_9450_n14109# a_10738_n13789# 0.01fF
C5220 a_10805_n11237# a_10738_n10301# 0.00fF
C5221 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_6941_n9525# 0.01fF
C5222 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VDD 0.86fF
C5223 a_9616_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C5224 a_5653_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C5225 a_797_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.12fF
C5226 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X a_5586_n9213# 0.03fF
C5227 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.32fF
C5228 a_1888_n5975# a_1978_n5405# 0.01fF
C5229 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkinv_4_4/A 0.08fF
C5230 a_8162_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.03fF
C5231 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_9450_n509# 0.00fF
C5232 a_501_n12325# a_501_n13413# 0.02fF
C5233 a_1978_n2685# VDD 0.44fF
C5234 a_8418_n509# a_8525_n509# 0.55fF
C5235 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X a_5752_n4887# 0.01fF
C5236 a_5752_n12503# a_7300_n12503# 0.01fF
C5237 a_6012_n12503# a_7040_n12503# 0.02fF
C5238 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_6941_n12325# 0.18fF
C5239 a_4464_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.03fF
C5240 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.02fF
C5241 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VDD 0.84fF
C5242 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkinv_4_3/A 0.70fF
C5243 a_4365_n10613# a_4554_n11933# 0.00fF
C5244 a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.01fF
C5245 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_4298_n5405# 0.03fF
C5246 a_9517_n11237# a_9616_n12503# 0.00fF
C5247 a_10738_n6173# VDD 0.13fF
C5248 a_8229_n4709# a_8229_n2997# 0.00fF
C5249 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8229_n13413# 0.01fF
C5250 a_5586_n11933# a_5586_n10301# 0.01fF
C5251 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.05fF
C5252 a_5842_n4317# a_4554_n4317# 0.01fF
C5253 a_5949_n4317# a_4298_n4317# 0.00fF
C5254 a_5586_n4317# a_4661_n4317# 0.02fF
C5255 p1d_b a_13765_n10301# 0.02fF
C5256 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_n428_n2167# 0.00fF
C5257 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C5258 a_8588_n8695# a_8588_n9783# 0.02fF
C5259 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X p2 0.02fF
C5260 a_3176_n3799# a_3266_n4317# 0.02fF
C5261 a_6941_n11237# a_8229_n11237# 0.01fF
C5262 a_6941_n3621# a_8328_n3799# 0.01fF
C5263 a_4365_n8437# a_5653_n8437# 0.01fF
C5264 a_7040_n3799# a_8229_n3621# 0.01fF
C5265 a_5752_n13591# a_5842_n11933# 0.00fF
C5266 a_501_n3621# a_1789_n3621# 0.01fF
C5267 a_5653_n4709# VDD 0.35fF
C5268 a_7237_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.12fF
C5269 a_5949_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C5270 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_7237_n10301# 0.02fF
C5271 a_8229_n13413# a_8328_n13591# 0.48fF
C5272 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C5273 a_8162_n9213# a_8418_n9213# 0.19fF
C5274 a_3077_n5797# a_3010_n4317# 0.00fF
C5275 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9876_n5975# 0.03fF
C5276 a_9813_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C5277 a_10738_n13789# a_11101_n13021# 0.01fF
C5278 a_1888_n3255# a_501_n2997# 0.01fF
C5279 a_10805_n8437# a_10738_n10301# 0.00fF
C5280 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1789_n3621# 0.01fF
C5281 a_11101_n11933# a_9450_n11933# 0.00fF
C5282 a_10994_n11933# a_9706_n11933# 0.01fF
C5283 a_11164_n13591# a_11164_n12503# 0.02fF
C5284 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.08fF
C5285 a_3176_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C5286 a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C5287 a_3077_n12325# a_3010_n13021# 0.01fF
C5288 a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.00fF
C5289 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_4298_n11933# 0.00fF
C5290 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.00fF
C5291 Bd_b sky130_fd_sc_hd__nand2_4_3/A 0.27fF
C5292 a_4298_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.03fF
C5293 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.02fF
C5294 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkinv_4_3/A 0.05fF
C5295 sky130_fd_sc_hd__nand2_4_3/B p2 0.06fF
C5296 sky130_fd_sc_hd__clkinv_4_3/Y a_11164_n4887# 0.01fF
C5297 a_5949_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.12fF
C5298 a_n688_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C5299 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_860_n9783# 0.00fF
C5300 a_4365_n12325# a_4724_n12503# 0.05fF
C5301 a_8162_n10301# a_8162_n11933# 0.01fF
C5302 a_8229_n12325# VDD 0.35fF
C5303 a_7130_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C5304 a_9517_n4709# a_9616_n3255# 0.00fF
C5305 sky130_fd_sc_hd__dfxbp_1_0/Q a_6658_n7363# 0.03fF
C5306 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkinv_1_4/Y 0.03fF
C5307 a_9517_n8437# a_9450_n9213# 0.01fF
C5308 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X a_6012_n4887# 0.03fF
C5309 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_8328_n12503# 0.01fF
C5310 a_4724_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C5311 a_7040_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.03fF
C5312 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.02fF
C5313 a_9813_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.01fF
C5314 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_9876_n1079# 0.03fF
C5315 Ad VDD 4.21fF
C5316 a_600_n9783# a_1789_n9525# 0.01fF
C5317 a_501_n9525# a_1888_n9783# 0.01fF
C5318 a_6941_n8437# a_6874_n9213# 0.01fF
C5319 a_4724_n5975# a_4661_n5405# 0.01fF
C5320 a_501_n12325# a_434_n11933# 0.01fF
C5321 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C5322 a_600_n8695# a_690_n9213# 0.01fF
C5323 sky130_fd_sc_hd__nand2_4_1/B a_10994_n5405# 0.00fF
C5324 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_4661_n9213# 0.00fF
C5325 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C5326 a_9517_n5797# a_10805_n5797# 0.01fF
C5327 a_3176_n11415# a_3373_n11933# 0.02fF
C5328 a_3436_n11415# a_3266_n11933# 0.04fF
C5329 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7300_n3255# 0.01fF
C5330 a_8229_n3621# a_8588_n3799# 0.05fF
C5331 a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C5332 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_4298_n4317# 0.03fF
C5333 a_7237_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5334 a_10904_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C5335 a_8229_n11237# a_8328_n11415# 0.49fF
C5336 a_6874_n5405# a_6941_n4709# 0.01fF
C5337 a_4365_n13413# a_5653_n13413# 0.01fF
C5338 a_3176_n1079# a_3266_n2685# 0.00fF
C5339 a_5653_n8437# a_5752_n8695# 0.49fF
C5340 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_4_4/A 0.04fF
C5341 a_7040_n4887# VDD 0.44fF
C5342 a_1789_n3621# a_1888_n3799# 0.49fF
C5343 a_8328_n13591# a_9616_n13591# 0.01fF
C5344 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.02fF
C5345 a_8229_n13413# a_9876_n13591# 0.00fF
C5346 a_8588_n13591# a_9517_n13413# 0.02fF
C5347 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6941_n821# 0.01fF
C5348 a_7130_n14109# a_7040_n12503# 0.00fF
C5349 a_6874_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.03fF
C5350 a_8525_n9213# a_9450_n9213# 0.02fF
C5351 a_8418_n9213# a_9706_n9213# 0.01fF
C5352 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_7300_n10871# 0.00fF
C5353 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C5354 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.08fF
C5355 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.83fF
C5356 sky130_fd_sc_hd__clkinv_1_0/A a_9616_n1079# 0.07fF
C5357 a_10805_n12325# a_10738_n13789# 0.01fF
C5358 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C5359 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_2085_n4317# 0.01fF
C5360 sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__nand2_4_2/A 0.26fF
C5361 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C5362 a_434_n1597# a_600_n3255# 0.00fF
C5363 a_690_n1597# a_501_n2997# 0.00fF
C5364 a_9450_n6493# a_9450_n8125# 0.01fF
C5365 a_5653_n10613# a_4365_n10613# 0.01fF
C5366 a_9616_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C5367 p1 p1d 0.20fF
C5368 a_9450_n2685# a_10738_n2685# 0.01fF
C5369 a_10994_n9213# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C5370 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C5371 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.29fF
C5372 a_7300_n4887# VDD 0.77fF
C5373 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_3436_n9783# 0.01fF
C5374 a_4464_n9783# a_4365_n10613# 0.00fF
C5375 a_11164_n8695# a_11101_n9213# 0.01fF
C5376 a_4724_n13591# a_4661_n11933# 0.00fF
C5377 a_7130_n2685# a_7130_n1597# 0.01fF
C5378 a_1888_n12503# a_3077_n12325# 0.01fF
C5379 a_1789_n12325# a_3176_n12503# 0.01fF
C5380 a_1888_n3255# a_1978_n4317# 0.01fF
C5381 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8418_n10301# 0.03fF
C5382 a_5752_n3799# a_5653_n1909# 0.00fF
C5383 a_2366_n8125# sky130_fd_sc_hd__clkinv_1_3/Y 0.34fF
C5384 a_5653_n3621# a_5752_n2167# 0.00fF
C5385 a_4298_n2685# a_5586_n2685# 0.01fF
C5386 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.02fF
C5387 a_4464_n12503# a_6012_n12503# 0.01fF
C5388 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.29fF
C5389 a_9450_n4317# a_9616_n3799# 0.04fF
C5390 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_5949_n2685# 0.01fF
C5391 a_9706_n4317# a_9517_n3621# 0.02fF
C5392 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.02fF
C5393 a_3010_n5405# a_3266_n5405# 0.19fF
C5394 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C5395 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_8588_n12503# 0.03fF
C5396 a_7237_n6493# a_7040_n5975# 0.02fF
C5397 a_7130_n6493# a_7300_n5975# 0.04fF
C5398 p1d_b a_13765_n12477# 0.12fF
C5399 a_13765_n11933# p1d 0.12fF
C5400 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.02fF
C5401 a_2148_n8695# VDD 0.80fF
C5402 a_9616_n9783# a_10805_n9525# 0.01fF
C5403 a_9517_n9525# a_10904_n9783# 0.01fF
C5404 a_9450_n2685# a_9616_n3799# 0.00fF
C5405 a_9706_n2685# a_9517_n3621# 0.00fF
C5406 a_1789_n9525# a_2148_n9783# 0.05fF
C5407 a_8162_n509# a_8162_n1597# 0.02fF
C5408 a_13765_n13565# p1 2.47fF
C5409 a_1978_n10301# a_2148_n8695# 0.00fF
C5410 a_2085_n10301# a_1888_n8695# 0.00fF
C5411 a_10805_n5797# a_10904_n5975# 0.48fF
C5412 a_9616_n10871# a_9616_n12503# 0.00fF
C5413 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_1722_n9213# 0.03fF
C5414 a_10738_n509# a_10805_n821# 0.03fF
C5415 a_9517_n1909# a_10805_n1909# 0.01fF
C5416 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__nand2_4_0/B 0.04fF
C5417 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_6874_n9213# 0.00fF
C5418 a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.00fF
C5419 a_4365_n3621# a_4365_n4709# 0.02fF
C5420 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_797_n2685# 0.01fF
C5421 a_2729_n8125# sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C5422 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.04fF
C5423 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_5949_n11933# 0.00fF
C5424 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C5425 a_11164_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.03fF
C5426 a_8525_n10301# a_8525_n9213# 0.02fF
C5427 a_8588_n11415# a_9517_n11237# 0.02fF
C5428 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_7/Y 0.02fF
C5429 a_4724_n3799# a_4661_n4317# 0.01fF
C5430 a_8588_n3799# a_9616_n3799# 0.02fF
C5431 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X a_9517_n3621# 0.18fF
C5432 a_4365_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C5433 a_2366_n509# a_2148_n1079# 0.03fF
C5434 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_4298_n2685# 0.00fF
C5435 a_5653_n13413# a_5752_n13591# 0.47fF
C5436 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C5437 sky130_fd_sc_hd__clkinv_1_5/A a_6101_n7254# 0.02fF
C5438 a_10738_n2685# a_11101_n2685# 0.05fF
C5439 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkinv_4_3/A 0.09fF
C5440 a_6794_n7203# p2 0.01fF
C5441 a_9517_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C5442 a_9616_n13591# a_9876_n13591# 0.28fF
C5443 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_10738_n8125# 0.02fF
C5444 a_10805_n11237# VDD 0.32fF
C5445 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VDD 0.90fF
C5446 a_7237_n509# a_7300_n1079# 0.01fF
C5447 a_11101_n11933# a_10994_n10301# 0.00fF
C5448 a_3077_n11237# a_4365_n11237# 0.01fF
C5449 a_2366_n6493# sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C5450 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.01fF
C5451 a_4464_n5975# a_4554_n4317# 0.00fF
C5452 a_10994_n11933# a_11101_n10301# 0.00fF
C5453 sky130_fd_sc_hd__clkinv_4_4/A A 0.01fF
C5454 sky130_fd_sc_hd__clkinv_1_0/A a_11164_n1079# 0.11fF
C5455 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_50/X 0.06fF
C5456 a_1789_n4709# a_3436_n4887# 0.00fF
C5457 a_8162_n6493# a_9706_n6493# 0.01fF
C5458 a_6941_n8437# a_5752_n8695# 0.01fF
C5459 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.33fF
C5460 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_600_n9783# 0.04fF
C5461 a_13765_n11933# a_13765_n13565# 0.01fF
C5462 a_13765_n2141# a_13765_n1597# 0.34fF
C5463 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_8588_n9783# 0.00fF
C5464 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VDD 0.85fF
C5465 a_8525_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.00fF
C5466 a_4464_n12503# a_4554_n13021# 0.02fF
C5467 a_5842_n13021# a_6012_n12503# 0.04fF
C5468 a_5949_n13021# a_5752_n12503# 0.02fF
C5469 a_6941_n10613# a_6874_n10301# 0.01fF
C5470 a_3077_n12325# a_3436_n12503# 0.05fF
C5471 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.04fF
C5472 a_9450_n13021# a_10738_n13021# 0.01fF
C5473 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n1597# 0.01fF
C5474 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C5475 a_8162_n10301# a_9706_n10301# 0.01fF
C5476 a_9876_n8695# a_9706_n10301# 0.00fF
C5477 a_4724_n9783# a_4724_n8695# 0.02fF
C5478 a_9616_n8695# a_9813_n10301# 0.00fF
C5479 a_5586_n2685# a_5842_n2685# 0.19fF
C5480 a_600_n1079# a_434_n2685# 0.00fF
C5481 a_860_n9783# sky130_fd_sc_hd__clkinv_1_3/A 0.00fF
C5482 a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.01fF
C5483 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.02fF
C5484 a_3176_n3255# a_3266_n1597# 0.00fF
C5485 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkinv_1_0/A 0.01fF
C5486 a_3373_n5405# a_4298_n5405# 0.02fF
C5487 a_3010_n5405# a_4661_n5405# 0.00fF
C5488 a_3266_n5405# a_4554_n5405# 0.01fF
C5489 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkinv_1_5/A 0.06fF
C5490 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A a_501_n2997# 0.17fF
C5491 a_3176_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C5492 a_6373_n7349# a_7212_n7203# 0.02fF
C5493 a_10805_n9525# a_11164_n9783# 0.05fF
C5494 a_9813_n6493# sky130_fd_sc_hd__clkinv_4_3/A 0.02fF
C5495 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X a_3077_n9525# 0.18fF
C5496 a_1888_n9783# a_3436_n9783# 0.01fF
C5497 a_2148_n9783# a_3176_n9783# 0.02fF
C5498 sky130_fd_sc_hd__dfxbp_1_0/Q_N a_5842_n9213# 0.00fF
C5499 a_5653_n11237# a_5842_n11933# 0.02fF
C5500 Bd VDD 4.20fF
C5501 a_7130_n2685# a_6941_n1909# 0.02fF
C5502 a_7130_n4317# a_6941_n4709# 0.02fF
C5503 a_6874_n4317# a_7040_n4887# 0.04fF
C5504 a_6874_n2685# a_7040_n2167# 0.04fF
C5505 a_10805_n1909# a_10904_n2167# 0.48fF
C5506 sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C5507 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.06fF
C5508 a_7300_n10871# a_7237_n9213# 0.00fF
C5509 a_7212_n7203# VDD 0.19fF
C5510 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X a_4661_n11933# 0.01fF
C5511 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.03fF
C5512 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VDD 2.54fF
C5513 a_10805_n8437# VDD 0.32fF
C5514 a_1789_n10613# VDD 0.35fF
C5515 a_n2436_n7037# VDD 0.79fF
C5516 a_434_n5405# a_690_n5405# 0.19fF
C5517 a_501_n11237# a_1888_n11415# 0.01fF
C5518 a_600_n11415# a_1789_n11237# 0.01fF
C5519 sky130_fd_sc_hd__nand2_4_1/A a_6665_n7459# 0.03fF
C5520 a_4724_n1079# a_4661_n2685# 0.00fF
C5521 a_501_n11237# a_501_n10613# 0.05fF
C5522 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C5523 a_4365_n11237# a_4464_n11415# 0.49fF
C5524 a_1789_n10613# a_1978_n10301# 0.02fF
C5525 a_1888_n10871# a_1722_n10301# 0.04fF
C5526 a_5842_n13021# a_4554_n13021# 0.01fF
C5527 a_434_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C5528 Ad_b a_6006_n7607# 0.01fF
C5529 a_5949_n13021# a_4298_n13021# 0.00fF
C5530 a_3176_n4887# a_3436_n4887# 0.28fF
C5531 a_3077_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.02fF
C5532 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_4365_n4709# 0.01fF
C5533 a_8328_n4887# a_8525_n5405# 0.02fF
C5534 a_8588_n4887# a_8418_n5405# 0.04fF
C5535 a_6874_n13021# VDD 0.75fF
C5536 a_3373_n5405# a_1722_n5405# 0.00fF
C5537 sky130_fd_sc_hd__dfxbp_1_1/D a_n1570_n6769# 0.15fF
C5538 a_8229_n9525# a_8328_n11415# 0.00fF
C5539 a_10994_n5405# a_10805_n3621# 0.00fF
C5540 a_3266_n5405# a_1978_n5405# 0.01fF
C5541 a_10738_n5405# a_10904_n3799# 0.00fF
C5542 a_3436_n12503# a_4464_n12503# 0.02fF
C5543 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_4365_n12325# 0.18fF
C5544 a_5586_n2685# a_5752_n3255# 0.04fF
C5545 a_8525_n2685# a_8525_n1597# 0.02fF
C5546 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.04fF
C5547 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C5548 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.08fF
C5549 a_2148_n13591# a_2085_n13021# 0.01fF
C5550 a_5949_n2685# a_5752_n1079# 0.00fF
C5551 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_5586_n5405# 0.00fF
C5552 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_8588_n5975# 0.03fF
C5553 a_9876_n3799# a_8229_n3621# 0.00fF
C5554 a_5842_n2685# a_6012_n1079# 0.00fF
C5555 a_4554_n5405# a_4661_n5405# 0.55fF
C5556 a_4298_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.03fF
C5557 a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C5558 a_2622_n6493# a_2622_n8125# 0.00fF
C5559 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_6658_n7363# 0.00fF
C5560 a_6874_n6493# a_6794_n7203# 0.01fF
C5561 a_9616_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C5562 a_7237_n6493# a_6665_n7459# 0.00fF
C5563 a_7130_n6493# a_6865_n7304# 0.01fF
C5564 a_4365_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C5565 a_3176_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.03fF
C5566 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.29fF
C5567 a_8162_n14109# a_8418_n14109# 0.19fF
C5568 a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C5569 a_9813_n11933# VDD 0.33fF
C5570 a_4623_n7349# a_4554_n9213# 0.00fF
C5571 a_9706_n6493# a_9517_n5797# 0.02fF
C5572 sky130_fd_sc_hd__nand2_4_2/A a_8418_n14109# 0.03fF
C5573 a_7040_n8695# a_6658_n7363# 0.00fF
C5574 a_4464_n5975# a_4623_n7349# 0.00fF
C5575 a_11164_n10871# a_11164_n12503# 0.01fF
C5576 a_7237_n6493# a_7130_n5405# 0.00fF
C5577 a_7130_n6493# a_7237_n5405# 0.00fF
C5578 a_5752_n3799# a_5752_n4887# 0.01fF
C5579 a_1888_n3255# a_1978_n2685# 0.02fF
C5580 a_3176_n10871# VDD 0.46fF
C5581 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VDD 0.78fF
C5582 a_797_n5405# a_1722_n5405# 0.02fF
C5583 a_690_n5405# a_1978_n5405# 0.01fF
C5584 a_5586_n10301# VDD 0.76fF
C5585 a_7300_n2167# a_7300_n3799# 0.01fF
C5586 a_7300_n8695# VDD 0.78fF
C5587 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__nand2_4_0/Y 0.44fF
C5588 sky130_fd_sc_hd__clkinv_4_3/Y Ad_b 0.07fF
C5589 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C5590 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_8162_n4317# 0.03fF
C5591 a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C5592 a_797_n10301# a_797_n9213# 0.02fF
C5593 a_3176_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.00fF
C5594 a_9616_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C5595 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_8328_n5975# 0.03fF
C5596 a_3010_n10301# a_4554_n10301# 0.01fF
C5597 a_3266_n10301# a_4298_n10301# 0.02fF
C5598 a_8418_n13021# VDD 0.46fF
C5599 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_9876_n9783# 0.00fF
C5600 a_10994_n9213# a_11164_n9783# 0.04fF
C5601 a_11101_n9213# a_10904_n9783# 0.02fF
C5602 a_9616_n8695# a_9813_n8125# 0.02fF
C5603 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7300_n12503# 0.03fF
C5604 a_7237_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C5605 a_n787_n12325# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C5606 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_1978_n1597# 0.01fF
C5607 a_3373_n1597# a_2085_n1597# 0.01fF
C5608 a_2366_n6493# a_2729_n6493# 0.05fF
C5609 a_7040_n13591# a_7237_n11933# 0.00fF
C5610 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6658_n7363# 0.00fF
C5611 a_7300_n13591# a_7130_n11933# 0.00fF
C5612 a_7130_n1597# a_6941_n821# 0.02fF
C5613 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_3176_n8695# 0.05fF
C5614 a_10994_n11933# a_10904_n13591# 0.00fF
C5615 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_4724_n11415# 0.00fF
C5616 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C5617 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C5618 a_3077_n1909# a_3266_n1597# 0.02fF
C5619 a_9876_n3799# a_9616_n3799# 0.28fF
C5620 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_9517_n3621# 0.02fF
C5621 a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C5622 a_3176_n2167# a_3010_n1597# 0.04fF
C5623 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5842_n5405# 0.03fF
C5624 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VDD 0.82fF
C5625 a_6941_n9525# a_8229_n9525# 0.01fF
C5626 a_8588_n2167# a_8525_n1597# 0.01fF
C5627 a_1789_n1909# a_2148_n2167# 0.05fF
C5628 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.01fF
C5629 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_3436_n3255# 0.01fF
C5630 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.03fF
C5631 a_6874_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C5632 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.00fF
C5633 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_11164_n11415# 0.03fF
C5634 a_5752_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C5635 a_1888_n5975# a_2148_n5975# 0.28fF
C5636 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.02fF
C5637 a_6012_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.29fF
C5638 a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C5639 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.02fF
C5640 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4365_n821# 0.01fF
C5641 a_10738_n9213# a_10738_n10301# 0.02fF
C5642 sky130_fd_sc_hd__clkinv_1_0/A a_434_n1597# 0.00fF
C5643 a_4298_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.03fF
C5644 a_8418_n14109# a_9706_n14109# 0.01fF
C5645 a_8525_n14109# a_9450_n14109# 0.02fF
C5646 sky130_fd_sc_hd__clkinv_4_8/A VDD 7.41fF
C5647 a_8162_n14109# a_9813_n14109# 0.00fF
C5648 a_7300_n11415# a_7130_n11933# 0.04fF
C5649 a_9813_n9213# a_10994_n9213# 0.01fF
C5650 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10738_n9213# 0.35fF
C5651 a_7237_n13021# a_7130_n14109# 0.00fF
C5652 a_7130_n13021# a_7237_n14109# 0.00fF
C5653 a_7040_n11415# a_7237_n11933# 0.02fF
C5654 sky130_fd_sc_hd__nand2_4_2/A a_9813_n14109# 0.03fF
C5655 a_9813_n1597# a_10994_n1597# 0.01fF
C5656 a_9706_n1597# a_11101_n1597# 0.01fF
C5657 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n1597# 0.35fF
C5658 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.04fF
C5659 a_5653_n12325# a_5586_n11933# 0.01fF
C5660 a_501_n4709# a_434_n5405# 0.01fF
C5661 a_10994_n5405# a_11164_n4887# 0.04fF
C5662 a_10738_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.02fF
C5663 a_434_n4317# a_501_n2997# 0.00fF
C5664 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_2085_n13021# 0.00fF
C5665 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C5666 a_9517_n4709# a_10805_n4709# 0.01fF
C5667 a_7130_n10301# VDD 0.44fF
C5668 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.01fF
C5669 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VDD 0.82fF
C5670 a_11164_n3799# a_10994_n2685# 0.00fF
C5671 a_10904_n3799# a_11101_n2685# 0.00fF
C5672 a_3176_n10871# a_3373_n10301# 0.02fF
C5673 a_3436_n10871# a_3266_n10301# 0.04fF
C5674 a_8588_n4887# a_8525_n4317# 0.01fF
C5675 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VDD 0.84fF
C5676 a_10904_n3799# a_10994_n4317# 0.02fF
C5677 a_8229_n1909# a_7300_n2167# 0.02fF
C5678 a_8588_n2167# a_6941_n1909# 0.00fF
C5679 a_8328_n2167# a_7040_n2167# 0.01fF
C5680 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_8588_n5975# 0.00fF
C5681 a_4464_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.03fF
C5682 a_6012_n3255# a_6941_n2997# 0.02fF
C5683 a_5752_n3255# a_7040_n3255# 0.01fF
C5684 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.03fF
C5685 a_5653_n11237# a_4365_n11237# 0.01fF
C5686 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.04fF
C5687 a_5752_n13591# a_6941_n13413# 0.01fF
C5688 a_5653_n13413# a_7040_n13591# 0.01fF
C5689 sky130_fd_sc_hd__clkinv_4_4/Y Bd_b 0.08fF
C5690 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A a_434_n2685# 0.03fF
C5691 a_9813_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.12fF
C5692 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkinv_1_5/A 0.21fF
C5693 a_7300_n9783# sky130_fd_sc_hd__nand2_4_3/Y 0.11fF
C5694 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_3436_n4887# 0.00fF
C5695 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.00fF
C5696 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.06fF
C5697 a_600_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.03fF
C5698 a_434_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.01fF
C5699 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.02fF
C5700 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_434_n5405# 0.04fF
C5701 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.04fF
C5702 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_9616_n3799# 0.00fF
C5703 a_2148_n2167# a_2148_n3799# 0.01fF
C5704 a_9813_n14109# a_9813_n13021# 0.02fF
C5705 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.08fF
C5706 a_8418_n8125# a_9813_n8125# 0.01fF
C5707 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C5708 a_8229_n12325# a_8162_n11933# 0.01fF
C5709 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3266_n9213# 0.03fF
C5710 a_2085_n9213# a_3373_n9213# 0.01fF
C5711 a_1722_n10301# a_1789_n9525# 0.01fF
C5712 a_1888_n2167# a_3436_n2167# 0.01fF
C5713 sky130_fd_sc_hd__nand2_4_0/Y a_7300_n2167# 0.11fF
C5714 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_3077_n1909# 0.18fF
C5715 a_2148_n2167# a_3176_n2167# 0.02fF
C5716 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.02fF
C5717 a_1888_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.00fF
C5718 a_2148_n5975# a_3436_n5975# 0.01fF
C5719 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_3176_n5975# 0.05fF
C5720 a_4661_n1597# a_4724_n1079# 0.01fF
C5721 a_9450_n14109# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C5722 a_9706_n14109# a_9813_n14109# 0.52fF
C5723 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C5724 a_2148_n13591# a_600_n13591# 0.01fF
C5725 a_10994_n9213# sky130_fd_sc_hd__clkinv_4_10/Y 0.01fF
C5726 a_1888_n13591# a_860_n13591# 0.02fF
C5727 a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.18fF
C5728 a_3176_n3255# VDD 0.46fF
C5729 a_6941_n1909# a_6941_n821# 0.02fF
C5730 a_1978_n1597# a_2085_n2685# 0.00fF
C5731 a_2085_n1597# a_1978_n2685# 0.00fF
C5732 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_4464_n2167# 0.05fF
C5733 a_3436_n2167# a_4724_n2167# 0.01fF
C5734 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_3436_n10871# 0.00fF
C5735 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.00fF
C5736 a_3176_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C5737 a_9517_n3621# VDD 0.34fF
C5738 a_5752_n5975# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C5739 a_10805_n4709# a_10904_n4887# 0.48fF
C5740 a_5842_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.05fF
C5741 a_8588_n10871# a_9876_n10871# 0.01fF
C5742 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_9616_n10871# 0.05fF
C5743 a_6012_n9783# a_5842_n9213# 0.04fF
C5744 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.06fF
C5745 a_690_n4317# a_1722_n4317# 0.02fF
C5746 a_434_n4317# a_1978_n4317# 0.01fF
C5747 a_5586_n1597# a_5752_n3255# 0.00fF
C5748 a_6941_n9525# a_6874_n9213# 0.01fF
C5749 a_8162_n1597# a_8328_n3255# 0.00fF
C5750 a_7237_n8125# a_6658_n7363# 0.00fF
C5751 sky130_fd_sc_hd__clkinv_1_0/A a_4365_n821# 0.06fF
C5752 a_8418_n1597# a_8229_n2997# 0.00fF
C5753 a_6874_n8125# a_6865_n7304# 0.02fF
C5754 a_7130_n8125# a_6665_n7459# 0.00fF
C5755 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.00fF
C5756 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_6012_n2167# 0.03fF
C5757 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C5758 sky130_fd_sc_hd__nand2_4_1/B VDD 1.40fF
C5759 a_7040_n3255# a_7300_n3255# 0.28fF
C5760 a_6941_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C5761 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X a_8229_n2997# 0.01fF
C5762 a_501_n3621# a_690_n5405# 0.00fF
C5763 a_6874_n6493# a_8162_n6493# 0.01fF
C5764 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C5765 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_2085_n10301# 0.00fF
C5766 a_600_n3799# a_434_n5405# 0.00fF
C5767 Bd_b a_6101_n7254# 0.01fF
C5768 a_5842_n1597# a_6012_n1079# 0.04fF
C5769 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5653_n5797# 0.00fF
C5770 a_5949_n1597# a_5752_n1079# 0.02fF
C5771 a_10738_n4317# sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C5772 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C5773 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X a_8525_n11933# 0.00fF
C5774 a_9616_n12503# a_9813_n13021# 0.02fF
C5775 a_8525_n1597# a_8328_n1079# 0.02fF
C5776 a_8418_n1597# a_8588_n1079# 0.04fF
C5777 a_3077_n9525# VDD 0.36fF
C5778 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C5779 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VDD 0.93fF
C5780 a_860_n3255# VDD 0.78fF
C5781 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_2148_n10871# 0.03fF
C5782 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C5783 a_797_n4317# a_797_n5405# 0.02fF
C5784 a_9616_n12503# a_9706_n14109# 0.00fF
C5785 a_501_n5797# a_860_n5975# 0.05fF
C5786 sky130_fd_sc_hd__nand2_4_2/A a_11164_n12503# 0.01fF
C5787 a_3373_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.12fF
C5788 a_3176_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.03fF
C5789 a_5653_n9525# a_5653_n8437# 0.02fF
C5790 a_9450_n6493# a_9616_n4887# 0.00fF
C5791 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.29fF
C5792 a_1789_n4709# a_2148_n4887# 0.05fF
C5793 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6865_n7304# 0.00fF
C5794 a_4365_n12325# a_4298_n11933# 0.01fF
C5795 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.03fF
C5796 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_8525_n11933# 0.01fF
C5797 a_3176_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C5798 a_9706_n1597# a_9616_n3255# 0.00fF
C5799 a_11101_n4317# a_11164_n4887# 0.01fF
C5800 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.04fF
C5801 a_4724_n3255# VDD 0.78fF
C5802 sky130_fd_sc_hd__nand2_1_4/Y Bd_b 0.01fF
C5803 a_n428_n4887# a_501_n4709# 0.02fF
C5804 a_9616_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C5805 a_1722_n9213# a_2085_n9213# 0.05fF
C5806 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8418_n14109# 0.03fF
C5807 a_5949_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C5808 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_7237_n13021# 0.02fF
C5809 a_6874_n1597# a_8162_n1597# 0.01fF
C5810 B_b Bd_b 0.20fF
C5811 a_4298_n1597# a_5586_n1597# 0.01fF
C5812 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.29fF
C5813 a_1722_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C5814 sky130_fd_sc_hd__clkinv_1_3/A VDD 6.20fF
C5815 a_3176_n8695# a_3266_n9213# 0.01fF
C5816 a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.00fF
C5817 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_10805_n3621# 0.17fF
C5818 a_9876_n3799# a_10904_n3799# 0.02fF
C5819 a_8418_n14109# a_8328_n13591# 0.02fF
C5820 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X a_8328_n3255# 0.05fF
C5821 a_9706_n8125# a_9517_n9525# 0.00fF
C5822 clk sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.04fF
C5823 a_9517_n4709# a_9517_n5797# 0.02fF
C5824 a_7300_n3255# a_8588_n3255# 0.01fF
C5825 a_7040_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C5826 a_8162_n6493# a_8418_n6493# 0.19fF
C5827 a_9517_n12325# a_9616_n12503# 0.49fF
C5828 a_5653_n5797# a_5653_n4709# 0.02fF
C5829 a_4661_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C5830 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5949_n5405# 0.02fF
C5831 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C5832 a_6941_n10613# a_6941_n12325# 0.00fF
C5833 a_10738_n9213# VDD 0.70fF
C5834 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.06fF
C5835 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.08fF
C5836 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkinv_4_4/A 0.02fF
C5837 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_n428_n4887# 0.02fF
C5838 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_860_n1079# 0.01fF
C5839 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.01fF
C5840 a_10805_n12325# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C5841 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.02fF
C5842 a_3266_n10301# a_3176_n9783# 0.01fF
C5843 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VDD 0.88fF
C5844 a_434_n2685# a_434_n4317# 0.01fF
C5845 a_4554_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.05fF
C5846 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VDD 0.88fF
C5847 a_9876_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.29fF
C5848 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_8525_n10301# 0.00fF
C5849 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C5850 a_5949_n9213# a_4554_n9213# 0.01fF
C5851 a_3436_n3799# a_3373_n2685# 0.00fF
C5852 a_2148_n4887# a_3176_n4887# 0.02fF
C5853 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_3077_n4709# 0.18fF
C5854 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkinv_1_4/Y 0.03fF
C5855 a_3077_n3621# a_3176_n3255# 0.01fF
C5856 sky130_fd_sc_hd__clkinv_1_0/A a_8229_n821# 0.06fF
C5857 a_3176_n3799# a_3077_n2997# 0.01fF
C5858 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10805_n2997# 0.00fF
C5859 a_8162_n4317# a_8229_n3621# 0.01fF
C5860 a_3077_n1909# VDD 0.36fF
C5861 a_8588_n10871# a_8418_n9213# 0.00fF
C5862 a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C5863 a_5653_n3621# a_6941_n3621# 0.01fF
C5864 a_9876_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C5865 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X a_8588_n3255# 0.00fF
C5866 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.06fF
C5867 a_1978_n9213# a_3373_n9213# 0.01fF
C5868 a_9706_n5405# a_9517_n3621# 0.00fF
C5869 a_1888_n13591# a_1978_n11933# 0.00fF
C5870 a_9450_n5405# a_9616_n3799# 0.00fF
C5871 a_4365_n10613# a_4554_n9213# 0.00fF
C5872 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.44fF
C5873 a_10904_n10871# a_10994_n11933# 0.01fF
C5874 a_7040_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C5875 a_5586_n1597# a_5842_n1597# 0.19fF
C5876 a_5586_n10301# a_5586_n9213# 0.02fF
C5877 a_4365_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C5878 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_4298_n9213# 0.03fF
C5879 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_8162_n8125# 0.00fF
C5880 a_5752_n2167# VDD 0.46fF
C5881 a_7130_n509# a_7237_n509# 0.55fF
C5882 a_6874_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.03fF
C5883 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_8162_n509# 0.00fF
C5884 a_10904_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.02fF
C5885 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_4_4/A 0.45fF
C5886 a_4724_n12503# a_5752_n12503# 0.02fF
C5887 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_5653_n12325# 0.18fF
C5888 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9517_n13413# 0.01fF
C5889 a_9450_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C5890 a_501_n8437# a_2148_n8695# 0.00fF
C5891 a_600_n8695# a_1888_n8695# 0.01fF
C5892 a_10904_n1079# a_10994_n2685# 0.00fF
C5893 a_8588_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.29fF
C5894 a_860_n8695# a_1789_n8437# 0.02fF
C5895 a_501_n4709# a_501_n3621# 0.02fF
C5896 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.05fF
C5897 a_8525_n6493# a_9450_n6493# 0.02fF
C5898 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C5899 a_434_n9213# a_1722_n9213# 0.01fF
C5900 a_9876_n12503# a_10805_n12325# 0.02fF
C5901 a_9517_n12325# a_11164_n12503# 0.00fF
C5902 a_9616_n12503# a_10904_n12503# 0.01fF
C5903 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_8525_n4317# 0.00fF
C5904 a_3077_n10613# a_3266_n11933# 0.00fF
C5905 a_3176_n10871# a_3010_n11933# 0.00fF
C5906 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_11101_n13021# 0.12fF
C5907 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkinv_4_3/A 0.70fF
C5908 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_3010_n5405# 0.03fF
C5909 a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C5910 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VDD 0.66fF
C5911 a_4298_n11933# a_4298_n10301# 0.01fF
C5912 a_690_n4317# a_860_n4887# 0.04fF
C5913 a_797_n4317# a_600_n4887# 0.02fF
C5914 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.01fF
C5915 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C5916 a_5653_n11237# a_6941_n11237# 0.01fF
C5917 a_5052_n7283# a_6101_n7254# 0.02fF
C5918 a_10805_n3621# VDD 0.32fF
C5919 a_3077_n8437# a_4365_n8437# 0.01fF
C5920 a_4661_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C5921 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5949_n10301# 0.02fF
C5922 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C5923 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_7300_n10871# 0.01fF
C5924 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_5842_n9213# 0.05fF
C5925 a_7130_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C5926 sky130_fd_sc_hd__clkinv_4_8/Y a_11164_n13591# 0.30fF
C5927 a_5949_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.12fF
C5928 a_6941_n13413# a_7040_n13591# 0.48fF
C5929 sky130_fd_sc_hd__nand2_4_0/A a_9706_n509# 0.10fF
C5930 a_1789_n5797# a_1722_n4317# 0.00fF
C5931 a_6874_n9213# a_7130_n9213# 0.19fF
C5932 a_9517_n1909# a_9450_n1597# 0.01fF
C5933 a_9813_n11933# a_8162_n11933# 0.00fF
C5934 a_7040_n9783# a_6941_n8437# 0.00fF
C5935 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_501_n3621# 0.01fF
C5936 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.03fF
C5937 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C5938 a_1789_n12325# a_1722_n13021# 0.01fF
C5939 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.02fF
C5940 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.03fF
C5941 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_3010_n11933# 0.00fF
C5942 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_797_n1597# 0.01fF
C5943 a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C5944 a_8229_n9525# a_8162_n8125# 0.00fF
C5945 a_4724_n9783# a_6012_n9783# 0.01fF
C5946 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_5752_n9783# 0.05fF
C5947 a_9876_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C5948 sky130_fd_sc_hd__clkinv_1_0/A B 0.01fF
C5949 a_5949_n1597# a_6874_n1597# 0.02fF
C5950 a_8588_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C5951 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X a_9813_n13021# 0.01fF
C5952 a_4464_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.00fF
C5953 a_6865_n7304# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C5954 a_9813_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C5955 a_4724_n8695# a_4661_n9213# 0.01fF
C5956 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C5957 a_6874_n10301# a_6874_n11933# 0.01fF
C5958 sky130_fd_sc_hd__nand2_1_4/Y a_5052_n7283# 0.01fF
C5959 a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C5960 a_5653_n12325# VDD 0.35fF
C5961 a_7300_n2167# VDD 0.78fF
C5962 a_7237_n509# a_8525_n509# 0.01fF
C5963 a_7130_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C5964 a_797_n2685# VDD 0.36fF
C5965 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.02fF
C5966 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8418_n509# 0.03fF
C5967 a_3436_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.00fF
C5968 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X a_4724_n4887# 0.03fF
C5969 a_9813_n14109# a_9876_n13591# 0.01fF
C5970 a_8229_n8437# a_8162_n9213# 0.01fF
C5971 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_7040_n12503# 0.01fF
C5972 a_5752_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.03fF
C5973 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.02fF
C5974 a_10904_n4887# a_10904_n5975# 0.01fF
C5975 a_13765_n1053# a_13765_n2685# 0.01fF
C5976 a_7040_n5975# a_7040_n4887# 0.01fF
C5977 a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C5978 a_10904_n12503# a_11164_n12503# 0.23fF
C5979 a_1722_n9213# a_1978_n9213# 0.19fF
C5980 a_8525_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.01fF
C5981 a_n2602_n7037# VDD 1.24fF
C5982 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkinv_4_3/A 0.01fF
C5983 a_n1654_n6671# VDD 0.02fF
C5984 a_8328_n10871# a_8328_n12503# 0.00fF
C5985 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.02fF
C5986 a_3436_n5975# a_3373_n5405# 0.01fF
C5987 a_5586_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C5988 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11164_n9783# 0.00fF
C5989 a_10738_n8125# a_10904_n8695# 0.03fF
C5990 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6012_n3255# 0.01fF
C5991 a_1888_n11415# a_2085_n11933# 0.02fF
C5992 a_2148_n11415# a_1978_n11933# 0.04fF
C5993 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C5994 a_6941_n11237# a_7040_n11415# 0.49fF
C5995 a_6941_n3621# a_7300_n3799# 0.05fF
C5996 a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C5997 a_4365_n8437# a_4464_n8695# 0.49fF
C5998 a_3077_n13413# a_4365_n13413# 0.01fF
C5999 a_4464_n4887# VDD 0.44fF
C6000 a_501_n3621# a_600_n3799# 0.49fF
C6001 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.02fF
C6002 a_7300_n13591# a_8229_n13413# 0.02fF
C6003 a_6941_n13413# a_8588_n13591# 0.00fF
C6004 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C6005 a_7040_n13591# a_8328_n13591# 0.01fF
C6006 a_6874_n9213# a_8525_n9213# 0.00fF
C6007 a_7130_n9213# a_8418_n9213# 0.01fF
C6008 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.08fF
C6009 a_n787_n4709# VDD 0.35fF
C6010 a_7237_n9213# a_8162_n9213# 0.02fF
C6011 a_3077_n1909# a_3077_n3621# 0.00fF
C6012 a_10738_n13789# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C6013 a_10805_n11237# a_10738_n13021# 0.00fF
C6014 a_8162_n6493# a_8162_n8125# 0.01fF
C6015 a_3266_n13021# a_4298_n13021# 0.02fF
C6016 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C6017 a_3010_n13021# a_4554_n13021# 0.01fF
C6018 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9450_n11933# 0.03fF
C6019 a_9813_n11933# a_9706_n11933# 0.55fF
C6020 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.04fF
C6021 a_797_n4317# a_860_n3799# 0.01fF
C6022 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_2148_n9783# 0.01fF
C6023 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C6024 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_860_n5975# 0.29fF
C6025 a_10904_n11415# a_10994_n10301# 0.01fF
C6026 a_9813_n14109# a_10738_n13789# 0.01fF
C6027 a_600_n12503# a_1789_n12325# 0.01fF
C6028 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_1888_n13591# 0.01fF
C6029 a_3436_n13591# a_3373_n11933# 0.00fF
C6030 a_4365_n9525# a_4298_n10301# 0.01fF
C6031 a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C6032 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkinv_4_7/A 0.81fF
C6033 a_3010_n2685# a_4298_n2685# 0.01fF
C6034 a_4365_n3621# a_4464_n2167# 0.00fF
C6035 a_3176_n12503# a_4724_n12503# 0.01fF
C6036 a_7040_n12503# VDD 0.44fF
C6037 a_8525_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.12fF
C6038 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A VDD 0.89fF
C6039 a_1888_n3255# a_3176_n3255# 0.01fF
C6040 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_7300_n12503# 0.03fF
C6041 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C6042 a_1888_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C6043 a_4365_n5797# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C6044 a_11164_n4887# VDD 0.67fF
C6045 a_8418_n2685# a_8229_n3621# 0.00fF
C6046 a_8328_n9783# a_9517_n9525# 0.01fF
C6047 a_8162_n2685# a_8328_n3799# 0.00fF
C6048 a_11164_n9783# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C6049 a_501_n9525# a_860_n9783# 0.05fF
C6050 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_11164_n9783# 0.01fF
C6051 a_n688_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C6052 a_13765_n2685# Ad_b 0.02fF
C6053 a_8328_n4887# a_8328_n3255# 0.00fF
C6054 a_5842_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C6055 a_5949_n4317# a_4661_n4317# 0.01fF
C6056 a_9517_n5797# a_9616_n5975# 0.49fF
C6057 a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.18fF
C6058 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_4554_n4317# 0.01fF
C6059 sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4317# 0.04fF
C6060 a_6941_n11237# a_8588_n11415# 0.00fF
C6061 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.04fF
C6062 a_7300_n11415# a_8229_n11237# 0.02fF
C6063 a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.17fF
C6064 a_3436_n3799# a_3373_n4317# 0.01fF
C6065 a_7040_n11415# a_8328_n11415# 0.01fF
C6066 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X a_8229_n3621# 0.18fF
C6067 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_3010_n2685# 0.00fF
C6068 a_7300_n3799# a_8328_n3799# 0.02fF
C6069 a_7040_n3799# a_8588_n3799# 0.01fF
C6070 a_4724_n8695# a_5653_n8437# 0.02fF
C6071 a_4464_n8695# a_5752_n8695# 0.01fF
C6072 a_4365_n13413# a_4464_n13591# 0.48fF
C6073 a_6012_n4887# VDD 0.77fF
C6074 a_4365_n8437# a_6012_n8695# 0.00fF
C6075 a_600_n3799# a_1888_n3799# 0.01fF
C6076 a_860_n3799# a_1789_n3621# 0.02fF
C6077 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C6078 a_1789_n11237# a_3077_n11237# 0.01fF
C6079 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_9517_n13413# 0.01fF
C6080 a_8328_n13591# a_8588_n13591# 0.28fF
C6081 a_8229_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.02fF
C6082 a_8162_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.03fF
C6083 a_8418_n9213# a_8525_n9213# 0.55fF
C6084 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6941_n12325# 0.00fF
C6085 a_6874_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C6086 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_9450_n9213# 0.00fF
C6087 a_3176_n5975# a_3266_n4317# 0.00fF
C6088 a_9813_n11933# a_9706_n10301# 0.00fF
C6089 a_n688_n4887# a_n787_n4709# 0.49fF
C6090 a_1888_n3255# a_860_n3255# 0.02fF
C6091 a_8328_n9783# a_8418_n10301# 0.01fF
C6092 a_10904_n8695# a_10994_n10301# 0.00fF
C6093 a_4464_n10871# a_4365_n10613# 0.49fF
C6094 a_4298_n13021# a_4661_n13021# 0.05fF
C6095 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.02fF
C6096 a_3176_n12503# a_3266_n13021# 0.02fF
C6097 a_6941_n8437# a_8229_n8437# 0.01fF
C6098 sky130_fd_sc_hd__clkinv_4_4/Y A_b 0.04fF
C6099 a_9450_n2685# a_9450_n4317# 0.01fF
C6100 a_5653_n10613# a_5586_n10301# 0.01fF
C6101 a_1789_n12325# a_2148_n12503# 0.05fF
C6102 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_7300_n10871# 0.01fF
C6103 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C6104 a_3077_n12325# VDD 0.36fF
C6105 a_8328_n8695# a_8525_n10301# 0.00fF
C6106 a_4298_n2685# a_4554_n2685# 0.19fF
C6107 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_5752_n12503# 0.01fF
C6108 a_4464_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.03fF
C6109 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.06fF
C6110 sky130_fd_sc_hd__dfxbp_1_0/Q a_6865_n7304# 0.02fF
C6111 a_8588_n12503# VDD 0.77fF
C6112 a_9616_n8695# a_9706_n9213# 0.01fF
C6113 a_2085_n5405# a_3010_n5405# 0.02fF
C6114 a_7040_n5975# a_7212_n7203# 0.00fF
C6115 a_9706_n6493# a_9616_n4887# 0.00fF
C6116 a_9517_n9525# a_9876_n9783# 0.05fF
C6117 a_600_n9783# a_2148_n9783# 0.01fF
C6118 a_860_n9783# a_1888_n9783# 0.02fF
C6119 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X a_1789_n9525# 0.18fF
C6120 a_5586_n13021# a_5653_n13413# 0.01fF
C6121 a_5586_n4317# a_5752_n4887# 0.04fF
C6122 a_5842_n4317# a_5653_n4709# 0.02fF
C6123 a_860_n8695# a_797_n9213# 0.01fF
C6124 a_9876_n5975# a_10805_n5797# 0.02fF
C6125 a_9616_n5975# a_10904_n5975# 0.01fF
C6126 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_4/A 0.11fF
C6127 a_9517_n5797# a_11164_n5975# 0.00fF
C6128 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.05fF
C6129 a_6012_n10871# a_5949_n9213# 0.00fF
C6130 a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.02fF
C6131 a_8328_n11415# a_8588_n11415# 0.28fF
C6132 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.03fF
C6133 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_3373_n11933# 0.01fF
C6134 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_9517_n11237# 0.01fF
C6135 a_9517_n1909# a_9616_n2167# 0.49fF
C6136 a_3436_n1079# a_3373_n2685# 0.00fF
C6137 a_8328_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.03fF
C6138 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_8588_n5975# 0.01fF
C6139 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X a_9616_n3799# 0.01fF
C6140 a_4464_n13591# a_5752_n13591# 0.01fF
C6141 a_7130_n5405# a_7040_n4887# 0.02fF
C6142 a_4724_n13591# a_5653_n13413# 0.02fF
C6143 a_5653_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.02fF
C6144 a_5752_n8695# a_6012_n8695# 0.28fF
C6145 a_1888_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.03fF
C6146 a_8229_n1909# a_8328_n3799# 0.00fF
C6147 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_3176_n8695# 0.01fF
C6148 a_8328_n2167# a_8229_n3621# 0.00fF
C6149 a_8328_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C6150 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X a_9616_n13591# 0.05fF
C6151 a_9616_n11415# VDD 0.42fF
C6152 a_3077_n11237# a_3176_n11415# 0.49fF
C6153 a_8588_n13591# a_9876_n13591# 0.01fF
C6154 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_9706_n9213# 0.03fF
C6155 a_9450_n4317# a_10994_n4317# 0.01fF
C6156 a_7237_n14109# a_7300_n12503# 0.00fF
C6157 a_9706_n4317# a_10738_n4317# 0.02fF
C6158 a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C6159 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_4298_n4317# 0.00fF
C6160 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.82fF
C6161 a_1888_n2167# a_1789_n821# 0.00fF
C6162 a_600_n10871# a_434_n10301# 0.04fF
C6163 a_11164_n12503# a_10738_n13789# 0.01fF
C6164 a_690_n1597# a_860_n3255# 0.00fF
C6165 a_797_n1597# a_600_n3255# 0.00fF
C6166 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C6167 a_13765_n8669# a_13765_n10301# 0.01fF
C6168 a_6012_n10871# a_4365_n10613# 0.00fF
C6169 a_7300_n4887# a_7130_n5405# 0.04fF
C6170 a_9706_n2685# a_10994_n2685# 0.01fF
C6171 a_2085_n5405# a_434_n5405# 0.00fF
C6172 a_6941_n9525# a_7040_n11415# 0.00fF
C6173 a_9813_n2685# a_10738_n2685# 0.02fF
C6174 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_4298_n13021# 0.03fF
C6175 a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C6176 a_7040_n9783# a_6941_n11237# 0.00fF
C6177 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C6178 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_2148_n4887# 0.01fF
C6179 a_9450_n2685# a_11101_n2685# 0.00fF
C6180 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__clkinv_4_10/Y 0.14fF
C6181 a_7237_n2685# a_7237_n1597# 0.02fF
C6182 a_8162_n10301# a_8525_n10301# 0.05fF
C6183 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C6184 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_3077_n12325# 0.18fF
C6185 a_2148_n12503# a_3176_n12503# 0.02fF
C6186 a_1888_n12503# a_3436_n12503# 0.01fF
C6187 a_9517_n8437# a_9450_n8125# 0.01fF
C6188 a_4464_n12503# VDD 0.44fF
C6189 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C6190 a_2729_n8125# sky130_fd_sc_hd__clkinv_1_3/Y 0.02fF
C6191 a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.00fF
C6192 a_4554_n2685# a_5842_n2685# 0.01fF
C6193 a_4661_n2685# a_5586_n2685# 0.02fF
C6194 a_4298_n2685# a_5949_n2685# 0.00fF
C6195 a_13765_n5405# VDD 2.23fF
C6196 a_9813_n4317# a_9616_n3799# 0.02fF
C6197 a_9450_n13021# a_9450_n14109# 0.02fF
C6198 a_3010_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.03fF
C6199 a_3266_n5405# a_3373_n5405# 0.55fF
C6200 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_7300_n5975# 0.03fF
C6201 a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.00fF
C6202 a_7237_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C6203 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_4298_n5405# 0.00fF
C6204 a_6874_n14109# a_7237_n14109# 0.05fF
C6205 a_6941_n8437# a_6874_n8125# 0.01fF
C6206 a_1789_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C6207 a_9616_n9783# a_11164_n9783# 0.01fF
C6208 a_9876_n9783# a_10904_n9783# 0.02fF
C6209 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X a_10805_n9525# 0.17fF
C6210 a_9813_n2685# a_9616_n3799# 0.00fF
C6211 a_1888_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C6212 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X a_3176_n9783# 0.01fF
C6213 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C6214 a_4365_n1909# a_4554_n2685# 0.02fF
C6215 a_8418_n509# a_8418_n1597# 0.01fF
C6216 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_2148_n8695# 0.00fF
C6217 a_10738_n8125# a_10805_n9525# 0.01fF
C6218 a_10738_n509# a_11164_n1079# 0.05fF
C6219 a_9876_n10871# a_9876_n12503# 0.01fF
C6220 a_10904_n5975# a_11164_n5975# 0.23fF
C6221 a_9517_n1909# a_11164_n2167# 0.00fF
C6222 a_501_n1909# a_600_n3799# 0.00fF
C6223 a_9876_n2167# a_10805_n1909# 0.02fF
C6224 sky130_fd_sc_hd__clkinv_4_8/A a_10738_n13021# 0.08fF
C6225 a_11101_n11933# a_10994_n13021# 0.00fF
C6226 a_10994_n11933# a_11101_n13021# 0.00fF
C6227 a_600_n2167# a_501_n3621# 0.00fF
C6228 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.08fF
C6229 a_9616_n2167# a_10904_n2167# 0.01fF
C6230 a_4464_n3799# a_4464_n4887# 0.01fF
C6231 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C6232 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.04fF
C6233 a_600_n10871# VDD 0.47fF
C6234 sky130_fd_sc_hd__clkinv_1_5/A a_6658_n7363# 0.23fF
C6235 a_10738_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.02fF
C6236 a_9876_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.29fF
C6237 sky130_fd_sc_hd__nand2_4_0/Y a_10994_n2685# 0.01fF
C6238 a_3436_n11415# a_4365_n11237# 0.02fF
C6239 a_10994_n2685# a_11101_n4317# 0.00fF
C6240 a_11101_n2685# a_10994_n4317# 0.00fF
C6241 a_3176_n11415# a_4464_n11415# 0.01fF
C6242 a_3077_n11237# a_4724_n11415# 0.00fF
C6243 a_11164_n11415# VDD 0.67fF
C6244 a_9813_n509# a_10738_n509# 0.01fF
C6245 a_10738_n4317# a_11101_n4317# 0.05fF
C6246 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.08fF
C6247 a_6012_n2167# a_6012_n3799# 0.01fF
C6248 a_4724_n5975# a_4661_n4317# 0.00fF
C6249 a_4365_n5797# a_4365_n4709# 0.02fF
C6250 a_13765_n1053# VDD 2.36fF
C6251 a_2148_n4887# a_3436_n4887# 0.01fF
C6252 a_1888_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.00fF
C6253 a_10738_n6173# sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C6254 a_8525_n6493# a_9706_n6493# 0.01fF
C6255 a_5842_n13021# VDD 0.45fF
C6256 a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.18fF
C6257 p1d_b p1 0.08fF
C6258 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C6259 a_3010_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C6260 a_5949_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.01fF
C6261 a_9813_n9213# a_9616_n9783# 0.02fF
C6262 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6012_n12503# 0.03fF
C6263 a_2085_n5405# a_1978_n5405# 0.55fF
C6264 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_1722_n5405# 0.03fF
C6265 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y 0.97fF
C6266 a_13765_n1597# Bd 0.15fF
C6267 a_9450_n13021# a_11101_n13021# 0.00fF
C6268 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_4464_n12503# 0.01fF
C6269 a_9706_n13021# a_10994_n13021# 0.01fF
C6270 a_3176_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.03fF
C6271 a_7040_n10871# a_7130_n10301# 0.02fF
C6272 a_6012_n13591# a_5842_n11933# 0.00fF
C6273 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.04fF
C6274 a_5586_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.03fF
C6275 a_5842_n2685# a_5949_n2685# 0.55fF
C6276 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C6277 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_9813_n10301# 0.00fF
C6278 a_860_n1079# a_690_n2685# 0.00fF
C6279 a_600_n1079# a_797_n2685# 0.00fF
C6280 a_5653_n2997# a_5586_n2685# 0.01fF
C6281 a_2366_n509# a_2622_n509# 0.19fF
C6282 a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C6283 a_10738_n5405# sky130_fd_sc_hd__clkinv_4_4/Y 0.00fF
C6284 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4554_n5405# 0.03fF
C6285 a_3266_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.01fF
C6286 a_1789_n1909# a_1978_n1597# 0.02fF
C6287 a_3373_n5405# a_4661_n5405# 0.01fF
C6288 a_1888_n2167# a_1722_n1597# 0.04fF
C6289 a_1789_n4709# VDD 0.36fF
C6290 a_13765_n11933# p1d_b 2.54fF
C6291 a_5653_n9525# a_6941_n9525# 0.01fF
C6292 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6665_n7459# 0.01fF
C6293 a_6865_n7304# a_7014_n7215# 0.00fF
C6294 a_6665_n7459# a_7212_n7203# 0.22fF
C6295 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A a_860_n3255# 0.02fF
C6296 a_3176_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C6297 a_8162_n8125# a_9450_n8125# 0.01fF
C6298 a_4464_n9783# a_3077_n9525# 0.01fF
C6299 a_4365_n9525# a_3176_n9783# 0.01fF
C6300 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X a_3436_n9783# 0.03fF
C6301 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C6302 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X 0.29fF
C6303 a_6874_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C6304 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6874_n1597# 0.01fF
C6305 a_9450_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C6306 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9450_n1597# 0.01fF
C6307 a_10738_n13789# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C6308 a_5752_n11415# a_5949_n11933# 0.02fF
C6309 a_6012_n11415# a_5842_n11933# 0.04fF
C6310 a_7237_n4317# a_7040_n4887# 0.02fF
C6311 a_7237_n2685# a_7040_n2167# 0.02fF
C6312 a_9616_n1079# a_10805_n821# 0.01fF
C6313 a_9517_n821# a_10904_n1079# 0.01fF
C6314 a_10994_n11933# a_10805_n12325# 0.02fF
C6315 a_10738_n11933# a_10904_n12503# 0.04fF
C6316 a_7130_n2685# a_7300_n2167# 0.04fF
C6317 a_10904_n2167# a_11164_n2167# 0.23fF
C6318 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C6319 a_11164_n8695# VDD 0.67fF
C6320 a_7041_n7581# VDD 0.00fF
C6321 a_434_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.03fF
C6322 a_690_n5405# a_797_n5405# 0.55fF
C6323 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_1722_n5405# 0.00fF
C6324 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C6325 a_860_n11415# a_1888_n11415# 0.02fF
C6326 a_600_n11415# a_2148_n11415# 0.01fF
C6327 a_2148_n10871# VDD 0.78fF
C6328 a_n2163_n6671# VDD 0.47fF
C6329 a_8588_n11415# a_8588_n10871# 0.09fF
C6330 sky130_fd_sc_hd__nand2_1_4/B VDD 2.93fF
C6331 a_3077_n1909# a_3077_n821# 0.02fF
C6332 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_797_n13021# 0.00fF
C6333 a_8229_n4709# a_9517_n4709# 0.01fF
C6334 a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C6335 a_4464_n11415# a_4724_n11415# 0.28fF
C6336 Bd_b sky130_fd_sc_hd__clkinv_4_3/A 0.22fF
C6337 a_9706_n509# a_9517_n821# 0.02fF
C6338 a_4554_n10301# VDD 0.44fF
C6339 a_5949_n13021# a_4661_n13021# 0.01fF
C6340 a_1888_n10871# a_2085_n10301# 0.02fF
C6341 a_7300_n4887# a_7237_n4317# 0.01fF
C6342 Ad_b a_6373_n7349# 0.00fF
C6343 a_2148_n10871# a_1978_n10301# 0.04fF
C6344 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_4554_n13021# 0.01fF
C6345 a_5842_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C6346 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_7300_n5975# 0.00fF
C6347 a_10904_n9783# a_10738_n10301# 0.04fF
C6348 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.02fF
C6349 a_10805_n9525# a_10994_n10301# 0.02fF
C6350 a_7237_n13021# VDD 0.35fF
C6351 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.03fF
C6352 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C6353 a_10994_n5405# a_11164_n3799# 0.00fF
C6354 a_11101_n5405# a_10904_n3799# 0.00fF
C6355 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_8525_n5405# 0.01fF
C6356 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_1978_n5405# 0.01fF
C6357 a_4365_n821# a_4464_n2167# 0.00fF
C6358 sky130_fd_sc_hd__clkinv_1_0/A a_860_n1079# 0.11fF
C6359 a_5949_n2685# a_5752_n3255# 0.02fF
C6360 a_5842_n2685# a_6012_n3255# 0.04fF
C6361 a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C6362 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.04fF
C6363 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_8162_n10301# 0.03fF
C6364 a_10738_n8125# a_10994_n9213# 0.01fF
C6365 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_4724_n11415# 0.01fF
C6366 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C6367 Ad_b VDD 8.08fF
C6368 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.06fF
C6369 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6012_n1079# 0.00fF
C6370 a_5949_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.00fF
C6371 a_4661_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.12fF
C6372 a_9876_n3799# a_8588_n3799# 0.01fF
C6373 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_8328_n3799# 0.00fF
C6374 a_3176_n4887# VDD 0.44fF
C6375 a_6941_n9525# a_7040_n9783# 0.49fF
C6376 a_434_n10301# a_501_n9525# 0.01fF
C6377 a_6941_n12325# a_6874_n11933# 0.01fF
C6378 a_2729_n6493# a_2729_n8125# 0.00fF
C6379 a_4623_n7349# a_4765_n7215# 0.01fF
C6380 a_4724_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C6381 a_8229_n10613# a_8418_n10301# 0.02fF
C6382 a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C6383 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C6384 a_3373_n1597# a_3436_n1079# 0.01fF
C6385 a_8162_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.03fF
C6386 a_8418_n14109# a_8525_n14109# 0.53fF
C6387 a_9706_n6493# a_9876_n5975# 0.04fF
C6388 a_4623_n7349# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C6389 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.41fF
C6390 a_n787_n9525# sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C6391 a_4724_n5975# sky130_fd_sc_hd__dfxbp_1_0/Q 0.00fF
C6392 sky130_fd_sc_hd__dfxbp_1_0/Q a_4661_n9213# 0.00fF
C6393 a_7300_n8695# a_6665_n7459# 0.00fF
C6394 a_797_n1597# a_690_n2685# 0.00fF
C6395 a_690_n1597# a_797_n2685# 0.00fF
C6396 a_7040_n8695# a_6865_n7304# 0.00fF
C6397 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_6658_n7363# 0.01fF
C6398 a_10805_n821# a_11164_n1079# 0.05fF
C6399 a_5653_n1909# a_5653_n821# 0.02fF
C6400 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_10994_n1597# 0.00fF
C6401 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C6402 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_2148_n10871# 0.00fF
C6403 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.10fF
C6404 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VDD 0.83fF
C6405 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_1978_n5405# 0.03fF
C6406 a_9517_n4709# a_9616_n4887# 0.49fF
C6407 a_6941_n3621# VDD 0.35fF
C6408 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.06fF
C6409 a_501_n821# a_1789_n821# 0.01fF
C6410 a_5949_n10301# VDD 0.35fF
C6411 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C6412 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.04fF
C6413 a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C6414 a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C6415 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_10738_n4317# 0.03fF
C6416 a_7130_n1597# a_6941_n2997# 0.00fF
C6417 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C6418 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A VDD 0.87fF
C6419 a_3266_n10301# a_4661_n10301# 0.01fF
C6420 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n10301# 0.35fF
C6421 a_3373_n10301# a_4554_n10301# 0.01fF
C6422 a_9876_n8695# sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C6423 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_797_n10301# 0.00fF
C6424 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_9813_n8125# 0.01fF
C6425 a_5752_n3255# a_6012_n3255# 0.28fF
C6426 a_5653_n13413# a_6012_n13591# 0.05fF
C6427 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.02fF
C6428 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C6429 a_7130_n1597# a_7300_n1079# 0.04fF
C6430 a_1888_n1079# a_1978_n2685# 0.00fF
C6431 a_7237_n1597# a_7040_n1079# 0.02fF
C6432 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10805_n3621# 0.00fF
C6433 a_9813_n6493# a_9813_n8125# 0.00fF
C6434 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6865_n7304# 0.00fF
C6435 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_7237_n11933# 0.00fF
C6436 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C6437 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.02fF
C6438 a_5653_n2997# a_7040_n3255# 0.01fF
C6439 a_501_n9525# VDD 0.36fF
C6440 a_11101_n11933# a_11164_n13591# 0.00fF
C6441 sky130_fd_sc_hd__clkinv_4_8/A a_10904_n13591# 0.15fF
C6442 a_434_n11933# a_600_n10871# 0.00fF
C6443 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_6012_n4887# 0.01fF
C6444 a_3436_n2167# a_3266_n1597# 0.04fF
C6445 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C6446 a_9517_n3621# a_9517_n2997# 0.05fF
C6447 a_4554_n1597# a_4365_n1909# 0.02fF
C6448 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.08fF
C6449 a_7300_n9783# a_8229_n9525# 0.02fF
C6450 a_2085_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.12fF
C6451 a_1888_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X 0.03fF
C6452 a_8418_n6493# a_8229_n4709# 0.00fF
C6453 a_8162_n6493# a_8328_n4887# 0.00fF
C6454 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.29fF
C6455 a_n787_n12325# a_n688_n12503# 0.49fF
C6456 a_4298_n13021# a_4298_n11933# 0.02fF
C6457 a_10994_n9213# a_10994_n10301# 0.01fF
C6458 a_501_n1909# a_600_n2167# 0.49fF
C6459 a_8418_n14109# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C6460 a_8525_n14109# a_9813_n14109# 0.01fF
C6461 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9706_n14109# 0.03fF
C6462 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C6463 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_7237_n11933# 0.01fF
C6464 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_11101_n9213# 0.02fF
C6465 a_3077_n12325# a_3010_n11933# 0.01fF
C6466 a_4661_n5405# a_4554_n4317# 0.00fF
C6467 a_4554_n5405# a_4661_n4317# 0.00fF
C6468 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_11101_n1597# 0.02fF
C6469 a_9517_n9525# VDD 0.34fF
C6470 a_690_n4317# a_600_n3255# 0.01fF
C6471 a_600_n4887# a_690_n5405# 0.02fF
C6472 a_11101_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.12fF
C6473 a_9450_n13021# a_9616_n13591# 0.04fF
C6474 a_9706_n13021# a_9517_n13413# 0.02fF
C6475 a_9616_n4887# a_10904_n4887# 0.01fF
C6476 a_9876_n4887# a_10805_n4709# 0.02fF
C6477 a_8328_n3799# VDD 0.44fF
C6478 a_8162_n1597# a_9450_n1597# 0.01fF
C6479 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VDD 0.89fF
C6480 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.29fF
C6481 a_1789_n8437# a_1722_n9213# 0.01fF
C6482 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11101_n2685# 0.00fF
C6483 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.06fF
C6484 a_8588_n2167# a_7300_n2167# 0.01fF
C6485 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.03fF
C6486 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_3373_n10301# 0.01fF
C6487 a_8328_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.05fF
C6488 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_7040_n2167# 0.00fF
C6489 a_11164_n3799# a_11101_n4317# 0.01fF
C6490 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_10994_n4317# 0.04fF
C6491 a_3010_n4317# a_4298_n4317# 0.01fF
C6492 sky130_fd_sc_hd__clkinv_1_0/A a_3176_n1079# 0.07fF
C6493 a_5949_n1597# a_5842_n2685# 0.00fF
C6494 a_5842_n1597# a_5949_n2685# 0.00fF
C6495 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_5842_n10301# 0.00fF
C6496 a_6012_n3255# a_7300_n3255# 0.01fF
C6497 a_8229_n11237# a_8162_n10301# 0.00fF
C6498 a_5752_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C6499 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X a_7040_n3255# 0.05fF
C6500 sky130_fd_sc_hd__nand2_4_3/Y a_10805_n8437# 0.02fF
C6501 a_6012_n11415# a_4365_n11237# 0.00fF
C6502 a_5653_n11237# a_4724_n11415# 0.02fF
C6503 a_6874_n6493# a_7130_n6493# 0.19fF
C6504 a_5752_n13591# a_7300_n13591# 0.01fF
C6505 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.02fF
C6506 a_5653_n2997# a_5586_n1597# 0.00fF
C6507 a_5752_n11415# a_4464_n11415# 0.01fF
C6508 a_3077_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.00fF
C6509 a_10904_n10871# a_10805_n11237# 0.01fF
C6510 a_10805_n10613# a_10904_n11415# 0.01fF
C6511 sky130_fd_sc_hd__clkinv_1_0/A a_10994_n1597# 0.01fF
C6512 a_8418_n10301# VDD 0.44fF
C6513 a_9706_n13021# a_9517_n11237# 0.00fF
C6514 a_5653_n10613# a_5653_n12325# 0.00fF
C6515 a_1888_n9783# VDD 0.47fF
C6516 a_3176_n3799# a_3077_n4709# 0.00fF
C6517 a_3077_n3621# a_3176_n4887# 0.00fF
C6518 B Bd_b 0.08fF
C6519 a_10994_n2685# VDD 0.42fF
C6520 a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C6521 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.00fF
C6522 a_10738_n4317# VDD 0.70fF
C6523 a_1978_n10301# a_1888_n9783# 0.01fF
C6524 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9813_n8125# 0.02fF
C6525 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.04fF
C6526 a_8328_n12503# a_8418_n11933# 0.01fF
C6527 a_8162_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C6528 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C6529 a_2085_n5405# a_1888_n3799# 0.00fF
C6530 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.02fF
C6531 a_8525_n8125# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C6532 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.00fF
C6533 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_3436_n2167# 0.03fF
C6534 a_10738_n5405# a_9450_n5405# 0.01fF
C6535 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.02fF
C6536 a_6941_n1909# a_6941_n2997# 0.02fF
C6537 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.06fF
C6538 a_13765_n9213# a_13765_n10301# 0.07fF
C6539 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_11101_n10301# 0.01fF
C6540 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.04fF
C6541 a_600_n11415# a_501_n12325# 0.00fF
C6542 sky130_fd_sc_hd__clkinv_1_0/A a_5653_n821# 0.06fF
C6543 a_9813_n14109# sky130_fd_sc_hd__nand2_4_2/B 0.13fF
C6544 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_860_n13591# 0.00fF
C6545 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.03fF
C6546 sky130_fd_sc_hd__nand2_4_0/A VDD 12.78fF
C6547 a_6874_n4317# a_6941_n3621# 0.01fF
C6548 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VDD 0.83fF
C6549 a_7040_n2167# a_7040_n1079# 0.01fF
C6550 a_10904_n9783# VDD 0.41fF
C6551 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1789_n2997# 0.00fF
C6552 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C6553 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_3010_n2685# 0.03fF
C6554 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_1722_n5405# 0.03fF
C6555 a_690_n9213# a_2085_n9213# 0.01fF
C6556 a_8162_n5405# a_8328_n3799# 0.00fF
C6557 a_8418_n5405# a_8229_n3621# 0.00fF
C6558 a_3176_n10871# a_3010_n9213# 0.00fF
C6559 a_3077_n10613# a_3266_n9213# 0.00fF
C6560 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkinv_1_0/A 0.02fF
C6561 a_4298_n1597# a_4554_n1597# 0.19fF
C6562 a_6874_n1597# a_7130_n1597# 0.19fF
C6563 a_690_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.02fF
C6564 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.02fF
C6565 a_9450_n1597# a_9706_n1597# 0.19fF
C6566 a_4298_n10301# a_4298_n9213# 0.02fF
C6567 a_690_n4317# a_2085_n4317# 0.01fF
C6568 a_797_n4317# a_1978_n4317# 0.01fF
C6569 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_7/Y 0.19fF
C6570 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_7/A 0.68fF
C6571 a_3077_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C6572 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1722_n4317# 0.35fF
C6573 a_8418_n1597# a_8588_n3255# 0.00fF
C6574 a_7040_n9783# a_7130_n9213# 0.02fF
C6575 a_8525_n1597# a_8328_n3255# 0.00fF
C6576 a_5949_n1597# a_5752_n3255# 0.00fF
C6577 a_5842_n1597# a_6012_n3255# 0.00fF
C6578 a_4298_n4317# a_4554_n4317# 0.19fF
C6579 sky130_fd_sc_hd__clkinv_1_0/A a_4724_n1079# 0.12fF
C6580 a_8162_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C6581 a_7300_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.29fF
C6582 a_6874_n6493# a_8525_n6493# 0.00fF
C6583 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.05fF
C6584 a_7237_n6493# a_8162_n6493# 0.02fF
C6585 a_11101_n4317# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C6586 a_7130_n6493# a_8418_n6493# 0.01fF
C6587 a_860_n3799# a_690_n5405# 0.00fF
C6588 Bd_b a_6658_n7363# 0.05fF
C6589 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C6590 a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C6591 a_600_n3799# a_797_n5405# 0.00fF
C6592 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_8588_n1079# 0.03fF
C6593 a_5949_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.01fF
C6594 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6012_n1079# 0.03fF
C6595 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C6596 a_1789_n10613# a_1978_n11933# 0.00fF
C6597 a_1888_n10871# a_1722_n11933# 0.00fF
C6598 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_9813_n13021# 0.01fF
C6599 a_3436_n9783# VDD 0.78fF
C6600 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.06fF
C6601 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.04fF
C6602 a_9450_n2685# a_9616_n1079# 0.00fF
C6603 a_9706_n2685# a_9517_n821# 0.00fF
C6604 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3077_n9525# 0.01fF
C6605 a_9876_n12503# a_9813_n14109# 0.00fF
C6606 a_3010_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C6607 a_9450_n5405# a_9450_n4317# 0.02fF
C6608 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X a_9450_n11933# 0.03fF
C6609 a_5752_n9783# a_5752_n8695# 0.01fF
C6610 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C6611 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_6012_n10871# 0.01fF
C6612 a_8229_n9525# a_8328_n8695# 0.00fF
C6613 a_1789_n2997# a_1888_n3799# 0.01fF
C6614 sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5405# 0.04fF
C6615 a_1888_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C6616 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.06fF
C6617 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.00fF
C6618 sky130_fd_sc_hd__clkinv_1_0/A a_7040_n1079# 0.07fF
C6619 a_4464_n12503# a_4554_n11933# 0.01fF
C6620 a_9813_n1597# a_9876_n3255# 0.00fF
C6621 a_5842_n5405# a_5653_n4709# 0.02fF
C6622 a_6665_n7459# sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C6623 a_5586_n5405# a_5752_n4887# 0.04fF
C6624 a_1888_n2167# VDD 0.47fF
C6625 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.16fF
C6626 a_1722_n4317# a_1888_n3799# 0.04fF
C6627 a_10805_n3621# a_10805_n2997# 0.05fF
C6628 a_n428_n4887# a_860_n4887# 0.01fF
C6629 a_501_n4709# a_600_n4887# 0.49fF
C6630 a_1978_n4317# a_1789_n3621# 0.02fF
C6631 a_600_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.04fF
C6632 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_3266_n9213# 0.00fF
C6633 a_1978_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.05fF
C6634 a_1888_n3255# a_1789_n4709# 0.00fF
C6635 a_6941_n9525# a_6874_n8125# 0.00fF
C6636 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.02fF
C6637 a_4554_n1597# a_5842_n1597# 0.01fF
C6638 a_6874_n1597# a_8525_n1597# 0.00fF
C6639 a_4661_n1597# a_5586_n1597# 0.02fF
C6640 a_4298_n1597# a_5949_n1597# 0.00fF
C6641 a_6012_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C6642 a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C6643 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_10738_n11933# 0.01fF
C6644 a_4623_n7349# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C6645 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_3266_n4317# 0.00fF
C6646 a_3436_n8695# a_3373_n9213# 0.01fF
C6647 a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C6648 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_8162_n9213# 0.03fF
C6649 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_3/Y 0.03fF
C6650 a_9616_n11415# a_9706_n11933# 0.02fF
C6651 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_7130_n509# 0.02fF
C6652 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_7130_n8125# 0.02fF
C6653 a_4724_n2167# VDD 0.78fF
C6654 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X a_11164_n3799# 0.03fF
C6655 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.00fF
C6656 a_8525_n14109# a_8588_n13591# 0.01fF
C6657 a_9616_n4887# a_9616_n5975# 0.01fF
C6658 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X a_10738_n2685# 0.00fF
C6659 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkinv_1_3/Y 0.06fF
C6660 a_9706_n8125# a_9876_n9783# 0.00fF
C6661 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C6662 a_5752_n5975# a_5752_n4887# 0.01fF
C6663 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_9450_n6493# 0.00fF
C6664 a_8162_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.03fF
C6665 a_8418_n6493# a_8525_n6493# 0.55fF
C6666 a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C6667 a_9616_n12503# a_9876_n12503# 0.28fF
C6668 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C6669 a_434_n9213# a_690_n9213# 0.19fF
C6670 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C6671 a_7040_n10871# a_7040_n12503# 0.00fF
C6672 a_2148_n5975# a_2085_n5405# 0.01fF
C6673 a_8162_n4317# a_9450_n4317# 0.01fF
C6674 a_11101_n9213# VDD 0.32fF
C6675 a_434_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.43fF
C6676 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_600_n4887# 0.04fF
C6677 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C6678 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C6679 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_9876_n9783# 0.00fF
C6680 a_3373_n10301# a_3436_n9783# 0.01fF
C6681 a_5653_n11237# a_5752_n11415# 0.49fF
C6682 a_6874_n1597# a_6941_n1909# 0.01fF
C6683 a_8229_n9525# a_8162_n10301# 0.01fF
C6684 a_1789_n13413# a_3077_n13413# 0.01fF
C6685 a_2148_n3255# a_1789_n2997# 0.05fF
C6686 a_3077_n8437# a_3176_n8695# 0.49fF
C6687 a_690_n2685# a_690_n4317# 0.01fF
C6688 a_6012_n13591# a_6941_n13413# 0.02fF
C6689 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_797_n11933# 0.01fF
C6690 a_5949_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.02fF
C6691 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_4661_n9213# 0.01fF
C6692 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C6693 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_5586_n4317# 0.01fF
C6694 a_5949_n9213# a_6874_n9213# 0.02fF
C6695 sky130_fd_sc_hd__clkinv_1_0/A a_8588_n1079# 0.12fF
C6696 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD 0.84fF
C6697 a_6874_n6493# a_6874_n8125# 0.01fF
C6698 a_n787_n9525# a_n688_n9783# 0.49fF
C6699 a_2622_n8125# sky130_fd_sc_hd__clkinv_1_3/A 0.01fF
C6700 a_2622_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.03fF
C6701 a_600_n5975# VDD 0.46fF
C6702 a_8418_n4317# a_8328_n3799# 0.02fF
C6703 a_1978_n13021# a_3010_n13021# 0.02fF
C6704 a_1722_n13021# a_3266_n13021# 0.01fF
C6705 a_3436_n2167# VDD 0.78fF
C6706 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.00fF
C6707 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8525_n9213# 0.00fF
C6708 a_5752_n3799# a_7040_n3799# 0.01fF
C6709 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_860_n9783# 0.01fF
C6710 a_5653_n3621# a_7300_n3799# 0.00fF
C6711 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C6712 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.40fF
C6713 a_2148_n13591# a_2085_n11933# 0.00fF
C6714 a_5842_n1597# a_5949_n1597# 0.55fF
C6715 a_5586_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.03fF
C6716 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_6874_n1597# 0.00fF
C6717 a_9616_n11415# a_9706_n10301# 0.01fF
C6718 a_11164_n10871# a_11101_n11933# 0.00fF
C6719 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C6720 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C6721 a_5842_n10301# a_5842_n9213# 0.01fF
C6722 a_1888_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.01fF
C6723 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.73fF
C6724 a_7237_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.12fF
C6725 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VDD 0.90fF
C6726 a_6941_n2997# a_7040_n4887# 0.00fF
C6727 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C6728 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_6012_n12503# 0.03fF
C6729 a_7040_n3255# a_6941_n4709# 0.00fF
C6730 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_1_4/B 0.14fF
C6731 a_11164_n1079# a_11101_n2685# 0.00fF
C6732 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_10994_n2685# 0.01fF
C6733 a_600_n4887# a_600_n3799# 0.01fF
C6734 a_860_n8695# a_2148_n8695# 0.01fF
C6735 sky130_fd_sc_hd__nand2_4_0/Y a_10904_n1079# 0.16fF
C6736 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_1888_n8695# 0.05fF
C6737 a_9876_n12503# a_11164_n12503# 0.01fF
C6738 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_10904_n12503# 0.05fF
C6739 a_9616_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.00fF
C6740 a_797_n9213# a_1722_n9213# 0.02fF
C6741 a_690_n9213# a_1978_n9213# 0.01fF
C6742 a_7130_n2685# a_6941_n3621# 0.00fF
C6743 a_3436_n10871# a_3266_n11933# 0.00fF
C6744 a_3176_n10871# a_3373_n11933# 0.00fF
C6745 a_6874_n2685# a_7040_n3799# 0.00fF
C6746 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.01fF
C6747 a_3077_n9525# a_3010_n9213# 0.01fF
C6748 sky130_fd_sc_hd__nand2_1_0/A a_n787_n1909# 0.07fF
C6749 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_860_n4887# 0.03fF
C6750 a_797_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C6751 a_1978_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.00fF
C6752 a_4554_n11933# a_4554_n10301# 0.01fF
C6753 a_9706_n509# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C6754 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.02fF
C6755 a_5653_n11237# a_7300_n11415# 0.00fF
C6756 a_6006_n7607# a_6373_n7349# 0.04fF
C6757 a_5052_n7283# a_6658_n7363# 0.00fF
C6758 a_6012_n11415# a_6941_n11237# 0.02fF
C6759 a_5752_n11415# a_7040_n11415# 0.01fF
C6760 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C6761 a_501_n10613# a_434_n9213# 0.00fF
C6762 a_6012_n3799# a_7040_n3799# 0.02fF
C6763 a_3077_n13413# a_3176_n13591# 0.48fF
C6764 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_6941_n3621# 0.18fF
C6765 sky130_fd_sc_hd__clkinv_4_4/A Ad_b 0.31fF
C6766 a_3077_n8437# a_4724_n8695# 0.00fF
C6767 a_3436_n8695# a_4365_n8437# 0.02fF
C6768 a_3176_n8695# a_4464_n8695# 0.01fF
C6769 a_3436_n4887# VDD 0.78fF
C6770 a_1722_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C6771 a_11164_n3799# VDD 0.67fF
C6772 a_7040_n8695# a_5653_n8437# 0.01fF
C6773 a_6941_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.02fF
C6774 a_7040_n13591# a_7300_n13591# 0.28fF
C6775 a_n688_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C6776 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_8229_n13413# 0.01fF
C6777 a_8229_n8437# a_9517_n8437# 0.01fF
C6778 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_8162_n9213# 0.00fF
C6779 a_1888_n5975# a_1978_n4317# 0.00fF
C6780 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/B 0.82fF
C6781 a_6874_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.03fF
C6782 a_7130_n9213# a_7237_n9213# 0.55fF
C6783 sky130_fd_sc_hd__clkinv_4_8/Y a_9876_n13591# 0.00fF
C6784 a_9616_n2167# a_9706_n1597# 0.02fF
C6785 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_3010_n4317# 0.01fF
C6786 a_6006_n7607# VDD 0.52fF
C6787 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_3/Y 0.05fF
C6788 a_3010_n13021# a_3373_n13021# 0.05fF
C6789 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_8418_n11933# 0.01fF
C6790 a_9813_n11933# a_8525_n11933# 0.01fF
C6791 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9517_n3621# 0.01fF
C6792 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9517_n5797# 0.01fF
C6793 a_9450_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.03fF
C6794 sky130_fd_sc_hd__clkinv_1_0/Y a_2366_n509# 0.34fF
C6795 a_1888_n12503# a_1978_n13021# 0.02fF
C6796 a_10738_n5405# a_11101_n5405# 0.05fF
C6797 a_3010_n13021# VDD 0.75fF
C6798 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_10738_n10301# 0.01fF
C6799 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6012_n10871# 0.01fF
C6800 a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C6801 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C6802 a_4724_n12503# a_4661_n13021# 0.01fF
C6803 sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# 0.58fF
C6804 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.02fF
C6805 a_3010_n2685# a_3266_n2685# 0.19fF
C6806 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C6807 p2 sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C6808 a_6012_n12503# VDD 0.77fF
C6809 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.06fF
C6810 a_7130_n10301# a_7130_n11933# 0.01fF
C6811 a_10805_n10613# a_10805_n9525# 0.02fF
C6812 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.02fF
C6813 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.02fF
C6814 a_5752_n8695# a_5949_n9213# 0.02fF
C6815 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.08fF
C6816 a_8328_n8695# a_8418_n9213# 0.01fF
C6817 a_8418_n13021# a_8525_n11933# 0.00fF
C6818 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.33fF
C6819 a_8525_n13021# a_8418_n11933# 0.00fF
C6820 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A a_501_n9525# 0.01fF
C6821 a_1722_n2685# a_1888_n3799# 0.00fF
C6822 a_1978_n2685# a_1789_n3621# 0.00fF
C6823 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.06fF
C6824 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.08fF
C6825 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5586_n10301# 0.00fF
C6826 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_1_3/A 0.73fF
C6827 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.12fF
C6828 a_5586_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C6829 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C6830 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_2085_n11933# 0.01fF
C6831 a_10738_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.01fF
C6832 sky130_fd_sc_hd__clkinv_4_8/Y a_10738_n13789# 0.01fF
C6833 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.05fF
C6834 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C6835 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_7300_n5975# 0.01fF
C6836 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C6837 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_8229_n11237# 0.01fF
C6838 a_7040_n11415# a_7300_n11415# 0.28fF
C6839 a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.02fF
C6840 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C6841 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_9876_n3255# 0.01fF
C6842 a_3077_n13413# a_4724_n13591# 0.00fF
C6843 a_7040_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C6844 a_3176_n13591# a_4464_n13591# 0.01fF
C6845 a_3436_n13591# a_4365_n13413# 0.02fF
C6846 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_8328_n3799# 0.01fF
C6847 a_2729_n509# a_2622_n509# 0.55fF
C6848 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_2366_n509# 0.02fF
C6849 a_9450_n6493# a_9813_n6493# 0.05fF
C6850 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD 0.86fF
C6851 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_5653_n8437# 0.01fF
C6852 a_4464_n8695# a_4724_n8695# 0.28fF
C6853 a_4365_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.02fF
C6854 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_8328_n13591# 0.05fF
C6855 a_7040_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C6856 a_2148_n3799# a_3176_n3799# 0.02fF
C6857 a_600_n3799# a_860_n3799# 0.28fF
C6858 a_501_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.02fF
C6859 a_7300_n13591# a_8588_n13591# 0.01fF
C6860 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_3077_n3621# 0.18fF
C6861 a_2366_n14109# VDD 0.77fF
C6862 a_1789_n11237# a_1888_n11415# 0.49fF
C6863 a_9517_n8437# a_9616_n8695# 0.49fF
C6864 a_1722_n1597# a_1789_n821# 0.01fF
C6865 a_7130_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C6866 a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C6867 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_3010_n4317# 0.00fF
C6868 a_7237_n9213# a_8525_n9213# 0.01fF
C6869 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8418_n9213# 0.03fF
C6870 a_3176_n2167# a_3176_n3799# 0.00fF
C6871 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_4724_n3255# 0.01fF
C6872 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C6873 a_501_n821# VDD 0.36fF
C6874 sky130_fd_sc_hd__clkinv_4_3/Y VDD 3.76fF
C6875 sky130_fd_sc_hd__nand2_4_3/Y a_10738_n9213# 0.08fF
C6876 a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C6877 a_8418_n6493# a_8418_n8125# 0.00fF
C6878 a_10904_n11415# a_10994_n13021# 0.00fF
C6879 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4298_n13021# 0.35fF
C6880 a_3266_n13021# a_4661_n13021# 0.01fF
C6881 a_3373_n13021# a_4554_n13021# 0.01fF
C6882 a_4724_n10871# a_3077_n10613# 0.00fF
C6883 a_4464_n10871# a_3176_n10871# 0.01fF
C6884 a_8229_n12325# a_8229_n13413# 0.02fF
C6885 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.08fF
C6886 a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C6887 a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C6888 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_3010_n13021# 0.03fF
C6889 a_5752_n9783# a_5653_n11237# 0.00fF
C6890 a_5653_n9525# a_5752_n11415# 0.00fF
C6891 a_6941_n8437# a_7040_n8695# 0.49fF
C6892 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.00fF
C6893 a_4554_n13021# VDD 0.47fF
C6894 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_9876_n13591# 0.01fF
C6895 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C6896 a_860_n12503# a_1888_n12503# 0.02fF
C6897 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_1789_n12325# 0.18fF
C6898 a_600_n12503# a_2148_n12503# 0.01fF
C6899 a_11164_n11415# a_11101_n10301# 0.00fF
C6900 a_4464_n9783# a_4554_n10301# 0.01fF
C6901 a_8229_n8437# a_8162_n8125# 0.01fF
C6902 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C6903 a_1888_n12503# VDD 0.44fF
C6904 a_3266_n2685# a_4554_n2685# 0.01fF
C6905 a_4623_n7349# sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C6906 a_3373_n2685# a_4298_n2685# 0.02fF
C6907 a_3010_n2685# a_4661_n2685# 0.00fF
C6908 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C6909 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_4724_n12503# 0.03fF
C6910 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VDD 0.86fF
C6911 a_8162_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C6912 a_8418_n2685# a_9450_n2685# 0.02fF
C6913 a_8162_n2685# a_9706_n2685# 0.01fF
C6914 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n11933# 0.00fF
C6915 a_8162_n13021# a_8162_n14109# 0.02fF
C6916 a_1888_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C6917 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_9450_n9213# 0.03fF
C6918 a_3010_n10301# VDD 0.76fF
C6919 a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C6920 a_2366_n14109# a_2729_n14109# 0.05fF
C6921 a_8328_n9783# a_9876_n9783# 0.01fF
C6922 a_8588_n9783# a_9616_n9783# 0.02fF
C6923 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_9517_n9525# 0.18fF
C6924 a_8229_n11237# a_8229_n12325# 0.02fF
C6925 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C6926 a_600_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C6927 a_8525_n2685# a_8328_n3799# 0.00fF
C6928 a_8418_n2685# a_8588_n3799# 0.00fF
C6929 a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C6930 a_1722_n10301# a_3266_n10301# 0.01fF
C6931 a_1978_n10301# a_3010_n10301# 0.02fF
C6932 a_8588_n4887# a_8588_n3255# 0.01fF
C6933 a_8229_n1909# a_8162_n2685# 0.01fF
C6934 a_7130_n509# a_7130_n1597# 0.01fF
C6935 a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.18fF
C6936 a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C6937 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_10805_n5797# 0.01fF
C6938 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.02fF
C6939 a_9616_n5975# a_9876_n5975# 0.28fF
C6940 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.02fF
C6941 a_4464_n11415# a_4365_n10613# 0.01fF
C6942 a_7040_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C6943 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.02fF
C6944 a_7300_n11415# a_8588_n11415# 0.01fF
C6945 sky130_fd_sc_hd__clkinv_1_5/A a_7300_n5975# 0.00fF
C6946 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.08fF
C6947 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_8328_n11415# 0.05fF
C6948 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_5653_n13413# 0.01fF
C6949 a_6874_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.03fF
C6950 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C6951 a_4464_n13591# a_4724_n13591# 0.28fF
C6952 a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.02fF
C6953 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X a_8588_n3799# 0.03fF
C6954 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6941_n4709# 0.01fF
C6955 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_2366_n14109# 0.00fF
C6956 a_4724_n8695# a_6012_n8695# 0.01fF
C6957 a_4464_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.00fF
C6958 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X a_5752_n8695# 0.05fF
C6959 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.29fF
C6960 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_4464_n3799# 0.01fF
C6961 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X a_1888_n3799# 0.05fF
C6962 a_7130_n14109# VDD 0.44fF
C6963 a_2148_n11415# a_3077_n11237# 0.02fF
C6964 a_1789_n11237# a_3436_n11415# 0.00fF
C6965 a_1888_n11415# a_3176_n11415# 0.01fF
C6966 a_8525_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.12fF
C6967 a_9450_n4317# a_9813_n4317# 0.05fF
C6968 a_3436_n5975# a_3373_n4317# 0.00fF
C6969 a_10805_n10613# a_10994_n9213# 0.00fF
C6970 a_10904_n10871# a_10738_n9213# 0.00fF
C6971 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.07fF
C6972 a_10805_n12325# a_10805_n11237# 0.02fF
C6973 a_9517_n821# VDD 0.34fF
C6974 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_10738_n13789# 0.00fF
C6975 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n8125# 0.00fF
C6976 a_9450_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C6977 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.15fF
C6978 a_11101_n5405# a_10994_n4317# 0.00fF
C6979 a_10738_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.08fF
C6980 a_4554_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.05fF
C6981 a_10994_n5405# a_11101_n4317# 0.00fF
C6982 a_6941_n8437# a_6874_n10301# 0.00fF
C6983 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_4365_n10613# 0.02fF
C6984 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_10738_n2685# 0.00fF
C6985 a_11164_n8695# a_11101_n10301# 0.00fF
C6986 a_6941_n8437# a_8588_n8695# 0.00fF
C6987 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_10994_n10301# 0.01fF
C6988 a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.01fF
C6989 a_3436_n12503# a_3373_n13021# 0.01fF
C6990 a_9706_n2685# a_9706_n4317# 0.01fF
C6991 a_5752_n10871# a_5842_n10301# 0.02fF
C6992 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_3176_n12503# 0.01fF
C6993 a_8162_n13021# a_9813_n13021# 0.00fF
C6994 a_7130_n10301# a_8525_n10301# 0.01fF
C6995 a_1888_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.03fF
C6996 a_501_n8437# a_501_n9525# 0.02fF
C6997 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_8525_n10301# 0.00fF
C6998 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C6999 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_5586_n10301# 0.03fF
C7000 a_3436_n12503# VDD 0.78fF
C7001 a_4554_n2685# a_4661_n2685# 0.55fF
C7002 a_4298_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C7003 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_5586_n2685# 0.00fF
C7004 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C7005 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_9876_n3255# 0.00fF
C7006 sky130_fd_sc_hd__dfxbp_1_0/Q p2 0.00fF
C7007 a_9450_n2685# a_9813_n2685# 0.05fF
C7008 a_4365_n2997# a_4298_n2685# 0.01fF
C7009 a_2085_n5405# a_3373_n5405# 0.01fF
C7010 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3266_n5405# 0.03fF
C7011 a_1888_n2167# a_1888_n3255# 0.01fF
C7012 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6874_n14109# 0.32fF
C7013 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.01fF
C7014 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_10904_n9783# 0.01fF
C7015 a_9616_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.03fF
C7016 a_860_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C7017 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X a_2148_n9783# 0.03fF
C7018 a_6874_n8125# a_8162_n8125# 0.01fF
C7019 a_3010_n10301# a_3373_n10301# 0.05fF
C7020 a_8162_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C7021 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8162_n1597# 0.01fF
C7022 a_9706_n8125# VDD 0.48fF
C7023 a_9876_n5975# a_11164_n5975# 0.01fF
C7024 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_10904_n5975# 0.05fF
C7025 a_10738_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.02fF
C7026 a_5949_n4317# a_5752_n4887# 0.02fF
C7027 a_5842_n4317# a_6012_n4887# 0.04fF
C7028 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.06fF
C7029 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.02fF
C7030 a_9616_n2167# a_9876_n2167# 0.28fF
C7031 a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C7032 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.05fF
C7033 a_8418_n8125# a_8525_n9213# 0.00fF
C7034 a_8525_n8125# a_8418_n9213# 0.00fF
C7035 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.29fF
C7036 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C7037 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_5752_n13591# 0.05fF
C7038 a_6012_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.29fF
C7039 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C7040 a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.02fF
C7041 a_3176_n11415# a_3436_n11415# 0.28fF
C7042 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_4365_n11237# 0.01fF
C7043 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD 0.79fF
C7044 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10738_n4317# 0.35fF
C7045 sky130_fd_sc_hd__nand2_4_3/B a_10805_n8437# 0.03fF
C7046 a_9706_n4317# a_11101_n4317# 0.01fF
C7047 a_9813_n4317# a_10994_n4317# 0.01fF
C7048 sky130_fd_sc_hd__clkinv_4_8/A a_9450_n14109# 0.01fF
C7049 a_600_n10871# a_797_n10301# 0.02fF
C7050 a_860_n10871# a_690_n10301# 0.04fF
C7051 a_10904_n1079# VDD 0.41fF
C7052 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_860_n3255# 0.00fF
C7053 a_4623_n7349# a_4765_n7542# 0.01fF
C7054 a_797_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C7055 a_9616_n9783# a_9450_n10301# 0.04fF
C7056 a_9517_n9525# a_9706_n10301# 0.02fF
C7057 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X a_600_n9783# 0.01fF
C7058 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_9706_n6493# 0.00fF
C7059 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.03fF
C7060 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_7237_n5405# 0.01fF
C7061 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_690_n5405# 0.01fF
C7062 a_2085_n5405# a_797_n5405# 0.01fF
C7063 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10994_n2685# 0.03fF
C7064 a_9813_n2685# a_11101_n2685# 0.01fF
C7065 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.04fF
C7066 a_7130_n509# a_6941_n1909# 0.00fF
C7067 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n4317# 0.00fF
C7068 a_6874_n509# a_7040_n2167# 0.00fF
C7069 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_9706_n10301# 0.00fF
C7070 a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C7071 a_9706_n509# VDD 0.48fF
C7072 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_6874_n10301# 0.03fF
C7073 a_9706_n13021# a_9813_n13021# 0.55fF
C7074 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_3436_n12503# 0.03fF
C7075 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.00fF
C7076 a_9450_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C7077 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_10738_n13021# 0.00fF
C7078 a_4554_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C7079 a_4661_n2685# a_5949_n2685# 0.01fF
C7080 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5842_n2685# 0.03fF
C7081 a_1722_n1597# a_3266_n1597# 0.01fF
C7082 a_1978_n1597# a_3010_n1597# 0.02fF
C7083 a_n787_n1909# a_n428_n2167# 0.05fF
C7084 a_9706_n13021# a_9706_n14109# 0.01fF
C7085 a_8229_n1909# sky130_fd_sc_hd__nand2_4_0/Y 0.08fF
C7086 a_10738_n6173# a_10805_n4709# 0.01fF
C7087 a_3373_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.12fF
C7088 a_5653_n9525# a_5752_n9783# 0.49fF
C7089 a_13765_n1597# a_13765_n1053# 0.31fF
C7090 a_8418_n10301# a_9706_n10301# 0.01fF
C7091 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X a_11164_n9783# 0.03fF
C7092 a_2148_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C7093 a_8162_n8125# a_8418_n8125# 0.19fF
C7094 a_8525_n509# a_8525_n1597# 0.02fF
C7095 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VDD 0.72fF
C7096 a_10738_n8125# a_11164_n9783# 0.01fF
C7097 a_4365_n2997# a_4365_n1909# 0.02fF
C7098 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_4/Y 0.13fF
C7099 a_9517_n821# a_9876_n1079# 0.05fF
C7100 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C7101 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__clkinv_4_3/Y 0.06fF
C7102 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_10904_n2167# 0.05fF
C7103 sky130_fd_sc_hd__clkinv_4_8/A a_11101_n13021# 0.10fF
C7104 a_9876_n2167# a_11164_n2167# 0.01fF
C7105 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_860_n10871# 0.00fF
C7106 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.00fF
C7107 a_10738_n9213# a_9450_n9213# 0.01fF
C7108 a_4724_n3799# a_4724_n4887# 0.02fF
C7109 a_600_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.03fF
C7110 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_690_n5405# 0.02fF
C7111 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VDD 0.90fF
C7112 sky130_fd_sc_hd__clkinv_1_5/A a_6865_n7304# 0.03fF
C7113 a_11101_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.12fF
C7114 a_8229_n4709# a_8328_n4887# 0.49fF
C7115 sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2685# 0.04fF
C7116 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C7117 a_3436_n11415# a_4724_n11415# 0.01fF
C7118 a_3176_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C7119 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_4464_n11415# 0.05fF
C7120 a_4464_n5975# a_4464_n4887# 0.01fF
C7121 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C7122 a_10994_n4317# sky130_fd_sc_hd__clkinv_4_3/A 0.01fF
C7123 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.02fF
C7124 a_8229_n10613# a_8328_n9783# 0.00fF
C7125 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A VDD 0.87fF
C7126 a_9517_n11237# a_10904_n11415# 0.01fF
C7127 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9876_n9783# 0.03fF
C7128 a_9450_n13021# a_9616_n12503# 0.04fF
C7129 a_9706_n13021# a_9517_n12325# 0.02fF
C7130 a_9813_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C7131 a_5653_n3621# VDD 0.35fF
C7132 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C7133 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_5949_n11933# 0.00fF
C7134 a_7300_n10871# a_7237_n10301# 0.01fF
C7135 a_6874_n6493# a_6941_n4709# 0.00fF
C7136 a_5949_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.12fF
C7137 a_4365_n2997# a_5752_n3255# 0.01fF
C7138 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_797_n2685# 0.00fF
C7139 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.00fF
C7140 a_2148_n2167# a_1978_n1597# 0.04fF
C7141 a_11101_n5405# sky130_fd_sc_hd__clkinv_4_4/Y 0.01fF
C7142 a_1888_n2167# a_2085_n1597# 0.02fF
C7143 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.02fF
C7144 a_8229_n3621# a_8229_n2997# 0.05fF
C7145 a_2148_n4887# VDD 0.78fF
C7146 a_5653_n9525# a_7300_n9783# 0.00fF
C7147 a_6012_n9783# a_6941_n9525# 0.02fF
C7148 a_5752_n9783# a_7040_n9783# 0.01fF
C7149 a_6658_n7363# sky130_fd_sc_hd__nand2_4_3/A 0.11fF
C7150 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6794_n7203# 0.00fF
C7151 a_6794_n7203# a_7212_n7203# 0.03fF
C7152 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C7153 a_1888_n8695# a_2085_n9213# 0.02fF
C7154 a_8525_n8125# a_9450_n8125# 0.02fF
C7155 a_3010_n13021# a_3010_n11933# 0.02fF
C7156 a_4724_n9783# a_3176_n9783# 0.01fF
C7157 a_4464_n9783# a_3436_n9783# 0.02fF
C7158 a_8162_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C7159 a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.18fF
C7160 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C7161 a_1722_n2685# a_3010_n2685# 0.01fF
C7162 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.03fF
C7163 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_5949_n11933# 0.01fF
C7164 a_5653_n1909# a_5586_n2685# 0.01fF
C7165 a_1789_n12325# a_1722_n11933# 0.01fF
C7166 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7300_n2167# 0.03fF
C7167 a_10994_n11933# a_11164_n12503# 0.04fF
C7168 a_3266_n5405# a_3373_n4317# 0.00fF
C7169 a_9616_n1079# a_11164_n1079# 0.01fF
C7170 a_11101_n11933# a_10904_n12503# 0.02fF
C7171 sky130_fd_sc_hd__clkinv_4_8/A a_10805_n12325# 0.07fF
C7172 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C7173 a_3373_n5405# a_3266_n4317# 0.00fF
C7174 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X a_10805_n821# 0.17fF
C7175 a_9876_n1079# a_10904_n1079# 0.02fF
C7176 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C7177 a_797_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.12fF
C7178 a_8418_n13021# a_8229_n13413# 0.02fF
C7179 a_8162_n13021# a_8328_n13591# 0.04fF
C7180 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.09fF
C7181 a_8328_n4887# a_9616_n4887# 0.01fF
C7182 a_8229_n4709# a_9876_n4887# 0.00fF
C7183 a_3176_n2167# a_3176_n1079# 0.01fF
C7184 a_8588_n4887# a_9517_n4709# 0.02fF
C7185 a_860_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.11fF
C7186 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.29fF
C7187 a_9813_n509# a_9616_n1079# 0.02fF
C7188 a_9706_n509# a_9876_n1079# 0.04fF
C7189 a_501_n821# a_600_n1079# 0.49fF
C7190 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VDD 0.89fF
C7191 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.02fF
C7192 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.06fF
C7193 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C7194 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_2085_n10301# 0.01fF
C7195 a_9876_n3799# a_9813_n4317# 0.01fF
C7196 Ad_b a_6665_n7459# 0.07fF
C7197 a_1722_n4317# a_3010_n4317# 0.01fF
C7198 a_10904_n9783# a_11101_n10301# 0.02fF
C7199 a_11164_n9783# a_10994_n10301# 0.04fF
C7200 a_6941_n11237# a_6874_n10301# 0.00fF
C7201 a_11101_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.00fF
C7202 a_4661_n1597# a_4554_n2685# 0.00fF
C7203 a_4554_n1597# a_4661_n2685# 0.00fF
C7204 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_4554_n10301# 0.00fF
C7205 a_9616_n3255# a_9517_n3621# 0.01fF
C7206 a_4554_n4317# a_4661_n2685# 0.00fF
C7207 a_4661_n4317# a_4554_n2685# 0.00fF
C7208 a_4365_n2997# a_4298_n1597# 0.00fF
C7209 a_4464_n13591# a_6012_n13591# 0.01fF
C7210 a_9517_n10613# a_9616_n11415# 0.01fF
C7211 a_5949_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C7212 a_9813_n2685# a_9876_n3799# 0.00fF
C7213 a_4365_n2997# a_4298_n4317# 0.00fF
C7214 a_1789_n821# VDD 0.36fF
C7215 a_501_n2997# a_501_n4709# 0.00fF
C7216 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6012_n3255# 0.03fF
C7217 a_5653_n2997# a_6012_n3255# 0.05fF
C7218 a_8162_n13021# a_8328_n11415# 0.00fF
C7219 a_8418_n13021# a_8229_n11237# 0.00fF
C7220 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C7221 a_9813_n11933# a_9616_n13591# 0.00fF
C7222 a_2085_n4317# a_1978_n5405# 0.00fF
C7223 a_9706_n6493# a_9813_n6493# 0.55fF
C7224 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C7225 a_690_n10301# a_600_n9783# 0.01fF
C7226 a_7040_n12503# a_7130_n11933# 0.01fF
C7227 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_8229_n9525# 0.01fF
C7228 a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.02fF
C7229 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C7230 a_7040_n9783# a_7300_n9783# 0.28fF
C7231 a_2366_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C7232 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A p2 0.02fF
C7233 a_5586_n13021# a_5752_n11415# 0.00fF
C7234 a_10994_n5405# VDD 0.43fF
C7235 a_13765_n8669# p2 2.54fF
C7236 a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C7237 a_10738_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C7238 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.06fF
C7239 a_690_n13021# a_1722_n13021# 0.02fF
C7240 a_434_n13021# a_1978_n13021# 0.01fF
C7241 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10738_n10301# 0.01fF
C7242 a_10994_n2685# a_10805_n2997# 0.02fF
C7243 a_8525_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.12fF
C7244 a_10738_n2685# a_10904_n3255# 0.04fF
C7245 a_8162_n2685# VDD 0.76fF
C7246 a_10738_n4317# a_10805_n2997# 0.00fF
C7247 a_10904_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.02fF
C7248 sky130_fd_sc_hd__clkinv_4_8/A p1d 0.01fF
C7249 a_8328_n9783# VDD 0.46fF
C7250 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_5586_n11933# 0.03fF
C7251 a_501_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.01fF
C7252 a_5752_n2167# a_5752_n1079# 0.01fF
C7253 a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C7254 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_501_n2997# 0.00fF
C7255 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C7256 a_9450_n509# a_10738_n509# 0.01fF
C7257 a_7130_n5405# a_6941_n3621# 0.00fF
C7258 a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C7259 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_10805_n4709# 0.01fF
C7260 a_9616_n4887# a_9876_n4887# 0.28fF
C7261 a_6874_n5405# a_7040_n3799# 0.00fF
C7262 a_3010_n10301# a_3010_n11933# 0.01fF
C7263 a_7300_n3799# VDD 0.77fF
C7264 sky130_fd_sc_hd__nand2_4_0/B a_10904_n1079# 0.02fF
C7265 a_8162_n1597# a_8418_n1597# 0.19fF
C7266 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_9813_n4317# 0.01fF
C7267 a_7237_n1597# a_7040_n3255# 0.00fF
C7268 a_3010_n4317# a_3266_n4317# 0.19fF
C7269 a_7130_n1597# a_7300_n3255# 0.00fF
C7270 a_1789_n8437# a_3176_n8695# 0.01fF
C7271 a_1888_n8695# a_3077_n8437# 0.01fF
C7272 sky130_fd_sc_hd__clkinv_1_0/A a_2148_n1079# 0.12fF
C7273 a_13765_n9757# p2d_b 0.12fF
C7274 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.02fF
C7275 a_3373_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C7276 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4661_n10301# 0.02fF
C7277 a_9706_n509# sky130_fd_sc_hd__nand2_4_0/B 0.05fF
C7278 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C7279 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.29fF
C7280 a_2148_n1079# a_2085_n2685# 0.00fF
C7281 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.02fF
C7282 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_7040_n13591# 0.01fF
C7283 a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C7284 a_4623_n7349# a_4724_n8695# 0.01fF
C7285 a_5752_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.03fF
C7286 sky130_fd_sc_hd__dfxbp_1_0/Q a_4464_n8695# 0.00fF
C7287 a_7237_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C7288 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7300_n1079# 0.03fF
C7289 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C7290 a_860_n9783# VDD 0.78fF
C7291 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_3/Y 0.64fF
C7292 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_3/A 0.19fF
C7293 a_690_n11933# a_860_n10871# 0.00fF
C7294 a_797_n11933# a_600_n10871# 0.00fF
C7295 a_690_n1597# a_501_n821# 0.02fF
C7296 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_434_n5405# 0.00fF
C7297 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.04fF
C7298 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_8162_n11933# 0.03fF
C7299 a_1722_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C7300 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1789_n9525# 0.01fF
C7301 a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C7302 a_9706_n4317# VDD 0.46fF
C7303 a_7130_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C7304 a_6941_n9525# a_7040_n8695# 0.00fF
C7305 a_8525_n6493# a_8328_n4887# 0.00fF
C7306 a_8418_n6493# a_8588_n4887# 0.00fF
C7307 a_n787_n12325# a_501_n12325# 0.01fF
C7308 a_n688_n12503# a_n428_n12503# 0.28fF
C7309 a_600_n3255# a_501_n3621# 0.01fF
C7310 a_501_n2997# a_600_n3799# 0.01fF
C7311 a_600_n2167# a_860_n2167# 0.28fF
C7312 a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X 0.02fF
C7313 a_11101_n9213# a_11101_n10301# 0.02fF
C7314 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__nand2_4_0/A 0.08fF
C7315 a_4554_n13021# a_4554_n11933# 0.01fF
C7316 a_1722_n1597# VDD 0.76fF
C7317 a_10738_n6173# a_10904_n5975# 0.03fF
C7318 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C7319 a_9706_n2685# VDD 0.43fF
C7320 a_4298_n5405# a_4464_n4887# 0.04fF
C7321 a_600_n12503# a_690_n13021# 0.02fF
C7322 a_3176_n12503# a_3266_n11933# 0.01fF
C7323 a_5586_n11933# VDD 0.76fF
C7324 a_4554_n5405# a_4365_n4709# 0.02fF
C7325 a_434_n13021# VDD 0.76fF
C7326 a_9876_n9783# VDD 0.74fF
C7327 a_860_n4887# a_797_n5405# 0.01fF
C7328 a_797_n4317# a_860_n3255# 0.00fF
C7329 a_9706_n13021# a_9876_n13591# 0.04fF
C7330 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_10904_n4887# 0.05fF
C7331 a_3373_n1597# a_4298_n1597# 0.02fF
C7332 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VDD 0.83fF
C7333 a_5842_n1597# a_7130_n1597# 0.01fF
C7334 a_8418_n1597# a_9706_n1597# 0.01fF
C7335 a_5586_n1597# a_7237_n1597# 0.00fF
C7336 a_8525_n1597# a_9450_n1597# 0.02fF
C7337 a_8162_n1597# a_9813_n1597# 0.00fF
C7338 a_10738_n509# a_10994_n1597# 0.01fF
C7339 a_8229_n1909# VDD 0.35fF
C7340 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.04fF
C7341 a_1888_n8695# a_1978_n9213# 0.01fF
C7342 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_1978_n4317# 0.00fF
C7343 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C7344 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A sky130_fd_sc_hd__clkinv_4_3/A 0.01fF
C7345 a_3010_n4317# a_4661_n4317# 0.00fF
C7346 a_3266_n4317# a_4554_n4317# 0.01fF
C7347 a_3373_n4317# a_4298_n4317# 0.02fF
C7348 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6874_n9213# 0.03fF
C7349 a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C7350 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.84fF
C7351 a_4365_n3621# a_5752_n3799# 0.01fF
C7352 a_4464_n3799# a_5653_n3621# 0.01fF
C7353 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X p2 0.02fF
C7354 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkinv_1_3/A 0.11fF
C7355 a_n860_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C7356 a_n688_n2167# VDD 0.51fF
C7357 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C7358 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_8162_n6493# 0.00fF
C7359 a_6012_n11415# a_4724_n11415# 0.01fF
C7360 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C7361 sky130_fd_sc_hd__dfxbp_1_0/Q a_6012_n8695# 0.01fF
C7362 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y 1.21fF
C7363 sky130_fd_sc_hd__nand2_4_3/Y a_11164_n8695# 0.12fF
C7364 a_5752_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.05fF
C7365 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_4464_n11415# 0.00fF
C7366 a_7130_n6493# a_7237_n6493# 0.55fF
C7367 a_6874_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.03fF
C7368 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VDD 0.90fF
C7369 a_2729_n509# sky130_fd_sc_hd__clkinv_1_0/Y 0.02fF
C7370 a_5752_n10871# a_5752_n12503# 0.00fF
C7371 a_13765_n2685# VDD 2.20fF
C7372 a_5586_n1597# a_5653_n1909# 0.01fF
C7373 a_8588_n12503# a_8525_n11933# 0.01fF
C7374 a_2085_n10301# a_2148_n9783# 0.01fF
C7375 a_11101_n4317# VDD 0.32fF
C7376 sky130_fd_sc_hd__nand2_4_0/Y VDD 7.70fF
C7377 a_8525_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C7378 a_6941_n9525# a_6874_n10301# 0.01fF
C7379 sky130_fd_sc_hd__nand2_4_3/B a_10738_n9213# 0.01fF
C7380 a_n1738_n6671# a_n1139_n6715# 0.04fF
C7381 a_11101_n5405# a_9450_n5405# 0.00fF
C7382 a_10994_n5405# a_9706_n5405# 0.01fF
C7383 a_3077_n5797# a_3176_n4887# 0.00fF
C7384 a_3176_n5975# a_3077_n4709# 0.00fF
C7385 a_7040_n2167# a_7040_n3255# 0.01fF
C7386 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_5586_n11933# 0.01fF
C7387 sky130_fd_sc_hd__nand2_4_3/Y Ad_b 0.00fF
C7388 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.04fF
C7389 a_3266_n1597# VDD 0.45fF
C7390 sky130_fd_sc_hd__clkinv_1_0/A a_6012_n1079# 0.12fF
C7391 a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C7392 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X p2 0.03fF
C7393 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_4298_n11933# 0.03fF
C7394 a_13765_n9757# VDD 2.19fF
C7395 a_7130_n4317# a_7040_n3799# 0.02fF
C7396 a_7300_n2167# a_7300_n1079# 0.02fF
C7397 a_4365_n3621# a_6012_n3799# 0.00fF
C7398 a_8418_n5405# a_8588_n3799# 0.00fF
C7399 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_2085_n9213# 0.02fF
C7400 a_797_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C7401 a_3176_n10871# a_3373_n9213# 0.00fF
C7402 a_3436_n10871# a_3266_n9213# 0.00fF
C7403 a_8525_n5405# a_8328_n3799# 0.00fF
C7404 a_2148_n3255# a_3077_n2997# 0.02fF
C7405 a_4298_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C7406 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_5586_n1597# 0.00fF
C7407 a_4554_n1597# a_4661_n1597# 0.55fF
C7408 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C7409 a_9450_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C7410 a_9706_n1597# a_9813_n1597# 0.55fF
C7411 a_6874_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C7412 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_8162_n1597# 0.00fF
C7413 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.02fF
C7414 a_9876_n10871# a_9813_n11933# 0.00fF
C7415 a_4554_n10301# a_4554_n9213# 0.01fF
C7416 a_434_n13021# a_501_n13413# 0.01fF
C7417 a_2366_n8125# a_2148_n9783# 0.00fF
C7418 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_2085_n4317# 0.02fF
C7419 a_797_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C7420 a_8525_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C7421 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6012_n3255# 0.00fF
C7422 a_4554_n4317# a_4661_n4317# 0.55fF
C7423 a_4298_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C7424 a_5949_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C7425 a_2729_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.12fF
C7426 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_8588_n3255# 0.00fF
C7427 a_7300_n9783# a_7237_n9213# 0.01fF
C7428 a_5752_n3255# a_5653_n4709# 0.00fF
C7429 a_7130_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C7430 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8418_n6493# 0.03fF
C7431 a_600_n5975# a_434_n4317# 0.00fF
C7432 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X a_797_n5405# 0.00fF
C7433 a_860_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C7434 a_501_n5797# a_690_n4317# 0.00fF
C7435 a_7237_n6493# a_8525_n6493# 0.01fF
C7436 a_2148_n10871# a_1978_n11933# 0.00fF
C7437 a_1789_n10613# a_1722_n9213# 0.00fF
C7438 a_10738_n10301# VDD 0.70fF
C7439 a_1888_n10871# a_2085_n11933# 0.00fF
C7440 a_8229_n12325# a_8418_n14109# 0.00fF
C7441 a_8328_n12503# a_8162_n14109# 0.00fF
C7442 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VDD 0.84fF
C7443 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_n428_n4887# 0.27fF
C7444 a_9706_n2685# a_9876_n1079# 0.00fF
C7445 a_9813_n2685# a_9616_n1079# 0.00fF
C7446 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C7447 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.05fF
C7448 a_9706_n5405# a_9706_n4317# 0.01fF
C7449 a_2148_n3255# a_600_n3255# 0.01fF
C7450 a_1789_n13413# a_1888_n13591# 0.48fF
C7451 a_6012_n9783# a_6012_n8695# 0.02fF
C7452 a_434_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.00fF
C7453 a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C7454 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.84fF
C7455 a_5842_n5405# a_6012_n4887# 0.04fF
C7456 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VDD 0.90fF
C7457 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8229_n3621# 0.01fF
C7458 a_8162_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C7459 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.02fF
C7460 a_1722_n13021# a_2085_n13021# 0.05fF
C7461 a_10904_n3799# a_10904_n3255# 0.07fF
C7462 a_2085_n4317# a_1888_n3799# 0.02fF
C7463 a_600_n4887# a_860_n4887# 0.28fF
C7464 a_501_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.02fF
C7465 a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.02fF
C7466 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_6941_n3621# 0.01fF
C7467 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C7468 a_5752_n3799# a_6012_n3799# 0.28fF
C7469 a_4365_n12325# a_4365_n11237# 0.02fF
C7470 a_7040_n9783# a_7130_n8125# 0.00fF
C7471 a_4661_n1597# a_5949_n1597# 0.01fF
C7472 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5842_n1597# 0.03fF
C7473 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_4365_n2997# 0.01fF
C7474 a_4554_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C7475 a_10738_n11933# a_10994_n11933# 0.19fF
C7476 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.04fF
C7477 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5586_n9213# 0.01fF
C7478 a_5586_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C7479 a_10994_n1597# a_10805_n821# 0.02fF
C7480 a_10738_n1597# a_10904_n1079# 0.04fF
C7481 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.06fF
C7482 a_9517_n10613# a_9517_n9525# 0.02fF
C7483 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C7484 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C7485 a_5842_n10301# a_5842_n11933# 0.01fF
C7486 a_7040_n8695# a_7130_n9213# 0.01fF
C7487 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A p2 0.05fF
C7488 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.08fF
C7489 a_9876_n4887# a_9876_n5975# 0.02fF
C7490 a_600_n1079# a_1789_n821# 0.01fF
C7491 sky130_fd_sc_hd__nand2_4_3/Y a_9517_n9525# 0.08fF
C7492 a_8525_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.12fF
C7493 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.29fF
C7494 a_6012_n5975# a_6012_n4887# 0.02fF
C7495 a_7237_n13021# a_7130_n11933# 0.00fF
C7496 a_7130_n13021# a_7237_n11933# 0.00fF
C7497 a_4464_n12503# a_4464_n10871# 0.00fF
C7498 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_1722_n9213# 0.00fF
C7499 a_434_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.03fF
C7500 a_690_n9213# a_797_n9213# 0.55fF
C7501 a_8229_n10613# VDD 0.35fF
C7502 p2d_b VDD 4.28fF
C7503 a_434_n2685# a_600_n3799# 0.00fF
C7504 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.06fF
C7505 a_8525_n4317# a_9450_n4317# 0.02fF
C7506 a_7300_n10871# a_7300_n12503# 0.01fF
C7507 a_434_n13021# a_434_n11933# 0.02fF
C7508 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.06fF
C7509 a_8418_n4317# a_9706_n4317# 0.01fF
C7510 a_8162_n4317# a_9813_n4317# 0.00fF
C7511 a_690_n2685# a_501_n3621# 0.00fF
C7512 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4298_n10301# 0.00fF
C7513 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C7514 a_797_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C7515 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.06fF
C7516 a_5752_n11415# a_6012_n11415# 0.28fF
C7517 a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.02fF
C7518 a_9450_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.08fF
C7519 a_2148_n13591# a_3077_n13413# 0.02fF
C7520 a_501_n1909# a_600_n3255# 0.00fF
C7521 a_600_n2167# a_501_n2997# 0.00fF
C7522 a_1888_n13591# a_3176_n13591# 0.01fF
C7523 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VDD 0.79fF
C7524 a_3176_n8695# a_3436_n8695# 0.28fF
C7525 a_3077_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.02fF
C7526 a_4623_n7349# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C7527 a_1789_n13413# a_3436_n13591# 0.00fF
C7528 a_797_n2685# a_797_n4317# 0.01fF
C7529 a_6012_n13591# a_7300_n13591# 0.01fF
C7530 a_8229_n8437# a_8328_n8695# 0.49fF
C7531 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X a_7040_n13591# 0.05fF
C7532 a_5949_n9213# a_7237_n9213# 0.01fF
C7533 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_7130_n9213# 0.03fF
C7534 a_8229_n5797# VDD 0.36fF
C7535 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.01fF
C7536 a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C7537 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_3436_n3255# 0.01fF
C7538 a_2148_n3255# a_2085_n4317# 0.00fF
C7539 a_7130_n6493# a_7130_n8125# 0.00fF
C7540 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkinv_1_3/A 0.45fF
C7541 a_n688_n9783# a_n428_n9783# 0.28fF
C7542 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.01fF
C7543 a_8525_n4317# a_8588_n3799# 0.01fF
C7544 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3010_n13021# 0.35fF
C7545 a_1978_n13021# a_3373_n13021# 0.01fF
C7546 a_2085_n13021# a_3266_n13021# 0.01fF
C7547 a_6941_n12325# a_6941_n13413# 0.02fF
C7548 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_501_n3621# 0.17fF
C7549 a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.01fF
C7550 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_1722_n13021# 0.03fF
C7551 a_5752_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C7552 a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C7553 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_8162_n8125# 0.00fF
C7554 sky130_fd_sc_hd__nand2_4_1/B a_10805_n4709# 0.01fF
C7555 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C7556 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10738_n5405# 0.35fF
C7557 a_9813_n5405# a_10994_n5405# 0.01fF
C7558 a_1978_n13021# VDD 0.46fF
C7559 a_5949_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.12fF
C7560 a_9876_n11415# a_9813_n10301# 0.00fF
C7561 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C7562 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VDD 0.86fF
C7563 a_6874_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C7564 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n11933# 0.00fF
C7565 a_6874_n2685# a_8418_n2685# 0.01fF
C7566 a_7130_n2685# a_8162_n2685# 0.02fF
C7567 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_8162_n9213# 0.03fF
C7568 a_13765_n9213# p2 0.12fF
C7569 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.00fF
C7570 a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C7571 a_9616_n12503# a_8229_n12325# 0.01fF
C7572 a_9517_n12325# a_8328_n12503# 0.01fF
C7573 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# 0.58fF
C7574 a_11164_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.00fF
C7575 a_434_n10301# VDD 0.76fF
C7576 a_860_n4887# a_860_n3799# 0.02fF
C7577 sky130_fd_sc_hd__nand2_4_3/Y a_10904_n9783# 0.05fF
C7578 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 1.54fF
C7579 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C7580 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1978_n9213# 0.03fF
C7581 a_6941_n11237# a_6941_n12325# 0.02fF
C7582 a_7130_n2685# a_7300_n3799# 0.00fF
C7583 a_7237_n2685# a_7040_n3799# 0.00fF
C7584 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C7585 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_3373_n11933# 0.00fF
C7586 a_434_n10301# a_1978_n10301# 0.01fF
C7587 a_690_n10301# a_1722_n10301# 0.02fF
C7588 a_3010_n5405# a_3077_n4709# 0.01fF
C7589 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_10738_n4317# 0.00fF
C7590 a_7300_n4887# a_7300_n3255# 0.01fF
C7591 a_3176_n9783# a_3266_n9213# 0.02fF
C7592 a_4661_n11933# a_4661_n10301# 0.01fF
C7593 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y 0.46fF
C7594 a_9616_n1079# a_8229_n821# 0.01fF
C7595 a_9517_n821# a_8328_n1079# 0.01fF
C7596 a_6012_n11415# a_7300_n11415# 0.01fF
C7597 a_6101_n7254# a_6658_n7363# 0.14fF
C7598 a_3077_n11237# a_3176_n10871# 0.01fF
C7599 a_3176_n11415# a_3077_n10613# 0.01fF
C7600 a_2366_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C7601 a_6006_n7607# a_6665_n7459# 0.03fF
C7602 a_5052_n7283# a_6865_n7304# 0.00fF
C7603 B B_b 0.47fF
C7604 a_5752_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C7605 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_7040_n11415# 0.05fF
C7606 a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.02fF
C7607 a_3176_n13591# a_3436_n13591# 0.28fF
C7608 a_11164_n3255# a_11164_n4887# 0.01fF
C7609 a_3436_n8695# a_4724_n8695# 0.01fF
C7610 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X a_7300_n3799# 0.03fF
C7611 a_3176_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C7612 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_4464_n8695# 0.05fF
C7613 a_5586_n10301# a_5752_n8695# 0.00fF
C7614 a_5842_n10301# a_5653_n8437# 0.00fF
C7615 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C7616 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_4365_n13413# 0.01fF
C7617 a_8229_n8437# a_8162_n10301# 0.00fF
C7618 a_8418_n6493# a_9813_n6493# 0.01fF
C7619 a_7040_n8695# a_6012_n8695# 0.02fF
C7620 a_7300_n8695# a_5752_n8695# 0.01fF
C7621 a_4365_n11237# a_4298_n10301# 0.00fF
C7622 a_8328_n8695# a_9616_n8695# 0.01fF
C7623 a_8588_n8695# a_9517_n8437# 0.02fF
C7624 a_8229_n8437# a_9876_n8695# 0.00fF
C7625 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.07fF
C7626 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.29fF
C7627 a_7237_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.12fF
C7628 a_8162_n5405# a_8229_n5797# 0.01fF
C7629 a_2148_n5975# a_2085_n4317# 0.00fF
C7630 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C7631 a_9876_n2167# a_9813_n1597# 0.01fF
C7632 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_10738_n13021# 0.00fF
C7633 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n8125# 0.00fF
C7634 a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C7635 a_10805_n1909# a_10805_n3621# 0.00fF
C7636 a_6373_n7349# VDD 0.43fF
C7637 a_8162_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C7638 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_4554_n13021# 0.00fF
C7639 a_9813_n5405# a_9706_n4317# 0.00fF
C7640 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.02fF
C7641 a_3266_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.05fF
C7642 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.06fF
C7643 a_1789_n5797# a_501_n5797# 0.01fF
C7644 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_1888_n3799# 0.01fF
C7645 a_2148_n12503# a_2085_n13021# 0.01fF
C7646 a_10994_n5405# sky130_fd_sc_hd__clkinv_4_4/A 0.01fF
C7647 a_4464_n10871# a_4554_n10301# 0.02fF
C7648 a_3373_n13021# VDD 0.34fF
C7649 a_600_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.03fF
C7650 a_860_n12503# VDD 0.78fF
C7651 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.08fF
C7652 a_3010_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C7653 a_3266_n2685# a_3373_n2685# 0.55fF
C7654 a_1789_n4709# a_1722_n5405# 0.01fF
C7655 a_1789_n821# a_3077_n821# 0.01fF
C7656 a_1888_n3255# a_1722_n1597# 0.00fF
C7657 a_8162_n2685# a_8525_n2685# 0.05fF
C7658 a_10904_n10871# a_10904_n9783# 0.01fF
C7659 a_6012_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.03fF
C7660 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_5949_n9213# 0.01fF
C7661 a_7237_n10301# a_7237_n11933# 0.01fF
C7662 a_3077_n2997# a_3010_n2685# 0.01fF
C7663 a_8588_n8695# a_8525_n9213# 0.01fF
C7664 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.06fF
C7665 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2366_n14109# 0.33fF
C7666 a_1978_n10301# VDD 0.44fF
C7667 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C7668 a_10738_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C7669 p2d a_13765_n9757# 2.55fF
C7670 a_8328_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.03fF
C7671 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A a_860_n9783# 0.00fF
C7672 a_2085_n2685# a_1888_n3799# 0.00fF
C7673 a_1722_n10301# a_2085_n10301# 0.05fF
C7674 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A a_4298_n9213# 0.03fF
C7675 a_600_n11415# a_600_n10871# 0.07fF
C7676 a_n688_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.02fF
C7677 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_9616_n5975# 0.05fF
C7678 a_7130_n8125# a_7237_n9213# 0.00fF
C7679 a_7237_n8125# a_7130_n9213# 0.00fF
C7680 Bd_b a_4661_n9213# 0.00fF
C7681 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.29fF
C7682 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.03fF
C7683 a_3176_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C7684 a_3436_n13591# a_4724_n13591# 0.01fF
C7685 a_5949_n5405# a_6012_n4887# 0.01fF
C7686 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.29fF
C7687 a_4724_n5975# Bd_b 0.00fF
C7688 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_4464_n13591# 0.05fF
C7689 a_8162_n509# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C7690 a_8328_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.01fF
C7691 a_2729_n14109# VDD 0.34fF
C7692 a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C7693 a_9616_n8695# a_9876_n8695# 0.28fF
C7694 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_3436_n3799# 0.03fF
C7695 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C7696 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.02fF
C7697 a_860_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.29fF
C7698 a_4623_n7349# sky130_fd_sc_hd__dfxbp_1_0/Q 0.55fF
C7699 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.02fF
C7700 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.05fF
C7701 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.02fF
C7702 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_3077_n11237# 0.01fF
C7703 a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.02fF
C7704 a_1888_n11415# a_2148_n11415# 0.28fF
C7705 a_3436_n2167# a_3436_n3799# 0.01fF
C7706 sky130_fd_sc_hd__nand2_4_3/Y a_11101_n9213# 0.10fF
C7707 a_8525_n6493# a_8525_n8125# 0.00fF
C7708 a_11164_n11415# a_11101_n13021# 0.00fF
C7709 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4661_n13021# 0.02fF
C7710 a_3373_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C7711 a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.02fF
C7712 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_3176_n10871# 0.00fF
C7713 a_4724_n10871# a_3436_n10871# 0.01fF
C7714 a_8328_n12503# a_8328_n13591# 0.01fF
C7715 a_4464_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.05fF
C7716 a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C7717 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n4317# 0.00fF
C7718 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VDD 0.87fF
C7719 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_5586_n10301# 0.03fF
C7720 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.02fF
C7721 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C7722 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_2148_n12503# 0.03fF
C7723 a_9517_n9525# a_9450_n9213# 0.01fF
C7724 a_8328_n8695# a_8418_n8125# 0.02fF
C7725 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD 0.86fF
C7726 a_4724_n9783# a_4661_n10301# 0.01fF
C7727 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_4724_n2167# 0.00fF
C7728 a_8162_n5405# VDD 0.76fF
C7729 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C7730 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4554_n2685# 0.03fF
C7731 a_10805_n13413# a_10994_n13021# 0.02fF
C7732 a_3266_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C7733 a_3373_n2685# a_4661_n2685# 0.01fF
C7734 a_690_n1597# a_1722_n1597# 0.02fF
C7735 a_434_n1597# a_1978_n1597# 0.01fF
C7736 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n2685# 0.35fF
C7737 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.04fF
C7738 a_8418_n2685# a_9813_n2685# 0.01fF
C7739 a_8525_n2685# a_9706_n2685# 0.01fF
C7740 a_n688_n4887# VDD 0.48fF
C7741 a_2085_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.12fF
C7742 a_8418_n13021# a_8418_n14109# 0.01fF
C7743 a_2622_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.04fF
C7744 a_9813_n6493# a_9616_n5975# 0.02fF
C7745 a_3373_n10301# VDD 0.35fF
C7746 a_4554_n11933# a_5586_n11933# 0.02fF
C7747 a_600_n12503# a_600_n13591# 0.01fF
C7748 a_2148_n3255# a_2085_n2685# 0.01fF
C7749 a_501_n1909# a_690_n2685# 0.02fF
C7750 a_600_n2167# a_434_n2685# 0.04fF
C7751 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_9876_n9783# 0.03fF
C7752 a_8328_n11415# a_8328_n12503# 0.01fF
C7753 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C7754 a_501_n13413# VDD 0.36fF
C7755 a_6874_n8125# a_7130_n8125# 0.19fF
C7756 a_8525_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C7757 a_10805_n4709# a_10805_n3621# 0.02fF
C7758 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8588_n3799# 0.01fF
C7759 a_2085_n10301# a_3266_n10301# 0.01fF
C7760 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n10301# 0.35fF
C7761 a_8328_n2167# a_8418_n2685# 0.01fF
C7762 a_1978_n10301# a_3373_n10301# 0.01fF
C7763 a_7237_n509# a_7237_n1597# 0.02fF
C7764 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C7765 a_8418_n10301# a_8525_n11933# 0.00fF
C7766 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.03fF
C7767 a_9876_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.29fF
C7768 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.02fF
C7769 a_3436_n3799# a_3436_n4887# 0.02fF
C7770 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.02fF
C7771 a_8162_n4317# a_8328_n5975# 0.00fF
C7772 a_8418_n4317# a_8229_n5797# 0.00fF
C7773 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.29fF
C7774 a_4365_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C7775 a_11164_n10871# a_10994_n9213# 0.00fF
C7776 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C7777 a_2148_n11415# a_3436_n11415# 0.01fF
C7778 a_1888_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C7779 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_3176_n11415# 0.05fF
C7780 a_10904_n10871# a_11101_n9213# 0.00fF
C7781 a_9706_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.05fF
C7782 sky130_fd_sc_hd__mux2_1_0/X a_4464_n8695# 0.00fF
C7783 a_434_n11933# a_434_n10301# 0.01fF
C7784 a_10904_n12503# a_10904_n11415# 0.01fF
C7785 a_9876_n1079# VDD 0.74fF
C7786 p2d p2d_b 0.47fF
C7787 a_11101_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.10fF
C7788 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C7789 a_13765_n8669# p2_b 0.12fF
C7790 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# 0.58fF
C7791 a_8229_n11237# a_9616_n11415# 0.01fF
C7792 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.08fF
C7793 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_434_n4317# 0.00fF
C7794 a_6874_n4317# VDD 0.76fF
C7795 a_6012_n10871# a_5949_n10301# 0.01fF
C7796 a_9813_n2685# a_9813_n4317# 0.01fF
C7797 a_8525_n13021# a_9813_n13021# 0.01fF
C7798 a_8418_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C7799 a_3077_n3621# VDD 0.35fF
C7800 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_9450_n8125# 0.03fF
C7801 a_7237_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C7802 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8525_n10301# 0.02fF
C7803 a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C7804 a_600_n8695# a_600_n9783# 0.01fF
C7805 a_3077_n11237# a_3077_n9525# 0.00fF
C7806 a_9706_n5405# VDD 0.45fF
C7807 a_4661_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.12fF
C7808 a_1722_n1597# a_2085_n1597# 0.05fF
C7809 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.02fF
C7810 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C7811 a_9706_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.05fF
C7812 a_4464_n3255# a_4554_n2685# 0.02fF
C7813 a_n860_n6173# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C7814 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.02fF
C7815 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n14109# 0.01fF
C7816 a_9450_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C7817 a_6941_n3621# a_6941_n2997# 0.05fF
C7818 sky130_fd_sc_hd__nand2_4_1/B a_10904_n5975# 0.02fF
C7819 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_7237_n14109# 0.01fF
C7820 a_10994_n11933# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C7821 a_8418_n10301# a_8525_n10301# 0.55fF
C7822 a_6874_n8125# a_8525_n8125# 0.00fF
C7823 a_8328_n4887# a_6941_n4709# 0.01fF
C7824 a_8229_n4709# a_7040_n4887# 0.01fF
C7825 a_7130_n8125# a_8418_n8125# 0.01fF
C7826 a_7237_n8125# a_8162_n8125# 0.02fF
C7827 a_3266_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.05fF
C7828 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_9450_n2685# 0.03fF
C7829 a_1722_n13021# a_1722_n11933# 0.02fF
C7830 a_501_n2997# a_1789_n2997# 0.01fF
C7831 a_5949_n9213# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C7832 a_1789_n8437# a_1888_n8695# 0.49fF
C7833 a_2085_n5405# a_1978_n4317# 0.00fF
C7834 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_9517_n821# 0.18fF
C7835 a_10738_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C7836 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6012_n4887# 0.03fF
C7837 a_9450_n10301# a_9450_n11933# 0.01fF
C7838 a_11101_n1597# a_10994_n2685# 0.00fF
C7839 a_10994_n1597# a_11101_n2685# 0.00fF
C7840 a_9813_n11933# a_9616_n12503# 0.02fF
C7841 sky130_fd_sc_hd__nand2_4_0/Y a_10738_n1597# 0.08fF
C7842 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C7843 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.29fF
C7844 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.43fF
C7845 a_600_n12503# a_690_n11933# 0.01fF
C7846 a_3010_n1597# a_3176_n1079# 0.04fF
C7847 a_3266_n1597# a_3077_n821# 0.02fF
C7848 a_434_n11933# VDD 0.77fF
C7849 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.02fF
C7850 a_7130_n13021# a_6941_n13413# 0.02fF
C7851 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_8588_n3799# 0.00fF
C7852 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C7853 a_7300_n4887# a_8229_n4709# 0.02fF
C7854 a_6874_n13021# a_7040_n13591# 0.04fF
C7855 a_1888_n2167# a_1888_n1079# 0.01fF
C7856 a_5752_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C7857 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Ad_b 0.02fF
C7858 a_8229_n1909# a_8588_n2167# 0.05fF
C7859 a_9813_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C7860 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.29fF
C7861 sky130_fd_sc_hd__clkinv_4_8/A a_9813_n14109# 0.02fF
C7862 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_11101_n4317# 0.02fF
C7863 sky130_fd_sc_hd__nand2_4_0/A a_11101_n1597# 0.00fF
C7864 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.03fF
C7865 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_797_n10301# 0.01fF
C7866 sky130_fd_sc_hd__dfxbp_1_0/Q a_5082_n7542# 0.01fF
C7867 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD 3.54fF
C7868 a_5653_n10613# a_5586_n11933# 0.00fF
C7869 a_9616_n9783# a_9813_n10301# 0.02fF
C7870 a_9876_n9783# a_9706_n10301# 0.04fF
C7871 a_3373_n1597# a_3266_n2685# 0.00fF
C7872 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkinv_1_5/A 0.02fF
C7873 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C7874 a_9813_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C7875 a_501_n11237# a_600_n9783# 0.00fF
C7876 a_600_n11415# a_501_n9525# 0.00fF
C7877 a_5653_n11237# a_5586_n10301# 0.00fF
C7878 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C7879 a_9517_n11237# a_9876_n11415# 0.05fF
C7880 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9876_n3799# 0.00fF
C7881 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_7300_n11415# 0.00fF
C7882 a_8418_n4317# VDD 0.47fF
C7883 a_9813_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.01fF
C7884 a_3373_n4317# a_3266_n2685# 0.00fF
C7885 a_3266_n4317# a_3373_n2685# 0.00fF
C7886 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__nand2_4_0/Y 0.06fF
C7887 a_7237_n509# a_7040_n2167# 0.00fF
C7888 a_4464_n3799# VDD 0.44fF
C7889 sky130_fd_sc_hd__nand2_4_0/B VDD 1.25fF
C7890 a_7130_n509# a_7300_n2167# 0.00fF
C7891 a_3077_n2997# a_3010_n4317# 0.00fF
C7892 a_8162_n5405# a_9706_n5405# 0.01fF
C7893 a_8418_n5405# a_9450_n5405# 0.02fF
C7894 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_3/Y 0.03fF
C7895 a_6874_n13021# a_7040_n11415# 0.00fF
C7896 a_10805_n4709# a_11164_n4887# 0.05fF
C7897 a_7130_n13021# a_6941_n11237# 0.00fF
C7898 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.02fF
C7899 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C7900 a_2085_n1597# a_3266_n1597# 0.01fF
C7901 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3010_n1597# 0.35fF
C7902 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_5586_n2685# 0.03fF
C7903 a_n688_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.02fF
C7904 a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C7905 a_8418_n2685# a_8229_n821# 0.00fF
C7906 a_10738_n8125# sky130_fd_sc_hd__clkinv_4_3/A 0.00fF
C7907 a_8162_n2685# a_8328_n1079# 0.00fF
C7908 a_8588_n2167# sky130_fd_sc_hd__nand2_4_0/Y 0.11fF
C7909 sky130_fd_sc_hd__nand2_4_3/B Ad_b 0.04fF
C7910 a_5752_n12503# a_5842_n11933# 0.01fF
C7911 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_1789_n5797# 0.18fF
C7912 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C7913 a_4365_n2997# a_5653_n2997# 0.01fF
C7914 a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.02fF
C7915 a_5752_n9783# a_6012_n9783# 0.28fF
C7916 a_3010_n10301# a_3010_n9213# 0.02fF
C7917 a_11164_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.00fF
C7918 a_8418_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C7919 a_8418_n8125# a_8525_n8125# 0.55fF
C7920 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_9450_n8125# 0.00fF
C7921 a_8162_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C7922 a_4464_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C7923 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.03fF
C7924 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.04fF
C7925 a_8229_n10613# a_8162_n11933# 0.00fF
C7926 a_9616_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.03fF
C7927 a_1789_n4709# a_1789_n3621# 0.02fF
C7928 sky130_fd_sc_hd__clkinv_4_8/A a_9616_n12503# 0.07fF
C7929 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_10904_n1079# 0.01fF
C7930 a_13765_n5949# A 2.52fF
C7931 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.00fF
C7932 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_860_n3799# 0.00fF
C7933 p2d VDD 4.20fF
C7934 a_501_n12325# a_501_n10613# 0.00fF
C7935 a_10994_n9213# a_9706_n9213# 0.01fF
C7936 a_11101_n9213# a_9450_n9213# 0.00fF
C7937 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.04fF
C7938 a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.01fF
C7939 a_10805_n13413# a_11164_n13591# 0.05fF
C7940 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C7941 a_1789_n2997# a_1978_n4317# 0.00fF
C7942 a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.02fF
C7943 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_9517_n4709# 0.01fF
C7944 a_8328_n4887# a_8588_n4887# 0.28fF
C7945 sky130_fd_sc_hd__clkinv_1_5/A p2 0.05fF
C7946 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.05fF
C7947 a_1722_n10301# a_1722_n11933# 0.01fF
C7948 a_10805_n13413# a_9517_n13413# 0.01fF
C7949 a_4724_n5975# a_4724_n4887# 0.02fF
C7950 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C7951 a_1722_n4317# a_1978_n4317# 0.19fF
C7952 a_6101_n7254# a_5842_n9213# 0.00fF
C7953 a_434_n11933# a_501_n13413# 0.00fF
C7954 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C7955 a_9706_n13021# a_9876_n12503# 0.04fF
C7956 a_600_n1079# VDD 0.49fF
C7957 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.08fF
C7958 sky130_fd_sc_hd__clkinv_4_4/A a_8229_n5797# 0.07fF
C7959 a_7130_n6493# a_7040_n4887# 0.00fF
C7960 a_4464_n3255# a_6012_n3255# 0.01fF
C7961 a_4724_n3255# a_5752_n3255# 0.02fF
C7962 VDD a_5586_n9213# 0.76fF
C7963 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_2085_n1597# 0.01fF
C7964 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.03fF
C7965 a_434_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.03fF
C7966 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_3176_n5975# 0.01fF
C7967 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_6874_n11933# 0.03fF
C7968 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkinv_1_4/Y 0.00fF
C7969 a_8328_n3799# a_8328_n3255# 0.07fF
C7970 a_6941_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C7971 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_7040_n9783# 0.05fF
C7972 a_5752_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.00fF
C7973 a_6012_n9783# a_7300_n9783# 0.01fF
C7974 a_7130_n6493# a_7300_n4887# 0.00fF
C7975 a_9450_n10301# a_10994_n10301# 0.01fF
C7976 a_9706_n10301# a_10738_n10301# 0.02fF
C7977 a_9813_n5405# VDD 0.33fF
C7978 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C7979 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_3436_n9783# 0.00fF
C7980 a_501_n5797# a_434_n5405# 0.01fF
C7981 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.03fF
C7982 a_434_n13021# a_797_n13021# 0.05fF
C7983 a_5752_n2167# a_5842_n2685# 0.01fF
C7984 a_3266_n13021# a_3266_n11933# 0.01fF
C7985 a_9813_n9213# a_9813_n10301# 0.02fF
C7986 a_1888_n3255# VDD 0.46fF
C7987 a_2085_n2685# a_3010_n2685# 0.02fF
C7988 a_8328_n2167# a_8229_n821# 0.00fF
C7989 a_8229_n1909# a_8328_n1079# 0.00fF
C7990 a_1888_n12503# a_1978_n11933# 0.01fF
C7991 a_1722_n2685# a_3373_n2685# 0.00fF
C7992 a_1978_n2685# a_3266_n2685# 0.01fF
C7993 a_7130_n2685# VDD 0.44fF
C7994 a_3077_n1909# a_4365_n1909# 0.01fF
C7995 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X a_11164_n1079# 0.03fF
C7996 a_9876_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.00fF
C7997 a_3010_n11933# VDD 0.76fF
C7998 a_11101_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C7999 sky130_fd_sc_hd__clkinv_4_8/A a_11164_n12503# 0.10fF
C8000 a_4724_n12503# a_4661_n11933# 0.01fF
C8001 a_8328_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C8002 a_3436_n2167# a_3436_n1079# 0.02fF
C8003 a_8418_n13021# a_8588_n13591# 0.04fF
C8004 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VDD 0.84fF
C8005 a_8525_n13021# a_8328_n13591# 0.02fF
C8006 a_8588_n4887# a_9876_n4887# 0.01fF
C8007 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_9616_n4887# 0.05fF
C8008 a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.02fF
C8009 a_7237_n1597# a_8162_n1597# 0.02fF
C8010 sky130_fd_sc_hd__nand2_4_0/B a_9876_n1079# 0.03fF
C8011 a_7130_n1597# a_8418_n1597# 0.01fF
C8012 a_9813_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.01fF
C8013 a_9813_n8125# a_9616_n9783# 0.00fF
C8014 a_9706_n4317# a_9517_n2997# 0.00fF
C8015 a_6874_n4317# a_8418_n4317# 0.01fF
C8016 a_7130_n4317# a_8162_n4317# 0.02fF
C8017 a_4365_n1909# a_5752_n2167# 0.01fF
C8018 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.08fF
C8019 a_1978_n4317# a_3266_n4317# 0.01fF
C8020 a_5752_n3799# a_5586_n4317# 0.04fF
C8021 a_9706_n8125# sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C8022 a_1722_n4317# a_3373_n4317# 0.00fF
C8023 a_5653_n3621# a_5842_n4317# 0.02fF
C8024 a_2085_n4317# a_3010_n4317# 0.02fF
C8025 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.03fF
C8026 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkinv_1_0/A 0.08fF
C8027 a_3077_n3621# a_4464_n3799# 0.01fF
C8028 a_3176_n3799# a_4365_n3621# 0.01fF
C8029 a_7040_n11415# a_7130_n10301# 0.01fF
C8030 a_2622_n6493# a_2729_n6493# 0.54fF
C8031 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C8032 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_4724_n2167# 0.01fF
C8033 a_9706_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C8034 a_4464_n3255# a_4554_n1597# 0.00fF
C8035 a_600_n3255# a_600_n4887# 0.00fF
C8036 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_6012_n13591# 0.03fF
C8037 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C8038 a_9706_n2685# a_9517_n2997# 0.02fF
C8039 a_4464_n3255# a_4554_n4317# 0.01fF
C8040 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.03fF
C8041 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD 1.18fF
C8042 a_8418_n13021# a_8588_n11415# 0.00fF
C8043 a_8525_n13021# a_8328_n11415# 0.00fF
C8044 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_7040_n3255# 0.01fF
C8045 VDD a_8162_n11933# 0.76fF
C8046 a_5752_n12503# a_5653_n13413# 0.00fF
C8047 a_5653_n12325# a_5752_n13591# 0.00fF
C8048 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9876_n13591# 0.00fF
C8049 a_9813_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C8050 a_7300_n12503# a_7237_n11933# 0.01fF
C8051 a_797_n10301# a_860_n9783# 0.01fF
C8052 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.29fF
C8053 a_2729_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C8054 a_2729_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C8055 a_5653_n9525# a_5586_n10301# 0.01fF
C8056 a_2148_n3799# a_1978_n5405# 0.00fF
C8057 a_9813_n5405# a_8162_n5405# 0.00fF
C8058 a_1888_n5975# a_1789_n4709# 0.00fF
C8059 a_1789_n5797# a_1888_n4887# 0.00fF
C8060 a_5752_n2167# a_5752_n3255# 0.01fF
C8061 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.04fF
C8062 a_10738_n10301# a_11101_n10301# 0.05fF
C8063 sky130_fd_sc_hd__clkinv_4_4/A VDD 5.98fF
C8064 a_4298_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C8065 a_690_n13021# a_2085_n13021# 0.01fF
C8066 a_6941_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C8067 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4298_n11933# 0.01fF
C8068 a_690_n1597# VDD 0.45fF
C8069 a_11101_n2685# a_10904_n3255# 0.02fF
C8070 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_4298_n2685# 0.00fF
C8071 a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C8072 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_3010_n11933# 0.03fF
C8073 a_10994_n2685# a_11164_n3255# 0.04fF
C8074 a_8525_n2685# VDD 0.35fF
C8075 a_10994_n4317# a_10904_n3255# 0.01fF
C8076 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X p2 0.02fF
C8077 a_4554_n11933# VDD 0.47fF
C8078 a_6012_n2167# a_6012_n1079# 0.02fF
C8079 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VDD 0.89fF
C8080 a_501_n821# a_1888_n1079# 0.01fF
C8081 a_7130_n5405# a_7300_n3799# 0.00fF
C8082 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.29fF
C8083 a_1888_n10871# a_2085_n9213# 0.00fF
C8084 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C8085 a_7237_n5405# a_7040_n3799# 0.00fF
C8086 a_2366_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C8087 p1_b VDD 4.25fF
C8088 a_3266_n10301# a_3266_n11933# 0.01fF
C8089 sky130_fd_sc_hd__nand2_4_3/B a_10904_n9783# 0.00fF
C8090 a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C8091 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_9450_n1597# 0.00fF
C8092 a_8162_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.03fF
C8093 a_8418_n1597# a_8525_n1597# 0.55fF
C8094 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Ad_b 0.09fF
C8095 a_8162_n4317# a_8525_n4317# 0.05fF
C8096 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_4298_n4317# 0.00fF
C8097 a_3010_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.03fF
C8098 a_7237_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C8099 a_3266_n4317# a_3373_n4317# 0.55fF
C8100 a_6012_n9783# a_5949_n9213# 0.01fF
C8101 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7300_n3255# 0.00fF
C8102 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.03fF
C8103 a_434_n10301# a_501_n8437# 0.00fF
C8104 a_1888_n8695# a_3436_n8695# 0.01fF
C8105 a_2148_n8695# a_3176_n8695# 0.02fF
C8106 a_3077_n821# VDD 0.36fF
C8107 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_8162_n10301# 0.01fF
C8108 a_4365_n3621# a_4724_n3799# 0.05fF
C8109 a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C8110 a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C8111 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_5586_n1597# 0.00fF
C8112 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_7130_n6493# 0.02fF
C8113 a_7130_n6493# a_7212_n7203# 0.00fF
C8114 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.02fF
C8115 a_10738_n11933# a_10805_n11237# 0.01fF
C8116 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkinv_1_5/A 0.03fF
C8117 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.00fF
C8118 a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C8119 a_10738_n1597# VDD 0.70fF
C8120 a_1978_n2685# a_1789_n2997# 0.02fF
C8121 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_860_n10871# 0.01fF
C8122 a_797_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.00fF
C8123 VDD a_9706_n11933# 0.46fF
C8124 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_1722_n4317# 0.03fF
C8125 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.09fF
C8126 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.05fF
C8127 a_8229_n11237# a_8418_n10301# 0.00fF
C8128 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VDD 0.84fF
C8129 a_9813_n8125# a_9813_n9213# 0.02fF
C8130 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_1/A 0.47fF
C8131 a_10738_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.00fF
C8132 a_8525_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.00fF
C8133 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_8588_n4887# 0.00fF
C8134 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9450_n5405# 0.03fF
C8135 a_9813_n5405# a_9706_n5405# 0.55fF
C8136 a_7040_n10871# a_8229_n10613# 0.01fF
C8137 a_6941_n10613# a_8328_n10871# 0.01fF
C8138 sky130_fd_sc_hd__clkinv_1_0/A a_2622_n509# 0.01fF
C8139 a_n428_n12503# a_501_n12325# 0.02fF
C8140 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkinv_1_0/Y 0.02fF
C8141 a_13765_n9213# p2_b 2.55fF
C8142 a_4661_n13021# a_4661_n11933# 0.02fF
C8143 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X 0.29fF
C8144 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_2148_n9783# 0.01fF
C8145 a_2085_n1597# VDD 0.35fF
C8146 a_11101_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C8147 a_3436_n12503# a_3373_n11933# 0.01fF
C8148 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VDD 0.85fF
C8149 a_4661_n5405# a_4464_n4887# 0.02fF
C8150 a_4554_n5405# a_4724_n4887# 0.04fF
C8151 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6941_n3621# 0.01fF
C8152 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.03fF
C8153 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.08fF
C8154 a_4365_n11237# a_4298_n13021# 0.00fF
C8155 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C8156 a_9450_n509# a_9616_n1079# 0.04fF
C8157 a_3077_n12325# a_3077_n11237# 0.02fF
C8158 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n11933# 0.00fF
C8159 a_5842_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C8160 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4554_n1597# 0.03fF
C8161 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_7130_n1597# 0.03fF
C8162 a_5949_n1597# a_7237_n1597# 0.01fF
C8163 a_501_n8437# VDD 0.37fF
C8164 a_3373_n1597# a_4661_n1597# 0.01fF
C8165 a_13765_n1597# a_13765_n2685# 0.07fF
C8166 a_8418_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C8167 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9706_n1597# 0.03fF
C8168 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11101_n2685# 0.01fF
C8169 a_8588_n2167# VDD 0.78fF
C8170 a_8525_n1597# a_9813_n1597# 0.01fF
C8171 a_9517_n11237# a_9616_n9783# 0.00fF
C8172 a_4298_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C8173 a_8162_n509# a_9706_n509# 0.01fF
C8174 a_3266_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C8175 a_3373_n4317# a_4661_n4317# 0.01fF
C8176 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4554_n4317# 0.03fF
C8177 a_9517_n1909# a_9616_n3799# 0.00fF
C8178 a_9616_n2167# a_9517_n3621# 0.00fF
C8179 a_4464_n1079# VDD 0.51fF
C8180 a_4724_n3799# a_5752_n3799# 0.02fF
C8181 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_5653_n3621# 0.18fF
C8182 a_7237_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.12fF
C8183 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VDD 1.21fF
C8184 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.02fF
C8185 a_5842_n13021# a_5949_n11933# 0.00fF
C8186 a_5949_n13021# a_5842_n11933# 0.00fF
C8187 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C8188 a_5653_n2997# a_5653_n4709# 0.00fF
C8189 sky130_fd_sc_hd__clkinv_1_5/A a_7130_n9213# 0.00fF
C8190 a_9706_n10301# VDD 0.43fF
C8191 a_5653_n10613# VDD 0.35fF
C8192 a_4464_n9783# VDD 0.47fF
C8193 a_6941_n5797# a_8328_n5975# 0.01fF
C8194 a_6012_n10871# a_6012_n12503# 0.01fF
C8195 sky130_fd_sc_hd__mux2_1_0/X a_4623_n7349# 0.22fF
C8196 a_4464_n12503# a_4365_n13413# 0.00fF
C8197 a_4365_n12325# a_4464_n13591# 0.00fF
C8198 a_7040_n5975# a_8229_n5797# 0.01fF
C8199 a_6012_n5975# a_6006_n7607# 0.00fF
C8200 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9450_n4317# 0.01fF
C8201 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.06fF
C8202 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.06fF
C8203 a_5842_n1597# a_5752_n2167# 0.02fF
C8204 a_7040_n9783# a_7130_n10301# 0.01fF
C8205 a_n1139_n6715# a_n2248_n7037# 0.01fF
C8206 A a_13765_n4861# 0.06fF
C8207 a_13765_n5949# Ad 0.06fF
C8208 a_7300_n2167# a_7300_n3255# 0.02fF
C8209 a_10805_n1909# a_10994_n2685# 0.02fF
C8210 a_10904_n2167# a_10738_n2685# 0.04fF
C8211 a_5653_n5797# VDD 0.36fF
C8212 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__clkinv_1_3/A 0.16fF
C8213 a_6941_n821# VDD 0.35fF
C8214 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1722_n13021# 0.35fF
C8215 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.04fF
C8216 a_7237_n4317# a_7300_n3799# 0.01fF
C8217 a_797_n13021# a_1978_n13021# 0.01fF
C8218 a_600_n12503# a_501_n11237# 0.00fF
C8219 a_4464_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C8220 a_4724_n3799# a_6012_n3799# 0.01fF
C8221 a_434_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C8222 a_6874_n14109# a_8162_n14109# 0.01fF
C8223 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_3373_n9213# 0.00fF
C8224 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.00fF
C8225 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_8588_n3799# 0.00fF
C8226 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6874_n8125# 0.00fF
C8227 a_8525_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C8228 a_7237_n9213# a_7212_n7203# 0.00fF
C8229 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_3176_n3255# 0.05fF
C8230 sky130_fd_sc_hd__nand2_4_2/A a_6874_n14109# 0.03fF
C8231 a_2148_n3255# a_3436_n3255# 0.01fF
C8232 a_2148_n3799# a_501_n3621# 0.00fF
C8233 a_4661_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.12fF
C8234 a_9813_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.12fF
C8235 a_9813_n11933# a_10738_n11933# 0.02fF
C8236 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.03fF
C8237 a_4661_n10301# a_4661_n9213# 0.02fF
C8238 a_1789_n1909# a_1888_n3799# 0.00fF
C8239 a_1888_n2167# a_1789_n3621# 0.00fF
C8240 a_690_n13021# a_600_n13591# 0.01fF
C8241 a_4554_n4317# a_4365_n4709# 0.02fF
C8242 a_4298_n4317# a_4464_n4887# 0.04fF
C8243 a_4661_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.12fF
C8244 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.08fF
C8245 a_9450_n509# a_9813_n509# 0.05fF
C8246 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C8247 a_434_n2685# a_1722_n2685# 0.01fF
C8248 a_10738_n13021# VDD 0.69fF
C8249 sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C8250 Bd_b p2 0.56fF
C8251 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.09fF
C8252 sky130_fd_sc_hd__nand2_4_3/Y a_8328_n9783# 0.05fF
C8253 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.02fF
C8254 a_600_n5975# a_797_n4317# 0.00fF
C8255 a_860_n5975# a_690_n4317# 0.00fF
C8256 a_5653_n11237# a_5653_n12325# 0.02fF
C8257 a_1888_n10871# a_1978_n9213# 0.00fF
C8258 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_690_n9213# 0.02fF
C8259 a_11101_n10301# VDD 0.32fF
C8260 a_7040_n10871# VDD 0.46fF
C8261 a_3077_n10613# a_4365_n10613# 0.01fF
C8262 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C8263 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_2085_n11933# 0.00fF
C8264 Ad_b sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C8265 a_8229_n5797# a_8588_n5975# 0.05fF
C8266 a_8229_n9525# a_9517_n9525# 0.01fF
C8267 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_9450_n4317# 0.00fF
C8268 a_8588_n12503# a_8418_n14109# 0.00fF
C8269 a_8328_n12503# a_8525_n14109# 0.00fF
C8270 a_6941_n5797# a_6658_n7363# 0.00fF
C8271 a_9813_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.00fF
C8272 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_600_n4887# 0.01fF
C8273 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9876_n1079# 0.00fF
C8274 a_9616_n8695# a_10805_n8437# 0.01fF
C8275 a_9517_n8437# a_10904_n8695# 0.01fF
C8276 a_8418_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.08fF
C8277 a_1888_n11415# a_1789_n10613# 0.01fF
C8278 a_1789_n11237# a_1888_n10871# 0.01fF
C8279 a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.01fF
C8280 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6941_n1909# 0.01fF
C8281 a_6874_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.03fF
C8282 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C8283 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_860_n3255# 0.00fF
C8284 a_501_n4709# a_n787_n4709# 0.01fF
C8285 a_501_n10613# a_1789_n10613# 0.01fF
C8286 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.04fF
C8287 a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C8288 a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.02fF
C8289 a_1888_n13591# a_2148_n13591# 0.28fF
C8290 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_8162_n10301# 0.03fF
C8291 a_4554_n10301# a_4365_n8437# 0.00fF
C8292 a_4298_n10301# a_4464_n8695# 0.00fF
C8293 a_8525_n2685# a_8418_n4317# 0.00fF
C8294 a_8418_n2685# a_8525_n4317# 0.00fF
C8295 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.28fF
C8296 a_7300_n8695# a_8229_n8437# 0.02fF
C8297 a_7040_n8695# a_8328_n8695# 0.01fF
C8298 a_6874_n5405# a_6941_n5797# 0.01fF
C8299 clk a_n1738_n6671# 0.01fF
C8300 a_7040_n5975# VDD 0.44fF
C8301 a_5949_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.12fF
C8302 a_9616_n4887# a_9517_n3621# 0.00fF
C8303 a_9517_n4709# a_9616_n3799# 0.00fF
C8304 a_8328_n1079# VDD 0.46fF
C8305 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n8125# 0.00fF
C8306 a_1978_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.05fF
C8307 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_3266_n13021# 0.00fF
C8308 a_11164_n3799# a_11164_n3255# 0.09fF
C8309 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.29fF
C8310 a_8162_n13021# a_9450_n13021# 0.01fF
C8311 a_860_n12503# a_797_n13021# 0.01fF
C8312 a_8229_n9525# a_8418_n10301# 0.02fF
C8313 a_797_n13021# VDD 0.35fF
C8314 a_9813_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.07fF
C8315 a_9813_n6493# a_9876_n4887# 0.00fF
C8316 a_7300_n9783# a_7237_n8125# 0.00fF
C8317 a_4464_n12503# a_4464_n11415# 0.01fF
C8318 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.02fF
C8319 a_2148_n3799# a_1888_n3799# 0.28fF
C8320 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_1789_n3621# 0.02fF
C8321 a_10738_n11933# sky130_fd_sc_hd__clkinv_4_8/A 0.00fF
C8322 a_10994_n11933# a_11101_n11933# 0.55fF
C8323 a_11101_n1597# a_10904_n1079# 0.02fF
C8324 a_10994_n1597# a_11164_n1079# 0.04fF
C8325 a_5586_n13021# a_6874_n13021# 0.01fF
C8326 a_5949_n10301# a_5949_n11933# 0.01fF
C8327 a_6874_n2685# a_7237_n2685# 0.05fF
C8328 a_9616_n10871# a_9616_n9783# 0.01fF
C8329 a_7300_n8695# a_7237_n9213# 0.01fF
C8330 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_n787_n4709# 0.01fF
C8331 a_1722_n2685# a_1978_n2685# 0.19fF
C8332 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_1789_n821# 0.18fF
C8333 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.04fF
C8334 sky130_fd_sc_hd__nand2_4_0/B a_10738_n1597# 0.01fF
C8335 a_5842_n13021# a_5752_n13591# 0.01fF
C8336 sky130_fd_sc_hd__nand2_4_3/Y a_9876_n9783# 0.11fF
C8337 a_10805_n4709# a_10738_n4317# 0.01fF
C8338 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.04fF
C8339 a_10805_n2997# VDD 0.32fF
C8340 a_797_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.12fF
C8341 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C8342 a_8525_n4317# a_9813_n4317# 0.01fF
C8343 a_690_n13021# a_690_n11933# 0.01fF
C8344 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9706_n4317# 0.03fF
C8345 a_797_n2685# a_600_n3799# 0.00fF
C8346 a_690_n2685# a_860_n3799# 0.00fF
C8347 a_8418_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C8348 a_434_n10301# a_797_n10301# 0.05fF
C8349 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X a_3010_n9213# 0.03fF
C8350 a_3077_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C8351 a_434_n4317# VDD 0.77fF
C8352 a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C8353 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.29fF
C8354 a_2148_n13591# a_3436_n13591# 0.01fF
C8355 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.29fF
C8356 a_1888_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.00fF
C8357 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X a_3176_n13591# 0.05fF
C8358 a_9517_n2997# VDD 0.34fF
C8359 a_7040_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C8360 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.02fF
C8361 a_n688_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.04fF
C8362 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.02fF
C8363 a_690_n1597# a_600_n1079# 0.01fF
C8364 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_9517_n8437# 0.01fF
C8365 a_8328_n8695# a_8588_n8695# 0.28fF
C8366 a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.02fF
C8367 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C8368 a_8588_n5975# VDD 0.78fF
C8369 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.03fF
C8370 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C8371 a_9876_n11415# a_9813_n13021# 0.00fF
C8372 a_7237_n6493# a_7237_n8125# 0.00fF
C8373 a_2085_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C8374 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.08fF
C8375 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3373_n13021# 0.02fF
C8376 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_860_n3799# 0.02fF
C8377 a_7040_n12503# a_7040_n13591# 0.01fF
C8378 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.08fF
C8379 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C8380 a_2148_n3799# a_2148_n3255# 0.09fF
C8381 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.08fF
C8382 a_9450_n13021# a_9706_n13021# 0.19fF
C8383 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_11101_n5405# 0.02fF
C8384 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VDD 0.87fF
C8385 a_501_n1909# a_1789_n1909# 0.01fF
C8386 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C8387 a_7040_n8695# a_7130_n8125# 0.02fF
C8388 sky130_fd_sc_hd__nand2_1_0/B VDD 1.53fF
C8389 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkinv_1_5/A 0.02fF
C8390 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C8391 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.00fF
C8392 a_7130_n10301# a_7237_n9213# 0.00fF
C8393 a_1789_n821# a_1888_n1079# 0.49fF
C8394 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.04fF
C8395 a_7237_n10301# a_7130_n9213# 0.00fF
C8396 a_7237_n2685# a_8418_n2685# 0.01fF
C8397 a_7130_n2685# a_8525_n2685# 0.01fF
C8398 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n2685# 0.35fF
C8399 a_9876_n12503# a_8328_n12503# 0.01fF
C8400 a_9616_n12503# a_8588_n12503# 0.02fF
C8401 a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.18fF
C8402 sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# 0.53fF
C8403 a_797_n10301# VDD 0.36fF
C8404 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C8405 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.04fF
C8406 a_3010_n11933# a_4554_n11933# 0.01fF
C8407 a_3266_n11933# a_4298_n11933# 0.02fF
C8408 a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C8409 a_7040_n11415# a_7040_n12503# 0.01fF
C8410 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7300_n3799# 0.01fF
C8411 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C8412 a_6874_n14109# a_6941_n13413# 0.01fF
C8413 a_3266_n5405# a_3176_n4887# 0.02fF
C8414 a_797_n10301# a_1978_n10301# 0.01fF
C8415 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n10301# 0.35fF
C8416 a_690_n10301# a_2085_n10301# 0.01fF
C8417 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C8418 a_4365_n9525# a_4298_n9213# 0.01fF
C8419 a_3436_n9783# a_3373_n9213# 0.01fF
C8420 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.02fF
C8421 a_9616_n1079# a_8588_n1079# 0.02fF
C8422 a_9876_n1079# a_8328_n1079# 0.01fF
C8423 a_6101_n7254# a_6865_n7304# 0.05fF
C8424 a_6373_n7349# a_6665_n7459# 0.39fF
C8425 a_13765_n1597# VDD 2.00fF
C8426 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.02fF
C8427 a_6006_n7607# a_6794_n7203# 0.02fF
C8428 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.29fF
C8429 a_6874_n10301# a_8162_n10301# 0.01fF
C8430 a_7130_n4317# a_6941_n5797# 0.00fF
C8431 a_5949_n10301# a_5752_n8695# 0.00fF
C8432 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9813_n6493# 0.02fF
C8433 a_8525_n6493# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C8434 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.02fF
C8435 a_5842_n10301# a_6012_n8695# 0.00fF
C8436 a_6874_n4317# a_7040_n5975# 0.00fF
C8437 a_7130_n509# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C8438 a_4464_n11415# a_4554_n10301# 0.01fF
C8439 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A VDD 1.13fF
C8440 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.03fF
C8441 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_6012_n8695# 0.00fF
C8442 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_9616_n8695# 0.05fF
C8443 a_8328_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C8444 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1789_n821# 0.01fF
C8445 a_8588_n8695# a_9876_n8695# 0.01fF
C8446 a_10738_n5405# a_10805_n5797# 0.01fF
C8447 a_1722_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.03fF
C8448 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.00fF
C8449 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_1888_n11415# 0.05fF
C8450 a_8418_n5405# a_8328_n5975# 0.01fF
C8451 a_9616_n10871# a_9813_n9213# 0.00fF
C8452 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C8453 a_10904_n13591# VDD 0.38fF
C8454 sky130_fd_sc_hd__nand2_4_3/Y a_10738_n10301# 0.00fF
C8455 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.08fF
C8456 a_9616_n12503# a_9616_n11415# 0.01fF
C8457 a_6665_n7459# VDD 0.89fF
C8458 a_1722_n9213# a_1888_n9783# 0.04fF
C8459 a_10904_n2167# a_10904_n3799# 0.00fF
C8460 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.44fF
C8461 a_1978_n9213# a_1789_n9525# 0.02fF
C8462 a_8229_n1909# a_8162_n509# 0.00fF
C8463 a_1789_n5797# a_860_n5975# 0.02fF
C8464 a_2148_n5975# a_501_n5797# 0.00fF
C8465 a_1888_n5975# a_600_n5975# 0.01fF
C8466 a_5586_n11933# a_7130_n11933# 0.01fF
C8467 a_3077_n8437# a_3176_n9783# 0.00fF
C8468 a_3176_n8695# a_3077_n9525# 0.00fF
C8469 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.08fF
C8470 a_4724_n10871# a_4661_n10301# 0.01fF
C8471 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_8162_n8125# 0.03fF
C8472 a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C8473 a_7130_n5405# VDD 0.47fF
C8474 a_1789_n11237# a_1789_n9525# 0.00fF
C8475 a_3373_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.12fF
C8476 a_1888_n3255# a_2085_n1597# 0.00fF
C8477 a_3176_n3255# a_3266_n2685# 0.02fF
C8478 a_434_n1597# a_797_n1597# 0.05fF
C8479 a_5653_n4709# a_6941_n4709# 0.01fF
C8480 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.02fF
C8481 a_1789_n821# a_3436_n1079# 0.00fF
C8482 a_1888_n4887# a_1978_n5405# 0.02fF
C8483 a_8418_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.05fF
C8484 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_9706_n2685# 0.00fF
C8485 a_5653_n3621# a_5842_n5405# 0.00fF
C8486 a_11164_n10871# a_11164_n9783# 0.02fF
C8487 a_n1738_n6671# sky130_fd_sc_hd__clkinv_1_5/A 0.11fF
C8488 a_5752_n3799# a_5586_n5405# 0.00fF
C8489 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n14109# 0.01fF
C8490 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.06fF
C8491 a_10904_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C8492 a_6874_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.03fF
C8493 a_1722_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.03fF
C8494 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VDD 0.89fF
C8495 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C8496 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2729_n14109# 0.02fF
C8497 a_4298_n11933# a_4661_n11933# 0.05fF
C8498 a_434_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C8499 a_n787_n12325# sky130_fd_sc_hd__nand2_1_4/B 0.28fF
C8500 a_5653_n10613# a_5586_n9213# 0.00fF
C8501 a_1978_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.05fF
C8502 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_3266_n10301# 0.00fF
C8503 a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C8504 a_860_n11415# a_860_n10871# 0.09fF
C8505 a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C8506 a_8162_n4317# a_8229_n2997# 0.00fF
C8507 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C8508 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C8509 a_8418_n10301# a_8418_n9213# 0.01fF
C8510 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.03fF
C8511 a_13765_n4861# Ad 2.55fF
C8512 a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C8513 a_1722_n1597# a_1888_n1079# 0.04fF
C8514 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.02fF
C8515 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.08fF
C8516 a_9706_n8125# sky130_fd_sc_hd__nand2_4_3/B 0.05fF
C8517 a_8418_n11933# a_9450_n11933# 0.02fF
C8518 a_8162_n11933# a_9706_n11933# 0.01fF
C8519 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_100/A 0.00fF
C8520 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C8521 a_10805_n10613# a_10994_n10301# 0.02fF
C8522 a_10904_n10871# a_10738_n10301# 0.04fF
C8523 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X a_5586_n10301# 0.01fF
C8524 a_8525_n509# sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C8525 a_9517_n10613# a_8229_n10613# 0.01fF
C8526 a_1888_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C8527 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.29fF
C8528 a_3176_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C8529 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Ad_b 0.03fF
C8530 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.29fF
C8531 a_3077_n4709# a_3010_n4317# 0.01fF
C8532 sky130_fd_sc_hd__dfxbp_1_0/Q_N a_7212_n7203# 0.01fF
C8533 a_8229_n8437# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C8534 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C8535 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VDD 0.82fF
C8536 a_2622_n8125# VDD 0.49fF
C8537 a_n1995_n6925# a_n1738_n6671# 0.10fF
C8538 a_n2436_n7037# a_n1139_n6715# 0.03fF
C8539 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkinv_4_3/A 0.44fF
C8540 a_8328_n9783# a_8525_n10301# 0.02fF
C8541 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C8542 a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.00fF
C8543 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.02fF
C8544 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.00fF
C8545 a_5842_n4317# VDD 0.47fF
C8546 a_8588_n12503# a_8588_n13591# 0.02fF
C8547 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6012_n11415# 0.00fF
C8548 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__nand2_4_0/Y 0.06fF
C8549 a_9616_n9783# a_9706_n9213# 0.02fF
C8550 a_10904_n2167# a_10738_n509# 0.00fF
C8551 a_8588_n8695# a_8525_n8125# 0.01fF
C8552 a_6874_n5405# a_8418_n5405# 0.01fF
C8553 a_7130_n5405# a_8162_n5405# 0.02fF
C8554 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.06fF
C8555 a_8525_n5405# VDD 0.35fF
C8556 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.02fF
C8557 a_5842_n13021# a_5653_n11237# 0.00fF
C8558 a_501_n4709# a_1789_n4709# 0.01fF
C8559 a_10805_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.05fF
C8560 sky130_fd_sc_hd__nand2_1_4/Y a_2729_n8125# 0.00fF
C8561 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_4298_n2685# 0.03fF
C8562 a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C8563 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1722_n1597# 0.35fF
C8564 a_6941_n4709# a_7040_n4887# 0.49fF
C8565 a_690_n1597# a_2085_n1597# 0.01fF
C8566 a_797_n1597# a_1978_n1597# 0.01fF
C8567 a_8525_n13021# a_8525_n14109# 0.02fF
C8568 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9813_n2685# 0.02fF
C8569 a_8525_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C8570 a_3077_n2997# a_4365_n2997# 0.01fF
C8571 a_7130_n2685# a_6941_n821# 0.00fF
C8572 a_6874_n2685# a_7040_n1079# 0.00fF
C8573 sky130_fd_sc_hd__nand2_4_1/B a_9876_n5975# 0.03fF
C8574 a_9813_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C8575 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5586_n11933# 0.35fF
C8576 a_860_n2167# a_690_n2685# 0.04fF
C8577 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.08fF
C8578 a_600_n2167# a_797_n2685# 0.02fF
C8579 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_434_n13021# 0.42fF
C8580 a_860_n12503# a_860_n13591# 0.02fF
C8581 a_7130_n8125# a_7237_n8125# 0.55fF
C8582 a_6874_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.03fF
C8583 a_8588_n11415# a_8588_n12503# 0.02fF
C8584 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_50/X 0.01fF
C8585 a_860_n13591# VDD 0.78fF
C8586 a_7300_n4887# a_6941_n4709# 0.05fF
C8587 a_10904_n4887# a_10904_n3799# 0.01fF
C8588 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.04fF
C8589 a_8588_n2167# a_8525_n2685# 0.01fF
C8590 sky130_fd_sc_hd__clkinv_4_7/Y VDD 2.22fF
C8591 a_501_n2997# a_600_n3255# 0.49fF
C8592 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3373_n10301# 0.02fF
C8593 a_2085_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.01fF
C8594 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.03fF
C8595 a_6941_n10613# a_6874_n11933# 0.00fF
C8596 a_2148_n8695# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C8597 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n13021# 0.01fF
C8598 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.04fF
C8599 a_10805_n5797# a_10994_n4317# 0.00fF
C8600 a_10904_n5975# a_10738_n4317# 0.00fF
C8601 a_9813_n9213# a_8162_n9213# 0.00fF
C8602 a_8418_n4317# a_8588_n5975# 0.00fF
C8603 a_8525_n4317# a_8328_n5975# 0.00fF
C8604 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.05fF
C8605 a_4724_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C8606 a_3436_n5975# a_3436_n4887# 0.02fF
C8607 a_9616_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C8608 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.02fF
C8609 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.05fF
C8610 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n1597# 0.01fF
C8611 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_1789_n4709# 0.01fF
C8612 a_690_n11933# a_690_n10301# 0.01fF
C8613 a_11164_n12503# a_11164_n11415# 0.02fF
C8614 a_9450_n8125# a_9517_n9525# 0.00fF
C8615 a_3176_n3255# a_1789_n2997# 0.01fF
C8616 a_8588_n11415# a_9616_n11415# 0.02fF
C8617 a_7237_n4317# VDD 0.35fF
C8618 a_8328_n11415# a_9876_n11415# 0.01fF
C8619 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.02fF
C8620 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C8621 a_860_n8695# a_860_n9783# 0.02fF
C8622 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.02fF
C8623 a_3436_n3799# VDD 0.77fF
C8624 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.08fF
C8625 sky130_fd_sc_hd__clkinv_4_4/A a_5653_n5797# 0.07fF
C8626 a_10805_n13413# a_10904_n12503# 0.00fF
C8627 a_3176_n11415# a_3176_n9783# 0.00fF
C8628 a_8162_n5405# a_8525_n5405# 0.05fF
C8629 a_3176_n1079# a_4365_n821# 0.01fF
C8630 a_3077_n821# a_4464_n1079# 0.01fF
C8631 a_9616_n4887# a_11164_n4887# 0.01fF
C8632 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_1_0/Y 0.63fF
C8633 sky130_fd_sc_hd__nand2_4_0/A a_2366_n509# 0.08fF
C8634 a_3077_n1909# a_3266_n2685# 0.02fF
C8635 VDD a_3010_n9213# 0.76fF
C8636 a_1978_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.05fF
C8637 a_3176_n2167# a_3010_n2685# 0.04fF
C8638 a_3077_n5797# VDD 0.36fF
C8639 a_4724_n3255# a_4661_n2685# 0.01fF
C8640 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_3266_n1597# 0.00fF
C8641 a_860_n2167# sky130_fd_sc_hd__clkinv_1_0/A 0.00fF
C8642 a_7040_n3799# a_7040_n3255# 0.07fF
C8643 a_10738_n6173# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C8644 a_2366_n6493# a_2366_n8125# 0.01fF
C8645 a_4365_n2997# a_4464_n3255# 0.49fF
C8646 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C8647 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y 1.53fF
C8648 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11164_n1079# 0.03fF
C8649 a_7237_n8125# a_8525_n8125# 0.01fF
C8650 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8418_n8125# 0.03fF
C8651 a_7130_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C8652 a_9517_n10613# VDD 0.34fF
C8653 a_1978_n13021# a_1978_n11933# 0.01fF
C8654 a_8588_n4887# a_7040_n4887# 0.01fF
C8655 a_4464_n2167# a_4554_n2685# 0.01fF
C8656 a_860_n3255# a_1789_n2997# 0.02fF
C8657 sky130_fd_sc_hd__nand2_4_3/Y VDD 7.72fF
C8658 a_1888_n8695# a_2148_n8695# 0.28fF
C8659 a_9706_n10301# a_9706_n11933# 0.01fF
C8660 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VDD 1.74fF
C8661 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9876_n12503# 0.03fF
C8662 a_9813_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C8663 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_9876_n1079# 0.03fF
C8664 sky130_fd_sc_hd__nand2_4_0/Y a_11101_n1597# 0.10fF
C8665 a_860_n12503# a_797_n11933# 0.01fF
C8666 a_10738_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.00fF
C8667 a_1888_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C8668 a_3266_n1597# a_3436_n1079# 0.04fF
C8669 a_9813_n9213# a_9706_n9213# 0.55fF
C8670 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9450_n9213# 0.03fF
C8671 a_501_n13413# a_860_n13591# 0.05fF
C8672 a_7130_n13021# a_7300_n13591# 0.04fF
C8673 a_797_n11933# VDD 0.35fF
C8674 a_7237_n13021# a_7040_n13591# 0.02fF
C8675 a_2148_n2167# a_2148_n1079# 0.02fF
C8676 a_4365_n821# a_5653_n821# 0.01fF
C8677 a_7300_n4887# a_8588_n4887# 0.01fF
C8678 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_8328_n4887# 0.05fF
C8679 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkinv_1_3/A 0.84fF
C8680 a_8328_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.03fF
C8681 a_5586_n4317# a_7130_n4317# 0.01fF
C8682 a_5842_n4317# a_6874_n4317# 0.02fF
C8683 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__dfxbp_1_0/Q 0.04fF
C8684 sky130_fd_sc_hd__dfxbp_1_0/Q a_7212_n7203# 0.01fF
C8685 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n10301# 0.00fF
C8686 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X a_9813_n10301# 0.01fF
C8687 a_9876_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C8688 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkinv_1_0/A 0.45fF
C8689 a_5752_n11415# a_5842_n10301# 0.01fF
C8690 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A VDD 0.88fF
C8691 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_10904_n11415# 0.01fF
C8692 a_10904_n2167# a_10805_n821# 0.00fF
C8693 a_10805_n1909# a_10904_n1079# 0.00fF
C8694 a_7237_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C8695 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD 0.84fF
C8696 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_7300_n2167# 0.00fF
C8697 a_3176_n3255# a_3266_n4317# 0.01fF
C8698 a_8162_n2685# a_8328_n3255# 0.04fF
C8699 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6941_n4709# 0.00fF
C8700 sky130_fd_sc_hd__clkinv_4_4/A a_7040_n5975# 0.07fF
C8701 a_6874_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C8702 a_8418_n2685# a_8229_n2997# 0.02fF
C8703 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9450_n5405# 0.35fF
C8704 a_8525_n5405# a_9706_n5405# 0.01fF
C8705 a_7237_n13021# a_7040_n11415# 0.00fF
C8706 a_4365_n821# a_4724_n1079# 0.05fF
C8707 a_7130_n13021# a_7300_n11415# 0.00fF
C8708 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_5752_n3255# 0.01fF
C8709 a_10904_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.02fF
C8710 VDD a_4554_n9213# 0.45fF
C8711 a_4464_n5975# VDD 0.49fF
C8712 a_8418_n2685# a_8588_n1079# 0.00fF
C8713 a_4724_n3255# a_5653_n2997# 0.02fF
C8714 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.05fF
C8715 a_8525_n2685# a_8328_n1079# 0.00fF
C8716 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.29fF
C8717 a_6012_n12503# a_5949_n11933# 0.01fF
C8718 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_2148_n5975# 0.03fF
C8719 a_3266_n10301# a_3266_n9213# 0.01fF
C8720 sky130_fd_sc_hd__nand2_1_4/Y a_3832_n7261# 0.01fF
C8721 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_4/Y 0.48fF
C8722 a_501_n11237# a_690_n13021# 0.00fF
C8723 a_9450_n10301# a_9813_n10301# 0.05fF
C8724 a_600_n11415# a_434_n13021# 0.00fF
C8725 a_8525_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.12fF
C8726 a_10904_n10871# VDD 0.41fF
C8727 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.04fF
C8728 a_4365_n9525# a_4724_n9783# 0.05fF
C8729 a_3010_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C8730 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3010_n11933# 0.01fF
C8731 a_5653_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C8732 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_5586_n2685# 0.03fF
C8733 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C8734 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8588_n12503# 0.00fF
C8735 a_8328_n10871# a_8418_n11933# 0.01fF
C8736 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_1722_n11933# 0.03fF
C8737 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_3010_n2685# 0.00fF
C8738 a_1888_n4887# a_1888_n3799# 0.01fF
C8739 a_9706_n4317# a_9616_n3255# 0.01fF
C8740 a_1978_n11933# VDD 0.47fF
C8741 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.70fF
C8742 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.29fF
C8743 a_1978_n10301# a_1978_n11933# 0.01fF
C8744 a_9706_n2685# a_9616_n3255# 0.02fF
C8745 a_7130_n1597# a_7237_n1597# 0.55fF
C8746 a_10805_n13413# a_9876_n13591# 0.02fF
C8747 a_6874_n4317# a_7237_n4317# 0.05fF
C8748 a_1722_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C8749 a_4365_n1909# a_4724_n2167# 0.05fF
C8750 a_1978_n4317# a_2085_n4317# 0.55fF
C8751 a_8162_n13021# a_8229_n12325# 0.01fF
C8752 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X a_6874_n10301# 0.01fF
C8753 a_8525_n4317# a_8418_n5405# 0.00fF
C8754 a_690_n11933# a_600_n13591# 0.00fF
C8755 a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.00fF
C8756 a_3077_n3621# a_3436_n3799# 0.05fF
C8757 a_8162_n509# VDD 0.79fF
C8758 a_8418_n4317# a_8525_n5405# 0.00fF
C8759 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_4298_n1597# 0.00fF
C8760 a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C8761 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VDD 0.83fF
C8762 a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C8763 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_4298_n4317# 0.01fF
C8764 sky130_fd_sc_hd__clkinv_4_4/A a_8588_n5975# 0.11fF
C8765 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_6012_n3255# 0.03fF
C8766 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C8767 a_5586_n13021# a_5653_n12325# 0.01fF
C8768 a_434_n2685# a_600_n3255# 0.04fF
C8769 a_690_n2685# a_501_n2997# 0.02fF
C8770 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.09fF
C8771 VDD a_7130_n11933# 0.47fF
C8772 a_8588_n3799# a_8588_n3255# 0.09fF
C8773 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.02fF
C8774 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n9213# 0.01fF
C8775 a_8229_n1909# a_8328_n3255# 0.00fF
C8776 a_8328_n2167# a_8229_n2997# 0.00fF
C8777 a_10738_n1597# a_10805_n2997# 0.00fF
C8778 p2 sky130_fd_sc_hd__nand2_4_3/A 0.34fF
C8779 a_5653_n10613# a_7040_n10871# 0.01fF
C8780 a_5752_n10871# a_6941_n10613# 0.01fF
C8781 a_7237_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C8782 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_7300_n4887# 0.00fF
C8783 a_9813_n10301# a_10994_n10301# 0.01fF
C8784 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_10738_n10301# 0.35fF
C8785 a_9706_n10301# a_11101_n10301# 0.01fF
C8786 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A p2 0.04fF
C8787 Bd_b a_4986_n7215# 0.01fF
C8788 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.04fF
C8789 a_3373_n13021# a_3373_n11933# 0.02fF
C8790 a_600_n5975# a_690_n5405# 0.01fF
C8791 a_690_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.05fF
C8792 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_1978_n13021# 0.00fF
C8793 a_6012_n2167# a_5949_n2685# 0.01fF
C8794 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VDD 0.89fF
C8795 a_2148_n12503# a_2085_n11933# 0.01fF
C8796 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3266_n2685# 0.03fF
C8797 a_2085_n2685# a_3373_n2685# 0.01fF
C8798 a_1978_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C8799 a_10805_n13413# a_10738_n13789# 0.03fF
C8800 a_10738_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C8801 a_5653_n2997# a_5752_n2167# 0.00fF
C8802 a_3266_n5405# a_3436_n4887# 0.04fF
C8803 a_3436_n2167# a_4365_n1909# 0.02fF
C8804 a_3373_n11933# VDD 0.35fF
C8805 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10805_n2997# 0.00fF
C8806 a_3077_n11237# a_3010_n13021# 0.00fF
C8807 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.06fF
C8808 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8588_n13591# 0.03fF
C8809 a_8525_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C8810 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkinv_4_8/A 0.02fF
C8811 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_5/A 1.46fF
C8812 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.04fF
C8813 a_1789_n12325# a_1789_n11237# 0.02fF
C8814 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C8815 a_3010_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C8816 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n11933# 0.00fF
C8817 a_9813_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C8818 sky130_fd_sc_hd__nand2_4_3/B a_9876_n9783# 0.00fF
C8819 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10805_n2997# 0.01fF
C8820 a_7130_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C8821 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8418_n1597# 0.03fF
C8822 a_1888_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C8823 a_7237_n1597# a_8525_n1597# 0.01fF
C8824 a_13765_n12477# a_13765_n13021# 0.34fF
C8825 a_8229_n11237# a_8328_n9783# 0.00fF
C8826 a_7130_n4317# a_8525_n4317# 0.01fF
C8827 a_7237_n4317# a_8418_n4317# 0.01fF
C8828 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8162_n4317# 0.35fF
C8829 a_1978_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C8830 a_2085_n4317# a_3373_n4317# 0.01fF
C8831 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3266_n4317# 0.03fF
C8832 a_9813_n8125# a_10738_n8125# 0.01fF
C8833 a_5752_n3799# a_5949_n4317# 0.02fF
C8834 a_1888_n1079# VDD 0.49fF
C8835 a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C8836 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_4365_n3621# 0.18fF
C8837 a_3436_n3799# a_4464_n3799# 0.02fF
C8838 a_3176_n3799# a_4724_n3799# 0.01fF
C8839 a_7300_n11415# a_7237_n10301# 0.00fF
C8840 a_4724_n3255# a_4661_n1597# 0.00fF
C8841 a_2729_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.12fF
C8842 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_9876_n11415# 0.01fF
C8843 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C8844 a_860_n3255# a_860_n4887# 0.01fF
C8845 a_4365_n2997# a_4365_n4709# 0.00fF
C8846 a_4365_n13413# a_4554_n13021# 0.02fF
C8847 a_4724_n3255# a_4661_n4317# 0.00fF
C8848 a_4464_n13591# a_4298_n13021# 0.04fF
C8849 a_8525_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C8850 a_5653_n5797# a_7040_n5975# 0.01fF
C8851 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8588_n11415# 0.00fF
C8852 a_5752_n5975# a_6941_n5797# 0.01fF
C8853 a_4724_n10871# a_4724_n12503# 0.01fF
C8854 a_3176_n12503# a_3077_n13413# 0.00fF
C8855 a_3077_n12325# a_3176_n13591# 0.00fF
C8856 sky130_fd_sc_hd__clkinv_4_4/A a_6665_n7459# 0.02fF
C8857 a_434_n11933# a_797_n11933# 0.05fF
C8858 a_9813_n6493# a_10738_n6173# 0.01fF
C8859 VDD a_8525_n11933# 0.35fF
C8860 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.00fF
C8861 a_9450_n9213# VDD 0.75fF
C8862 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.06fF
C8863 a_7040_n1079# a_8229_n821# 0.01fF
C8864 a_6941_n821# a_8328_n1079# 0.01fF
C8865 a_7130_n1597# a_7040_n2167# 0.02fF
C8866 a_4554_n1597# a_4464_n2167# 0.02fF
C8867 a_5752_n9783# a_5842_n10301# 0.01fF
C8868 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.06fF
C8869 a_7237_n6493# sky130_fd_sc_hd__clkinv_1_5/A 0.00fF
C8870 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_8418_n5405# 0.01fF
C8871 a_10738_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.02fF
C8872 a_6941_n10613# a_7300_n10871# 0.05fF
C8873 a_9813_n5405# a_8525_n5405# 0.01fF
C8874 a_6012_n2167# a_6012_n3255# 0.02fF
C8875 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A a_434_n4317# 0.01fF
C8876 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A VDD 0.89fF
C8877 a_9450_n6493# a_9450_n5405# 0.02fF
C8878 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_10904_n3255# 0.02fF
C8879 a_5949_n4317# a_6012_n3799# 0.01fF
C8880 a_11101_n4317# a_11164_n3255# 0.00fF
C8881 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VDD 0.88fF
C8882 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VDD 0.83fF
C8883 a_4365_n12325# a_4365_n10613# 0.00fF
C8884 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.04fF
C8885 a_9517_n1909# a_9450_n2685# 0.01fF
C8886 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_7300_n3799# 0.00fF
C8887 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_2085_n9213# 0.00fF
C8888 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C8889 a_7237_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C8890 a_3373_n10301# a_3373_n11933# 0.01fF
C8891 a_3373_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.12fF
C8892 a_8525_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.12fF
C8893 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C8894 a_8418_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.05fF
C8895 a_3373_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.12fF
C8896 a_5653_n1909# a_6941_n1909# 0.01fF
C8897 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.08fF
C8898 a_10904_n5975# sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C8899 a_690_n10301# a_600_n8695# 0.00fF
C8900 a_3077_n11237# a_3010_n10301# 0.00fF
C8901 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.00fF
C8902 a_3436_n1079# VDD 0.79fF
C8903 a_4464_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.03fF
C8904 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.03fF
C8905 p2d sky130_fd_sc_hd__nand2_4_3/Y 0.01fF
C8906 a_4298_n5405# VDD 0.76fF
C8907 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_5752_n3799# 0.01fF
C8908 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C8909 a_9517_n13413# a_9450_n11933# 0.00fF
C8910 a_10994_n11933# a_10904_n11415# 0.02fF
C8911 a_600_n10871# a_690_n9213# 0.00fF
C8912 a_4464_n10871# VDD 0.46fF
C8913 a_11101_n1597# VDD 0.32fF
C8914 a_8525_n10301# VDD 0.35fF
C8915 a_6941_n5797# a_7300_n5975# 0.05fF
C8916 a_434_n11933# a_1978_n11933# 0.01fF
C8917 a_690_n11933# a_1722_n11933# 0.02fF
C8918 a_1789_n10613# a_3077_n10613# 0.01fF
C8919 a_7040_n8695# a_7212_n7203# 0.00fF
C8920 a_8525_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.00fF
C8921 a_1789_n8437# a_1789_n9525# 0.02fF
C8922 a_8588_n11415# a_8418_n10301# 0.00fF
C8923 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X a_6874_n10301# 0.03fF
C8924 a_8229_n821# a_8588_n1079# 0.05fF
C8925 a_8162_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C8926 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5653_n1909# 0.01fF
C8927 a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C8928 a_5586_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.03fF
C8929 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_7300_n8695# 0.01fF
C8930 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.01fF
C8931 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.04fF
C8932 a_7130_n2685# a_7237_n4317# 0.00fF
C8933 a_7237_n2685# a_7130_n4317# 0.00fF
C8934 a_7300_n10871# a_8328_n10871# 0.02fF
C8935 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_8229_n10613# 0.18fF
C8936 a_1978_n2685# a_2085_n4317# 0.00fF
C8937 a_2085_n2685# a_1978_n4317# 0.00fF
C8938 a_501_n5797# a_600_n4887# 0.00fF
C8939 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C8940 a_600_n5975# a_501_n4709# 0.00fF
C8941 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X a_860_n3799# 0.01fF
C8942 a_11164_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.03fF
C8943 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.04fF
C8944 a_9517_n11237# a_9450_n11933# 0.01fF
C8945 a_8328_n4887# a_8229_n3621# 0.00fF
C8946 a_4623_n7349# Bd_b 0.43fF
C8947 a_8229_n4709# a_8328_n3799# 0.00fF
C8948 a_5752_n1079# VDD 0.46fF
C8949 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.06fF
C8950 a_4661_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C8951 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_4724_n4887# 0.03fF
C8952 sky130_fd_sc_hd__clkinv_4_1/Y B_b 0.04fF
C8953 a_9876_n3799# a_9876_n3255# 0.09fF
C8954 a_4464_n11415# a_4554_n13021# 0.00fF
C8955 a_6874_n13021# a_8162_n13021# 0.01fF
C8956 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.02fF
C8957 a_1722_n5405# VDD 0.76fF
C8958 a_3176_n12503# a_3176_n11415# 0.01fF
C8959 a_860_n8695# VDD 0.81fF
C8960 sky130_fd_sc_hd__nand2_4_2/A a_2622_n14109# 0.03fF
C8961 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.02fF
C8962 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/X 0.04fF
C8963 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C8964 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.02fF
C8965 a_600_n11415# a_434_n10301# 0.00fF
C8966 a_501_n11237# a_690_n10301# 0.00fF
C8967 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.02fF
C8968 a_6941_n1909# a_7040_n2167# 0.49fF
C8969 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_501_n13413# 0.18fF
C8970 a_8525_n509# a_9706_n509# 0.01fF
C8971 a_8418_n509# a_9813_n509# 0.01fF
C8972 a_434_n2685# a_690_n2685# 0.19fF
C8973 a_1722_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.00fF
C8974 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD 0.84fF
C8975 a_5586_n5405# a_6874_n5405# 0.01fF
C8976 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.04fF
C8977 a_5842_n5405# VDD 0.47fF
C8978 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.63fF
C8979 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.04fF
C8980 a_9517_n4709# a_9450_n4317# 0.01fF
C8981 sky130_fd_sc_hd__clkinv_4_7/Y p1_b 0.04fF
C8982 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_1722_n9213# 0.00fF
C8983 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C8984 a_6012_n10871# VDD 0.78fF
C8985 a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C8986 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VDD 0.85fF
C8987 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X a_8229_n5797# 0.18fF
C8988 a_9450_n14109# VDD 0.75fF
C8989 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD 0.91fF
C8990 a_7040_n5975# a_8588_n5975# 0.01fF
C8991 a_7300_n5975# a_8328_n5975# 0.02fF
C8992 a_3077_n10613# a_3176_n10871# 0.49fF
C8993 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C8994 a_8229_n9525# a_8328_n9783# 0.49fF
C8995 a_10904_n4887# a_10738_n5405# 0.04fF
C8996 a_10805_n4709# a_10994_n5405# 0.02fF
C8997 a_4365_n10613# a_4298_n10301# 0.01fF
C8998 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6101_n7254# 0.00fF
C8999 a_4554_n9213# a_5586_n9213# 0.02fF
C9000 a_4298_n9213# a_5842_n9213# 0.01fF
C9001 a_7237_n5405# sky130_fd_sc_hd__clkinv_4_3/A 0.05fF
C9002 a_n787_n9525# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C9003 a_7300_n9783# a_7237_n10301# 0.01fF
C9004 a_9517_n11237# a_9450_n10301# 0.00fF
C9005 a_5949_n1597# a_6012_n2167# 0.01fF
C9006 sky130_fd_sc_hd__dfxbp_1_1/D a_n1738_n6671# 0.10fF
C9007 a_6941_n2997# VDD 0.35fF
C9008 a_501_n10613# a_600_n10871# 0.49fF
C9009 a_n2602_n7037# a_n1139_n6715# 0.03fF
C9010 a_434_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X 0.01fF
C9011 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C9012 a_7040_n8695# a_7300_n8695# 0.28fF
C9013 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.04fF
C9014 a_10904_n2167# a_11101_n2685# 0.02fF
C9015 a_11164_n2167# a_10994_n2685# 0.04fF
C9016 a_6012_n5975# VDD 0.77fF
C9017 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.01fF
C9018 a_10805_n1909# sky130_fd_sc_hd__nand2_4_0/Y 0.08fF
C9019 a_3077_n5797# sky130_fd_sc_hd__clkinv_4_4/A 0.07fF
C9020 a_7300_n1079# VDD 0.78fF
C9021 a_10904_n13591# a_10738_n13021# 0.04fF
C9022 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.08fF
C9023 a_10805_n2997# a_9517_n2997# 0.01fF
C9024 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_2085_n13021# 0.02fF
C9025 a_797_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C9026 a_8162_n13021# a_8418_n13021# 0.19fF
C9027 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.02fF
C9028 a_600_n11415# VDD 0.44fF
C9029 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.02fF
C9030 a_7130_n14109# a_8418_n14109# 0.01fF
C9031 a_7237_n14109# a_8162_n14109# 0.02fF
C9032 a_6874_n14109# a_8525_n14109# 0.00fF
C9033 a_11164_n2167# sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C9034 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_600_n3799# 0.00fF
C9035 a_2148_n3799# a_860_n3799# 0.01fF
C9036 a_9813_n11933# a_11101_n11933# 0.01fF
C9037 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10994_n11933# 0.03fF
C9038 sky130_fd_sc_hd__nand2_4_2/A a_7237_n14109# 0.02fF
C9039 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_797_n5405# 0.01fF
C9040 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.00fF
C9041 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.04fF
C9042 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C9043 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_1_5/A 0.02fF
C9044 a_5586_n13021# a_5842_n13021# 0.19fF
C9045 a_4554_n4317# a_4724_n4887# 0.04fF
C9046 a_4661_n4317# a_4464_n4887# 0.02fF
C9047 a_5586_n5405# a_5586_n4317# 0.02fF
C9048 a_7130_n8125# sky130_fd_sc_hd__clkinv_1_5/A 0.02fF
C9049 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X a_6012_n4887# 0.00fF
C9050 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C9051 a_797_n2685# a_1722_n2685# 0.02fF
C9052 a_434_n2685# a_2085_n2685# 0.00fF
C9053 a_5842_n10301# a_5949_n9213# 0.00fF
C9054 a_11101_n13021# VDD 0.32fF
C9055 a_690_n2685# a_1978_n2685# 0.01fF
C9056 a_600_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.03fF
C9057 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C9058 a_1888_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C9059 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.69fF
C9060 a_1722_n11933# a_3266_n11933# 0.01fF
C9061 a_1978_n11933# a_3010_n11933# 0.02fF
C9062 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C9063 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C9064 a_5752_n11415# a_5752_n12503# 0.01fF
C9065 a_9616_n3255# VDD 0.45fF
C9066 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A VDD 0.66fF
C9067 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VDD 0.83fF
C9068 a_3436_n10871# a_4365_n10613# 0.02fF
C9069 a_434_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.04fF
C9070 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_434_n11933# 0.01fF
C9071 a_501_n1909# a_n787_n1909# 0.01fF
C9072 a_2148_n9783# a_2085_n9213# 0.01fF
C9073 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X a_8525_n14109# 0.00fF
C9074 a_8229_n9525# a_9876_n9783# 0.00fF
C9075 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C9076 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.04fF
C9077 a_9706_n13021# a_9813_n11933# 0.00fF
C9078 a_8162_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.07fF
C9079 a_13765_n5405# a_13765_n5949# 0.31fF
C9080 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.04fF
C9081 a_9876_n8695# a_10904_n8695# 0.02fF
C9082 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_10805_n8437# 0.17fF
C9083 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C9084 a_6941_n5797# a_6865_n7304# 0.01fF
C9085 a_7300_n5975# a_6658_n7363# 0.00fF
C9086 a_9616_n8695# a_11164_n8695# 0.01fF
C9087 a_7040_n5975# a_6665_n7459# 0.00fF
C9088 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkinv_4_3/A 0.44fF
C9089 a_860_n4887# a_n787_n4709# 0.00fF
C9090 a_8229_n11237# a_8229_n10613# 0.05fF
C9091 a_5842_n4317# a_5653_n5797# 0.00fF
C9092 a_5586_n4317# a_5752_n5975# 0.00fF
C9093 a_5586_n10301# a_6874_n10301# 0.01fF
C9094 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.29fF
C9095 a_4554_n10301# a_4724_n8695# 0.00fF
C9096 a_4661_n10301# a_4464_n8695# 0.00fF
C9097 a_8328_n3255# VDD 0.46fF
C9098 a_501_n10613# a_2148_n10871# 0.00fF
C9099 a_7040_n8695# a_7130_n10301# 0.00fF
C9100 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_8328_n8695# 0.05fF
C9101 a_7300_n8695# a_8588_n8695# 0.01fF
C9102 a_7040_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.00fF
C9103 clk a_n2248_n7037# 0.01fF
C9104 a_9450_n8125# a_9706_n8125# 0.19fF
C9105 a_7130_n5405# a_7040_n5975# 0.01fF
C9106 a_13765_n2141# Bd_b 0.12fF
C9107 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD 0.84fF
C9108 a_2622_n14109# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C9109 a_4464_n5975# sky130_fd_sc_hd__clkinv_4_4/A 0.07fF
C9110 a_9517_n10613# a_9706_n11933# 0.00fF
C9111 a_9616_n10871# a_9450_n11933# 0.00fF
C9112 a_434_n9213# a_600_n9783# 0.04fF
C9113 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.00fF
C9114 a_690_n9213# a_501_n9525# 0.02fF
C9115 a_7237_n8125# a_7212_n7203# 0.02fF
C9116 a_8525_n13021# a_9450_n13021# 0.02fF
C9117 a_8418_n13021# a_9706_n13021# 0.01fF
C9118 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.08fF
C9119 a_4724_n8695# Ad_b 0.00fF
C9120 a_4298_n11933# a_5842_n11933# 0.01fF
C9121 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C9122 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.02fF
C9123 a_2148_n2167# a_2148_n3255# 0.02fF
C9124 a_11101_n11933# sky130_fd_sc_hd__clkinv_4_8/A 0.01fF
C9125 a_n688_n9783# a_501_n9525# 0.01fF
C9126 a_4623_n7349# a_5052_n7283# 0.04fF
C9127 a_n787_n9525# a_600_n9783# 0.01fF
C9128 a_11101_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.01fF
C9129 a_5586_n13021# a_7237_n13021# 0.00fF
C9130 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.02fF
C9131 a_600_n1079# a_1888_n1079# 0.01fF
C9132 a_4365_n4709# a_5653_n4709# 0.01fF
C9133 a_10805_n12325# VDD 0.32fF
C9134 a_9876_n10871# a_9876_n9783# 0.02fF
C9135 a_7130_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.05fF
C9136 a_4365_n3621# a_4554_n5405# 0.00fF
C9137 a_1722_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.03fF
C9138 a_4464_n3799# a_4298_n5405# 0.00fF
C9139 a_1978_n2685# a_2085_n2685# 0.55fF
C9140 sky130_fd_sc_hd__nand2_4_3/B VDD 1.28fF
C9141 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.06fF
C9142 a_9616_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C9143 sky130_fd_sc_hd__nand2_4_1/A Bd_b 0.66fF
C9144 a_9450_n1597# a_9517_n821# 0.01fF
C9145 a_3010_n11933# a_3373_n11933# 0.05fF
C9146 a_10904_n4887# a_10994_n4317# 0.01fF
C9147 a_11164_n3255# VDD 0.67fF
C9148 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.02fF
C9149 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkinv_4_3/A 0.06fF
C9150 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3077_n4709# 0.01fF
C9151 a_797_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.00fF
C9152 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_860_n3799# 0.01fF
C9153 a_690_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.05fF
C9154 a_3010_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C9155 a_6874_n4317# a_6941_n2997# 0.00fF
C9156 a_9706_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.07fF
C9157 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A a_2148_n4887# 0.00fF
C9158 a_6874_n1597# VDD 0.76fF
C9159 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_8328_n1079# 0.03fF
C9160 a_1789_n2997# a_1789_n4709# 0.00fF
C9161 a_9616_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C9162 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C9163 a_10738_n13021# sky130_fd_sc_hd__clkinv_4_7/Y 0.00fF
C9164 a_797_n4317# VDD 0.35fF
C9165 a_6874_n10301# a_7130_n10301# 0.19fF
C9166 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C9167 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_860_n3255# 0.01fF
C9168 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C9169 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.02fF
C9170 a_6874_n11933# a_8418_n11933# 0.01fF
C9171 a_7130_n11933# a_8162_n11933# 0.02fF
C9172 a_5653_n3621# a_5842_n2685# 0.00fF
C9173 a_5752_n3799# a_5586_n2685# 0.00fF
C9174 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.07fF
C9175 a_2729_n509# sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C9176 a_9517_n10613# a_9706_n10301# 0.02fF
C9177 a_9616_n10871# a_9450_n10301# 0.04fF
C9178 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C9179 a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C9180 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_4298_n10301# 0.01fF
C9181 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X a_8162_n10301# 0.00fF
C9182 a_797_n1597# a_860_n1079# 0.01fF
C9183 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.29fF
C9184 a_8162_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.03fF
C9185 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8229_n5797# 0.01fF
C9186 a_1789_n4709# a_1722_n4317# 0.01fF
C9187 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.02fF
C9188 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C9189 a_3077_n10613# a_3077_n9525# 0.02fF
C9190 a_8229_n13413# VDD 0.35fF
C9191 a_8162_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C9192 a_7300_n12503# a_7300_n13591# 0.02fF
C9193 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/X 0.09fF
C9194 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X Ad_b 0.02fF
C9195 a_5586_n11933# a_5949_n11933# 0.05fF
C9196 a_501_n1909# a_2148_n2167# 0.00fF
C9197 a_600_n2167# a_1888_n2167# 0.01fF
C9198 a_8229_n8437# a_8418_n10301# 0.00fF
C9199 a_8328_n9783# a_8418_n9213# 0.02fF
C9200 a_860_n2167# a_1789_n1909# 0.02fF
C9201 a_7300_n8695# a_7237_n8125# 0.01fF
C9202 a_5949_n5405# VDD 0.34fF
C9203 a_501_n10613# a_501_n9525# 0.02fF
C9204 a_6874_n2685# a_5586_n2685# 0.01fF
C9205 a_6941_n12325# a_8229_n12325# 0.01fF
C9206 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C9207 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_3077_n821# 0.01fF
C9208 a_5653_n4709# a_5752_n4887# 0.49fF
C9209 a_1789_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C9210 a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.02fF
C9211 p1d VDD 4.21fF
C9212 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C9213 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8525_n2685# 0.02fF
C9214 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_8588_n12503# 0.00fF
C9215 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C9216 a_797_n13021# a_860_n13591# 0.01fF
C9217 a_3373_n11933# a_4554_n11933# 0.01fF
C9218 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4298_n11933# 0.35fF
C9219 a_8229_n11237# VDD 0.35fF
C9220 a_3266_n11933# a_4661_n11933# 0.01fF
C9221 a_7300_n11415# a_7300_n12503# 0.02fF
C9222 a_1789_n3621# VDD 0.35fF
C9223 A a_13765_n4317# 0.02fF
C9224 a_13765_n5949# Ad_b 0.12fF
C9225 a_797_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C9226 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_2085_n10301# 0.02fF
C9227 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.08fF
C9228 a_7130_n14109# a_7040_n13591# 0.02fF
C9229 a_501_n11237# a_690_n11933# 0.02fF
C9230 a_600_n11415# a_434_n11933# 0.04fF
C9231 a_9616_n8695# a_9517_n9525# 0.00fF
C9232 a_9517_n8437# a_9616_n9783# 0.00fF
C9233 a_4464_n9783# a_4554_n9213# 0.02fF
C9234 a_5653_n3621# a_5752_n3255# 0.01fF
C9235 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X a_8588_n1079# 0.00fF
C9236 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_3436_n10871# 0.01fF
C9237 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.01fF
C9238 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A 0.53fF
C9239 a_6658_n7363# a_6865_n7304# 0.54fF
C9240 a_9517_n5797# a_9706_n4317# 0.00fF
C9241 a_2085_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C9242 a_6101_n7254# p2 0.01fF
C9243 a_6373_n7349# a_6794_n7203# 0.10fF
C9244 a_7237_n10301# a_8162_n10301# 0.02fF
C9245 a_7237_n4317# a_7040_n5975# 0.00fF
C9246 a_7130_n4317# a_7300_n5975# 0.00fF
C9247 a_9616_n5975# a_9450_n4317# 0.00fF
C9248 a_8162_n11933# a_8525_n11933# 0.05fF
C9249 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6012_n8695# 0.00fF
C9250 a_5949_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.00fF
C9251 a_4724_n11415# a_4661_n10301# 0.00fF
C9252 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/A 0.47fF
C9253 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.02fF
C9254 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C9255 a_7040_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.07fF
C9256 a_10994_n5405# a_10904_n5975# 0.01fF
C9257 a_8525_n5405# a_8588_n5975# 0.01fF
C9258 a_13765_n13565# VDD 2.05fF
C9259 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C9260 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_9813_n9213# 0.00fF
C9261 a_9876_n12503# a_9876_n11415# 0.02fF
C9262 sky130_fd_sc_hd__nand2_4_3/Y a_11101_n10301# 0.01fF
C9263 a_11164_n2167# a_11164_n3799# 0.01fF
C9264 a_6794_n7203# VDD 0.33fF
C9265 a_1978_n9213# a_2148_n9783# 0.04fF
C9266 a_4464_n5975# a_5653_n5797# 0.01fF
C9267 a_4365_n5797# a_5752_n5975# 0.01fF
C9268 a_9616_n13591# VDD 0.42fF
C9269 a_8328_n2167# a_8418_n509# 0.00fF
C9270 a_8229_n9525# a_8229_n10613# 0.02fF
C9271 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Bd_b 0.05fF
C9272 a_2148_n5975# a_860_n5975# 0.01fF
C9273 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_600_n5975# 0.00fF
C9274 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_9450_n9213# 0.03fF
C9275 a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C9276 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.08fF
C9277 a_9450_n6493# sky130_fd_sc_hd__clkinv_4_3/A 0.01fF
C9278 a_1888_n11415# a_1888_n9783# 0.00fF
C9279 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_3077_n1909# 0.01fF
C9280 a_1888_n1079# a_3077_n821# 0.01fF
C9281 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VDD 0.88fF
C9282 a_6874_n5405# a_7237_n5405# 0.05fF
C9283 a_3010_n1597# a_3010_n2685# 0.02fF
C9284 a_8229_n12325# a_8328_n12503# 0.49fF
C9285 sky130_fd_sc_hd__nand2_1_0/A a_n428_n4887# 0.02fF
C9286 a_2366_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C9287 a_6012_n4887# a_6941_n4709# 0.02fF
C9288 a_n2248_n7037# sky130_fd_sc_hd__clkinv_1_5/A 0.01fF
C9289 a_5752_n4887# a_7040_n4887# 0.01fF
C9290 a_690_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_43/A 0.05fF
C9291 a_3436_n3255# a_3373_n2685# 0.01fF
C9292 a_7237_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.12fF
C9293 a_3077_n2997# a_3176_n3255# 0.49fF
C9294 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C9295 a_10805_n1909# VDD 0.32fF
C9296 a_10805_n13413# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C9297 a_4554_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.05fF
C9298 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6941_n3621# 0.00fF
C9299 a_5752_n10871# a_5842_n9213# 0.00fF
C9300 a_n428_n12503# sky130_fd_sc_hd__nand2_1_4/B 0.14fF
C9301 a_7300_n4887# a_5752_n4887# 0.01fF
C9302 a_4365_n11237# a_4298_n11933# 0.01fF
C9303 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_5586_n9213# 0.03fF
C9304 a_8418_n4317# a_8328_n3255# 0.01fF
C9305 a_797_n11933# a_797_n13021# 0.02fF
C9306 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkinv_1_3/A 0.05fF
C9307 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.02fF
C9308 a_2085_n1597# a_1888_n1079# 0.02fF
C9309 a_1978_n1597# a_2148_n1079# 0.04fF
C9310 a_8525_n11933# a_9706_n11933# 0.01fF
C9311 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_9450_n11933# 0.35fF
C9312 a_9616_n10871# a_8328_n10871# 0.01fF
C9313 a_9876_n10871# a_8229_n10613# 0.00fF
C9314 a_5842_n13021# a_6012_n13591# 0.04fF
C9315 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkinv_1_3/A 0.84fF
C9316 a_10904_n10871# a_11101_n10301# 0.02fF
C9317 a_11164_n10871# a_10994_n10301# 0.04fF
C9318 a_8588_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.12fF
C9319 a_3176_n4887# a_3266_n4317# 0.01fF
C9320 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VDD 2.18fF
C9321 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_434_n10301# 0.00fF
C9322 a_4464_n10871# a_4554_n11933# 0.01fF
C9323 a_n2163_n6671# a_n1139_n6715# 0.02fF
C9324 a_n1995_n6925# a_n2248_n7037# 0.03fF
C9325 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.03fF
C9326 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X a_8525_n10301# 0.01fF
C9327 a_n1570_n6769# a_n1738_n6671# 0.53fF
C9328 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.04fF
C9329 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_9450_n509# 0.00fF
C9330 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_9616_n11415# 0.01fF
C9331 a_5752_n13591# a_5586_n11933# 0.00fF
C9332 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A VDD 0.88fF
C9333 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.01fF
C9334 a_9813_n6493# sky130_fd_sc_hd__nand2_4_1/B 0.13fF
C9335 a_9616_n2167# a_9517_n821# 0.00fF
C9336 a_9517_n1909# a_9616_n1079# 0.00fF
C9337 a_6874_n2685# a_7040_n3255# 0.04fF
C9338 a_7130_n2685# a_6941_n2997# 0.02fF
C9339 a_7237_n5405# a_8418_n5405# 0.01fF
C9340 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8162_n5405# 0.35fF
C9341 a_3077_n821# a_3436_n1079# 0.05fF
C9342 a_7130_n5405# a_8525_n5405# 0.01fF
C9343 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C9344 a_5949_n13021# a_5752_n11415# 0.00fF
C9345 a_5842_n13021# a_6012_n11415# 0.00fF
C9346 Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.02fF
C9347 a_860_n4887# a_1789_n4709# 0.02fF
C9348 a_600_n4887# a_1888_n4887# 0.01fF
C9349 a_501_n4709# a_2148_n4887# 0.00fF
C9350 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_2085_n1597# 0.02fF
C9351 a_8162_n6493# a_8229_n5797# 0.01fF
C9352 a_1888_n5975# VDD 0.47fF
C9353 a_797_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.01fF
C9354 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.04fF
C9355 a_7237_n2685# a_7040_n1079# 0.00fF
C9356 a_7130_n2685# a_7300_n1079# 0.00fF
C9357 a_3077_n2997# a_4724_n3255# 0.00fF
C9358 a_3436_n3255# a_4365_n2997# 0.02fF
C9359 Ad_b sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C9360 a_3176_n3255# a_4464_n3255# 0.01fF
C9361 a_3077_n3621# a_1789_n3621# 0.01fF
C9362 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.04fF
C9363 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_797_n2685# 0.01fF
C9364 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.03fF
C9365 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.04fF
C9366 a_13765_n5405# a_13765_n4861# 0.34fF
C9367 a_10738_n1597# a_11101_n1597# 0.05fF
C9368 a_7237_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.12fF
C9369 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1722_n11933# 0.01fF
C9370 a_8328_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C9371 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_7040_n4887# 0.03fF
C9372 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.06fF
C9373 a_600_n3255# a_860_n3255# 0.28fF
C9374 a_501_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.02fF
C9375 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.06fF
C9376 a_9450_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C9377 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9517_n2997# 0.00fF
C9378 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n11933# 0.00fF
C9379 a_7040_n10871# a_7130_n11933# 0.01fF
C9380 a_2366_n8125# a_2729_n8125# 0.05fF
C9381 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Bd_b 0.03fF
C9382 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_8418_n9213# 0.01fF
C9383 a_9813_n9213# a_8525_n9213# 0.01fF
C9384 a_11164_n5975# a_10994_n4317# 0.00fF
C9385 a_10904_n5975# a_11101_n4317# 0.00fF
C9386 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8588_n5975# 0.00fF
C9387 a_10805_n5797# sky130_fd_sc_hd__clkinv_4_3/A 0.02fF
C9388 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.02fF
C9389 a_8229_n9525# VDD 0.35fF
C9390 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VDD 0.73fF
C9391 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.29fF
C9392 a_8418_n509# a_8229_n821# 0.02fF
C9393 a_8162_n509# a_8328_n1079# 0.04fF
C9394 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkinv_1_3/A 0.82fF
C9395 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.04fF
C9396 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.04fF
C9397 a_5586_n4317# a_5949_n4317# 0.05fF
C9398 a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C9399 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_5586_n11933# 0.01fF
C9400 a_10805_n4709# VDD 0.32fF
C9401 a_797_n11933# a_797_n10301# 0.01fF
C9402 a_6874_n13021# a_6941_n12325# 0.01fF
C9403 a_7237_n4317# a_7130_n5405# 0.00fF
C9404 a_7130_n4317# a_7237_n5405# 0.00fF
C9405 clk a_n2436_n7037# 0.07fF
C9406 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C9407 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_9876_n11415# 0.03fF
C9408 a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C9409 a_600_n2167# a_501_n821# 0.00fF
C9410 a_3436_n11415# a_3436_n9783# 0.01fF
C9411 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.04fF
C9412 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_9706_n5405# 0.00fF
C9413 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C9414 a_4365_n9525# a_4365_n11237# 0.00fF
C9415 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_10738_n9213# 0.03fF
C9416 sky130_fd_sc_hd__clkinv_4_4/A a_6012_n5975# 0.11fF
C9417 a_3176_n1079# a_4724_n1079# 0.01fF
C9418 a_8418_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.05fF
C9419 a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C9420 a_3436_n1079# a_4464_n1079# 0.02fF
C9421 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_4365_n821# 0.18fF
C9422 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_11164_n4887# 0.03fF
C9423 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.00fF
C9424 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_3077_n4709# 0.01fF
C9425 VDD a_3373_n9213# 0.35fF
C9426 a_3176_n2167# a_3373_n2685# 0.02fF
C9427 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.08fF
C9428 a_3436_n5975# VDD 0.79fF
C9429 a_3436_n2167# a_3266_n2685# 0.04fF
C9430 a_9616_n2167# a_9706_n509# 0.00fF
C9431 a_4464_n3255# a_4724_n3255# 0.28fF
C9432 a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.02fF
C9433 a_7300_n3799# a_7300_n3255# 0.09fF
C9434 a_3077_n1909# a_3077_n2997# 0.02fF
C9435 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_5653_n2997# 0.01fF
C9436 sky130_fd_sc_hd__nand2_4_3/Y a_6665_n7459# 0.01fF
C9437 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n9213# 0.01fF
C9438 a_3010_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C9439 a_4464_n10871# a_5653_n10613# 0.01fF
C9440 a_8525_n10301# a_9706_n10301# 0.01fF
C9441 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n10301# 0.35fF
C9442 a_9876_n10871# VDD 0.74fF
C9443 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C9444 a_4464_n9783# a_4464_n10871# 0.01fF
C9445 a_2085_n13021# a_2085_n11933# 0.02fF
C9446 a_4724_n2167# a_4661_n2685# 0.01fF
C9447 a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C9448 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C9449 a_8328_n10871# a_8162_n9213# 0.00fF
C9450 a_8229_n10613# a_8418_n9213# 0.00fF
C9451 a_8162_n6493# VDD 0.78fF
C9452 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X a_8162_n11933# 0.01fF
C9453 a_4365_n2997# a_4464_n2167# 0.00fF
C9454 a_1789_n11237# a_1722_n13021# 0.00fF
C9455 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.06fF
C9456 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7300_n13591# 0.03fF
C9457 a_4365_n821# a_6012_n1079# 0.00fF
C9458 a_4724_n1079# a_5653_n821# 0.02fF
C9459 a_7237_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C9460 a_501_n8437# a_860_n8695# 0.05fF
C9461 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_2085_n5405# 0.00fF
C9462 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C9463 a_4464_n1079# a_5752_n1079# 0.01fF
C9464 a_600_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.03fF
C9465 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.04fF
C9466 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.02fF
C9467 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n11933# 0.00fF
C9468 a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C9469 a_9517_n5797# a_8229_n5797# 0.01fF
C9470 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6874_n4317# 0.35fF
C9471 sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13021# 0.04fF
C9472 a_5842_n4317# a_7237_n4317# 0.01fF
C9473 a_5949_n4317# a_7130_n4317# 0.01fF
C9474 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C9475 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_3/Y 0.05fF
C9476 a_9517_n4709# a_9450_n5405# 0.01fF
C9477 a_1888_n2167# a_1789_n2997# 0.00fF
C9478 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_501_n13413# 0.00fF
C9479 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__dfxbp_1_0/Q 0.01fF
C9480 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C9481 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C9482 a_6012_n11415# a_5949_n10301# 0.00fF
C9483 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.08fF
C9484 a_7130_n509# VDD 0.46fF
C9485 sky130_fd_sc_hd__nand2_1_4/Y a_3077_n8437# 0.00fF
C9486 a_3436_n3255# a_3373_n1597# 0.00fF
C9487 a_8418_n2685# a_8588_n3255# 0.04fF
C9488 a_8525_n2685# a_8328_n3255# 0.02fF
C9489 a_4464_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.03fF
C9490 a_3176_n13591# a_3010_n13021# 0.04fF
C9491 a_3436_n3255# a_3373_n4317# 0.00fF
C9492 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.85fF
C9493 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkinv_1_3/A 0.08fF
C9494 a_3077_n13413# a_3266_n13021# 0.02fF
C9495 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7300_n11415# 0.00fF
C9496 a_7237_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C9497 a_1888_n12503# a_1789_n13413# 0.00fF
C9498 a_1789_n12325# a_1888_n13591# 0.00fF
C9499 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.89fF
C9500 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_2366_n509# 0.00fF
C9501 a_10805_n1909# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C9502 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8588_n1079# 0.00fF
C9503 a_6874_n9213# VDD 0.76fF
C9504 VDD a_5949_n11933# 0.35fF
C9505 Ad_b a_13765_n4861# 0.22fF
C9506 a_5653_n821# a_7040_n1079# 0.01fF
C9507 a_5752_n1079# a_6941_n821# 0.01fF
C9508 a_13765_n4317# Ad 0.12fF
C9509 a_9517_n12325# a_9450_n11933# 0.01fF
C9510 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.06fF
C9511 a_10805_n11237# a_10904_n11415# 0.48fF
C9512 a_3373_n10301# a_3373_n9213# 0.02fF
C9513 sky130_fd_sc_hd__dfxbp_1_0/Q Ad_b 0.26fF
C9514 a_5653_n10613# a_6012_n10871# 0.05fF
C9515 a_9706_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.05fF
C9516 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_10994_n10301# 0.00fF
C9517 sky130_fd_sc_hd__clkinv_1_6/Y VDD 2.06fF
C9518 a_860_n11415# a_690_n13021# 0.00fF
C9519 a_501_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.18fF
C9520 a_4464_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.03fF
C9521 sky130_fd_sc_hd__clkinv_4_8/A a_6941_n12325# 0.08fF
C9522 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_797_n13021# 0.01fF
C9523 a_8162_n6493# a_8162_n5405# 0.02fF
C9524 a_3077_n12325# a_3077_n10613# 0.00fF
C9525 a_1722_n9213# VDD 0.76fF
C9526 a_9813_n4317# a_9876_n3255# 0.00fF
C9527 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VDD 0.88fF
C9528 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_4365_n1909# 0.01fF
C9529 a_5586_n5405# a_5752_n5975# 0.04fF
C9530 a_5842_n5405# a_5653_n5797# 0.02fF
C9531 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_6941_n821# 0.01fF
C9532 a_5949_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C9533 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6012_n3799# 0.00fF
C9534 a_4365_n8437# VDD 0.36fF
C9535 a_9450_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.07fF
C9536 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n2685# 0.01fF
C9537 a_9813_n2685# a_9876_n3255# 0.01fF
C9538 a_1888_n3255# a_1789_n3621# 0.01fF
C9539 a_2085_n10301# a_2085_n11933# 0.01fF
C9540 a_5653_n11237# a_5586_n11933# 0.01fF
C9541 a_7237_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.12fF
C9542 a_7130_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.05fF
C9543 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_8418_n4317# 0.00fF
C9544 a_2085_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.12fF
C9545 a_3010_n10301# a_3176_n8695# 0.00fF
C9546 a_3266_n10301# a_3077_n8437# 0.00fF
C9547 a_8418_n13021# a_8328_n12503# 0.02fF
C9548 a_1789_n11237# a_1722_n10301# 0.00fF
C9549 a_4554_n1597# a_3010_n1597# 0.01fF
C9550 a_4298_n1597# a_3266_n1597# 0.02fF
C9551 a_797_n11933# a_860_n13591# 0.00fF
C9552 a_3176_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.03fF
C9553 a_2148_n3799# a_1978_n4317# 0.04fF
C9554 a_8525_n509# VDD 0.35fF
C9555 a_8229_n13413# a_8162_n11933# 0.00fF
C9556 a_13765_n9213# sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C9557 a_5653_n5797# a_6012_n5975# 0.05fF
C9558 a_9517_n5797# VDD 0.34fF
C9559 a_797_n2685# a_600_n3255# 0.02fF
C9560 a_690_n2685# a_860_n3255# 0.04fF
C9561 a_6941_n3621# a_6941_n4709# 0.02fF
C9562 a_4365_n13413# VDD 0.35fF
C9563 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_434_n11933# 0.44fF
C9564 a_8418_n9213# VDD 0.44fF
C9565 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.88fF
C9566 a_6941_n821# a_7300_n1079# 0.05fF
C9567 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.09fF
C9568 a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C9569 a_6012_n10871# a_7040_n10871# 0.02fF
C9570 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_6941_n10613# 0.18fF
C9571 a_10994_n1597# a_10904_n3255# 0.00fF
C9572 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_1_5/A 0.37fF
C9573 a_5752_n10871# a_7300_n10871# 0.01fF
C9574 sky130_fd_sc_hd__clkinv_1_5/A a_7212_n7203# 0.28fF
C9575 a_9706_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.01fF
C9576 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_11101_n10301# 0.02fF
C9577 a_n2436_n7037# sky130_fd_sc_hd__clkinv_1_5/A 0.16fF
C9578 a_4298_n2685# VDD 0.76fF
C9579 sky130_fd_sc_hd__clkinv_4_8/A a_8328_n12503# 0.07fF
C9580 a_6012_n8695# a_6101_n7254# 0.00fF
C9581 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6006_n7607# 0.00fF
C9582 a_860_n5975# a_797_n5405# 0.01fF
C9583 a_8229_n11237# a_8162_n11933# 0.01fF
C9584 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C9585 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_2148_n4887# 0.00fF
C9586 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.04fF
C9587 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_9876_n3255# 0.00fF
C9588 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.06fF
C9589 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.06fF
C9590 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_8588_n1079# 0.01fF
C9591 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.02fF
C9592 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.02fF
C9593 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_3436_n4887# 0.03fF
C9594 a_3373_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C9595 a_9706_n6493# sky130_fd_sc_hd__clkinv_4_3/A 0.02fF
C9596 a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.01fF
C9597 a_600_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C9598 a_3176_n11415# a_3266_n13021# 0.00fF
C9599 a_11164_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.00fF
C9600 a_5752_n8695# VDD 0.47fF
C9601 a_1888_n12503# a_1888_n11415# 0.01fF
C9602 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.00fF
C9603 a_3077_n11237# VDD 0.35fF
C9604 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.02fF
C9605 p1d p1_b 0.53fF
C9606 a_4724_n11415# a_4724_n12503# 0.02fF
C9607 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X a_1722_n11933# 0.00fF
C9608 a_7237_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C9609 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8525_n4317# 0.02fF
C9610 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C9611 a_5653_n1909# a_5752_n2167# 0.49fF
C9612 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.02fF
C9613 a_9876_n5975# sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C9614 a_9450_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C9615 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VDD 0.83fF
C9616 a_5586_n13021# a_4554_n13021# 0.02fF
C9617 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C9618 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.03fF
C9619 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.02fF
C9620 a_3266_n5405# VDD 0.47fF
C9621 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_4724_n3799# 0.03fF
C9622 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C9623 a_3176_n2167# a_3373_n1597# 0.02fF
C9624 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C9625 a_4464_n3255# a_4464_n4887# 0.00fF
C9626 a_10738_n13021# a_11101_n13021# 0.05fF
C9627 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A VDD 1.32fF
C9628 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10805_n11237# 0.01fF
C9629 a_10805_n8437# a_10904_n8695# 0.48fF
C9630 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C9631 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C9632 a_n2436_n7037# a_n1995_n6925# 0.22fF
C9633 a_4724_n13591# a_4554_n13021# 0.04fF
C9634 a_4464_n13591# a_4661_n13021# 0.02fF
C9635 a_1789_n10613# a_1888_n10871# 0.49fF
C9636 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C9637 a_5752_n5975# a_7300_n5975# 0.01fF
C9638 a_6012_n5975# a_7040_n5975# 0.02fF
C9639 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6941_n5797# 0.18fF
C9640 a_10904_n5975# VDD 0.39fF
C9641 a_5752_n13591# VDD 0.43fF
C9642 a_690_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.05fF
C9643 a_3010_n9213# a_4554_n9213# 0.01fF
C9644 a_3266_n9213# a_4298_n9213# 0.02fF
C9645 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.11fF
C9646 a_7040_n1079# a_8588_n1079# 0.01fF
C9647 a_7300_n1079# a_8328_n1079# 0.02fF
C9648 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A a_8229_n821# 0.18fF
C9649 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_3/A 0.32fF
C9650 a_4661_n1597# a_4724_n2167# 0.01fF
C9651 a_6012_n9783# a_5949_n10301# 0.01fF
C9652 a_7237_n1597# a_7300_n2167# 0.01fF
C9653 a_3176_n5975# a_4365_n5797# 0.01fF
C9654 a_3077_n5797# a_4464_n5975# 0.01fF
C9655 a_7040_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C9656 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_8328_n10871# 0.01fF
C9657 a_13765_n13565# p1_b 0.12fF
C9658 p1 a_13765_n13021# 0.12fF
C9659 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C9660 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_2148_n4887# 0.01fF
C9661 a_11101_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.12fF
C9662 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.02fF
C9663 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.04fF
C9664 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.04fF
C9665 a_5842_n2685# VDD 0.44fF
C9666 a_9706_n13021# a_9616_n11415# 0.00fF
C9667 sky130_fd_sc_hd__clkinv_4_10/Y p2_b 0.04fF
C9668 a_2366_n509# VDD 0.81fF
C9669 a_600_n11415# a_797_n13021# 0.00fF
C9670 a_7300_n8695# sky130_fd_sc_hd__clkinv_1_5/A 0.00fF
C9671 a_1888_n2167# a_1722_n2685# 0.04fF
C9672 a_1789_n1909# a_1978_n2685# 0.02fF
C9673 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.08fF
C9674 a_10994_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.04fF
C9675 a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C9676 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_4298_n13021# 0.00fF
C9677 a_6874_n13021# a_7130_n13021# 0.19fF
C9678 a_9517_n10613# a_10904_n10871# 0.01fF
C9679 a_9616_n10871# a_10805_n10613# 0.01fF
C9680 a_690_n5405# VDD 0.48fF
C9681 a_9616_n2167# a_9706_n2685# 0.01fF
C9682 a_6941_n8437# a_6658_n7363# 0.01fF
C9683 a_4464_n11415# VDD 0.44fF
C9684 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.02fF
C9685 a_13765_n11933# a_13765_n13021# 0.07fF
C9686 a_4365_n1909# VDD 0.36fF
C9687 a_5752_n2167# a_7040_n2167# 0.01fF
C9688 a_6012_n2167# a_6941_n1909# 0.02fF
C9689 a_5653_n1909# a_7300_n2167# 0.00fF
C9690 a_3266_n4317# a_3436_n4887# 0.04fF
C9691 a_3176_n11415# a_3266_n10301# 0.01fF
C9692 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_9706_n509# 0.00fF
C9693 a_797_n10301# a_860_n8695# 0.00fF
C9694 a_10805_n12325# a_10738_n13021# 0.01fF
C9695 a_4661_n5405# VDD 0.35fF
C9696 a_6874_n1597# a_6941_n821# 0.01fF
C9697 a_8229_n1909# a_9616_n2167# 0.01fF
C9698 a_8328_n2167# a_9517_n1909# 0.01fF
C9699 a_9616_n13591# a_9706_n11933# 0.00fF
C9700 a_9450_n8125# VDD 0.80fF
C9701 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.02fF
C9702 a_10994_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.04fF
C9703 a_11101_n11933# a_11164_n11415# 0.01fF
C9704 a_860_n10871# a_797_n9213# 0.00fF
C9705 a_9616_n5975# a_9450_n5405# 0.04fF
C9706 a_2148_n10871# a_3077_n10613# 0.02fF
C9707 a_9517_n5797# a_9706_n5405# 0.02fF
C9708 a_1888_n10871# a_3176_n10871# 0.01fF
C9709 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VDD 0.83fF
C9710 a_1789_n10613# a_3436_n10871# 0.00fF
C9711 a_8418_n14109# VDD 0.45fF
C9712 a_600_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C9713 a_9616_n8695# a_9706_n8125# 0.02fF
C9714 a_7040_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.03fF
C9715 a_797_n11933# a_1978_n11933# 0.01fF
C9716 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n11933# 0.35fF
C9717 clk sky130_fd_sc_hd__clkinv_1_3/A 0.00fF
C9718 a_690_n11933# a_2085_n11933# 0.01fF
C9719 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_8328_n5975# 0.01fF
C9720 a_6941_n9525# a_8588_n9783# 0.00fF
C9721 a_7040_n9783# a_8328_n9783# 0.01fF
C9722 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.04fF
C9723 a_4298_n9213# a_4661_n9213# 0.05fF
C9724 a_6941_n11237# a_6941_n10613# 0.05fF
C9725 a_1888_n8695# a_1888_n9783# 0.01fF
C9726 a_10994_n11933# a_10805_n13413# 0.00fF
C9727 a_5586_n4317# a_5586_n2685# 0.01fF
C9728 a_10805_n1909# a_10738_n1597# 0.01fF
C9729 a_4298_n10301# a_5586_n10301# 0.01fF
C9730 a_9616_n3255# a_10805_n2997# 0.01fF
C9731 a_4365_n5797# a_4724_n5975# 0.05fF
C9732 a_5752_n3255# VDD 0.46fF
C9733 a_9616_n2167# sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C9734 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD 0.86fF
C9735 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Ad_b 0.04fF
C9736 a_1888_n5975# sky130_fd_sc_hd__clkinv_4_4/A 0.07fF
C9737 a_2148_n3799# a_1978_n2685# 0.00fF
C9738 a_860_n12503# a_n787_n12325# 0.00fF
C9739 a_600_n12503# a_n688_n12503# 0.01fF
C9740 a_n787_n12325# VDD 0.35fF
C9741 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VDD 0.83fF
C9742 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.09fF
C9743 a_501_n1909# a_434_n1597# 0.01fF
C9744 a_9616_n3255# a_9517_n2997# 0.49fF
C9745 a_7237_n13021# a_8162_n13021# 0.02fF
C9746 a_6874_n13021# a_8525_n13021# 0.00fF
C9747 a_2148_n3255# a_1978_n1597# 0.00fF
C9748 a_7130_n13021# a_8418_n13021# 0.01fF
C9749 a_4724_n11415# a_4661_n13021# 0.00fF
C9750 a_10805_n10613# a_11164_n10871# 0.05fF
C9751 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_8162_n14109# 0.00fF
C9752 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C9753 a_3436_n12503# a_3436_n11415# 0.02fF
C9754 a_6006_n7607# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.19fF
C9755 a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C9756 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.01fF
C9757 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 2.12fF
C9758 a_9813_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.12fF
C9759 a_860_n11415# a_690_n10301# 0.00fF
C9760 a_600_n11415# a_797_n10301# 0.00fF
C9761 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_860_n13591# 0.02fF
C9762 a_8588_n10871# a_8588_n9783# 0.02fF
C9763 a_7040_n2167# a_7300_n2167# 0.28fF
C9764 a_6941_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C9765 a_8525_n509# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C9766 a_3176_n3799# a_3010_n5405# 0.00fF
C9767 a_434_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.03fF
C9768 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9813_n509# 0.02fF
C9769 a_690_n2685# a_797_n2685# 0.55fF
C9770 a_8328_n3255# a_9517_n2997# 0.01fF
C9771 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VDD 0.84fF
C9772 a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.00fF
C9773 a_3077_n3621# a_3266_n5405# 0.00fF
C9774 a_5586_n5405# a_7237_n5405# 0.00fF
C9775 a_5842_n5405# a_7130_n5405# 0.01fF
C9776 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C9777 a_1722_n11933# a_2085_n11933# 0.05fF
C9778 sky130_fd_sc_hd__clkinv_4_3/A p2 0.00fF
C9779 a_9616_n4887# a_9706_n4317# 0.01fF
C9780 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_4365_n10613# 0.01fF
C9781 a_9813_n14109# VDD 0.33fF
C9782 a_3176_n10871# a_3436_n10871# 0.28fF
C9783 a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.02fF
C9784 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_3266_n11933# 0.00fF
C9785 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X a_8588_n5975# 0.03fF
C9786 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_9517_n9525# 0.01fF
C9787 a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.02fF
C9788 a_10904_n4887# a_11101_n5405# 0.02fF
C9789 a_10805_n11237# a_10805_n9525# 0.00fF
C9790 a_7130_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.23fF
C9791 a_4298_n1597# VDD 0.76fF
C9792 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_10904_n8695# 0.01fF
C9793 a_4661_n9213# a_5842_n9213# 0.01fF
C9794 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_5586_n9213# 0.35fF
C9795 a_9450_n1597# VDD 0.75fF
C9796 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.01fF
C9797 a_4298_n4317# VDD 0.76fF
C9798 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.08fF
C9799 a_6874_n9213# a_5586_n9213# 0.01fF
C9800 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.06fF
C9801 a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.02fF
C9802 a_10805_n2997# a_11164_n3255# 0.05fF
C9803 a_5586_n10301# a_5842_n10301# 0.19fF
C9804 a_5842_n11933# a_6874_n11933# 0.02fF
C9805 sky130_fd_sc_hd__dfxbp_1_1/D a_n2248_n7037# 0.25fF
C9806 a_4365_n3621# a_4554_n2685# 0.00fF
C9807 a_7300_n3255# VDD 0.78fF
C9808 a_4464_n3799# a_4298_n2685# 0.00fF
C9809 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.29fF
C9810 a_6874_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.03fF
C9811 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6941_n5797# 0.01fF
C9812 a_8418_n8125# a_9706_n8125# 0.01fF
C9813 a_11164_n2167# sky130_fd_sc_hd__nand2_4_0/Y 0.11fF
C9814 a_3436_n5975# sky130_fd_sc_hd__clkinv_4_4/A 0.11fF
C9815 a_1789_n12325# a_501_n12325# 0.01fF
C9816 a_9517_n10613# a_9450_n9213# 0.00fF
C9817 a_10904_n13591# a_11101_n13021# 0.02fF
C9818 a_11164_n13591# a_10994_n13021# 0.04fF
C9819 a_1789_n10613# a_1789_n9525# 0.02fF
C9820 a_6012_n12503# a_6012_n13591# 0.02fF
C9821 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_860_n11415# 0.01fF
C9822 a_11164_n3255# a_9517_n2997# 0.00fF
C9823 a_8418_n13021# a_8525_n13021# 0.55fF
C9824 a_8162_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.03fF
C9825 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_9450_n13021# 0.00fF
C9826 a_501_n4709# VDD 0.36fF
C9827 sky130_fd_sc_hd__nand2_4_3/Y a_9450_n9213# 0.07fF
C9828 a_5752_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C9829 a_7237_n14109# a_8525_n14109# 0.01fF
C9830 a_7130_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C9831 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C9832 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkinv_4_8/A 0.06fF
C9833 a_434_n4317# a_797_n4317# 0.05fF
C9834 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.02fF
C9835 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C9836 a_4365_n4709# a_4464_n4887# 0.49fF
C9837 a_5842_n5405# a_5842_n4317# 0.01fF
C9838 a_5653_n12325# a_6941_n12325# 0.01fF
C9839 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X a_501_n2997# 0.00fF
C9840 a_4661_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C9841 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_4724_n4887# 0.03fF
C9842 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkinv_4_7/A 0.03fF
C9843 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.03fF
C9844 a_9616_n12503# VDD 0.42fF
C9845 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_n787_n4709# 0.01fF
C9846 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1978_n2685# 0.03fF
C9847 a_690_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.01fF
C9848 a_797_n2685# a_2085_n2685# 0.01fF
C9849 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n509# 0.00fF
C9850 a_5653_n11237# VDD 0.35fF
C9851 a_2085_n11933# a_3266_n11933# 0.01fF
C9852 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3010_n11933# 0.35fF
C9853 a_1978_n11933# a_3373_n11933# 0.01fF
C9854 a_10805_n8437# a_10805_n9525# 0.02fF
C9855 a_6012_n11415# a_6012_n12503# 0.02fF
C9856 a_9517_n4709# sky130_fd_sc_hd__clkinv_4_3/A 0.07fF
C9857 a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C9858 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_10738_n4317# 0.03fF
C9859 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VDD 0.84fF
C9860 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X Ad_b 0.02fF
C9861 a_501_n1909# a_n428_n2167# 0.02fF
C9862 a_860_n2167# a_n787_n1909# 0.00fF
C9863 a_600_n2167# a_n688_n2167# 0.01fF
C9864 a_2085_n5405# a_2148_n4887# 0.01fF
C9865 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.08fF
C9866 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C9867 A_b A 0.47fF
C9868 a_7040_n5975# a_6794_n7203# 0.00fF
C9869 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X a_6665_n7459# 0.00fF
C9870 a_8525_n13021# sky130_fd_sc_hd__clkinv_4_8/A 0.05fF
C9871 a_8229_n8437# a_8328_n9783# 0.00fF
C9872 a_5842_n1597# VDD 0.44fF
C9873 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X a_7300_n1079# 0.00fF
C9874 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_11164_n8695# 0.03fF
C9875 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.00fF
C9876 a_8328_n11415# a_8328_n10871# 0.07fF
C9877 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A VDD 0.73fF
C9878 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_2148_n10871# 0.01fF
C9879 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C9880 a_5842_n4317# a_6012_n5975# 0.00fF
C9881 a_5949_n4317# a_5752_n5975# 0.00fF
C9882 a_4661_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C9883 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_4724_n8695# 0.00fF
C9884 a_5586_n10301# a_7237_n10301# 0.00fF
C9885 a_5842_n10301# a_7130_n10301# 0.01fF
C9886 a_5949_n10301# a_6874_n10301# 0.02fF
C9887 a_7300_n8695# a_7237_n10301# 0.00fF
C9888 a_6874_n11933# a_7237_n11933# 0.05fF
C9889 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VDD 0.82fF
C9890 sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C9891 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.02fF
C9892 clk a_n2602_n7037# 0.39fF
C9893 a_7237_n5405# a_7300_n5975# 0.01fF
C9894 a_9876_n10871# a_9706_n11933# 0.00fF
C9895 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkinv_4_7/A 0.45fF
C9896 a_7130_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C9897 a_690_n9213# a_860_n9783# 0.04fF
C9898 a_10904_n13591# a_10805_n12325# 0.00fF
C9899 a_9876_n2167# a_9876_n3799# 0.01fF
C9900 a_797_n9213# a_600_n9783# 0.02fF
C9901 a_7040_n13591# VDD 0.43fF
C9902 Bd Bd_b 0.47fF
C9903 sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__clkinv_1_3/A 0.18fF
C9904 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Bd_b 0.14fF
C9905 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9706_n13021# 0.03fF
C9906 a_3077_n2997# a_3176_n4887# 0.00fF
C9907 a_3176_n3255# a_3077_n4709# 0.00fF
C9908 a_6941_n9525# a_6941_n10613# 0.02fF
C9909 a_4554_n11933# a_5949_n11933# 0.01fF
C9910 a_4464_n3799# a_4365_n1909# 0.00fF
C9911 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Ad_b 0.02fF
C9912 a_4661_n11933# a_5842_n11933# 0.01fF
C9913 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/X 0.04fF
C9914 a_n688_n4887# a_501_n4709# 0.01fF
C9915 a_5752_n8695# a_5586_n9213# 0.04fF
C9916 a_5653_n8437# a_5842_n9213# 0.02fF
C9917 sky130_fd_sc_hd__dfxbp_1_0/Q a_6006_n7607# 0.37fF
C9918 a_8418_n509# a_9450_n509# 0.02fF
C9919 a_n688_n9783# a_860_n9783# 0.01fF
C9920 a_n428_n9783# a_600_n9783# 0.02fF
C9921 a_4623_n7349# a_6101_n7254# 0.01fF
C9922 a_4464_n4887# a_5752_n4887# 0.01fF
C9923 a_6941_n12325# a_7040_n12503# 0.49fF
C9924 a_4724_n4887# a_5653_n4709# 0.02fF
C9925 a_4365_n4709# a_6012_n4887# 0.00fF
C9926 a_860_n1079# a_2148_n1079# 0.01fF
C9927 a_600_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.00fF
C9928 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X a_1888_n1079# 0.05fF
C9929 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.04fF
C9930 a_11164_n12503# VDD 0.67fF
C9931 a_4464_n3799# a_4661_n5405# 0.00fF
C9932 a_2085_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.12fF
C9933 a_4724_n3799# a_4554_n5405# 0.00fF
C9934 a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C9935 a_9706_n1597# a_9616_n1079# 0.01fF
C9936 a_7040_n11415# VDD 0.44fF
C9937 a_3266_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.05fF
C9938 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_4554_n11933# 0.00fF
C9939 a_600_n3799# VDD 0.44fF
C9940 a_10904_n4887# sky130_fd_sc_hd__clkinv_4_3/A 0.07fF
C9941 a_4365_n5797# a_4554_n5405# 0.02fF
C9942 a_4464_n5975# a_4298_n5405# 0.04fF
C9943 a_6874_n14109# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.03fF
C9944 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6941_n13413# 0.01fF
C9945 a_4464_n10871# a_4554_n9213# 0.00fF
C9946 a_3077_n11237# a_3010_n11933# 0.01fF
C9947 a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C9948 p1d_b p2d_b 0.11fF
C9949 a_7130_n4317# a_7040_n3255# 0.01fF
C9950 a_8229_n4709# a_8229_n5797# 0.02fF
C9951 a_10904_n8695# sky130_fd_sc_hd__clkinv_1_3/A 0.06fF
C9952 a_10805_n1909# a_10805_n2997# 0.02fF
C9953 a_11101_n13021# sky130_fd_sc_hd__clkinv_4_7/Y 0.01fF
C9954 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_3010_n1597# 0.00fF
C9955 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_8162_n10301# 0.00fF
C9956 a_6874_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.03fF
C9957 a_7130_n10301# a_7237_n10301# 0.55fF
C9958 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_n688_n4887# 0.01fF
C9959 a_7237_n11933# a_8418_n11933# 0.01fF
C9960 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8162_n11933# 0.35fF
C9961 a_5752_n3799# a_5949_n2685# 0.00fF
C9962 a_8588_n10871# a_6941_n10613# 0.00fF
C9963 a_7130_n11933# a_8525_n11933# 0.01fF
C9964 a_10738_n6173# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C9965 a_9616_n10871# a_9813_n10301# 0.02fF
C9966 a_9876_n10871# a_9706_n10301# 0.04fF
C9967 sky130_fd_sc_hd__nand2_1_4/Y a_4623_n7349# 0.02fF
C9968 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/X 0.09fF
C9969 sky130_fd_sc_hd__clkinv_4_4/A a_9517_n5797# 0.07fF
C9970 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10805_n5797# 0.01fF
C9971 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/X 0.06fF
C9972 a_10738_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.03fF
C9973 a_5653_n3621# a_5653_n2997# 0.05fF
C9974 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.06fF
C9975 sky130_fd_sc_hd__clkinv_1_4/Y VDD 4.78fF
C9976 a_1888_n4887# a_1978_n4317# 0.01fF
C9977 a_8525_n8125# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C9978 a_8588_n13591# VDD 0.76fF
C9979 a_10904_n8695# a_10738_n9213# 0.04fF
C9980 a_10805_n8437# a_10994_n9213# 0.02fF
C9981 a_3176_n10871# a_3176_n9783# 0.01fF
C9982 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.04fF
C9983 a_4365_n13413# a_4554_n11933# 0.00fF
C9984 a_4464_n13591# a_4298_n11933# 0.00fF
C9985 a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.00fF
C9986 a_2148_n2167# sky130_fd_sc_hd__clkinv_1_0/Y 0.00fF
C9987 a_6874_n10301# a_8418_n10301# 0.01fF
C9988 a_600_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X 0.00fF
C9989 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_7130_n11933# 0.00fF
C9990 a_860_n2167# a_2148_n2167# 0.01fF
C9991 a_8588_n8695# a_8418_n10301# 0.00fF
C9992 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_1888_n2167# 0.05fF
C9993 a_8588_n9783# a_8525_n9213# 0.01fF
C9994 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6874_n5405# 0.35fF
C9995 a_5949_n5405# a_7130_n5405# 0.01fF
C9996 sky130_fd_sc_hd__mux2_1_0/X Ad_b 0.02fF
C9997 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.08fF
C9998 a_4365_n12325# a_5653_n12325# 0.01fF
C9999 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.04fF
C10000 a_6874_n2685# a_5949_n2685# 0.02fF
C10001 a_7237_n2685# a_5586_n2685# 0.00fF
C10002 a_7130_n2685# a_5842_n2685# 0.01fF
C10003 a_7040_n12503# a_8328_n12503# 0.01fF
C10004 a_5653_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.02fF
C10005 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X a_6941_n4709# 0.01fF
C10006 a_7300_n12503# a_8229_n12325# 0.02fF
C10007 a_5752_n4887# a_6012_n4887# 0.28fF
C10008 a_6941_n12325# a_8588_n12503# 0.00fF
C10009 a_6874_n6493# a_6941_n5797# 0.01fF
C10010 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C10011 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.06fF
C10012 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10805_n821# 0.01fF
C10013 a_8588_n11415# VDD 0.77fF
C10014 a_9616_n2167# VDD 0.45fF
C10015 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C10016 a_5949_n2685# a_6012_n3799# 0.00fF
C10017 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Ad_b 0.03fF
C10018 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4661_n11933# 0.02fF
C10019 a_3373_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C10020 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.04fF
C10021 a_9876_n4887# a_9876_n3799# 0.02fF
C10022 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_5586_n9213# 0.00fF
C10023 a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C10024 a_1722_n10301# a_1789_n8437# 0.00fF
C10025 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C10026 a_7237_n14109# a_7300_n13591# 0.01fF
C10027 a_4724_n9783# a_4661_n9213# 0.01fF
C10028 a_860_n11415# a_690_n11933# 0.04fF
C10029 a_5752_n10871# a_5842_n11933# 0.01fF
C10030 a_600_n11415# a_797_n11933# 0.02fF
C10031 a_9813_n1597# a_9706_n509# 0.00fF
C10032 a_9706_n1597# a_9813_n509# 0.00fF
C10033 a_4365_n3621# a_4554_n4317# 0.02fF
C10034 a_10904_n13591# a_9616_n13591# 0.01fF
C10035 a_11164_n13591# a_9517_n13413# 0.00fF
C10036 a_4464_n3799# a_4298_n4317# 0.04fF
C10037 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8229_n2997# 0.00fF
C10038 a_8162_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C10039 a_8229_n3621# a_9517_n3621# 0.01fF
C10040 a_6665_n7459# a_6794_n7203# 0.23fF
C10041 a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.17fF
C10042 a_6658_n7363# p2 0.35fF
C10043 a_7237_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C10044 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7300_n5975# 0.00fF
C10045 a_9616_n5975# a_9813_n4317# 0.00fF
C10046 a_9876_n5975# a_9706_n4317# 0.00fF
C10047 a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C10048 a_10738_n11933# a_10738_n10301# 0.01fF
C10049 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A 0.63fF
C10050 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8229_n10613# 0.02fF
C10051 a_8588_n10871# a_8328_n10871# 0.28fF
C10052 a_5653_n9525# VDD 0.35fF
C10053 a_8418_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.05fF
C10054 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_9706_n11933# 0.00fF
C10055 a_7130_n509# a_6941_n821# 0.02fF
C10056 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C10057 a_6874_n509# a_7040_n1079# 0.04fF
C10058 sky130_fd_sc_hd__clkinv_4_4/A a_10904_n5975# 0.07fF
C10059 a_11101_n5405# a_11164_n5975# 0.01fF
C10060 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkinv_1_3/A 0.84fF
C10061 a_3077_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C10062 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X a_3010_n4317# 0.03fF
C10063 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C10064 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.01fF
C10065 a_5586_n13021# a_5586_n11933# 0.02fF
C10066 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.04fF
C10067 a_434_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C10068 a_8418_n8125# a_8328_n9783# 0.00fF
C10069 a_8229_n4709# VDD 0.35fF
C10070 a_4464_n5975# a_6012_n5975# 0.01fF
C10071 a_4724_n5975# a_5752_n5975# 0.02fF
C10072 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VDD 0.76fF
C10073 a_5842_n4317# a_5949_n5405# 0.00fF
C10074 a_8588_n2167# a_8525_n509# 0.00fF
C10075 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C10076 a_9517_n8437# a_9450_n10301# 0.00fF
C10077 a_4365_n9525# a_4464_n8695# 0.00fF
C10078 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C10079 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A a_3436_n9783# 0.01fF
C10080 a_4464_n9783# a_4365_n8437# 0.00fF
C10081 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_8418_n5405# 0.00fF
C10082 a_2148_n11415# a_2148_n9783# 0.01fF
C10083 a_7130_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.05fF
C10084 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_3077_n821# 0.18fF
C10085 a_2148_n1079# a_3176_n1079# 0.02fF
C10086 a_1888_n1079# a_3436_n1079# 0.01fF
C10087 a_8162_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C10088 a_10805_n4709# a_10805_n2997# 0.00fF
C10089 a_3266_n1597# a_3266_n2685# 0.01fF
C10090 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X Bd_b 0.02fF
C10091 a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.02fF
C10092 a_8328_n12503# a_8588_n12503# 0.28fF
C10093 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X a_7040_n4887# 0.05fF
C10094 a_n2602_n7037# sky130_fd_sc_hd__clkinv_1_5/A 0.11fF
C10095 p1d_b VDD 4.28fF
C10096 sky130_fd_sc_hd__nand2_1_0/A a_600_n4887# 0.01fF
C10097 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.08fF
C10098 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VDD 0.83fF
C10099 a_3176_n3255# a_3436_n3255# 0.28fF
C10100 a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.02fF
C10101 a_6012_n3799# a_6012_n3255# 0.09fF
C10102 a_11164_n2167# VDD 0.67fF
C10103 a_1789_n9525# a_3077_n9525# 0.01fF
C10104 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.03fF
C10105 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_6012_n4887# 0.00fF
C10106 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_6874_n11933# 0.01fF
C10107 a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C10108 a_4464_n11415# a_4554_n11933# 0.02fF
C10109 a_7040_n10871# a_6874_n9213# 0.00fF
C10110 a_6941_n10613# a_7130_n9213# 0.00fF
C10111 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_1722_n2685# 0.00fF
C10112 a_8525_n10301# a_8525_n11933# 0.01fF
C10113 a_8525_n4317# a_8588_n3255# 0.00fF
C10114 sky130_fd_sc_hd__clkinv_1_5/A a_n787_n4709# 0.00fF
C10115 a_9517_n3621# a_9616_n3799# 0.49fF
C10116 a_4464_n1079# a_4298_n2685# 0.00fF
C10117 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.04fF
C10118 a_4365_n821# a_4554_n2685# 0.00fF
C10119 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6665_n7459# 0.02fF
C10120 a_2085_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.01fF
C10121 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_2148_n1079# 0.03fF
C10122 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/Y 0.46fF
C10123 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6012_n13591# 0.03fF
C10124 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_8328_n10871# 0.00fF
C10125 a_7040_n9783# VDD 0.46fF
C10126 a_5949_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C10127 a_10904_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.02fF
C10128 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.02fF
C10129 sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# 0.53fF
C10130 a_1722_n1597# a_1789_n2997# 0.00fF
C10131 a_13765_n2141# B_b 0.15fF
C10132 a_8229_n4709# a_8162_n5405# 0.01fF
C10133 a_4724_n10871# a_4661_n11933# 0.00fF
C10134 a_3176_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C10135 sky130_fd_sc_hd__dfxbp_1_1/D a_n2436_n7037# 0.73fF
C10136 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9517_n9525# 0.00fF
C10137 a_9450_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.00fF
C10138 a_9616_n4887# VDD 0.42fF
C10139 a_n2602_n7037# a_n1995_n6925# 0.30fF
C10140 a_n1570_n6769# a_n2248_n7037# 0.01fF
C10141 a_n2163_n6671# a_n2068_n6671# 0.02fF
C10142 a_3077_n12325# a_4365_n12325# 0.01fF
C10143 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.85fF
C10144 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8525_n5405# 0.02fF
C10145 a_7237_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C10146 a_7237_n2685# a_7040_n3255# 0.02fF
C10147 a_7130_n2685# a_7300_n3255# 0.04fF
C10148 a_1789_n13413# a_1978_n13021# 0.02fF
C10149 a_3176_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.03fF
C10150 a_1888_n13591# a_1722_n13021# 0.04fF
C10151 a_9876_n8695# a_9813_n9213# 0.01fF
C10152 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_4464_n1079# 0.01fF
C10153 a_5949_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.00fF
C10154 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6012_n11415# 0.00fF
C10155 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X a_1888_n4887# 0.05fF
C10156 a_860_n4887# a_2148_n4887# 0.01fF
C10157 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_4_1/A 0.04fF
C10158 a_5586_n2685# a_5653_n821# 0.00fF
C10159 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.89fF
C10160 a_600_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C10161 a_8418_n6493# a_8328_n5975# 0.02fF
C10162 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD 0.85fF
C10163 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7300_n1079# 0.00fF
C10164 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.00fF
C10165 a_600_n2167# VDD 0.47fF
C10166 a_3176_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C10167 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X a_4464_n3255# 0.05fF
C10168 a_3436_n3255# a_4724_n3255# 0.01fF
C10169 a_6874_n6493# a_6658_n7363# 0.00fF
C10170 sky130_fd_sc_hd__nand2_4_1/B Bd_b 0.07fF
C10171 a_3436_n3799# a_1789_n3621# 0.00fF
C10172 a_3176_n3799# a_1888_n3799# 0.01fF
C10173 a_2085_n10301# a_2085_n9213# 0.02fF
C10174 A_b Ad 0.53fF
C10175 a_10994_n1597# sky130_fd_sc_hd__clkinv_4_1/Y 0.01fF
C10176 a_3077_n9525# a_3176_n9783# 0.49fF
C10177 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VDD 0.82fF
C10178 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.29fF
C10179 a_10805_n10613# a_10904_n12503# 0.00fF
C10180 a_10904_n10871# a_10805_n12325# 0.00fF
C10181 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X a_5586_n11933# 0.03fF
C10182 a_6874_n6493# a_6874_n5405# 0.02fF
C10183 a_7300_n10871# a_7237_n11933# 0.00fF
C10184 a_1789_n12325# a_1789_n10613# 0.00fF
C10185 a_9813_n10301# a_9706_n9213# 0.00fF
C10186 a_7130_n6493# VDD 0.46fF
C10187 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Bd_b 0.03fF
C10188 a_2622_n8125# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.04fF
C10189 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.02fF
C10190 a_11164_n5975# sky130_fd_sc_hd__clkinv_4_3/A 0.12fF
C10191 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_5653_n821# 0.01fF
C10192 a_8525_n509# a_8328_n1079# 0.02fF
C10193 a_6941_n1909# a_7040_n3799# 0.00fF
C10194 a_8418_n509# a_8588_n1079# 0.04fF
C10195 a_7040_n2167# a_6941_n3621# 0.00fF
C10196 a_3176_n4887# a_4365_n4709# 0.01fF
C10197 a_3077_n4709# a_4464_n4887# 0.01fF
C10198 a_5842_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.05fF
C10199 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.02fF
C10200 a_10738_n9213# a_10805_n9525# 0.01fF
C10201 a_7130_n13021# a_7040_n12503# 0.02fF
C10202 a_4464_n1079# a_4365_n1909# 0.00fF
C10203 clk a_n2163_n6671# 0.01fF
C10204 a_2729_n509# VDD 0.36fF
C10205 a_6941_n13413# a_6874_n11933# 0.00fF
C10206 a_5949_n9213# a_6101_n7254# 0.00fF
C10207 clk sky130_fd_sc_hd__nand2_1_4/B 0.07fF
C10208 a_4365_n12325# a_4464_n12503# 0.49fF
C10209 a_4464_n9783# a_4464_n11415# 0.00fF
C10210 a_1789_n821# a_1722_n2685# 0.00fF
C10211 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C10212 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A a_4724_n1079# 0.03fF
C10213 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C10214 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.02fF
C10215 a_4298_n5405# a_5842_n5405# 0.01fF
C10216 a_4554_n5405# a_5586_n5405# 0.02fF
C10217 a_1789_n13413# VDD 0.35fF
C10218 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C10219 Bd_b sky130_fd_sc_hd__clkinv_1_3/A 0.22fF
C10220 a_8328_n2167# a_8162_n1597# 0.04fF
C10221 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_3373_n2685# 0.01fF
C10222 a_8229_n1909# a_8418_n1597# 0.02fF
C10223 a_9876_n2167# a_9813_n509# 0.00fF
C10224 a_3176_n2167# a_3176_n3255# 0.01fF
C10225 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.29fF
C10226 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.09fF
C10227 a_5653_n821# a_6012_n1079# 0.05fF
C10228 a_9876_n11415# a_10805_n11237# 0.02fF
C10229 a_9616_n11415# a_10904_n11415# 0.01fF
C10230 a_4464_n10871# a_6012_n10871# 0.01fF
C10231 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_5653_n10613# 0.18fF
C10232 a_4724_n10871# a_5752_n10871# 0.02fF
C10233 a_8525_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C10234 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9813_n10301# 0.02fF
C10235 a_4724_n9783# a_4724_n10871# 0.02fF
C10236 a_10738_n11933# VDD 0.70fF
C10237 a_6941_n11237# a_6874_n11933# 0.01fF
C10238 a_6874_n13021# a_6874_n14109# 0.02fF
C10239 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.04fF
C10240 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.06fF
C10241 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkinv_1_3/A 0.00fF
C10242 a_9450_n1597# a_10738_n1597# 0.01fF
C10243 a_8328_n10871# a_8525_n9213# 0.00fF
C10244 a_690_n9213# VDD 0.46fF
C10245 a_8525_n6493# VDD 0.35fF
C10246 a_2366_n6493# a_2148_n5975# 0.03fF
C10247 a_9517_n11237# a_9616_n10871# 0.01fF
C10248 a_600_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.03fF
C10249 a_1888_n11415# a_1978_n13021# 0.00fF
C10250 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X a_5752_n1079# 0.05fF
C10251 a_10738_n6173# a_10738_n5405# 0.01fF
C10252 a_4724_n1079# a_6012_n1079# 0.01fF
C10253 a_4464_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.00fF
C10254 a_3176_n8695# VDD 0.49fF
C10255 a_10805_n3621# a_10738_n2685# 0.00fF
C10256 a_8328_n4887# a_8162_n4317# 0.04fF
C10257 a_8418_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.08fF
C10258 a_8229_n8437# VDD 0.36fF
C10259 a_8229_n4709# a_8418_n4317# 0.02fF
C10260 a_3077_n10613# a_3010_n10301# 0.01fF
C10261 a_2366_n14109# a_2148_n13591# 0.03fF
C10262 a_9517_n5797# a_8588_n5975# 0.02fF
C10263 a_9876_n5975# a_8229_n5797# 0.00fF
C10264 a_9616_n5975# a_8328_n5975# 0.01fF
C10265 a_n688_n9783# VDD 0.51fF
C10266 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C10267 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_7237_n4317# 0.02fF
C10268 a_9616_n4887# a_9706_n5405# 0.02fF
C10269 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.00fF
C10270 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_10805_n9525# 0.01fF
C10271 a_3373_n1597# a_3010_n1597# 0.05fF
C10272 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_3010_n9213# 0.00fF
C10273 a_8162_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.03fF
C10274 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8229_n12325# 0.01fF
C10275 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.03fF
C10276 a_9706_n2685# a_9813_n1597# 0.00fF
C10277 a_9813_n2685# a_9706_n1597# 0.00fF
C10278 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.02fF
C10279 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VDD 0.92fF
C10280 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.02fF
C10281 a_501_n10613# a_434_n10301# 0.01fF
C10282 a_7130_n9213# a_6658_n7363# 0.00fF
C10283 a_6874_n9213# a_6665_n7459# 0.00fF
C10284 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.02fF
C10285 a_8525_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C10286 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.03fF
C10287 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A 0.01fF
C10288 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8588_n3255# 0.03fF
C10289 a_3436_n13591# a_3266_n13021# 0.04fF
C10290 a_3176_n13591# a_3373_n13021# 0.02fF
C10291 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X a_5653_n5797# 0.18fF
C10292 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.03fF
C10293 a_10994_n9213# sky130_fd_sc_hd__clkinv_1_3/A 0.01fF
C10294 a_3176_n13591# VDD 0.45fF
C10295 a_10904_n3799# a_9517_n3621# 0.01fF
C10296 a_10805_n3621# a_9616_n3799# 0.01fF
C10297 a_1789_n1909# a_3077_n1909# 0.01fF
C10298 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C10299 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_4724_n13591# 0.01fF
C10300 a_7237_n9213# VDD 0.35fF
C10301 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X a_6941_n821# 0.18fF
C10302 a_6012_n1079# a_7040_n1079# 0.02fF
C10303 a_1888_n5975# a_3077_n5797# 0.01fF
C10304 sky130_fd_sc_hd__nand2_4_2/A a_10994_n13021# 0.00fF
C10305 a_5752_n1079# a_7300_n1079# 0.01fF
C10306 a_1789_n5797# a_3176_n5975# 0.01fF
C10307 a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C10308 a_10904_n11415# a_11164_n11415# 0.23fF
C10309 a_9616_n12503# a_9706_n11933# 0.01fF
C10310 a_10738_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C10311 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.04fF
C10312 a_5752_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.03fF
C10313 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_7040_n10871# 0.01fF
C10314 a_4554_n1597# a_4365_n821# 0.02fF
C10315 a_4298_n1597# a_4464_n1079# 0.04fF
C10316 a_9813_n8125# a_9706_n9213# 0.00fF
C10317 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A 0.02fF
C10318 a_3266_n2685# VDD 0.44fF
C10319 a_10738_n9213# a_10994_n9213# 0.19fF
C10320 a_1789_n13413# a_501_n13413# 0.01fF
C10321 sky130_fd_sc_hd__clkinv_4_8/A a_7300_n12503# 0.10fF
C10322 a_8418_n6493# a_8418_n5405# 0.01fF
C10323 a_1722_n1597# a_1722_n2685# 0.02fF
C10324 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C10325 a_3176_n12503# a_3176_n10871# 0.00fF
C10326 a_3077_n1909# a_4464_n2167# 0.01fF
C10327 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_3010_n13021# 0.00fF
C10328 a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C10329 a_5842_n5405# a_6012_n5975# 0.04fF
C10330 a_4724_n8695# VDD 0.84fF
C10331 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.02fF
C10332 a_9813_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C10333 a_1888_n11415# VDD 0.44fF
C10334 a_9616_n8695# VDD 0.45fF
C10335 a_5653_n9525# a_5586_n9213# 0.01fF
C10336 a_2085_n10301# a_1978_n9213# 0.00fF
C10337 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.08fF
C10338 a_501_n10613# VDD 0.36fF
C10339 a_4464_n2167# a_5752_n2167# 0.01fF
C10340 a_4724_n2167# a_5653_n1909# 0.02fF
C10341 a_3266_n10301# a_3436_n8695# 0.00fF
C10342 a_3373_n10301# a_3176_n8695# 0.00fF
C10343 a_4661_n1597# a_3266_n1597# 0.01fF
C10344 a_1888_n11415# a_1978_n10301# 0.01fF
C10345 a_8525_n13021# a_8588_n12503# 0.01fF
C10346 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.00fF
C10347 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C10348 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_2085_n4317# 0.01fF
C10349 a_5586_n1597# a_5653_n821# 0.01fF
C10350 a_8162_n1597# a_8229_n821# 0.01fF
C10351 a_2085_n5405# VDD 0.35fF
C10352 a_8328_n13591# a_8418_n11933# 0.00fF
C10353 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_10738_n13021# 0.35fF
C10354 a_9813_n11933# a_9876_n11415# 0.01fF
C10355 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C10356 a_9813_n13021# a_10994_n13021# 0.01fF
C10357 a_8229_n9525# sky130_fd_sc_hd__nand2_4_3/Y 0.08fF
C10358 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.02fF
C10359 a_13765_n5405# a_13765_n4317# 0.07fF
C10360 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_1_4/Y 0.07fF
C10361 a_6874_n8125# VDD 0.76fF
C10362 a_5586_n13021# VDD 0.74fF
C10363 a_860_n10871# a_1789_n10613# 0.02fF
C10364 a_600_n10871# a_1888_n10871# 0.01fF
C10365 a_5752_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.03fF
C10366 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X a_7040_n5975# 0.01fF
C10367 a_9876_n5975# VDD 0.73fF
C10368 a_9517_n1909# a_9450_n509# 0.00fF
C10369 a_4724_n13591# VDD 0.81fF
C10370 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_860_n3255# 0.03fF
C10371 a_797_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C10372 a_7040_n3799# a_7040_n4887# 0.01fF
C10373 a_3077_n1909# a_3176_n2167# 0.49fF
C10374 a_3010_n9213# a_3373_n9213# 0.05fF
C10375 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A VDD 0.88fF
C10376 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_797_n11933# 0.01fF
C10377 a_7040_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.03fF
C10378 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X a_8328_n1079# 0.01fF
C10379 a_5653_n11237# a_5653_n10613# 0.05fF
C10380 a_3077_n5797# a_3436_n5975# 0.05fF
C10381 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C10382 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_8588_n3255# 0.01fF
C10383 a_11101_n1597# a_11164_n3255# 0.00fF
C10384 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C10385 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X a_7300_n10871# 0.03fF
C10386 a_n2163_n6671# sky130_fd_sc_hd__clkinv_1_5/A 0.08fF
C10387 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.01fF
C10388 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A 2.37fF
C10389 a_8328_n11415# a_8418_n11933# 0.02fF
C10390 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_5/A 0.92fF
C10391 a_4661_n2685# VDD 0.35fF
C10392 a_10994_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.04fF
C10393 a_501_n11237# a_860_n11415# 0.05fF
C10394 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.01fF
C10395 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.70fF
C10396 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n5405# 0.01fF
C10397 a_9450_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C10398 sky130_fd_sc_hd__mux2_1_0/X a_6006_n7607# 0.01fF
C10399 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C10400 a_5949_n13021# a_6874_n13021# 0.02fF
C10401 a_1888_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X 0.03fF
C10402 a_3436_n11415# a_3373_n13021# 0.00fF
C10403 a_5842_n13021# a_7130_n13021# 0.01fF
C10404 a_8525_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.01fF
C10405 a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C10406 a_9517_n10613# a_9876_n10871# 0.05fF
C10407 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VDD 0.83fF
C10408 a_2148_n12503# a_2148_n11415# 0.02fF
C10409 a_3436_n11415# VDD 0.77fF
C10410 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_8588_n9783# 0.00fF
C10411 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.04fF
C10412 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.00fF
C10413 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_6941_n1909# 0.01fF
C10414 a_5752_n2167# a_6012_n2167# 0.28fF
C10415 a_5653_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C10416 sky130_fd_sc_hd__clkinv_1_5/A Ad_b 0.55fF
C10417 a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C10418 a_7040_n3255# a_8229_n2997# 0.01fF
C10419 a_6941_n2997# a_8328_n3255# 0.01fF
C10420 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_3010_n10301# 0.01fF
C10421 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.35fF
C10422 a_4298_n5405# a_5949_n5405# 0.00fF
C10423 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.03fF
C10424 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_3373_n1597# 0.01fF
C10425 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X a_9450_n11933# 0.00fF
C10426 a_9517_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C10427 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A VDD 0.88fF
C10428 a_9813_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C10429 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C10430 a_10994_n13021# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C10431 a_4724_n3255# a_4724_n4887# 0.01fF
C10432 a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.01fF
C10433 a_10904_n8695# a_11164_n8695# 0.23fF
C10434 a_8418_n8125# VDD 0.45fF
C10435 a_n2436_n7037# a_n1570_n6769# 0.13fF
C10436 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_3077_n10613# 0.01fF
C10437 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C10438 a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.02fF
C10439 a_1888_n10871# a_2148_n10871# 0.28fF
C10440 a_n1995_n6925# a_n2163_n6671# 0.38fF
C10441 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_4661_n13021# 0.01fF
C10442 a_1789_n2997# VDD 0.35fF
C10443 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_7300_n5975# 0.03fF
C10444 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_3436_n13591# 0.01fF
C10445 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X 0.01fF
C10446 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_1978_n11933# 0.00fF
C10447 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C10448 a_13765_n5949# VDD 2.07fF
C10449 a_9616_n4887# a_9813_n5405# 0.02fF
C10450 a_600_n2167# a_600_n1079# 0.01fF
C10451 a_3266_n9213# a_4661_n9213# 0.01fF
C10452 a_3373_n9213# a_4554_n9213# 0.01fF
C10453 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4298_n9213# 0.35fF
C10454 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A a_8588_n1079# 0.03fF
C10455 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_4365_n5797# 0.18fF
C10456 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.08fF
C10457 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C10458 a_3176_n5975# a_4724_n5975# 0.01fF
C10459 a_3436_n5975# a_4464_n5975# 0.02fF
C10460 a_1722_n4317# VDD 0.76fF
C10461 a_4298_n10301# a_4554_n10301# 0.19fF
C10462 a_3077_n3621# a_3266_n2685# 0.00fF
C10463 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.08fF
C10464 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.06fF
C10465 a_3176_n3799# a_3010_n2685# 0.00fF
C10466 a_1789_n4709# a_3077_n4709# 0.01fF
C10467 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_9450_n11933# 0.03fF
C10468 a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C10469 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A VDD 0.89fF
C10470 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.00fF
C10471 a_5653_n2997# VDD 0.35fF
C10472 a_2148_n2167# a_1978_n2685# 0.04fF
C10473 a_1888_n2167# a_2085_n2685# 0.02fF
C10474 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.02fF
C10475 a_9876_n3255# a_8229_n2997# 0.00fF
C10476 a_9616_n3255# a_8328_n3255# 0.01fF
C10477 a_1722_n9213# a_3010_n9213# 0.01fF
C10478 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_8162_n13021# 0.00fF
C10479 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.03fF
C10480 a_7130_n13021# a_7237_n13021# 0.55fF
C10481 a_9876_n10871# a_10904_n10871# 0.02fF
C10482 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_10805_n10613# 0.17fF
C10483 a_9616_n10871# a_11164_n10871# 0.01fF
C10484 a_9876_n2167# a_9813_n2685# 0.01fF
C10485 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A VDD 0.88fF
C10486 a_6941_n8437# a_6865_n7304# 0.02fF
C10487 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VDD 0.84fF
C10488 p1d_b p1_b 0.20fF
C10489 a_6874_n1597# a_6941_n2997# 0.00fF
C10490 a_9450_n1597# a_9517_n2997# 0.00fF
C10491 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkinv_4_7/A 0.05fF
C10492 a_11164_n13591# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C10493 a_10805_n3621# a_10904_n3799# 0.48fF
C10494 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X a_7040_n2167# 0.05fF
C10495 a_5752_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C10496 a_6012_n2167# a_7300_n2167# 0.01fF
C10497 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_3436_n4887# 0.03fF
C10498 a_3373_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C10499 a_8229_n2997# a_8588_n3255# 0.05fF
C10500 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.00fF
C10501 a_3436_n11415# a_3373_n10301# 0.00fF
C10502 a_8328_n2167# a_9876_n2167# 0.01fF
C10503 a_1789_n3621# a_1722_n5405# 0.00fF
C10504 a_13765_n4317# Ad_b 2.86fF
C10505 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_6874_n5405# 0.00fF
C10506 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_9517_n1909# 0.18fF
C10507 a_8588_n2167# a_9616_n2167# 0.02fF
C10508 a_5842_n5405# a_5949_n5405# 0.55fF
C10509 a_5586_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.03fF
C10510 a_10904_n12503# a_10994_n13021# 0.02fF
C10511 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C10512 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C10513 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_9450_n4317# 0.03fF
C10514 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C10515 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.02fF
C10516 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X a_3176_n10871# 0.05fF
C10517 a_2148_n10871# a_3436_n10871# 0.01fF
C10518 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VDD 0.87fF
C10519 a_11101_n5405# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C10520 a_1888_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.00fF
C10521 a_9876_n5975# a_9706_n5405# 0.04fF
C10522 a_434_n4317# a_501_n4709# 0.01fF
C10523 a_7300_n9783# a_8588_n9783# 0.01fF
C10524 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A a_8328_n9783# 0.05fF
C10525 a_797_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C10526 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_2085_n11933# 0.02fF
C10527 a_7040_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.00fF
C10528 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X a_4298_n10301# 0.03fF
C10529 a_9813_n6493# a_9706_n8125# 0.00fF
C10530 a_8418_n1597# VDD 0.44fF
C10531 a_4554_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.05fF
C10532 a_9706_n6493# a_9813_n8125# 0.00fF
C10533 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_5842_n9213# 0.00fF
C10534 a_2148_n8695# a_2148_n9783# 0.02fF
C10535 a_7040_n11415# a_7040_n10871# 0.07fF
C10536 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_860_n10871# 0.01fF
C10537 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X a_9450_n10301# 0.01fF
C10538 sky130_fd_sc_hd__clkinv_4_8/A a_10805_n13413# 0.02fF
C10539 a_5842_n4317# a_5842_n2685# 0.01fF
C10540 a_10904_n2167# a_10994_n1597# 0.02fF
C10541 a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C10542 a_3266_n4317# VDD 0.47fF
C10543 a_9616_n3255# a_11164_n3255# 0.01fF
C10544 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X a_10805_n2997# 0.17fF
C10545 a_9876_n3255# a_10904_n3255# 0.02fF
C10546 a_4298_n10301# a_5949_n10301# 0.00fF
C10547 a_4554_n10301# a_5842_n10301# 0.01fF
C10548 a_4661_n10301# a_5586_n10301# 0.02fF
C10549 a_434_n11933# a_501_n10613# 0.00fF
C10550 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VDD 0.83fF
C10551 a_3077_n4709# a_3176_n4887# 0.49fF
C10552 a_5949_n5405# a_6012_n5975# 0.01fF
C10553 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C10554 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C10555 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_4_4/A 0.85fF
C10556 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_8588_n3799# 0.01fF
C10557 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__nand2_4_0/Y 0.69fF
C10558 a_8588_n10871# a_8418_n11933# 0.00fF
C10559 a_600_n12503# a_501_n12325# 0.49fF
C10560 a_860_n12503# a_n428_n12503# 0.01fF
C10561 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_n688_n12503# 0.00fF
C10562 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.01fF
C10563 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X a_2085_n2685# 0.00fF
C10564 a_n428_n12503# VDD 0.83fF
C10565 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X a_9517_n2997# 0.02fF
C10566 a_10805_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C10567 sky130_fd_sc_hd__nand2_4_3/Y a_8418_n9213# 0.08fF
C10568 a_600_n2167# a_690_n1597# 0.02fF
C10569 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.02fF
C10570 sky130_fd_sc_hd__clkinv_4_8/Y VDD 3.54fF
C10571 a_5653_n9525# a_5653_n10613# 0.02fF
C10572 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.00fF
C10573 a_7237_n13021# a_8525_n13021# 0.01fF
C10574 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8418_n13021# 0.03fF
C10575 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X a_2085_n1597# 0.00fF
C10576 a_7130_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C10577 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.04fF
C10578 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Ad_b 0.02fF
C10579 a_4365_n9525# a_5752_n9783# 0.01fF
C10580 a_4464_n9783# a_5653_n9525# 0.01fF
C10581 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C10582 a_6373_n7349# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.02fF
C10583 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_434_n4317# 0.44fF
C10584 a_4464_n8695# a_4298_n9213# 0.04fF
C10585 a_4365_n8437# a_4554_n9213# 0.02fF
C10586 a_7130_n509# a_8162_n509# 0.02fF
C10587 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C10588 a_6874_n509# a_8418_n509# 0.01fF
C10589 a_5653_n12325# a_5752_n12503# 0.49fF
C10590 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.29fF
C10591 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5586_n4317# 0.01fF
C10592 a_3436_n4887# a_4365_n4709# 0.02fF
C10593 a_9706_n14109# a_9517_n13413# 0.02fF
C10594 a_9450_n14109# a_9616_n13591# 0.04fF
C10595 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.04fF
C10596 a_3436_n3799# a_3266_n5405# 0.00fF
C10597 a_797_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_45/A 0.12fF
C10598 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X a_9517_n2997# 0.18fF
C10599 a_3176_n3799# a_3373_n5405# 0.00fF
C10600 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.02fF
C10601 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_10904_n2167# 0.01fF
C10602 a_5842_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C10603 sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD 0.50fF
C10604 a_1978_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.05fF
C10605 a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C10606 a_n1139_n6715# VDD 0.47fF
C10607 a_3176_n5975# a_3010_n5405# 0.04fF
C10608 a_3077_n5797# a_3266_n5405# 0.02fF
C10609 a_9876_n4887# a_9813_n4317# 0.01fF
C10610 a_8328_n4887# sky130_fd_sc_hd__clkinv_4_3/A 0.07fF
C10611 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.29fF
C10612 a_434_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.00fF
C10613 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.04fF
C10614 a_10904_n11415# a_10904_n9783# 0.00fF
C10615 a_1789_n11237# a_1722_n11933# 0.01fF
C10616 a_5842_n4317# a_5752_n3255# 0.01fF
C10617 a_13765_n5405# Bd_b 0.10fF
C10618 a_4661_n1597# VDD 0.35fF
C10619 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkinv_4_8/A 0.44fF
C10620 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X a_6865_n7304# 0.00fF
C10621 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C10622 a_9813_n1597# VDD 0.33fF
C10623 a_7130_n9213# a_5842_n9213# 0.01fF
C10624 a_7237_n9213# a_5586_n9213# 0.00fF
C10625 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C10626 a_4661_n4317# VDD 0.35fF
C10627 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_6874_n10301# 0.00fF
C10628 a_4724_n3799# a_4554_n2685# 0.00fF
C10629 a_4464_n3799# a_4661_n2685# 0.00fF
C10630 a_n2602_n7037# sky130_fd_sc_hd__dfxbp_1_1/D 0.41fF
C10631 a_5586_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.03fF
C10632 a_5842_n10301# a_5949_n10301# 0.55fF
C10633 a_5949_n11933# a_7130_n11933# 0.01fF
C10634 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_6874_n11933# 0.35fF
C10635 a_5842_n11933# a_7237_n11933# 0.01fF
C10636 a_4365_n3621# a_4365_n2997# 0.05fF
C10637 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.05fF
C10638 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9706_n8125# 0.03fF
C10639 a_690_n4317# a_501_n3621# 0.02fF
C10640 a_434_n4317# a_600_n3799# 0.04fF
C10641 a_501_n821# a_690_n2685# 0.00fF
C10642 a_2148_n12503# a_501_n12325# 0.00fF
C10643 a_9616_n10871# a_9706_n9213# 0.00fF
C10644 a_6012_n13591# VDD 0.76fF
C10645 a_11164_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C10646 a_1888_n10871# a_1888_n9783# 0.01fF
C10647 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.04fF
C10648 a_9517_n12325# a_9517_n13413# 0.02fF
C10649 a_3176_n13591# a_3010_n11933# 0.00fF
C10650 a_3077_n13413# a_3266_n11933# 0.00fF
C10651 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_1722_n1597# 0.03fF
C10652 a_8525_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.12fF
C10653 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_5842_n11933# 0.00fF
C10654 a_860_n4887# VDD 0.78fF
C10655 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X a_10738_n13021# 0.03fF
C10656 a_9517_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C10657 a_690_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.05fF
C10658 a_1888_n5975# a_1722_n5405# 0.04fF
C10659 a_n688_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.02fF
C10660 a_1789_n5797# a_1978_n5405# 0.02fF
C10661 a_8162_n509# a_8525_n509# 0.05fF
C10662 a_1722_n2685# VDD 0.76fF
C10663 a_5653_n12325# a_7300_n12503# 0.00fF
C10664 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C10665 a_4365_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.02fF
C10666 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X a_5653_n4709# 0.01fF
C10667 a_6012_n12503# a_6941_n12325# 0.02fF
C10668 a_4464_n4887# a_4724_n4887# 0.28fF
C10669 a_5752_n12503# a_7040_n12503# 0.01fF
C10670 a_13765_n10301# p2 0.02fF
C10671 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VDD 0.79fF
C10672 a_13765_n1053# Bd_b 0.02fF
C10673 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.02fF
C10674 a_9450_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X 0.03fF
C10675 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9517_n821# 0.01fF
C10676 a_2085_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C10677 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3373_n11933# 0.02fF
C10678 a_6012_n11415# VDD 0.77fF
C10679 a_4365_n10613# a_4298_n11933# 0.00fF
C10680 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A 0.97fF
C10681 a_10904_n8695# a_10904_n9783# 0.01fF
C10682 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.04fF
C10683 a_9517_n11237# a_9517_n12325# 0.02fF
C10684 a_9876_n4887# sky130_fd_sc_hd__clkinv_4_3/A 0.10fF
C10685 a_5842_n4317# a_4298_n4317# 0.01fF
C10686 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X a_n688_n2167# 0.00fF
C10687 a_5586_n4317# a_4554_n4317# 0.02fF
C10688 a_860_n2167# a_n428_n2167# 0.01fF
C10689 a_600_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C10690 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.08fF
C10691 a_13765_n11933# a_13765_n10301# 0.04fF
C10692 a_3176_n3799# a_3010_n4317# 0.04fF
C10693 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6941_n2997# 0.00fF
C10694 a_3077_n3621# a_3266_n4317# 0.02fF
C10695 a_6874_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C10696 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A VDD 0.89fF
C10697 a_6941_n3621# a_8229_n3621# 0.01fF
C10698 a_5653_n13413# a_5842_n11933# 0.00fF
C10699 a_5842_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C10700 a_5949_n10301# a_7237_n10301# 0.01fF
C10701 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_7130_n10301# 0.03fF
C10702 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6012_n5975# 0.00fF
C10703 a_7130_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.05fF
C10704 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_8418_n11933# 0.00fF
C10705 a_5949_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C10706 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C10707 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C10708 a_9813_n5405# a_9876_n5975# 0.01fF
C10709 a_9450_n8125# sky130_fd_sc_hd__nand2_4_3/Y 0.01fF
C10710 a_10738_n13789# a_10994_n13021# 0.01fF
C10711 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.06fF
C10712 a_10738_n11933# a_9706_n11933# 0.02fF
C10713 a_10994_n11933# a_9450_n11933# 0.01fF
C10714 a_797_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C10715 a_9616_n2167# a_9517_n2997# 0.00fF
C10716 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C10717 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_3/A 0.47fF
C10718 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_860_n9783# 0.03fF
C10719 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VDD 0.82fF
C10720 a_7040_n9783# a_7040_n10871# 0.01fF
C10721 a_4661_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C10722 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5949_n11933# 0.02fF
C10723 a_6012_n8695# a_5842_n9213# 0.04fF
C10724 sky130_fd_sc_hd__nand2_1_4/B Bd_b 0.02fF
C10725 a_n688_n4887# a_860_n4887# 0.01fF
C10726 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C10727 a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.17fF
C10728 a_6874_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C10729 sky130_fd_sc_hd__dfxbp_1_0/Q a_6373_n7349# 0.04fF
C10730 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9450_n509# 0.35fF
C10731 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_8229_n12325# 0.01fF
C10732 a_4464_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C10733 a_6941_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C10734 a_7040_n12503# a_7300_n12503# 0.28fF
C10735 a_4724_n4887# a_6012_n4887# 0.01fF
C10736 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X a_5752_n4887# 0.05fF
C10737 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.02fF
C10738 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.00fF
C10739 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_4661_n5405# 0.00fF
C10740 a_9450_n13021# a_9450_n11933# 0.02fF
C10741 a_9813_n1597# a_9876_n1079# 0.01fF
C10742 sky130_fd_sc_hd__clkinv_1_3/Y VDD 1.20fF
C10743 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD 0.84fF
C10744 a_13765_n4861# VDD 1.90fF
C10745 a_13765_n8669# a_13765_n9757# 0.07fF
C10746 sky130_fd_sc_hd__dfxbp_1_0/Q VDD 2.09fF
C10747 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VDD 0.84fF
C10748 a_501_n9525# a_1789_n9525# 0.01fF
C10749 a_4464_n5975# a_4661_n5405# 0.02fF
C10750 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C10751 a_4724_n5975# a_4554_n5405# 0.04fF
C10752 sky130_fd_sc_hd__nand2_4_1/B a_10738_n5405# 0.01fF
C10753 a_4724_n10871# a_4661_n9213# 0.00fF
C10754 Bd_b Ad_b 5.22fF
C10755 a_501_n8437# a_690_n9213# 0.02fF
C10756 a_600_n8695# a_434_n9213# 0.04fF
C10757 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.87fF
C10758 a_3176_n11415# a_3266_n11933# 0.02fF
C10759 a_7237_n4317# a_7300_n3255# 0.00fF
C10760 a_8328_n4887# a_8328_n5975# 0.01fF
C10761 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A 2.37fF
C10762 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__clkinv_1_3/A 0.68fF
C10763 a_3176_n1079# a_3010_n2685# 0.00fF
C10764 a_10904_n2167# a_10904_n3255# 0.01fF
C10765 a_11164_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.33fF
C10766 a_3077_n821# a_3266_n2685# 0.00fF
C10767 a_8229_n3621# a_8328_n3799# 0.49fF
C10768 a_6941_n4709# VDD 0.35fF
C10769 a_7237_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.12fF
C10770 a_8229_n13413# a_9616_n13591# 0.01fF
C10771 a_8328_n13591# a_9517_n13413# 0.01fF
C10772 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8525_n11933# 0.02fF
C10773 a_7237_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C10774 a_6874_n14109# a_7040_n12503# 0.00fF
C10775 a_8588_n10871# a_7300_n10871# 0.01fF
C10776 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C10777 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_9813_n10301# 0.01fF
C10778 a_7130_n14109# a_6941_n12325# 0.00fF
C10779 a_8418_n9213# a_9450_n9213# 0.02fF
C10780 a_8162_n9213# a_9706_n9213# 0.01fF
C10781 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_7040_n10871# 0.00fF
C10782 sky130_fd_sc_hd__clkinv_4_4/A a_9876_n5975# 0.11fF
C10783 sky130_fd_sc_hd__clkinv_1_0/A a_9517_n821# 0.06fF
C10784 a_1888_n3255# a_1789_n2997# 0.49fF
C10785 a_434_n1597# a_501_n2997# 0.00fF
C10786 a_2148_n4887# a_2085_n4317# 0.01fF
C10787 a_4464_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.03fF
C10788 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_5752_n5975# 0.01fF
C10789 p1 a_13765_n12477# 0.06fF
C10790 a_13765_n13565# p1d 0.06fF
C10791 a_10904_n8695# a_11101_n9213# 0.02fF
C10792 a_3436_n10871# a_3436_n9783# 0.02fF
C10793 a_4365_n9525# a_4365_n10613# 0.02fF
C10794 a_11164_n8695# a_10994_n9213# 0.04fF
C10795 a_4464_n13591# a_4661_n11933# 0.00fF
C10796 a_4724_n13591# a_4554_n11933# 0.00fF
C10797 a_1888_n3255# a_1722_n4317# 0.00fF
C10798 a_7237_n10301# a_8418_n10301# 0.01fF
C10799 a_1789_n12325# a_3077_n12325# 0.01fF
C10800 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkinv_4_3/A 0.05fF
C10801 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/X 0.02fF
C10802 a_5653_n3621# a_5653_n1909# 0.00fF
C10803 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C10804 a_4365_n12325# a_6012_n12503# 0.00fF
C10805 a_4464_n12503# a_5752_n12503# 0.01fF
C10806 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.08fF
C10807 a_5949_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C10808 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_7237_n5405# 0.02fF
C10809 a_1888_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X 0.03fF
C10810 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3010_n2685# 0.01fF
C10811 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_5842_n2685# 0.01fF
C10812 a_9450_n4317# a_9517_n3621# 0.01fF
C10813 a_7130_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.03fF
C10814 a_7237_n2685# a_5949_n2685# 0.01fF
C10815 a_7300_n12503# a_8588_n12503# 0.01fF
C10816 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X a_8328_n12503# 0.05fF
C10817 a_7040_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C10818 a_6012_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.29fF
C10819 a_7130_n6493# a_7040_n5975# 0.02fF
C10820 a_13765_n11933# a_13765_n12477# 0.31fF
C10821 a_1888_n8695# VDD 0.49fF
C10822 a_13765_n2141# B 0.06fF
C10823 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VDD 0.83fF
C10824 a_9517_n9525# a_10805_n9525# 0.01fF
C10825 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.03fF
C10826 a_1789_n9525# a_1888_n9783# 0.49fF
C10827 a_9450_n2685# a_9517_n3621# 0.00fF
C10828 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.04fF
C10829 a_9616_n4887# a_9517_n2997# 0.00fF
C10830 a_1978_n10301# a_1888_n8695# 0.00fF
C10831 a_9517_n10613# a_9616_n12503# 0.00fF
C10832 a_9616_n10871# a_9517_n12325# 0.00fF
C10833 a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C10834 a_10738_n11933# a_10738_n13021# 0.02fF
C10835 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.03fF
C10836 a_6012_n10871# a_5949_n11933# 0.00fF
C10837 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.08fF
C10838 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X a_4298_n11933# 0.03fF
C10839 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_9876_n9783# 0.01fF
C10840 a_8328_n11415# a_9517_n11237# 0.01fF
C10841 a_4724_n3799# a_4554_n4317# 0.04fF
C10842 a_4464_n3799# a_4661_n4317# 0.02fF
C10843 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C10844 a_11164_n13591# a_9876_n13591# 0.01fF
C10845 a_10904_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.05fF
C10846 a_8525_n10301# a_8418_n9213# 0.00fF
C10847 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_690_n2685# 0.02fF
C10848 a_8588_n3799# a_9517_n3621# 0.02fF
C10849 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkinv_4_4/A 0.04fF
C10850 a_8328_n3799# a_9616_n3799# 0.01fF
C10851 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X 0.02fF
C10852 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_9813_n4317# 0.00fF
C10853 a_9876_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C10854 a_10738_n2685# a_10994_n2685# 0.19fF
C10855 a_6865_n7304# p2 0.01fF
C10856 sky130_fd_sc_hd__clkinv_1_5/A a_6006_n7607# 0.01fF
C10857 a_10738_n2685# a_10738_n4317# 0.01fF
C10858 a_9517_n13413# a_9876_n13591# 0.05fF
C10859 a_6012_n9783# VDD 0.78fF
C10860 a_7237_n509# a_7040_n1079# 0.02fF
C10861 a_10994_n11933# a_10994_n10301# 0.01fF
C10862 a_4365_n5797# a_4554_n4317# 0.00fF
C10863 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C10864 a_4464_n5975# a_4298_n4317# 0.00fF
C10865 a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C10866 a_7130_n509# a_7300_n1079# 0.04fF
C10867 sky130_fd_sc_hd__clkinv_1_0/A a_10904_n1079# 0.06fF
C10868 sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# 0.52fF
C10869 a_13765_n8669# p2d_b 0.02fF
C10870 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_501_n9525# 0.18fF
C10871 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X a_434_n10301# 0.01fF
C10872 a_6941_n8437# a_5653_n8437# 0.01fF
C10873 a_10904_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.02fF
C10874 a_8525_n8125# a_8588_n9783# 0.00fF
C10875 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C10876 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C10877 a_8588_n4887# VDD 0.77fF
C10878 a_4365_n12325# a_4554_n13021# 0.02fF
C10879 a_5842_n13021# a_5752_n12503# 0.02fF
C10880 a_4464_n12503# a_4298_n13021# 0.04fF
C10881 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.04fF
C10882 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.02fF
C10883 a_8162_n10301# a_9450_n10301# 0.01fF
C10884 a_3077_n12325# a_3176_n12503# 0.49fF
C10885 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/A 0.02fF
C10886 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_50/X 0.01fF
C10887 a_9616_n8695# a_9706_n10301# 0.00fF
C10888 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C10889 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A 0.00fF
C10890 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X a_3436_n1079# 0.03fF
C10891 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.02fF
C10892 a_10904_n4887# a_10904_n3255# 0.00fF
C10893 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.29fF
C10894 a_3010_n5405# a_4554_n5405# 0.01fF
C10895 a_3266_n5405# a_4298_n5405# 0.02fF
C10896 a_3176_n3255# a_3010_n1597# 0.00fF
C10897 a_3077_n2997# a_3266_n1597# 0.00fF
C10898 a_8162_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.03fF
C10899 a_n1612_n7037# sky130_fd_sc_hd__clkinv_1_5/A 0.01fF
C10900 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8229_n5797# 0.01fF
C10901 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.29fF
C10902 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.05fF
C10903 a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C10904 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.09fF
C10905 a_6101_n7254# a_7212_n7203# 0.01fF
C10906 a_11164_n13591# a_10738_n13789# 0.05fF
C10907 a_10805_n9525# a_10904_n9783# 0.48fF
C10908 a_1888_n9783# a_3176_n9783# 0.01fF
C10909 sky130_fd_sc_hd__nand2_1_4/B a_5052_n7283# 0.00fF
C10910 a_1789_n9525# a_3436_n9783# 0.00fF
C10911 a_2148_n9783# a_3077_n9525# 0.02fF
C10912 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C10913 a_6874_n4317# a_6941_n4709# 0.01fF
C10914 a_6874_n2685# a_6941_n1909# 0.01fF
C10915 a_4724_n11415# a_4661_n11933# 0.01fF
C10916 a_9450_n8125# a_9450_n9213# 0.02fF
C10917 a_2729_n6493# VDD 0.35fF
C10918 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_2085_n9213# 0.01fF
C10919 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.02fF
C10920 a_7300_n10871# a_7130_n9213# 0.00fF
C10921 a_7040_n10871# a_7237_n9213# 0.00fF
C10922 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C10923 a_4724_n1079# a_4554_n2685# 0.00fF
C10924 a_4464_n1079# a_4661_n2685# 0.00fF
C10925 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6794_n7203# 0.00fF
C10926 a_501_n11237# a_1789_n11237# 0.01fF
C10927 sky130_fd_sc_hd__nand2_4_1/A a_6658_n7363# 0.03fF
C10928 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkinv_4_3/A 0.09fF
C10929 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.00fF
C10930 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VDD 0.90fF
C10931 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD 1.18fF
C10932 a_5842_n13021# a_4298_n13021# 0.01fF
C10933 Ad_b a_5052_n7283# 0.08fF
C10934 a_1789_n10613# a_1722_n10301# 0.01fF
C10935 a_3077_n4709# a_3436_n4887# 0.05fF
C10936 a_9450_n6493# a_9706_n6493# 0.19fF
C10937 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C10938 a_8328_n4887# a_8418_n5405# 0.02fF
C10939 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.03fF
C10940 sky130_fd_sc_hd__clkinv_1_4/Y a_3010_n9213# 0.00fF
C10941 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_1888_n9783# 0.01fF
C10942 sky130_fd_sc_hd__dfxbp_1_1/D a_n2163_n6671# 0.07fF
C10943 a_3266_n5405# a_1722_n5405# 0.01fF
C10944 a_3010_n5405# a_1978_n5405# 0.02fF
C10945 a_10738_n5405# a_10805_n3621# 0.00fF
C10946 a_8229_n9525# a_8229_n11237# 0.00fF
C10947 a_n2602_n7037# a_n1570_n6769# 0.14fF
C10948 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD 0.79fF
C10949 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6941_n12325# 0.01fF
C10950 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C10951 a_n2163_n6671# a_n2037_n7037# 0.02fF
C10952 a_6874_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.03fF
C10953 a_8418_n2685# a_8525_n1597# 0.00fF
C10954 a_8525_n2685# a_8418_n1597# 0.00fF
C10955 B_b Bd 0.53fF
C10956 a_3436_n12503# a_4365_n12325# 0.02fF
C10957 a_3176_n12503# a_4464_n12503# 0.01fF
C10958 a_4464_n10871# a_4464_n11415# 0.07fF
C10959 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X a_10738_n10301# 0.00fF
C10960 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.01fF
C10961 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_9876_n1079# 0.01fF
C10962 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7300_n3255# 0.03fF
C10963 a_2148_n13591# a_1978_n13021# 0.04fF
C10964 a_7237_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C10965 a_1888_n13591# a_2085_n13021# 0.02fF
C10966 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.06fF
C10967 a_4298_n5405# a_4661_n5405# 0.05fF
C10968 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.02fF
C10969 a_5842_n2685# a_5752_n1079# 0.00fF
C10970 a_8525_n6493# a_8588_n5975# 0.01fF
C10971 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VDD 0.91fF
C10972 a_7130_n6493# a_6665_n7459# 0.00fF
C10973 a_6874_n6493# a_6865_n7304# 0.01fF
C10974 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.02fF
C10975 a_7237_n6493# a_6658_n7363# 0.00fF
C10976 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_1888_n3799# 0.00fF
C10977 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A a_1789_n2997# 0.01fF
C10978 a_9616_n11415# a_9876_n11415# 0.28fF
C10979 a_3077_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C10980 a_3176_n9783# a_3436_n9783# 0.28fF
C10981 a_4464_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.03fF
C10982 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.04fF
C10983 sky130_fd_sc_hd__nand2_4_2/A a_8162_n14109# 0.03fF
C10984 a_434_n1597# a_434_n2685# 0.02fF
C10985 a_1888_n3255# a_1722_n2685# 0.04fF
C10986 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VDD 0.99fF
C10987 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C10988 a_7130_n6493# a_7130_n5405# 0.01fF
C10989 a_5752_n3799# a_5653_n4709# 0.00fF
C10990 a_5653_n3621# a_5752_n4887# 0.00fF
C10991 a_13765_n8669# VDD 2.36fF
C10992 a_1888_n12503# a_1888_n10871# 0.00fF
C10993 a_434_n5405# a_1978_n5405# 0.01fF
C10994 a_690_n5405# a_1722_n5405# 0.02fF
C10995 a_3077_n10613# VDD 0.35fF
C10996 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_1722_n13021# 0.00fF
C10997 a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.00fF
C10998 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_8588_n1079# 0.03fF
C10999 a_797_n10301# a_690_n9213# 0.00fF
C11000 sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# 0.58fF
C11001 a_7237_n1597# sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C11002 a_690_n10301# a_797_n9213# 0.00fF
C11003 a_7040_n8695# VDD 0.47fF
C11004 a_3176_n4887# a_4724_n4887# 0.01fF
C11005 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X a_8229_n5797# 0.02fF
C11006 a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C11007 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X a_9450_n5405# 0.03fF
C11008 a_3010_n10301# a_4298_n10301# 0.01fF
C11009 a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C11010 a_8162_n13021# VDD 0.75fF
C11011 a_10994_n9213# a_10904_n9783# 0.02fF
C11012 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_9616_n9783# 0.00fF
C11013 a_2366_n6493# a_2622_n6493# 0.19fF
C11014 a_7237_n13021# a_7300_n12503# 0.01fF
C11015 a_3373_n1597# a_1978_n1597# 0.01fF
C11016 sky130_fd_sc_hd__clkinv_1_0/A a_1789_n821# 0.06fF
C11017 a_8328_n10871# a_8162_n10301# 0.04fF
C11018 a_7040_n13591# a_7130_n11933# 0.00fF
C11019 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_3077_n8437# 0.18fF
C11020 a_4724_n9783# a_4724_n11415# 0.01fF
C11021 a_10738_n11933# a_10904_n13591# 0.00fF
C11022 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C11023 a_13765_n5405# A_b 2.54fF
C11024 a_4661_n5405# a_5842_n5405# 0.01fF
C11025 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5586_n5405# 0.35fF
C11026 a_3077_n1909# a_3010_n1597# 0.01fF
C11027 a_9876_n3799# a_9517_n3621# 0.05fF
C11028 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6941_n821# 0.00fF
C11029 a_2148_n13591# VDD 0.78fF
C11030 a_8588_n2167# a_8418_n1597# 0.04fF
C11031 a_8328_n2167# a_8525_n1597# 0.02fF
C11032 a_1789_n1909# a_1888_n2167# 0.49fF
C11033 a_3436_n2167# a_3436_n3255# 0.02fF
C11034 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__nand2_4_0/B 0.02fF
C11035 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A VDD 0.89fF
C11036 sky130_fd_sc_hd__clkinv_4_4/A a_860_n4887# 0.00fF
C11037 a_2366_n6493# sky130_fd_sc_hd__nand2_4_1/A 0.08fF
C11038 a_1789_n5797# a_2148_n5975# 0.05fF
C11039 a_5752_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.03fF
C11040 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X a_10904_n11415# 0.05fF
C11041 a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C11042 a_9876_n11415# a_11164_n11415# 0.01fF
C11043 a_9616_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.00fF
C11044 a_5653_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C11045 a_501_n12325# a_690_n13021# 0.02fF
C11046 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C11047 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X a_6012_n10871# 0.03fF
C11048 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.04fF
C11049 a_11101_n11933# VDD 0.32fF
C11050 a_9813_n9213# a_10738_n9213# 0.02fF
C11051 a_8162_n14109# a_9706_n14109# 0.01fF
C11052 a_8418_n14109# a_9450_n14109# 0.02fF
C11053 a_7040_n11415# a_7130_n11933# 0.02fF
C11054 a_7130_n13021# a_7130_n14109# 0.01fF
C11055 sky130_fd_sc_hd__nand2_4_2/A a_9706_n14109# 0.04fF
C11056 a_4298_n5405# a_4298_n4317# 0.02fF
C11057 a_8162_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C11058 a_9450_n1597# a_11101_n1597# 0.00fF
C11059 a_9813_n1597# a_10738_n1597# 0.02fF
C11060 a_9706_n1597# a_10994_n1597# 0.01fF
C11061 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n5405# 0.01fF
C11062 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X a_4724_n2167# 0.01fF
C11063 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C11064 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A VDD 0.89fF
C11065 a_2148_n11415# a_2085_n13021# 0.00fF
C11066 a_6874_n10301# VDD 0.76fF
C11067 a_10738_n6173# a_11101_n5405# 0.01fF
C11068 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.02fF
C11069 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VDD 0.83fF
C11070 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C11071 a_8588_n4887# a_8418_n4317# 0.04fF
C11072 a_8328_n4887# a_8525_n4317# 0.02fF
C11073 a_10904_n3799# a_10994_n2685# 0.01fF
C11074 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__nand2_4_0/Y 0.44fF
C11075 a_8588_n8695# VDD 0.79fF
C11076 a_3176_n10871# a_3266_n10301# 0.02fF
C11077 a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C11078 a_8229_n1909# a_7040_n2167# 0.01fF
C11079 a_8328_n2167# a_6941_n1909# 0.01fF
C11080 a_10805_n3621# a_10994_n4317# 0.02fF
C11081 a_10904_n3799# a_10738_n4317# 0.04fF
C11082 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X a_8328_n5975# 0.00fF
C11083 a_9876_n5975# a_8588_n5975# 0.01fF
C11084 a_4464_n2167# a_4724_n2167# 0.28fF
C11085 a_5586_n1597# a_5586_n2685# 0.02fF
C11086 a_9706_n13021# VDD 0.45fF
C11087 a_13765_n9213# a_13765_n9757# 0.34fF
C11088 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_11164_n9783# 0.33fF
C11089 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3266_n1597# 0.05fF
C11090 a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C11091 a_5752_n3255# a_6941_n2997# 0.01fF
C11092 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X a_1722_n10301# 0.01fF
C11093 a_4554_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.00fF
C11094 a_5653_n13413# a_6941_n13413# 0.01fF
C11095 a_6874_n9213# a_6794_n7203# 0.00fF
C11096 a_7237_n9213# a_6665_n7459# 0.00fF
C11097 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X a_8162_n11933# 0.00fF
C11098 a_7130_n9213# a_6865_n7304# 0.00fF
C11099 a_8229_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C11100 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_6658_n7363# 0.00fF
C11101 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X a_4464_n8695# 0.01fF
C11102 a_3436_n3255# a_3436_n4887# 0.01fF
C11103 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.03fF
C11104 a_7040_n9783# sky130_fd_sc_hd__nand2_4_3/Y 0.04fF
C11105 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X a_3373_n13021# 0.01fF
C11106 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A 1.21fF
C11107 a_600_n10871# a_860_n10871# 0.28fF
C11108 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X a_6012_n5975# 0.03fF
C11109 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X a_2148_n13591# 0.01fF
C11110 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C11111 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VDD 0.84fF
C11112 a_11164_n3799# a_9616_n3799# 0.01fF
C11113 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VDD 0.82fF
C11114 a_2085_n9213# a_3266_n9213# 0.01fF
C11115 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3010_n9213# 0.35fF
C11116 a_9706_n14109# a_9813_n13021# 0.00fF
C11117 a_8162_n8125# a_9813_n8125# 0.00fF
C11118 sky130_fd_sc_hd__nand2_4_0/Y a_7040_n2167# 0.04fF
C11119 a_1789_n1909# a_3436_n2167# 0.00fF
C11120 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X a_434_n11933# 0.03fF
C11121 a_1888_n2167# a_3176_n2167# 0.01fF
C11122 a_2148_n2167# a_3077_n1909# 0.02fF
C11123 a_1888_n5975# a_3436_n5975# 0.01fF
C11124 a_2148_n5975# a_3176_n5975# 0.02fF
C11125 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_3077_n5797# 0.18fF
C11126 a_6012_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.00fF
C11127 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X a_7300_n1079# 0.03fF
C11128 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A 2.26fF
C11129 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.37fF
C11130 a_4554_n1597# a_4724_n1079# 0.04fF
C11131 a_4661_n1597# a_4464_n1079# 0.02fF
C11132 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A VDD 0.89fF
C11133 a_2148_n13591# a_501_n13413# 0.00fF
C11134 a_10994_n9213# a_11101_n9213# 0.55fF
C11135 a_10738_n9213# sky130_fd_sc_hd__clkinv_4_10/Y 0.00fF
C11136 a_1789_n13413# a_860_n13591# 0.02fF
C11137 a_1888_n13591# a_600_n13591# 0.01fF
C11138 a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C11139 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X a_8162_n11933# 0.03fF
C11140 a_9813_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C11141 a_9450_n14109# a_9813_n14109# 0.05fF
C11142 a_3077_n2997# VDD 0.35fF
C11143 a_8525_n6493# a_8525_n5405# 0.02fF
C11144 a_1978_n1597# a_1978_n2685# 0.01fF
C11145 a_3436_n2167# a_4464_n2167# 0.02fF
C11146 a_3436_n12503# a_3436_n10871# 0.01fF
C11147 a_3176_n2167# a_4724_n2167# 0.01fF
C11148 a_5842_n13021# a_5949_n13021# 0.55fF
C11149 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__dfxbp_1_0/Q 0.03fF
C11150 a_600_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X 0.01fF
C11151 a_8588_n10871# a_9616_n10871# 0.02fF
C11152 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_9517_n10613# 0.18fF
C11153 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD 0.76fF
C11154 a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.01fF
C11155 a_5752_n9783# a_5842_n9213# 0.02fF
C11156 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD 0.84fF
C11157 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C11158 a_434_n4317# a_1722_n4317# 0.01fF
C11159 a_6874_n8125# a_6665_n7459# 0.00fF
C11160 a_8162_n1597# a_8229_n2997# 0.00fF
C11161 a_7130_n8125# a_6658_n7363# 0.01fF
C11162 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X a_5752_n2167# 0.05fF
C11163 a_3373_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.00fF
C11164 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_3436_n8695# 0.00fF
C11165 a_4464_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C11166 a_4724_n2167# a_6012_n2167# 0.01fF
C11167 a_9813_n6493# VDD 0.35fF
C11168 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.03fF
C11169 a_2148_n11415# a_2085_n10301# 0.00fF
C11170 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.08fF
C11171 Bd_b a_6006_n7607# 0.01fF
C11172 a_6941_n2997# a_7300_n3255# 0.05fF
C11173 a_501_n3621# a_434_n5405# 0.00fF
C11174 a_5842_n1597# a_5752_n1079# 0.01fF
C11175 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6874_n9213# 0.01fF
C11176 a_8418_n1597# a_8328_n1079# 0.01fF
C11177 a_8588_n13591# a_8525_n11933# 0.00fF
C11178 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.08fF
C11179 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_11101_n13021# 0.02fF
C11180 A_b Ad_b 0.33fF
C11181 a_7237_n8125# VDD 0.34fF
C11182 a_860_n10871# a_2148_n10871# 0.01fF
C11183 a_600_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C11184 a_600_n3255# VDD 0.47fF
C11185 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X a_1888_n10871# 0.05fF
C11186 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.29fF
C11187 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/Y 0.73fF
C11188 sky130_fd_sc_hd__nand2_4_0/A a_10738_n509# 0.12fF
C11189 a_690_n4317# a_797_n5405# 0.00fF
C11190 a_797_n4317# a_690_n5405# 0.00fF
C11191 a_9517_n12325# a_9706_n14109# 0.00fF
C11192 a_9616_n12503# a_9450_n14109# 0.00fF
C11193 a_501_n5797# a_600_n5975# 0.49fF
C11194 sky130_fd_sc_hd__nand2_4_2/B a_10994_n13021# 0.00fF
C11195 a_3266_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.05fF
C11196 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_4554_n9213# 0.00fF
C11197 a_9450_n8125# sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C11198 a_3176_n2167# a_3436_n2167# 0.28fF
C11199 a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.02fF
C11200 a_5752_n11415# a_5752_n10871# 0.07fF
C11201 a_3176_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.03fF
C11202 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X a_4464_n5975# 0.01fF
C11203 a_9450_n6493# a_9517_n4709# 0.00fF
C11204 a_1789_n4709# a_1888_n4887# 0.49fF
C11205 p2_b a_13765_n10301# 0.06fF
C11206 a_13765_n9213# p2d_b 0.06fF
C11207 a_8588_n11415# a_8525_n11933# 0.01fF
C11208 a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C11209 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X a_6665_n7459# 0.01fF
C11210 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.02fF
C11211 a_10994_n4317# a_11164_n4887# 0.04fF
C11212 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C11213 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X a_7300_n3799# 0.01fF
C11214 a_4464_n3255# VDD 0.46fF
C11215 a_9450_n1597# a_9616_n3255# 0.00fF
C11216 a_3010_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.01fF
C11217 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X a_5752_n2167# 0.01fF
C11218 a_10738_n6173# sky130_fd_sc_hd__clkinv_4_3/A 0.49fF
C11219 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.02fF
C11220 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_7130_n13021# 0.03fF
C11221 a_5842_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C11222 a_5949_n13021# a_7237_n13021# 0.01fF
C11223 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8162_n14109# 0.34fF
C11224 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C11225 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_10904_n10871# 0.01fF
C11226 a_9616_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.03fF
C11227 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.04fF
C11228 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.42fF
C11229 a_3176_n8695# a_3010_n9213# 0.04fF
C11230 a_3077_n8437# a_3266_n9213# 0.02fF
C11231 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.06fF
C11232 a_9876_n3799# a_10805_n3621# 0.02fF
C11233 sky130_fd_sc_hd__mux2_1_0/X VDD 1.02fF
C11234 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.29fF
C11235 a_8418_n14109# a_8229_n13413# 0.02fF
C11236 a_8162_n14109# a_8328_n13591# 0.04fF
C11237 Bd_b sky130_fd_sc_hd__clkinv_4_3/Y 0.18fF
C11238 a_7040_n3255# a_8588_n3255# 0.01fF
C11239 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X a_8229_n2997# 0.18fF
C11240 a_7300_n3255# a_8328_n3255# 0.02fF
C11241 a_4661_n5405# a_5949_n5405# 0.01fF
C11242 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6941_n821# 0.01fF
C11243 a_6874_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X 0.03fF
C11244 a_4554_n5405# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C11245 a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C11246 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X a_10738_n13021# 0.03fF
C11247 p2d a_13765_n8669# 0.06fF
C11248 a_11164_n8695# sky130_fd_sc_hd__nand2_4_3/A 0.04fF
C11249 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.00fF
C11250 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A 0.32fF
C11251 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VDD 0.94fF
C11252 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C11253 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_3/A 0.26fF
C11254 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C11255 a_n2163_n6671# a_n1570_n6769# 0.05fF
C11256 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.29fF
C11257 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.03fF
C11258 a_9616_n11415# a_9616_n9783# 0.00fF
C11259 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X a_9813_n5405# 0.01fF
C11260 a_860_n2167# a_860_n1079# 0.02fF
C11261 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4661_n9213# 0.02fF
C11262 a_3373_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C11263 a_3266_n10301# a_3077_n9525# 0.02fF
C11264 a_3010_n10301# a_3176_n9783# 0.04fF
C11265 a_7237_n1597# VDD 0.35fF
C11266 a_5586_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C11267 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X a_4724_n5975# 0.03fF
C11268 a_5949_n9213# a_4298_n9213# 0.00fF
C11269 a_8588_n11415# a_8525_n10301# 0.00fF
C11270 a_9616_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C11271 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X a_10738_n1597# 0.03fF
C11272 a_2085_n4317# VDD 0.35fF
C11273 a_3436_n3799# a_3266_n2685# 0.00fF
C11274 a_3176_n3799# a_3373_n2685# 0.00fF
C11275 a_4554_n10301# a_4661_n10301# 0.55fF
C11276 a_4298_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C11277 a_1888_n4887# a_3176_n4887# 0.01fF
C11278 a_2148_n4887# a_3077_n4709# 0.02fF
C11279 a_2366_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C11280 a_3077_n3621# a_3077_n2997# 0.05fF
C11281 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X sky130_fd_sc_hd__clkinv_1_0/A 0.02fF
C11282 Ad_b sky130_fd_sc_hd__nand2_4_3/A 0.32fF
C11283 sky130_fd_sc_hd__clkinv_4_3/A Ad 0.01fF
C11284 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A Ad_b 0.03fF
C11285 a_600_n10871# a_600_n9783# 0.01fF
C11286 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_25/A 0.03fF
C11287 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X a_2085_n2685# 0.01fF
C11288 a_1978_n9213# a_3266_n9213# 0.01fF
C11289 a_1722_n9213# a_3373_n9213# 0.00fF
C11290 a_9616_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.05fF
C11291 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X a_8328_n3255# 0.00fF
C11292 a_9876_n3255# a_8588_n3255# 0.01fF
C11293 a_4365_n10613# a_4298_n9213# 0.00fF
C11294 sky130_fd_sc_hd__nand2_4_3/Y a_7237_n9213# 0.05fF
C11295 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_9706_n14109# 0.00fF
C11296 a_7237_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.12fF
C11297 a_9450_n5405# a_9517_n3621# 0.00fF
C11298 a_1888_n13591# a_1722_n11933# 0.00fF
C11299 a_1789_n13413# a_1978_n11933# 0.00fF
C11300 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.06fF
C11301 a_6941_n13413# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C11302 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X a_11164_n10871# 0.03fF
C11303 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.06fF
C11304 a_10904_n10871# a_10738_n11933# 0.00fF
C11305 a_10805_n10613# a_10994_n11933# 0.00fF
C11306 sky130_fd_sc_hd__clkinv_4_3/A a_7040_n4887# 0.04fF
C11307 a_5653_n1909# VDD 0.35fF
C11308 a_8229_n9525# a_8418_n9213# 0.02fF
C11309 a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A 0.01fF
C11310 a_6874_n509# a_7237_n509# 0.05fF
C11311 a_10904_n3799# a_11164_n3799# 0.23fF
C11312 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C11313 a_4724_n12503# a_5653_n12325# 0.02fF
C11314 a_9813_n6493# a_9706_n5405# 0.00fF
C11315 a_10904_n1079# a_10738_n2685# 0.00fF
C11316 a_10805_n821# a_10994_n2685# 0.00fF
C11317 a_600_n8695# a_1789_n8437# 0.01fF
C11318 a_501_n8437# a_1888_n8695# 0.01fF
C11319 a_8328_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C11320 a_8418_n6493# a_9450_n6493# 0.02fF
C11321 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_161/A 0.03fF
C11322 a_1888_n3799# a_1978_n5405# 0.00fF
C11323 a_9517_n12325# a_10904_n12503# 0.01fF
C11324 a_9616_n12503# a_10805_n12325# 0.01fF
C11325 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X a_9876_n2167# 0.03fF
C11326 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C11327 a_11164_n12503# a_11101_n13021# 0.01fF
C11328 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_10994_n13021# 0.04fF
C11329 a_3077_n10613# a_3010_n11933# 0.00fF
C11330 a_7300_n4887# sky130_fd_sc_hd__clkinv_4_3/A 0.10fF
C11331 a_13765_n9213# VDD 2.00fF
C11332 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/X 0.02fF
C11333 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkinv_4_4/A 0.02fF
C11334 a_690_n4317# a_600_n4887# 0.01fF
C11335 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.02fF
C11336 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A 0.00fF
C11337 a_5052_n7283# a_6006_n7607# 0.02fF
C11338 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A VDD 0.89fF
C11339 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A VDD 0.88fF
C11340 a_5949_n4317# a_5949_n2685# 0.01fF
C11341 a_6874_n9213# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C11342 sky130_fd_sc_hd__clkinv_4_8/Y a_10904_n13591# 0.02fF
C11343 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A VDD 0.88fF
C11344 a_11164_n2167# a_11101_n1597# 0.01fF
C11345 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X a_11164_n3255# 0.03fF
C11346 a_5949_n9213# a_5842_n9213# 0.55fF
C11347 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_5586_n9213# 0.03fF
C11348 a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.01fF
C11349 a_7300_n11415# a_7300_n10871# 0.09fF
C11350 a_5842_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.05fF
C11351 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5842_n10301# 0.03fF
C11352 a_4661_n10301# a_5949_n10301# 0.01fF
C11353 a_4554_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C11354 a_5653_n2997# a_5842_n4317# 0.00fF
C11355 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C11356 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.06fF
C11357 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C11358 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8525_n11933# 0.00fF
C11359 a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.00fF
C11360 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X a_501_n12325# 0.02fF
C11361 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_9450_n9213# 0.00fF
C11362 a_6941_n9525# a_6941_n8437# 0.02fF
C11363 a_860_n2167# a_797_n1597# 0.01fF
C11364 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.44fF
C11365 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.02fF
C11366 a_5752_n9783# a_5752_n10871# 0.01fF
C11367 a_5842_n1597# a_6874_n1597# 0.02fF
C11368 a_9876_n13591# a_9813_n13021# 0.01fF
C11369 a_8328_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C11370 a_4464_n9783# a_6012_n9783# 0.01fF
C11371 a_4724_n9783# a_5752_n9783# 0.02fF
C11372 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_5653_n9525# 0.18fF
C11373 sky130_fd_sc_hd__nand2_4_2/A a_10738_n13789# 0.11fF
C11374 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_797_n4317# 0.01fF
C11375 a_4724_n8695# a_4554_n9213# 0.04fF
C11376 a_4464_n8695# a_4661_n9213# 0.02fF
C11377 a_9706_n1597# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C11378 a_6665_n7459# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.02fF
C11379 a_7040_n2167# VDD 0.46fF
C11380 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkinv_4_4/A 0.08fF
C11381 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8162_n509# 0.35fF
C11382 a_7130_n509# a_8525_n509# 0.01fF
C11383 a_7237_n509# a_8418_n509# 0.01fF
C11384 a_690_n2685# VDD 0.45fF
C11385 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X a_6941_n12325# 0.01fF
C11386 a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.02fF
C11387 a_5752_n12503# a_6012_n12503# 0.28fF
C11388 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X a_4464_n4887# 0.05fF
C11389 a_3436_n4887# a_4724_n4887# 0.01fF
C11390 a_10805_n4709# a_10904_n5975# 0.00fF
C11391 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.00fF
C11392 a_9813_n14109# a_9616_n13591# 0.02fF
C11393 a_9706_n14109# a_9876_n13591# 0.04fF
C11394 a_10904_n4887# a_10805_n5797# 0.00fF
C11395 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X a_3373_n5405# 0.00fF
C11396 a_6941_n5797# a_7040_n4887# 0.00fF
C11397 a_7040_n5975# a_6941_n4709# 0.00fF
C11398 a_8162_n13021# a_8162_n11933# 0.02fF
C11399 a_10805_n12325# a_11164_n12503# 0.05fF
C11400 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkinv_4_3/A 0.70fF
C11401 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.06fF
C11402 a_n2068_n6671# VDD 0.02fF
C11403 a_3176_n5975# a_3373_n5405# 0.02fF
C11404 a_8229_n10613# a_8328_n12503# 0.00fF
C11405 a_8328_n10871# a_8229_n12325# 0.00fF
C11406 a_3436_n5975# a_3266_n5405# 0.04fF
C11407 a_11164_n11415# a_11164_n9783# 0.01fF
C11408 a_10738_n8125# a_10805_n8437# 0.03fF
C11409 a_1888_n11415# a_1978_n11933# 0.02fF
C11410 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/X 0.01fF
C11411 a_5949_n4317# a_6012_n3255# 0.00fF
C11412 a_6941_n3621# a_7040_n3799# 0.49fF
C11413 a_9616_n2167# a_9616_n3255# 0.01fF
C11414 a_4365_n4709# VDD 0.36fF
C11415 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VDD 1.23fF
C11416 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_5842_n9213# 0.01fF
C11417 a_5949_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.12fF
C11418 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X a_4661_n2685# 0.00fF
C11419 a_6941_n13413# a_8328_n13591# 0.01fF
C11420 a_7040_n13591# a_8229_n13413# 0.01fF
C11421 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C11422 a_5949_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C11423 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_7237_n11933# 0.02fF
C11424 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.03fF
C11425 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X a_8525_n10301# 0.01fF
C11426 a_7130_n9213# a_8162_n9213# 0.02fF
C11427 a_6874_n9213# a_8418_n9213# 0.01fF
C11428 a_4464_n3799# a_4464_n3255# 0.07fF
C11429 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.01fF
C11430 a_9813_n11933# a_9450_n11933# 0.05fF
C11431 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11164_n4887# 0.03fF
C11432 a_690_n4317# a_860_n3799# 0.04fF
C11433 a_797_n4317# a_600_n3799# 0.02fF
C11434 a_3010_n13021# a_4298_n13021# 0.01fF
C11435 a_2148_n10871# a_2148_n9783# 0.02fF
C11436 a_9450_n6493# a_9616_n5975# 0.04fF
C11437 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X a_600_n5975# 0.03fF
C11438 p1 sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C11439 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.01fF
C11440 a_3176_n13591# a_3373_n11933# 0.00fF
C11441 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_1789_n13413# 0.01fF
C11442 a_3436_n13591# a_3266_n11933# 0.00fF
C11443 a_9706_n14109# a_10738_n13789# 0.01fF
C11444 a_10805_n11237# a_10994_n10301# 0.00fF
C11445 a_10904_n11415# a_10738_n10301# 0.00fF
C11446 a_9616_n12503# a_9616_n13591# 0.01fF
C11447 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X a_7040_n9783# 0.01fF
C11448 a_9876_n13591# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C11449 sky130_fd_sc_hd__clkinv_1_0/A VDD 6.18fF
C11450 a_3077_n12325# a_4724_n12503# 0.00fF
C11451 a_2148_n5975# a_1978_n5405# 0.04fF
C11452 a_6941_n12325# VDD 0.35fF
C11453 a_8418_n509# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.05fF
C11454 a_2085_n2685# VDD 0.35fF
C11455 a_501_n12325# a_600_n13591# 0.00fF
C11456 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X a_7040_n12503# 0.05fF
C11457 a_4724_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.29fF
C11458 a_6012_n12503# a_7300_n12503# 0.01fF
C11459 a_5752_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C11460 a_1888_n3255# a_3077_n2997# 0.01fF
C11461 a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C11462 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_7/Y 0.14fF
C11463 a_501_n9525# a_600_n9783# 0.49fF
C11464 a_8162_n2685# a_8229_n3621# 0.00fF
C11465 a_11164_n8695# a_11164_n9783# 0.02fF
C11466 clk VDD 2.76fF
C11467 a_n787_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C11468 a_8229_n4709# a_8328_n3255# 0.00fF
C11469 a_8328_n4887# a_8229_n2997# 0.00fF
C11470 a_13765_n2685# a_13765_n4317# 0.04fF
C11471 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C11472 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.07fF
C11473 a_9813_n6493# a_9813_n5405# 0.02fF
C11474 a_5586_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.35fF
C11475 a_5842_n4317# a_4661_n4317# 0.01fF
C11476 a_5949_n4317# a_4554_n4317# 0.01fF
C11477 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.01fF
C11478 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X a_3010_n11933# 0.03fF
C11479 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_8588_n9783# 0.01fF
C11480 a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C11481 a_7040_n3799# a_8328_n3799# 0.01fF
C11482 a_7300_n3799# a_8229_n3621# 0.02fF
C11483 a_6941_n11237# a_8328_n11415# 0.01fF
C11484 a_7040_n11415# a_8229_n11237# 0.01fF
C11485 a_3436_n3799# a_3266_n4317# 0.04fF
C11486 a_3176_n3799# a_3373_n4317# 0.02fF
C11487 a_6941_n3621# a_8588_n3799# 0.00fF
C11488 a_4464_n8695# a_5653_n8437# 0.01fF
C11489 a_4365_n8437# a_5752_n8695# 0.01fF
C11490 a_5752_n4887# VDD 0.44fF
C11491 a_5752_n13591# a_5949_n11933# 0.00fF
C11492 a_501_n3621# a_1888_n3799# 0.01fF
C11493 a_600_n3799# a_1789_n3621# 0.01fF
C11494 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.02fF
C11495 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/A 0.01fF
C11496 a_8229_n13413# a_8588_n13591# 0.05fF
C11497 a_3176_n5975# a_3010_n4317# 0.00fF
C11498 a_3077_n5797# a_3266_n4317# 0.00fF
C11499 a_8162_n9213# a_8525_n9213# 0.05fF
C11500 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X a_n688_n4887# 0.02fF
C11501 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.06fF
C11502 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.85fF
C11503 a_10738_n5405# a_10738_n4317# 0.02fF
C11504 a_1888_n3255# a_600_n3255# 0.01fF
C11505 a_4298_n13021# a_4554_n13021# 0.19fF
C11506 a_11164_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.03fF
C11507 a_10904_n8695# a_10738_n10301# 0.00fF
C11508 a_10805_n8437# a_10994_n10301# 0.00fF
C11509 a_11101_n11933# a_9706_n11933# 0.01fF
C11510 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C11511 a_3077_n12325# a_3266_n13021# 0.02fF
C11512 sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# 0.58fF
C11513 a_3176_n12503# a_3010_n13021# 0.04fF
C11514 a_1789_n12325# a_1888_n12503# 0.49fF
C11515 a_7300_n9783# a_7300_n10871# 0.02fF
C11516 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_8418_n10301# 0.00fF
C11517 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/A 0.04fF
C11518 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C11519 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X a_5653_n12325# 0.01fF
C11520 a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.02fF
C11521 a_4464_n12503# a_4724_n12503# 0.28fF
C11522 a_8328_n12503# VDD 0.44fF
C11523 a_9616_n4887# a_9616_n3255# 0.00fF
C11524 sky130_fd_sc_hd__dfxbp_1_0/Q a_6665_n7459# 0.04fF
C11525 a_9706_n6493# a_9517_n4709# 0.00fF
C11526 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6941_n5797# 0.01fF
C11527 a_6874_n6493# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.03fF
C11528 a_9616_n8695# a_9450_n9213# 0.04fF
C11529 a_9517_n8437# a_9706_n9213# 0.02fF
C11530 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.29fF
C11531 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.02fF
C11532 a_9706_n13021# a_9706_n11933# 0.01fF
C11533 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.06fF
C11534 a_9517_n9525# a_9616_n9783# 0.49fF
C11535 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C11536 a_860_n9783# a_1789_n9525# 0.02fF
C11537 a_600_n9783# a_1888_n9783# 0.01fF
C11538 a_501_n9525# a_2148_n9783# 0.00fF
C11539 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.03fF
C11540 a_6941_n8437# a_7130_n9213# 0.02fF
C11541 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1789_n8437# 0.00fF
C11542 a_501_n12325# a_690_n11933# 0.02fF
C11543 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.02fF
C11544 a_5586_n4317# a_5653_n4709# 0.01fF
C11545 a_9517_n5797# a_10904_n5975# 0.01fF
C11546 a_860_n8695# a_690_n9213# 0.04fF
C11547 a_7130_n4317# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C11548 a_9616_n5975# a_10805_n5797# 0.01fF
C11549 a_600_n8695# a_797_n9213# 0.02fF
C11550 a_3436_n11415# a_3373_n11933# 0.01fF
C11551 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C11552 a_8162_n8125# a_8162_n9213# 0.02fF
C11553 a_5752_n10871# a_5949_n9213# 0.00fF
C11554 a_8229_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C11555 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X a_9517_n3621# 0.01fF
C11556 a_8588_n4887# a_8588_n5975# 0.02fF
C11557 a_3436_n1079# a_3266_n2685# 0.00fF
C11558 a_8328_n3799# a_8588_n3799# 0.28fF
C11559 a_3176_n1079# a_3373_n2685# 0.00fF
C11560 a_8229_n11237# a_8588_n11415# 0.05fF
C11561 a_5653_n8437# a_6012_n8695# 0.05fF
C11562 a_7130_n5405# a_6941_n4709# 0.02fF
C11563 a_4365_n13413# a_5752_n13591# 0.01fF
C11564 a_4464_n13591# a_5653_n13413# 0.01fF
C11565 a_6874_n5405# a_7040_n4887# 0.04fF
C11566 a_11164_n2167# a_11164_n3255# 0.02fF
C11567 a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C11568 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X a_3077_n8437# 0.01fF
C11569 a_8229_n1909# a_8229_n3621# 0.00fF
C11570 a_8588_n13591# a_9616_n13591# 0.02fF
C11571 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X a_9517_n13413# 0.18fF
C11572 a_8328_n13591# a_9876_n13591# 0.01fF
C11573 a_7130_n14109# a_7300_n12503# 0.00fF
C11574 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C11575 sky130_fd_sc_hd__clkinv_1_0/A a_9876_n1079# 0.12fF
C11576 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n10301# 0.00fF
C11577 a_7237_n14109# a_7040_n12503# 0.00fF
C11578 a_8525_n9213# a_9706_n9213# 0.01fF
C11579 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_9450_n9213# 0.35fF
C11580 a_10738_n11933# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C11581 a_1789_n1909# a_1789_n821# 0.02fF
C11582 a_10904_n12503# a_10738_n13789# 0.00fF
C11583 a_9450_n4317# a_10738_n4317# 0.01fF
C11584 a_690_n1597# a_600_n3255# 0.00fF
C11585 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.06fF
C11586 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C11587 a_5586_n13021# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C11588 a_5752_n10871# a_4365_n10613# 0.01fF
C11589 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD 0.86fF
C11590 a_9450_n2685# a_10994_n2685# 0.01fF
C11591 a_11101_n9213# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C11592 p2d a_13765_n9213# 0.15fF
C11593 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.04fF
C11594 a_9706_n2685# a_10738_n2685# 0.02fF
C11595 a_6941_n9525# a_6941_n11237# 0.00fF
C11596 a_2148_n3799# a_2148_n4887# 0.02fF
C11597 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_11101_n9213# 0.01fF
C11598 a_1888_n12503# a_3176_n12503# 0.01fF
C11599 a_1789_n12325# a_3436_n12503# 0.00fF
C11600 a_2148_n12503# a_3077_n12325# 0.02fF
C11601 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C11602 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X a_4661_n11933# 0.00fF
C11603 a_7237_n2685# a_7130_n1597# 0.00fF
C11604 a_7130_n2685# a_7237_n1597# 0.00fF
C11605 a_1888_n3255# a_2085_n4317# 0.00fF
C11606 a_4365_n12325# VDD 0.36fF
C11607 a_4554_n2685# a_5586_n2685# 0.02fF
C11608 a_4298_n2685# a_5842_n2685# 0.01fF
C11609 a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C11610 a_5752_n3799# a_5752_n2167# 0.00fF
C11611 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X a_9450_n10301# 0.00fF
C11612 a_2622_n8125# sky130_fd_sc_hd__clkinv_1_3/Y 0.03fF
C11613 a_4464_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C11614 sky130_fd_sc_hd__clkinv_1_6/Y a_n787_n12325# 0.00fF
C11615 a_9706_n4317# a_9616_n3799# 0.02fF
C11616 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.02fF
C11617 a_3010_n5405# a_3373_n5405# 0.05fF
C11618 a_7237_n6493# a_7300_n5975# 0.01fF
C11619 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.02fF
C11620 a_6874_n14109# a_7130_n14109# 0.19fF
C11621 p1d_b p1d 0.47fF
C11622 a_9876_n9783# a_10805_n9525# 0.02fF
C11623 a_9517_n9525# a_11164_n9783# 0.00fF
C11624 a_9616_n9783# a_10904_n9783# 0.01fF
C11625 a_1789_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.02fF
C11626 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X a_3077_n9525# 0.01fF
C11627 a_1888_n9783# a_2148_n9783# 0.28fF
C11628 a_9706_n2685# a_9616_n3799# 0.01fF
C11629 a_10738_n13789# VSS 1.09fF
C11630 a_n860_n13789# VSS 0.01fF
C11631 sky130_fd_sc_hd__nand2_4_2/B VSS 1.06fF
C11632 a_9813_n14109# VSS 0.32fF
C11633 a_9706_n14109# VSS 0.41fF
C11634 a_9450_n14109# VSS 0.58fF
C11635 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS 0.81fF
C11636 a_8525_n14109# VSS 0.32fF
C11637 a_8418_n14109# VSS 0.41fF
C11638 a_8162_n14109# VSS 0.58fF
C11639 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS 0.81fF
C11640 a_7237_n14109# VSS 0.32fF
C11641 a_7130_n14109# VSS 0.41fF
C11642 a_6874_n14109# VSS 0.57fF
C11643 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS 2.07fF
C11644 a_2729_n14109# VSS 0.33fF
C11645 a_2622_n14109# VSS 0.41fF
C11646 a_2366_n14109# VSS 0.58fF
C11647 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A VSS 1.03fF
C11648 sky130_fd_sc_hd__nand2_4_2/A VSS 4.02fF
C11649 p1 VSS 2.96fF
C11650 a_13765_n13565# VSS 2.07fF
C11651 a_11164_n13591# VSS 0.52fF
C11652 a_10904_n13591# VSS 0.37fF
C11653 a_10805_n13413# VSS 0.31fF
C11654 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS 0.87fF
C11655 a_9876_n13591# VSS 0.59fF
C11656 a_9616_n13591# VSS 0.41fF
C11657 a_9517_n13413# VSS 0.33fF
C11658 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS 0.83fF
C11659 a_8588_n13591# VSS 0.61fF
C11660 a_8328_n13591# VSS 0.41fF
C11661 a_8229_n13413# VSS 0.33fF
C11662 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS 0.84fF
C11663 a_7300_n13591# VSS 0.61fF
C11664 a_7040_n13591# VSS 0.41fF
C11665 a_6941_n13413# VSS 0.33fF
C11666 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS 0.85fF
C11667 a_6012_n13591# VSS 0.62fF
C11668 a_5752_n13591# VSS 0.43fF
C11669 a_5653_n13413# VSS 0.34fF
C11670 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS 0.84fF
C11671 a_4724_n13591# VSS 0.61fF
C11672 a_4464_n13591# VSS 0.42fF
C11673 a_4365_n13413# VSS 0.34fF
C11674 sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VSS 0.85fF
C11675 a_3436_n13591# VSS 0.60fF
C11676 a_3176_n13591# VSS 0.41fF
C11677 a_3077_n13413# VSS 0.34fF
C11678 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS 0.84fF
C11679 a_2148_n13591# VSS 0.60fF
C11680 a_1888_n13591# VSS 0.41fF
C11681 a_1789_n13413# VSS 0.34fF
C11682 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS 0.84fF
C11683 a_860_n13591# VSS 0.61fF
C11684 a_600_n13591# VSS 0.42fF
C11685 a_501_n13413# VSS 0.35fF
C11686 p1_b VSS 3.36fF
C11687 a_13765_n13021# VSS 2.12fF
C11688 sky130_fd_sc_hd__clkinv_4_7/Y VSS 1.92fF
C11689 sky130_fd_sc_hd__clkinv_4_7/A VSS 12.47fF
C11690 a_11101_n13021# VSS 0.33fF
C11691 a_10994_n13021# VSS 0.43fF
C11692 a_10738_n13021# VSS 0.61fF
C11693 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS 0.91fF
C11694 a_9813_n13021# VSS 0.33fF
C11695 a_9706_n13021# VSS 0.43fF
C11696 a_9450_n13021# VSS 0.62fF
C11697 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A VSS 0.91fF
C11698 a_8525_n13021# VSS 0.34fF
C11699 a_8418_n13021# VSS 0.44fF
C11700 a_8162_n13021# VSS 0.63fF
C11701 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X VSS 0.91fF
C11702 a_7237_n13021# VSS 0.34fF
C11703 a_7130_n13021# VSS 0.44fF
C11704 a_6874_n13021# VSS 0.63fF
C11705 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A VSS 0.91fF
C11706 a_5949_n13021# VSS 0.34fF
C11707 a_5842_n13021# VSS 0.44fF
C11708 a_5586_n13021# VSS 0.63fF
C11709 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS 0.91fF
C11710 a_4661_n13021# VSS 0.34fF
C11711 a_4554_n13021# VSS 0.44fF
C11712 a_4298_n13021# VSS 0.63fF
C11713 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X VSS 0.91fF
C11714 a_3373_n13021# VSS 0.34fF
C11715 a_3266_n13021# VSS 0.44fF
C11716 a_3010_n13021# VSS 0.63fF
C11717 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS 0.91fF
C11718 a_2085_n13021# VSS 0.34fF
C11719 a_1978_n13021# VSS 0.44fF
C11720 a_1722_n13021# VSS 0.63fF
C11721 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A VSS 0.91fF
C11722 a_797_n13021# VSS 0.34fF
C11723 a_690_n13021# VSS 0.44fF
C11724 a_434_n13021# VSS 0.63fF
C11725 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS 0.59fF
C11726 p1d VSS 3.18fF
C11727 a_13765_n12477# VSS 2.24fF
C11728 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS 0.71fF
C11729 a_11164_n12503# VSS 0.57fF
C11730 a_10904_n12503# VSS 0.41fF
C11731 a_10805_n12325# VSS 0.34fF
C11732 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS 0.91fF
C11733 a_9876_n12503# VSS 0.62fF
C11734 a_9616_n12503# VSS 0.43fF
C11735 a_9517_n12325# VSS 0.35fF
C11736 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS 0.88fF
C11737 a_8588_n12503# VSS 0.64fF
C11738 a_8328_n12503# VSS 0.44fF
C11739 a_8229_n12325# VSS 0.35fF
C11740 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS 0.88fF
C11741 a_7300_n12503# VSS 0.64fF
C11742 a_7040_n12503# VSS 0.44fF
C11743 a_6941_n12325# VSS 0.35fF
C11744 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS 0.88fF
C11745 a_6012_n12503# VSS 0.63fF
C11746 a_5752_n12503# VSS 0.43fF
C11747 a_5653_n12325# VSS 0.35fF
C11748 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS 0.89fF
C11749 a_4724_n12503# VSS 0.64fF
C11750 a_4464_n12503# VSS 0.44fF
C11751 a_4365_n12325# VSS 0.35fF
C11752 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS 0.88fF
C11753 a_3436_n12503# VSS 0.64fF
C11754 a_3176_n12503# VSS 0.44fF
C11755 a_3077_n12325# VSS 0.35fF
C11756 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS 0.88fF
C11757 a_2148_n12503# VSS 0.64fF
C11758 a_1888_n12503# VSS 0.44fF
C11759 a_1789_n12325# VSS 0.35fF
C11760 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS 0.89fF
C11761 a_860_n12503# VSS 0.64fF
C11762 a_600_n12503# VSS 0.44fF
C11763 a_501_n12325# VSS 0.35fF
C11764 a_n428_n12503# VSS 0.70fF
C11765 a_n688_n12503# VSS 0.48fF
C11766 a_n787_n12325# VSS 0.38fF
C11767 p1d_b VSS 3.37fF
C11768 a_13765_n11933# VSS 2.19fF
C11769 sky130_fd_sc_hd__clkinv_4_8/Y VSS 2.71fF
C11770 sky130_fd_sc_hd__clkinv_4_8/A VSS 8.50fF
C11771 a_11101_n11933# VSS 0.33fF
C11772 a_10994_n11933# VSS 0.43fF
C11773 a_10738_n11933# VSS 0.61fF
C11774 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS 0.92fF
C11775 a_9813_n11933# VSS 0.33fF
C11776 a_9706_n11933# VSS 0.43fF
C11777 a_9450_n11933# VSS 0.62fF
C11778 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A VSS 0.91fF
C11779 a_8525_n11933# VSS 0.34fF
C11780 a_8418_n11933# VSS 0.44fF
C11781 a_8162_n11933# VSS 0.63fF
C11782 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS 0.92fF
C11783 a_7237_n11933# VSS 0.34fF
C11784 a_7130_n11933# VSS 0.44fF
C11785 a_6874_n11933# VSS 0.63fF
C11786 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A VSS 0.92fF
C11787 a_5949_n11933# VSS 0.34fF
C11788 a_5842_n11933# VSS 0.44fF
C11789 a_5586_n11933# VSS 0.63fF
C11790 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS 0.92fF
C11791 a_4661_n11933# VSS 0.34fF
C11792 a_4554_n11933# VSS 0.44fF
C11793 a_4298_n11933# VSS 0.63fF
C11794 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A VSS 0.92fF
C11795 a_3373_n11933# VSS 0.34fF
C11796 a_3266_n11933# VSS 0.44fF
C11797 a_3010_n11933# VSS 0.63fF
C11798 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS 0.92fF
C11799 a_2085_n11933# VSS 0.34fF
C11800 a_1978_n11933# VSS 0.44fF
C11801 a_1722_n11933# VSS 0.63fF
C11802 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A VSS 0.92fF
C11803 a_797_n11933# VSS 0.35fF
C11804 a_690_n11933# VSS 0.44fF
C11805 a_434_n11933# VSS 0.63fF
C11806 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS 0.60fF
C11807 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS 1.20fF
C11808 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS 0.66fF
C11809 a_11164_n11415# VSS 0.57fF
C11810 a_10904_n11415# VSS 0.40fF
C11811 a_10805_n11237# VSS 0.34fF
C11812 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS 0.93fF
C11813 a_9876_n11415# VSS 0.62fF
C11814 a_9616_n11415# VSS 0.43fF
C11815 a_9517_n11237# VSS 0.35fF
C11816 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS 0.90fF
C11817 a_8588_n11415# VSS 0.64fF
C11818 a_8328_n11415# VSS 0.44fF
C11819 a_8229_n11237# VSS 0.36fF
C11820 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS 0.90fF
C11821 a_7300_n11415# VSS 0.64fF
C11822 a_7040_n11415# VSS 0.44fF
C11823 a_6941_n11237# VSS 0.36fF
C11824 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS 0.90fF
C11825 a_6012_n11415# VSS 0.64fF
C11826 a_5752_n11415# VSS 0.44fF
C11827 a_5653_n11237# VSS 0.36fF
C11828 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS 0.90fF
C11829 a_4724_n11415# VSS 0.64fF
C11830 a_4464_n11415# VSS 0.44fF
C11831 a_4365_n11237# VSS 0.36fF
C11832 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS 0.90fF
C11833 a_3436_n11415# VSS 0.64fF
C11834 a_3176_n11415# VSS 0.44fF
C11835 a_3077_n11237# VSS 0.36fF
C11836 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS 0.90fF
C11837 a_2148_n11415# VSS 0.64fF
C11838 a_1888_n11415# VSS 0.44fF
C11839 a_1789_n11237# VSS 0.36fF
C11840 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS 0.92fF
C11841 a_860_n11415# VSS 0.65fF
C11842 a_600_n11415# VSS 0.44fF
C11843 a_501_n11237# VSS 0.36fF
C11844 sky130_fd_sc_hd__clkinv_1_6/Y VSS 1.44fF
C11845 a_11164_n10871# VSS 0.56fF
C11846 a_10904_n10871# VSS 0.39fF
C11847 a_10805_n10613# VSS 0.34fF
C11848 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS 0.88fF
C11849 a_9876_n10871# VSS 0.62fF
C11850 a_9616_n10871# VSS 0.41fF
C11851 a_9517_n10613# VSS 0.35fF
C11852 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS 0.90fF
C11853 a_8588_n10871# VSS 0.64fF
C11854 a_8328_n10871# VSS 0.42fF
C11855 a_8229_n10613# VSS 0.36fF
C11856 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS 0.90fF
C11857 a_7300_n10871# VSS 0.64fF
C11858 a_7040_n10871# VSS 0.42fF
C11859 a_6941_n10613# VSS 0.36fF
C11860 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS 0.90fF
C11861 a_6012_n10871# VSS 0.64fF
C11862 a_5752_n10871# VSS 0.42fF
C11863 a_5653_n10613# VSS 0.36fF
C11864 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS 0.90fF
C11865 a_4724_n10871# VSS 0.64fF
C11866 a_4464_n10871# VSS 0.42fF
C11867 a_4365_n10613# VSS 0.36fF
C11868 sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VSS 0.90fF
C11869 a_3436_n10871# VSS 0.64fF
C11870 a_3176_n10871# VSS 0.42fF
C11871 a_3077_n10613# VSS 0.36fF
C11872 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS 0.90fF
C11873 a_2148_n10871# VSS 0.64fF
C11874 a_1888_n10871# VSS 0.42fF
C11875 a_1789_n10613# VSS 0.36fF
C11876 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS 0.85fF
C11877 a_860_n10871# VSS 0.64fF
C11878 a_600_n10871# VSS 0.43fF
C11879 a_501_n10613# VSS 0.37fF
C11880 p2d_b VSS 3.24fF
C11881 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A VSS 0.71fF
C11882 a_13765_n10301# VSS 2.38fF
C11883 a_11101_n10301# VSS 0.33fF
C11884 a_10994_n10301# VSS 0.44fF
C11885 a_10738_n10301# VSS 0.62fF
C11886 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS 0.92fF
C11887 a_9813_n10301# VSS 0.33fF
C11888 a_9706_n10301# VSS 0.45fF
C11889 a_9450_n10301# VSS 0.63fF
C11890 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A VSS 0.92fF
C11891 a_8525_n10301# VSS 0.34fF
C11892 a_8418_n10301# VSS 0.45fF
C11893 a_8162_n10301# VSS 0.63fF
C11894 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS 0.92fF
C11895 a_7237_n10301# VSS 0.34fF
C11896 a_7130_n10301# VSS 0.45fF
C11897 a_6874_n10301# VSS 0.63fF
C11898 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A VSS 0.92fF
C11899 a_5949_n10301# VSS 0.34fF
C11900 a_5842_n10301# VSS 0.45fF
C11901 a_5586_n10301# VSS 0.63fF
C11902 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS 0.92fF
C11903 a_4661_n10301# VSS 0.34fF
C11904 a_4554_n10301# VSS 0.45fF
C11905 a_4298_n10301# VSS 0.63fF
C11906 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A VSS 0.92fF
C11907 a_3373_n10301# VSS 0.34fF
C11908 a_3266_n10301# VSS 0.45fF
C11909 a_3010_n10301# VSS 0.63fF
C11910 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS 0.92fF
C11911 a_2085_n10301# VSS 0.34fF
C11912 a_1978_n10301# VSS 0.45fF
C11913 a_1722_n10301# VSS 0.63fF
C11914 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A VSS 0.92fF
C11915 a_797_n10301# VSS 0.34fF
C11916 a_690_n10301# VSS 0.46fF
C11917 a_434_n10301# VSS 0.63fF
C11918 p2d VSS 3.33fF
C11919 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS 0.61fF
C11920 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VSS 1.80fF
C11921 a_13765_n9757# VSS 2.05fF
C11922 a_11164_n9783# VSS 0.57fF
C11923 a_10904_n9783# VSS 0.39fF
C11924 a_10805_n9525# VSS 0.34fF
C11925 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS 0.86fF
C11926 a_9876_n9783# VSS 0.62fF
C11927 a_9616_n9783# VSS 0.42fF
C11928 a_9517_n9525# VSS 0.35fF
C11929 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS 0.82fF
C11930 a_8588_n9783# VSS 0.64fF
C11931 a_8328_n9783# VSS 0.43fF
C11932 a_8229_n9525# VSS 0.36fF
C11933 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS 0.83fF
C11934 a_7300_n9783# VSS 0.64fF
C11935 a_7040_n9783# VSS 0.43fF
C11936 a_6941_n9525# VSS 0.36fF
C11937 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS 0.84fF
C11938 a_6012_n9783# VSS 0.64fF
C11939 a_5752_n9783# VSS 0.43fF
C11940 a_5653_n9525# VSS 0.36fF
C11941 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS 0.84fF
C11942 a_4724_n9783# VSS 0.64fF
C11943 a_4464_n9783# VSS 0.43fF
C11944 a_4365_n9525# VSS 0.36fF
C11945 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS 0.84fF
C11946 a_3436_n9783# VSS 0.64fF
C11947 a_3176_n9783# VSS 0.43fF
C11948 a_3077_n9525# VSS 0.36fF
C11949 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS 0.84fF
C11950 a_2148_n9783# VSS 0.64fF
C11951 a_1888_n9783# VSS 0.43fF
C11952 a_1789_n9525# VSS 0.36fF
C11953 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS 0.84fF
C11954 a_860_n9783# VSS 0.64fF
C11955 a_600_n9783# VSS 0.43fF
C11956 a_501_n9525# VSS 0.36fF
C11957 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS 1.11fF
C11958 a_n428_n9783# VSS 0.69fF
C11959 a_n688_n9783# VSS 0.47fF
C11960 a_n787_n9525# VSS 0.38fF
C11961 p2_b VSS 3.22fF
C11962 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS 0.69fF
C11963 a_13765_n9213# VSS 2.32fF
C11964 sky130_fd_sc_hd__clkinv_4_10/Y VSS 2.03fF
C11965 a_11101_n9213# VSS 0.33fF
C11966 a_10994_n9213# VSS 0.44fF
C11967 a_10738_n9213# VSS 0.62fF
C11968 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS 0.89fF
C11969 a_9813_n9213# VSS 0.33fF
C11970 a_9706_n9213# VSS 0.44fF
C11971 a_9450_n9213# VSS 0.63fF
C11972 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A VSS 0.89fF
C11973 a_8525_n9213# VSS 0.34fF
C11974 a_8418_n9213# VSS 0.45fF
C11975 a_8162_n9213# VSS 0.63fF
C11976 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS 0.90fF
C11977 a_7237_n9213# VSS 0.34fF
C11978 a_7130_n9213# VSS 0.45fF
C11979 a_6874_n9213# VSS 0.63fF
C11980 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A VSS 0.91fF
C11981 a_5949_n9213# VSS 0.34fF
C11982 a_5842_n9213# VSS 0.45fF
C11983 a_5586_n9213# VSS 0.63fF
C11984 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS 0.91fF
C11985 a_4661_n9213# VSS 0.34fF
C11986 a_4554_n9213# VSS 0.45fF
C11987 a_4298_n9213# VSS 0.63fF
C11988 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A VSS 0.91fF
C11989 a_3373_n9213# VSS 0.34fF
C11990 a_3266_n9213# VSS 0.45fF
C11991 a_3010_n9213# VSS 0.63fF
C11992 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS 0.91fF
C11993 a_2085_n9213# VSS 0.34fF
C11994 a_1978_n9213# VSS 0.45fF
C11995 a_1722_n9213# VSS 0.64fF
C11996 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A VSS 0.91fF
C11997 a_797_n9213# VSS 0.35fF
C11998 a_690_n9213# VSS 0.46fF
C11999 a_434_n9213# VSS 0.64fF
C12000 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS 0.62fF
C12001 a_13765_n8669# VSS 2.08fF
C12002 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS 2.89fF
C12003 a_11164_n8695# VSS 0.57fF
C12004 a_10904_n8695# VSS 0.39fF
C12005 a_10805_n8437# VSS 0.34fF
C12006 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS 0.92fF
C12007 a_9876_n8695# VSS 0.62fF
C12008 a_9616_n8695# VSS 0.42fF
C12009 a_9517_n8437# VSS 0.35fF
C12010 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS 0.89fF
C12011 a_8588_n8695# VSS 0.64fF
C12012 a_8328_n8695# VSS 0.43fF
C12013 a_8229_n8437# VSS 0.36fF
C12014 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS 0.89fF
C12015 a_7300_n8695# VSS 0.64fF
C12016 a_7040_n8695# VSS 0.43fF
C12017 a_6941_n8437# VSS 0.36fF
C12018 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS 0.90fF
C12019 a_6012_n8695# VSS 0.66fF
C12020 a_5752_n8695# VSS 0.46fF
C12021 a_5653_n8437# VSS 0.36fF
C12022 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS 0.89fF
C12023 a_4724_n8695# VSS 0.65fF
C12024 a_4464_n8695# VSS 0.42fF
C12025 a_4365_n8437# VSS 0.36fF
C12026 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS 0.90fF
C12027 a_3436_n8695# VSS 0.65fF
C12028 a_3176_n8695# VSS 0.43fF
C12029 a_3077_n8437# VSS 0.36fF
C12030 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS 0.90fF
C12031 a_2148_n8695# VSS 0.65fF
C12032 a_1888_n8695# VSS 0.43fF
C12033 a_1789_n8437# VSS 0.36fF
C12034 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS 0.90fF
C12035 a_860_n8695# VSS 0.66fF
C12036 a_600_n8695# VSS 0.44fF
C12037 a_501_n8437# VSS 0.37fF
C12038 a_10738_n8125# VSS 1.10fF
C12039 sky130_fd_sc_hd__nand2_4_3/Y VSS 8.33fF
C12040 a_n860_n8125# VSS 0.00fF
C12041 sky130_fd_sc_hd__nand2_4_3/B VSS 1.25fF
C12042 a_9813_n8125# VSS 0.34fF
C12043 a_9706_n8125# VSS 0.45fF
C12044 a_9450_n8125# VSS 0.62fF
C12045 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS 0.96fF
C12046 a_8525_n8125# VSS 0.37fF
C12047 a_8418_n8125# VSS 0.50fF
C12048 a_8162_n8125# VSS 0.67fF
C12049 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS 0.98fF
C12050 a_7237_n8125# VSS 0.34fF
C12051 a_7130_n8125# VSS 0.44fF
C12052 a_6874_n8125# VSS 0.61fF
C12053 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS 2.83fF
C12054 a_2729_n8125# VSS 0.35fF
C12055 a_2622_n8125# VSS 0.46fF
C12056 a_2366_n8125# VSS 0.64fF
C12057 sky130_fd_sc_hd__clkinv_1_3/Y VSS 1.28fF
C12058 sky130_fd_sc_hd__clkinv_1_3/A VSS 13.93fF
C12059 sky130_fd_sc_hd__nand2_4_3/A VSS 5.08fF
C12060 a_7212_n7203# VSS 0.14fF
C12061 a_7014_n7215# VSS 0.01fF
C12062 a_6593_n7215# VSS 0.01fF
C12063 sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS 0.31fF
C12064 a_4986_n7215# VSS 0.01fF
C12065 a_4765_n7215# VSS 0.01fF
C12066 a_3832_n7261# VSS 0.01fF
C12067 sky130_fd_sc_hd__clkinv_1_4/Y VSS 1.60fF
C12068 p2 VSS 9.17fF
C12069 a_6794_n7203# VSS 0.39fF
C12070 a_6865_n7304# VSS 0.32fF
C12071 a_6665_n7459# VSS 0.61fF
C12072 a_6658_n7363# VSS 0.82fF
C12073 a_6373_n7349# VSS 0.39fF
C12074 a_6101_n7254# VSS 0.65fF
C12075 a_6006_n7607# VSS 0.31fF
C12076 a_5052_n7283# VSS 0.50fF
C12077 sky130_fd_sc_hd__dfxbp_1_0/Q VSS 1.48fF
C12078 a_4623_n7349# VSS 0.54fF
C12079 sky130_fd_sc_hd__mux2_1_0/X VSS 0.76fF
C12080 sky130_fd_sc_hd__nand2_1_4/B VSS 6.41fF
C12081 sky130_fd_sc_hd__nand2_1_4/Y VSS 1.85fF
C12082 a_n1612_n7037# VSS 0.00fF
C12083 a_n2037_n7037# VSS 0.00fF
C12084 a_n2248_n7037# VSS 0.14fF
C12085 a_n1139_n6715# VSS 0.29fF
C12086 a_n1738_n6671# VSS 0.41fF
C12087 a_n1570_n6769# VSS 0.64fF
C12088 a_n2163_n6671# VSS 0.32fF
C12089 a_n1995_n6925# VSS 0.36fF
C12090 a_n2436_n7037# VSS 0.60fF
C12091 sky130_fd_sc_hd__dfxbp_1_1/D VSS 1.16fF
C12092 a_n2602_n7037# VSS 0.85fF
C12093 clk VSS 3.84fF
C12094 a_10738_n6173# VSS 1.19fF
C12095 a_n860_n6173# VSS 0.01fF
C12096 sky130_fd_sc_hd__nand2_4_1/B VSS 1.19fF
C12097 a_9813_n6493# VSS 0.34fF
C12098 a_9706_n6493# VSS 0.44fF
C12099 a_9450_n6493# VSS 0.62fF
C12100 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS 0.90fF
C12101 a_8525_n6493# VSS 0.37fF
C12102 a_8418_n6493# VSS 0.48fF
C12103 a_8162_n6493# VSS 0.67fF
C12104 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS 0.91fF
C12105 a_7237_n6493# VSS 0.36fF
C12106 a_7130_n6493# VSS 0.48fF
C12107 a_6874_n6493# VSS 0.66fF
C12108 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS 2.46fF
C12109 a_2729_n6493# VSS 0.37fF
C12110 a_2622_n6493# VSS 0.48fF
C12111 a_2366_n6493# VSS 0.67fF
C12112 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A VSS 1.20fF
C12113 sky130_fd_sc_hd__nand2_4_1/A VSS 5.01fF
C12114 A VSS 3.15fF
C12115 a_13765_n5949# VSS 2.10fF
C12116 a_11164_n5975# VSS 0.54fF
C12117 a_10904_n5975# VSS 0.37fF
C12118 a_10805_n5797# VSS 0.32fF
C12119 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS 0.93fF
C12120 a_9876_n5975# VSS 0.60fF
C12121 a_9616_n5975# VSS 0.41fF
C12122 a_9517_n5797# VSS 0.34fF
C12123 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS 0.90fF
C12124 a_8588_n5975# VSS 0.65fF
C12125 a_8328_n5975# VSS 0.44fF
C12126 a_8229_n5797# VSS 0.36fF
C12127 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS 0.91fF
C12128 a_7300_n5975# VSS 0.65fF
C12129 a_7040_n5975# VSS 0.44fF
C12130 a_6941_n5797# VSS 0.35fF
C12131 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS 0.91fF
C12132 a_6012_n5975# VSS 0.64fF
C12133 a_5752_n5975# VSS 0.44fF
C12134 a_5653_n5797# VSS 0.36fF
C12135 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS 0.91fF
C12136 a_4724_n5975# VSS 0.65fF
C12137 a_4464_n5975# VSS 0.43fF
C12138 a_4365_n5797# VSS 0.36fF
C12139 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS 0.91fF
C12140 a_3436_n5975# VSS 0.65fF
C12141 a_3176_n5975# VSS 0.45fF
C12142 a_3077_n5797# VSS 0.35fF
C12143 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS 0.91fF
C12144 a_2148_n5975# VSS 0.64fF
C12145 a_1888_n5975# VSS 0.45fF
C12146 a_1789_n5797# VSS 0.36fF
C12147 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS 0.91fF
C12148 a_860_n5975# VSS 0.65fF
C12149 a_600_n5975# VSS 0.43fF
C12150 a_501_n5797# VSS 0.37fF
C12151 A_b VSS 3.36fF
C12152 a_13765_n5405# VSS 2.12fF
C12153 sky130_fd_sc_hd__clkinv_4_4/Y VSS 1.92fF
C12154 sky130_fd_sc_hd__clkinv_4_4/A VSS 13.93fF
C12155 a_11101_n5405# VSS 0.33fF
C12156 a_10994_n5405# VSS 0.43fF
C12157 a_10738_n5405# VSS 0.61fF
C12158 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS 0.91fF
C12159 a_9813_n5405# VSS 0.33fF
C12160 a_9706_n5405# VSS 0.43fF
C12161 a_9450_n5405# VSS 0.62fF
C12162 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A VSS 0.91fF
C12163 a_8525_n5405# VSS 0.34fF
C12164 a_8418_n5405# VSS 0.44fF
C12165 a_8162_n5405# VSS 0.63fF
C12166 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS 0.91fF
C12167 a_7237_n5405# VSS 0.34fF
C12168 a_7130_n5405# VSS 0.44fF
C12169 a_6874_n5405# VSS 0.63fF
C12170 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A VSS 0.91fF
C12171 a_5949_n5405# VSS 0.34fF
C12172 a_5842_n5405# VSS 0.44fF
C12173 a_5586_n5405# VSS 0.63fF
C12174 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS 0.91fF
C12175 a_4661_n5405# VSS 0.34fF
C12176 a_4554_n5405# VSS 0.44fF
C12177 a_4298_n5405# VSS 0.63fF
C12178 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A VSS 0.92fF
C12179 a_3373_n5405# VSS 0.34fF
C12180 a_3266_n5405# VSS 0.44fF
C12181 a_3010_n5405# VSS 0.63fF
C12182 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS 0.91fF
C12183 a_2085_n5405# VSS 0.34fF
C12184 a_1978_n5405# VSS 0.44fF
C12185 a_1722_n5405# VSS 0.63fF
C12186 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A VSS 0.92fF
C12187 a_797_n5405# VSS 0.35fF
C12188 a_690_n5405# VSS 0.45fF
C12189 a_434_n5405# VSS 0.64fF
C12190 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A VSS 0.60fF
C12191 Ad VSS 3.18fF
C12192 a_13765_n4861# VSS 2.24fF
C12193 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A VSS 0.71fF
C12194 a_11164_n4887# VSS 0.57fF
C12195 a_10904_n4887# VSS 0.41fF
C12196 a_10805_n4709# VSS 0.34fF
C12197 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS 0.91fF
C12198 a_9876_n4887# VSS 0.62fF
C12199 a_9616_n4887# VSS 0.43fF
C12200 a_9517_n4709# VSS 0.35fF
C12201 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS 0.88fF
C12202 a_8588_n4887# VSS 0.64fF
C12203 a_8328_n4887# VSS 0.44fF
C12204 a_8229_n4709# VSS 0.35fF
C12205 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS 0.88fF
C12206 a_7300_n4887# VSS 0.64fF
C12207 a_7040_n4887# VSS 0.44fF
C12208 a_6941_n4709# VSS 0.35fF
C12209 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS 0.88fF
C12210 a_6012_n4887# VSS 0.63fF
C12211 a_5752_n4887# VSS 0.43fF
C12212 a_5653_n4709# VSS 0.35fF
C12213 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS 0.89fF
C12214 a_4724_n4887# VSS 0.64fF
C12215 a_4464_n4887# VSS 0.44fF
C12216 a_4365_n4709# VSS 0.35fF
C12217 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS 0.88fF
C12218 a_3436_n4887# VSS 0.64fF
C12219 a_3176_n4887# VSS 0.44fF
C12220 a_3077_n4709# VSS 0.35fF
C12221 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS 0.88fF
C12222 a_2148_n4887# VSS 0.64fF
C12223 a_1888_n4887# VSS 0.44fF
C12224 a_1789_n4709# VSS 0.35fF
C12225 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS 0.89fF
C12226 a_860_n4887# VSS 0.64fF
C12227 a_600_n4887# VSS 0.44fF
C12228 a_501_n4709# VSS 0.35fF
C12229 a_n428_n4887# VSS 0.70fF
C12230 a_n688_n4887# VSS 0.48fF
C12231 a_n787_n4709# VSS 0.38fF
C12232 Ad_b VSS 16.44fF
C12233 a_13765_n4317# VSS 2.19fF
C12234 sky130_fd_sc_hd__clkinv_4_3/Y VSS 2.74fF
C12235 sky130_fd_sc_hd__clkinv_4_3/A VSS 8.56fF
C12236 a_11101_n4317# VSS 0.33fF
C12237 a_10994_n4317# VSS 0.43fF
C12238 a_10738_n4317# VSS 0.61fF
C12239 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS 0.92fF
C12240 a_9813_n4317# VSS 0.33fF
C12241 a_9706_n4317# VSS 0.43fF
C12242 a_9450_n4317# VSS 0.62fF
C12243 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A VSS 0.91fF
C12244 a_8525_n4317# VSS 0.34fF
C12245 a_8418_n4317# VSS 0.44fF
C12246 a_8162_n4317# VSS 0.63fF
C12247 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS 0.92fF
C12248 a_7237_n4317# VSS 0.34fF
C12249 a_7130_n4317# VSS 0.44fF
C12250 a_6874_n4317# VSS 0.63fF
C12251 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A VSS 0.92fF
C12252 a_5949_n4317# VSS 0.34fF
C12253 a_5842_n4317# VSS 0.44fF
C12254 a_5586_n4317# VSS 0.63fF
C12255 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS 0.92fF
C12256 a_4661_n4317# VSS 0.34fF
C12257 a_4554_n4317# VSS 0.44fF
C12258 a_4298_n4317# VSS 0.63fF
C12259 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A VSS 0.92fF
C12260 a_3373_n4317# VSS 0.34fF
C12261 a_3266_n4317# VSS 0.44fF
C12262 a_3010_n4317# VSS 0.63fF
C12263 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS 0.92fF
C12264 a_2085_n4317# VSS 0.34fF
C12265 a_1978_n4317# VSS 0.44fF
C12266 a_1722_n4317# VSS 0.63fF
C12267 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A VSS 0.92fF
C12268 a_797_n4317# VSS 0.35fF
C12269 a_690_n4317# VSS 0.44fF
C12270 a_434_n4317# VSS 0.63fF
C12271 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A VSS 0.60fF
C12272 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VSS 1.23fF
C12273 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A VSS 0.66fF
C12274 a_11164_n3799# VSS 0.57fF
C12275 a_10904_n3799# VSS 0.40fF
C12276 a_10805_n3621# VSS 0.34fF
C12277 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS 0.93fF
C12278 a_9876_n3799# VSS 0.62fF
C12279 a_9616_n3799# VSS 0.43fF
C12280 a_9517_n3621# VSS 0.35fF
C12281 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS 0.90fF
C12282 a_8588_n3799# VSS 0.64fF
C12283 a_8328_n3799# VSS 0.44fF
C12284 a_8229_n3621# VSS 0.36fF
C12285 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS 0.90fF
C12286 a_7300_n3799# VSS 0.64fF
C12287 a_7040_n3799# VSS 0.44fF
C12288 a_6941_n3621# VSS 0.36fF
C12289 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS 0.90fF
C12290 a_6012_n3799# VSS 0.64fF
C12291 a_5752_n3799# VSS 0.44fF
C12292 a_5653_n3621# VSS 0.36fF
C12293 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS 0.90fF
C12294 a_4724_n3799# VSS 0.64fF
C12295 a_4464_n3799# VSS 0.44fF
C12296 a_4365_n3621# VSS 0.36fF
C12297 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS 0.90fF
C12298 a_3436_n3799# VSS 0.64fF
C12299 a_3176_n3799# VSS 0.44fF
C12300 a_3077_n3621# VSS 0.36fF
C12301 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS 0.90fF
C12302 a_2148_n3799# VSS 0.64fF
C12303 a_1888_n3799# VSS 0.44fF
C12304 a_1789_n3621# VSS 0.36fF
C12305 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS 0.92fF
C12306 a_860_n3799# VSS 0.65fF
C12307 a_600_n3799# VSS 0.44fF
C12308 a_501_n3621# VSS 0.36fF
C12309 a_11164_n3255# VSS 0.56fF
C12310 a_10904_n3255# VSS 0.39fF
C12311 a_10805_n2997# VSS 0.34fF
C12312 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS 0.88fF
C12313 a_9876_n3255# VSS 0.62fF
C12314 a_9616_n3255# VSS 0.41fF
C12315 a_9517_n2997# VSS 0.35fF
C12316 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS 0.90fF
C12317 a_8588_n3255# VSS 0.64fF
C12318 a_8328_n3255# VSS 0.42fF
C12319 a_8229_n2997# VSS 0.36fF
C12320 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS 0.90fF
C12321 a_7300_n3255# VSS 0.64fF
C12322 a_7040_n3255# VSS 0.42fF
C12323 a_6941_n2997# VSS 0.36fF
C12324 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS 0.90fF
C12325 a_6012_n3255# VSS 0.64fF
C12326 a_5752_n3255# VSS 0.42fF
C12327 a_5653_n2997# VSS 0.36fF
C12328 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS 0.90fF
C12329 a_4724_n3255# VSS 0.64fF
C12330 a_4464_n3255# VSS 0.42fF
C12331 a_4365_n2997# VSS 0.36fF
C12332 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS 0.90fF
C12333 a_3436_n3255# VSS 0.64fF
C12334 a_3176_n3255# VSS 0.42fF
C12335 a_3077_n2997# VSS 0.36fF
C12336 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VSS 0.90fF
C12337 a_2148_n3255# VSS 0.64fF
C12338 a_1888_n3255# VSS 0.42fF
C12339 a_1789_n2997# VSS 0.36fF
C12340 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS 0.85fF
C12341 a_860_n3255# VSS 0.64fF
C12342 a_600_n3255# VSS 0.43fF
C12343 a_501_n2997# VSS 0.37fF
C12344 sky130_fd_sc_hd__clkinv_1_5/A VSS 5.66fF
C12345 Bd_b VSS 9.24fF
C12346 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X VSS 0.71fF
C12347 a_13765_n2685# VSS 2.38fF
C12348 a_11101_n2685# VSS 0.33fF
C12349 a_10994_n2685# VSS 0.44fF
C12350 a_10738_n2685# VSS 0.62fF
C12351 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS 0.92fF
C12352 a_9813_n2685# VSS 0.33fF
C12353 a_9706_n2685# VSS 0.45fF
C12354 a_9450_n2685# VSS 0.63fF
C12355 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A VSS 0.92fF
C12356 a_8525_n2685# VSS 0.34fF
C12357 a_8418_n2685# VSS 0.45fF
C12358 a_8162_n2685# VSS 0.63fF
C12359 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS 0.92fF
C12360 a_7237_n2685# VSS 0.34fF
C12361 a_7130_n2685# VSS 0.45fF
C12362 a_6874_n2685# VSS 0.63fF
C12363 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A VSS 0.92fF
C12364 a_5949_n2685# VSS 0.34fF
C12365 a_5842_n2685# VSS 0.45fF
C12366 a_5586_n2685# VSS 0.63fF
C12367 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS 0.92fF
C12368 a_4661_n2685# VSS 0.34fF
C12369 a_4554_n2685# VSS 0.45fF
C12370 a_4298_n2685# VSS 0.63fF
C12371 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A VSS 0.92fF
C12372 a_3373_n2685# VSS 0.34fF
C12373 a_3266_n2685# VSS 0.45fF
C12374 a_3010_n2685# VSS 0.63fF
C12375 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A VSS 0.92fF
C12376 a_2085_n2685# VSS 0.34fF
C12377 a_1978_n2685# VSS 0.45fF
C12378 a_1722_n2685# VSS 0.63fF
C12379 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A VSS 0.92fF
C12380 a_797_n2685# VSS 0.34fF
C12381 a_690_n2685# VSS 0.46fF
C12382 a_434_n2685# VSS 0.63fF
C12383 Bd VSS 3.33fF
C12384 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS 0.61fF
C12385 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VSS 1.63fF
C12386 a_13765_n2141# VSS 2.05fF
C12387 a_11164_n2167# VSS 0.57fF
C12388 a_10904_n2167# VSS 0.39fF
C12389 a_10805_n1909# VSS 0.34fF
C12390 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS 0.86fF
C12391 a_9876_n2167# VSS 0.62fF
C12392 a_9616_n2167# VSS 0.42fF
C12393 a_9517_n1909# VSS 0.35fF
C12394 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS 0.82fF
C12395 a_8588_n2167# VSS 0.64fF
C12396 a_8328_n2167# VSS 0.43fF
C12397 a_8229_n1909# VSS 0.36fF
C12398 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS 0.83fF
C12399 a_7300_n2167# VSS 0.64fF
C12400 a_7040_n2167# VSS 0.43fF
C12401 a_6941_n1909# VSS 0.36fF
C12402 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS 0.84fF
C12403 a_6012_n2167# VSS 0.64fF
C12404 a_5752_n2167# VSS 0.43fF
C12405 a_5653_n1909# VSS 0.36fF
C12406 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS 0.84fF
C12407 a_4724_n2167# VSS 0.64fF
C12408 a_4464_n2167# VSS 0.43fF
C12409 a_4365_n1909# VSS 0.36fF
C12410 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS 0.84fF
C12411 a_3436_n2167# VSS 0.64fF
C12412 a_3176_n2167# VSS 0.43fF
C12413 a_3077_n1909# VSS 0.36fF
C12414 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VSS 0.84fF
C12415 a_2148_n2167# VSS 0.64fF
C12416 a_1888_n2167# VSS 0.43fF
C12417 a_1789_n1909# VSS 0.36fF
C12418 sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VSS 0.84fF
C12419 a_860_n2167# VSS 0.64fF
C12420 a_600_n2167# VSS 0.43fF
C12421 a_501_n1909# VSS 0.36fF
C12422 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS 1.15fF
C12423 a_n428_n2167# VSS 0.69fF
C12424 a_n688_n2167# VSS 0.47fF
C12425 a_n787_n1909# VSS 0.38fF
C12426 B_b VSS 3.22fF
C12427 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS 0.69fF
C12428 a_13765_n1597# VSS 2.32fF
C12429 sky130_fd_sc_hd__clkinv_4_1/Y VSS 2.03fF
C12430 a_11101_n1597# VSS 0.33fF
C12431 a_10994_n1597# VSS 0.44fF
C12432 a_10738_n1597# VSS 0.62fF
C12433 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS 0.89fF
C12434 a_9813_n1597# VSS 0.33fF
C12435 a_9706_n1597# VSS 0.44fF
C12436 a_9450_n1597# VSS 0.63fF
C12437 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A VSS 0.89fF
C12438 a_8525_n1597# VSS 0.34fF
C12439 a_8418_n1597# VSS 0.45fF
C12440 a_8162_n1597# VSS 0.63fF
C12441 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS 0.90fF
C12442 a_7237_n1597# VSS 0.34fF
C12443 a_7130_n1597# VSS 0.45fF
C12444 a_6874_n1597# VSS 0.63fF
C12445 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A VSS 0.91fF
C12446 a_5949_n1597# VSS 0.34fF
C12447 a_5842_n1597# VSS 0.45fF
C12448 a_5586_n1597# VSS 0.63fF
C12449 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS 0.91fF
C12450 a_4661_n1597# VSS 0.34fF
C12451 a_4554_n1597# VSS 0.45fF
C12452 a_4298_n1597# VSS 0.63fF
C12453 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A VSS 0.91fF
C12454 a_3373_n1597# VSS 0.34fF
C12455 a_3266_n1597# VSS 0.45fF
C12456 a_3010_n1597# VSS 0.63fF
C12457 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A VSS 0.91fF
C12458 a_2085_n1597# VSS 0.34fF
C12459 a_1978_n1597# VSS 0.45fF
C12460 a_1722_n1597# VSS 0.63fF
C12461 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A VSS 0.91fF
C12462 a_797_n1597# VSS 0.34fF
C12463 a_690_n1597# VSS 0.45fF
C12464 a_434_n1597# VSS 0.63fF
C12465 B VSS 3.21fF
C12466 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X VSS 0.62fF
C12467 a_13765_n1053# VSS 2.05fF
C12468 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS 2.86fF
C12469 a_11164_n1079# VSS 0.56fF
C12470 a_10904_n1079# VSS 0.39fF
C12471 a_10805_n821# VSS 0.33fF
C12472 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS 0.89fF
C12473 a_9876_n1079# VSS 0.61fF
C12474 a_9616_n1079# VSS 0.42fF
C12475 a_9517_n821# VSS 0.35fF
C12476 sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VSS 0.86fF
C12477 a_8588_n1079# VSS 0.63fF
C12478 a_8328_n1079# VSS 0.42fF
C12479 a_8229_n821# VSS 0.35fF
C12480 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS 0.87fF
C12481 a_7300_n1079# VSS 0.63fF
C12482 a_7040_n1079# VSS 0.42fF
C12483 a_6941_n821# VSS 0.35fF
C12484 sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VSS 0.88fF
C12485 a_6012_n1079# VSS 0.67fF
C12486 a_5752_n1079# VSS 0.46fF
C12487 a_5653_n821# VSS 0.36fF
C12488 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS 0.86fF
C12489 a_4724_n1079# VSS 0.64fF
C12490 a_4464_n1079# VSS 0.42fF
C12491 a_4365_n821# VSS 0.36fF
C12492 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VSS 0.88fF
C12493 a_3436_n1079# VSS 0.64fF
C12494 a_3176_n1079# VSS 0.42fF
C12495 a_3077_n821# VSS 0.36fF
C12496 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VSS 0.87fF
C12497 a_2148_n1079# VSS 0.64fF
C12498 a_1888_n1079# VSS 0.42fF
C12499 a_1789_n821# VSS 0.36fF
C12500 sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VSS 0.87fF
C12501 a_860_n1079# VSS 0.64fF
C12502 a_600_n1079# VSS 0.43fF
C12503 a_501_n821# VSS 0.37fF
C12504 a_10738_n509# VSS 1.08fF
C12505 sky130_fd_sc_hd__nand2_4_0/Y VSS 8.30fF
C12506 a_n860_n509# VSS 0.00fF
C12507 sky130_fd_sc_hd__nand2_4_0/B VSS 1.19fF
C12508 a_9813_n509# VSS 0.33fF
C12509 a_9706_n509# VSS 0.45fF
C12510 a_9450_n509# VSS 0.61fF
C12511 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS 0.91fF
C12512 a_8525_n509# VSS 0.33fF
C12513 a_8418_n509# VSS 0.45fF
C12514 a_8162_n509# VSS 0.61fF
C12515 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS 0.92fF
C12516 a_7237_n509# VSS 0.33fF
C12517 a_7130_n509# VSS 0.44fF
C12518 a_6874_n509# VSS 0.60fF
C12519 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS 2.63fF
C12520 a_2729_n509# VSS 0.34fF
C12521 a_2622_n509# VSS 0.46fF
C12522 a_2366_n509# VSS 0.61fF
C12523 sky130_fd_sc_hd__clkinv_1_0/Y VSS 1.19fF
C12524 sky130_fd_sc_hd__clkinv_1_0/A VSS 13.40fF
C12525 sky130_fd_sc_hd__nand2_4_0/A VSS 4.31fF
C12526 sky130_fd_sc_hd__nand2_1_0/A VSS 1.38fF
C12527 sky130_fd_sc_hd__nand2_1_0/B VSS 1.68fF
C12528 VDD VSS 1347.57fF
.ends

