magic
tech sky130A
magscale 1 2
timestamp 1654656593
<< nmos >>
rect -2374 -140 -2254 140
rect -2196 -140 -2076 140
rect -2018 -140 -1898 140
rect -1840 -140 -1720 140
rect -1662 -140 -1542 140
rect -1484 -140 -1364 140
rect -1306 -140 -1186 140
rect -1128 -140 -1008 140
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
rect 1008 -140 1128 140
rect 1186 -140 1306 140
rect 1364 -140 1484 140
rect 1542 -140 1662 140
rect 1720 -140 1840 140
rect 1898 -140 2018 140
rect 2076 -140 2196 140
rect 2254 -140 2374 140
<< ndiff >>
rect -2432 128 -2374 140
rect -2432 -128 -2420 128
rect -2386 -128 -2374 128
rect -2432 -140 -2374 -128
rect -2254 128 -2196 140
rect -2254 -128 -2242 128
rect -2208 -128 -2196 128
rect -2254 -140 -2196 -128
rect -2076 128 -2018 140
rect -2076 -128 -2064 128
rect -2030 -128 -2018 128
rect -2076 -140 -2018 -128
rect -1898 128 -1840 140
rect -1898 -128 -1886 128
rect -1852 -128 -1840 128
rect -1898 -140 -1840 -128
rect -1720 128 -1662 140
rect -1720 -128 -1708 128
rect -1674 -128 -1662 128
rect -1720 -140 -1662 -128
rect -1542 128 -1484 140
rect -1542 -128 -1530 128
rect -1496 -128 -1484 128
rect -1542 -140 -1484 -128
rect -1364 128 -1306 140
rect -1364 -128 -1352 128
rect -1318 -128 -1306 128
rect -1364 -140 -1306 -128
rect -1186 128 -1128 140
rect -1186 -128 -1174 128
rect -1140 -128 -1128 128
rect -1186 -140 -1128 -128
rect -1008 128 -950 140
rect -1008 -128 -996 128
rect -962 -128 -950 128
rect -1008 -140 -950 -128
rect -830 128 -772 140
rect -830 -128 -818 128
rect -784 -128 -772 128
rect -830 -140 -772 -128
rect -652 128 -594 140
rect -652 -128 -640 128
rect -606 -128 -594 128
rect -652 -140 -594 -128
rect -474 128 -416 140
rect -474 -128 -462 128
rect -428 -128 -416 128
rect -474 -140 -416 -128
rect -296 128 -238 140
rect -296 -128 -284 128
rect -250 -128 -238 128
rect -296 -140 -238 -128
rect -118 128 -60 140
rect -118 -128 -106 128
rect -72 -128 -60 128
rect -118 -140 -60 -128
rect 60 128 118 140
rect 60 -128 72 128
rect 106 -128 118 128
rect 60 -140 118 -128
rect 238 128 296 140
rect 238 -128 250 128
rect 284 -128 296 128
rect 238 -140 296 -128
rect 416 128 474 140
rect 416 -128 428 128
rect 462 -128 474 128
rect 416 -140 474 -128
rect 594 128 652 140
rect 594 -128 606 128
rect 640 -128 652 128
rect 594 -140 652 -128
rect 772 128 830 140
rect 772 -128 784 128
rect 818 -128 830 128
rect 772 -140 830 -128
rect 950 128 1008 140
rect 950 -128 962 128
rect 996 -128 1008 128
rect 950 -140 1008 -128
rect 1128 128 1186 140
rect 1128 -128 1140 128
rect 1174 -128 1186 128
rect 1128 -140 1186 -128
rect 1306 128 1364 140
rect 1306 -128 1318 128
rect 1352 -128 1364 128
rect 1306 -140 1364 -128
rect 1484 128 1542 140
rect 1484 -128 1496 128
rect 1530 -128 1542 128
rect 1484 -140 1542 -128
rect 1662 128 1720 140
rect 1662 -128 1674 128
rect 1708 -128 1720 128
rect 1662 -140 1720 -128
rect 1840 128 1898 140
rect 1840 -128 1852 128
rect 1886 -128 1898 128
rect 1840 -140 1898 -128
rect 2018 128 2076 140
rect 2018 -128 2030 128
rect 2064 -128 2076 128
rect 2018 -140 2076 -128
rect 2196 128 2254 140
rect 2196 -128 2208 128
rect 2242 -128 2254 128
rect 2196 -140 2254 -128
rect 2374 128 2432 140
rect 2374 -128 2386 128
rect 2420 -128 2432 128
rect 2374 -140 2432 -128
<< ndiffc >>
rect -2420 -128 -2386 128
rect -2242 -128 -2208 128
rect -2064 -128 -2030 128
rect -1886 -128 -1852 128
rect -1708 -128 -1674 128
rect -1530 -128 -1496 128
rect -1352 -128 -1318 128
rect -1174 -128 -1140 128
rect -996 -128 -962 128
rect -818 -128 -784 128
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect 784 -128 818 128
rect 962 -128 996 128
rect 1140 -128 1174 128
rect 1318 -128 1352 128
rect 1496 -128 1530 128
rect 1674 -128 1708 128
rect 1852 -128 1886 128
rect 2030 -128 2064 128
rect 2208 -128 2242 128
rect 2386 -128 2420 128
<< poly >>
rect -2356 212 -2272 228
rect -2356 195 -2340 212
rect -2374 178 -2340 195
rect -2288 195 -2272 212
rect -2178 212 -2094 228
rect -2178 195 -2162 212
rect -2288 178 -2254 195
rect -2374 140 -2254 178
rect -2196 178 -2162 195
rect -2110 195 -2094 212
rect -2000 212 -1916 228
rect -2000 195 -1984 212
rect -2110 178 -2076 195
rect -2196 140 -2076 178
rect -2018 178 -1984 195
rect -1932 195 -1916 212
rect -1822 212 -1738 228
rect -1822 195 -1806 212
rect -1932 178 -1898 195
rect -2018 140 -1898 178
rect -1840 178 -1806 195
rect -1754 195 -1738 212
rect -1644 212 -1560 228
rect -1644 195 -1628 212
rect -1754 178 -1720 195
rect -1840 140 -1720 178
rect -1662 178 -1628 195
rect -1576 195 -1560 212
rect -1466 212 -1382 228
rect -1466 195 -1450 212
rect -1576 178 -1542 195
rect -1662 140 -1542 178
rect -1484 178 -1450 195
rect -1398 195 -1382 212
rect -1288 212 -1204 228
rect -1288 195 -1272 212
rect -1398 178 -1364 195
rect -1484 140 -1364 178
rect -1306 178 -1272 195
rect -1220 195 -1204 212
rect -1110 212 -1026 228
rect -1110 195 -1094 212
rect -1220 178 -1186 195
rect -1306 140 -1186 178
rect -1128 178 -1094 195
rect -1042 195 -1026 212
rect -932 212 -848 228
rect -932 195 -916 212
rect -1042 178 -1008 195
rect -1128 140 -1008 178
rect -950 178 -916 195
rect -864 195 -848 212
rect -754 212 -670 228
rect -754 195 -738 212
rect -864 178 -830 195
rect -950 140 -830 178
rect -772 178 -738 195
rect -686 195 -670 212
rect -576 212 -492 228
rect -576 195 -560 212
rect -686 178 -652 195
rect -772 140 -652 178
rect -594 178 -560 195
rect -508 195 -492 212
rect -398 212 -314 228
rect -398 195 -382 212
rect -508 178 -474 195
rect -594 140 -474 178
rect -416 178 -382 195
rect -330 195 -314 212
rect -220 212 -136 228
rect -220 195 -204 212
rect -330 178 -296 195
rect -416 140 -296 178
rect -238 178 -204 195
rect -152 195 -136 212
rect -42 212 42 228
rect -42 195 -26 212
rect -152 178 -118 195
rect -238 140 -118 178
rect -60 178 -26 195
rect 26 195 42 212
rect 136 212 220 228
rect 136 195 152 212
rect 26 178 60 195
rect -60 140 60 178
rect 118 178 152 195
rect 204 195 220 212
rect 314 212 398 228
rect 314 195 330 212
rect 204 178 238 195
rect 118 140 238 178
rect 296 178 330 195
rect 382 195 398 212
rect 492 212 576 228
rect 492 195 508 212
rect 382 178 416 195
rect 296 140 416 178
rect 474 178 508 195
rect 560 195 576 212
rect 670 212 754 228
rect 670 195 686 212
rect 560 178 594 195
rect 474 140 594 178
rect 652 178 686 195
rect 738 195 754 212
rect 848 212 932 228
rect 848 195 864 212
rect 738 178 772 195
rect 652 140 772 178
rect 830 178 864 195
rect 916 195 932 212
rect 1026 212 1110 228
rect 1026 195 1042 212
rect 916 178 950 195
rect 830 140 950 178
rect 1008 178 1042 195
rect 1094 195 1110 212
rect 1204 212 1288 228
rect 1204 195 1220 212
rect 1094 178 1128 195
rect 1008 140 1128 178
rect 1186 178 1220 195
rect 1272 195 1288 212
rect 1382 212 1466 228
rect 1382 195 1398 212
rect 1272 178 1306 195
rect 1186 140 1306 178
rect 1364 178 1398 195
rect 1450 195 1466 212
rect 1560 212 1644 228
rect 1560 195 1576 212
rect 1450 178 1484 195
rect 1364 140 1484 178
rect 1542 178 1576 195
rect 1628 195 1644 212
rect 1738 212 1822 228
rect 1738 195 1754 212
rect 1628 178 1662 195
rect 1542 140 1662 178
rect 1720 178 1754 195
rect 1806 195 1822 212
rect 1916 212 2000 228
rect 1916 195 1932 212
rect 1806 178 1840 195
rect 1720 140 1840 178
rect 1898 178 1932 195
rect 1984 195 2000 212
rect 2094 212 2178 228
rect 2094 195 2110 212
rect 1984 178 2018 195
rect 1898 140 2018 178
rect 2076 178 2110 195
rect 2162 195 2178 212
rect 2272 212 2356 228
rect 2272 195 2288 212
rect 2162 178 2196 195
rect 2076 140 2196 178
rect 2254 178 2288 195
rect 2340 195 2356 212
rect 2340 178 2374 195
rect 2254 140 2374 178
rect -2374 -178 -2254 -140
rect -2374 -195 -2340 -178
rect -2356 -212 -2340 -195
rect -2288 -195 -2254 -178
rect -2196 -178 -2076 -140
rect -2196 -195 -2162 -178
rect -2288 -212 -2272 -195
rect -2356 -228 -2272 -212
rect -2178 -212 -2162 -195
rect -2110 -195 -2076 -178
rect -2018 -178 -1898 -140
rect -2018 -195 -1984 -178
rect -2110 -212 -2094 -195
rect -2178 -228 -2094 -212
rect -2000 -212 -1984 -195
rect -1932 -195 -1898 -178
rect -1840 -178 -1720 -140
rect -1840 -195 -1806 -178
rect -1932 -212 -1916 -195
rect -2000 -228 -1916 -212
rect -1822 -212 -1806 -195
rect -1754 -195 -1720 -178
rect -1662 -178 -1542 -140
rect -1662 -195 -1628 -178
rect -1754 -212 -1738 -195
rect -1822 -228 -1738 -212
rect -1644 -212 -1628 -195
rect -1576 -195 -1542 -178
rect -1484 -178 -1364 -140
rect -1484 -195 -1450 -178
rect -1576 -212 -1560 -195
rect -1644 -228 -1560 -212
rect -1466 -212 -1450 -195
rect -1398 -195 -1364 -178
rect -1306 -178 -1186 -140
rect -1306 -195 -1272 -178
rect -1398 -212 -1382 -195
rect -1466 -228 -1382 -212
rect -1288 -212 -1272 -195
rect -1220 -195 -1186 -178
rect -1128 -178 -1008 -140
rect -1128 -195 -1094 -178
rect -1220 -212 -1204 -195
rect -1288 -228 -1204 -212
rect -1110 -212 -1094 -195
rect -1042 -195 -1008 -178
rect -950 -178 -830 -140
rect -950 -195 -916 -178
rect -1042 -212 -1026 -195
rect -1110 -228 -1026 -212
rect -932 -212 -916 -195
rect -864 -195 -830 -178
rect -772 -178 -652 -140
rect -772 -195 -738 -178
rect -864 -212 -848 -195
rect -932 -228 -848 -212
rect -754 -212 -738 -195
rect -686 -195 -652 -178
rect -594 -178 -474 -140
rect -594 -195 -560 -178
rect -686 -212 -670 -195
rect -754 -228 -670 -212
rect -576 -212 -560 -195
rect -508 -195 -474 -178
rect -416 -178 -296 -140
rect -416 -195 -382 -178
rect -508 -212 -492 -195
rect -576 -228 -492 -212
rect -398 -212 -382 -195
rect -330 -195 -296 -178
rect -238 -178 -118 -140
rect -238 -195 -204 -178
rect -330 -212 -314 -195
rect -398 -228 -314 -212
rect -220 -212 -204 -195
rect -152 -195 -118 -178
rect -60 -178 60 -140
rect -60 -195 -26 -178
rect -152 -212 -136 -195
rect -220 -228 -136 -212
rect -42 -212 -26 -195
rect 26 -195 60 -178
rect 118 -178 238 -140
rect 118 -195 152 -178
rect 26 -212 42 -195
rect -42 -228 42 -212
rect 136 -212 152 -195
rect 204 -195 238 -178
rect 296 -178 416 -140
rect 296 -195 330 -178
rect 204 -212 220 -195
rect 136 -228 220 -212
rect 314 -212 330 -195
rect 382 -195 416 -178
rect 474 -178 594 -140
rect 474 -195 508 -178
rect 382 -212 398 -195
rect 314 -228 398 -212
rect 492 -212 508 -195
rect 560 -195 594 -178
rect 652 -178 772 -140
rect 652 -195 686 -178
rect 560 -212 576 -195
rect 492 -228 576 -212
rect 670 -212 686 -195
rect 738 -195 772 -178
rect 830 -178 950 -140
rect 830 -195 864 -178
rect 738 -212 754 -195
rect 670 -228 754 -212
rect 848 -212 864 -195
rect 916 -195 950 -178
rect 1008 -178 1128 -140
rect 1008 -195 1042 -178
rect 916 -212 932 -195
rect 848 -228 932 -212
rect 1026 -212 1042 -195
rect 1094 -195 1128 -178
rect 1186 -178 1306 -140
rect 1186 -195 1220 -178
rect 1094 -212 1110 -195
rect 1026 -228 1110 -212
rect 1204 -212 1220 -195
rect 1272 -195 1306 -178
rect 1364 -178 1484 -140
rect 1364 -195 1398 -178
rect 1272 -212 1288 -195
rect 1204 -228 1288 -212
rect 1382 -212 1398 -195
rect 1450 -195 1484 -178
rect 1542 -178 1662 -140
rect 1542 -195 1576 -178
rect 1450 -212 1466 -195
rect 1382 -228 1466 -212
rect 1560 -212 1576 -195
rect 1628 -195 1662 -178
rect 1720 -178 1840 -140
rect 1720 -195 1754 -178
rect 1628 -212 1644 -195
rect 1560 -228 1644 -212
rect 1738 -212 1754 -195
rect 1806 -195 1840 -178
rect 1898 -178 2018 -140
rect 1898 -195 1932 -178
rect 1806 -212 1822 -195
rect 1738 -228 1822 -212
rect 1916 -212 1932 -195
rect 1984 -195 2018 -178
rect 2076 -178 2196 -140
rect 2076 -195 2110 -178
rect 1984 -212 2000 -195
rect 1916 -228 2000 -212
rect 2094 -212 2110 -195
rect 2162 -195 2196 -178
rect 2254 -178 2374 -140
rect 2254 -195 2288 -178
rect 2162 -212 2178 -195
rect 2094 -228 2178 -212
rect 2272 -212 2288 -195
rect 2340 -195 2374 -178
rect 2340 -212 2356 -195
rect 2272 -228 2356 -212
<< polycont >>
rect -2340 178 -2288 212
rect -2162 178 -2110 212
rect -1984 178 -1932 212
rect -1806 178 -1754 212
rect -1628 178 -1576 212
rect -1450 178 -1398 212
rect -1272 178 -1220 212
rect -1094 178 -1042 212
rect -916 178 -864 212
rect -738 178 -686 212
rect -560 178 -508 212
rect -382 178 -330 212
rect -204 178 -152 212
rect -26 178 26 212
rect 152 178 204 212
rect 330 178 382 212
rect 508 178 560 212
rect 686 178 738 212
rect 864 178 916 212
rect 1042 178 1094 212
rect 1220 178 1272 212
rect 1398 178 1450 212
rect 1576 178 1628 212
rect 1754 178 1806 212
rect 1932 178 1984 212
rect 2110 178 2162 212
rect 2288 178 2340 212
rect -2340 -212 -2288 -178
rect -2162 -212 -2110 -178
rect -1984 -212 -1932 -178
rect -1806 -212 -1754 -178
rect -1628 -212 -1576 -178
rect -1450 -212 -1398 -178
rect -1272 -212 -1220 -178
rect -1094 -212 -1042 -178
rect -916 -212 -864 -178
rect -738 -212 -686 -178
rect -560 -212 -508 -178
rect -382 -212 -330 -178
rect -204 -212 -152 -178
rect -26 -212 26 -178
rect 152 -212 204 -178
rect 330 -212 382 -178
rect 508 -212 560 -178
rect 686 -212 738 -178
rect 864 -212 916 -178
rect 1042 -212 1094 -178
rect 1220 -212 1272 -178
rect 1398 -212 1450 -178
rect 1576 -212 1628 -178
rect 1754 -212 1806 -178
rect 1932 -212 1984 -178
rect 2110 -212 2162 -178
rect 2288 -212 2340 -178
<< locali >>
rect -2420 178 -2340 212
rect -2288 178 -2272 212
rect -2178 178 -2162 212
rect -2110 178 -2094 212
rect -2000 178 -1984 212
rect -1932 178 -1916 212
rect -1822 178 -1806 212
rect -1754 178 -1738 212
rect -1644 178 -1628 212
rect -1576 178 -1560 212
rect -1466 178 -1450 212
rect -1398 178 -1382 212
rect -1288 178 -1272 212
rect -1220 178 -1204 212
rect -1110 178 -1094 212
rect -1042 178 -1026 212
rect -932 178 -916 212
rect -864 178 -848 212
rect -754 178 -738 212
rect -686 178 -670 212
rect -576 178 -560 212
rect -508 178 -492 212
rect -398 178 -382 212
rect -330 178 -314 212
rect -220 178 -204 212
rect -152 178 -136 212
rect -42 178 -26 212
rect 26 178 42 212
rect 136 178 152 212
rect 204 178 220 212
rect 314 178 330 212
rect 382 178 398 212
rect 492 178 508 212
rect 560 178 576 212
rect 670 178 686 212
rect 738 178 754 212
rect 848 178 864 212
rect 916 178 932 212
rect 1026 178 1042 212
rect 1094 178 1110 212
rect 1204 178 1220 212
rect 1272 178 1288 212
rect 1382 178 1398 212
rect 1450 178 1466 212
rect 1560 178 1576 212
rect 1628 178 1644 212
rect 1738 178 1754 212
rect 1806 178 1822 212
rect 1916 178 1932 212
rect 1984 178 2000 212
rect 2094 178 2110 212
rect 2162 178 2178 212
rect 2272 178 2288 212
rect 2340 178 2420 212
rect -2420 128 -2386 178
rect -2420 -178 -2386 -128
rect -2242 128 -2208 144
rect -2242 -144 -2208 -128
rect -2064 128 -2030 144
rect -2064 -144 -2030 -128
rect -1886 128 -1852 144
rect -1886 -144 -1852 -128
rect -1708 128 -1674 144
rect -1708 -144 -1674 -128
rect -1530 128 -1496 144
rect -1530 -144 -1496 -128
rect -1352 128 -1318 144
rect -1352 -144 -1318 -128
rect -1174 128 -1140 144
rect -1174 -144 -1140 -128
rect -996 128 -962 144
rect -996 -144 -962 -128
rect -818 128 -784 144
rect -818 -144 -784 -128
rect -640 128 -606 144
rect -640 -144 -606 -128
rect -462 128 -428 144
rect -462 -144 -428 -128
rect -284 128 -250 144
rect -284 -144 -250 -128
rect -106 128 -72 144
rect -106 -144 -72 -128
rect 72 128 106 144
rect 72 -144 106 -128
rect 250 128 284 144
rect 250 -144 284 -128
rect 428 128 462 144
rect 428 -144 462 -128
rect 606 128 640 144
rect 606 -144 640 -128
rect 784 128 818 144
rect 784 -144 818 -128
rect 962 128 996 144
rect 962 -144 996 -128
rect 1140 128 1174 144
rect 1140 -144 1174 -128
rect 1318 128 1352 144
rect 1318 -144 1352 -128
rect 1496 128 1530 144
rect 1496 -144 1530 -128
rect 1674 128 1708 144
rect 1674 -144 1708 -128
rect 1852 128 1886 144
rect 1852 -144 1886 -128
rect 2030 128 2064 144
rect 2030 -144 2064 -128
rect 2208 128 2242 144
rect 2208 -144 2242 -128
rect 2386 128 2420 178
rect 2386 -178 2420 -128
rect -2420 -212 -2340 -178
rect -2288 -212 -2272 -178
rect -2178 -212 -2162 -178
rect -2110 -212 -2094 -178
rect -2000 -212 -1984 -178
rect -1932 -212 -1916 -178
rect -1822 -212 -1806 -178
rect -1754 -212 -1738 -178
rect -1644 -212 -1628 -178
rect -1576 -212 -1560 -178
rect -1466 -212 -1450 -178
rect -1398 -212 -1382 -178
rect -1288 -212 -1272 -178
rect -1220 -212 -1204 -178
rect -1110 -212 -1094 -178
rect -1042 -212 -1026 -178
rect -932 -212 -916 -178
rect -864 -212 -848 -178
rect -754 -212 -738 -178
rect -686 -212 -670 -178
rect -576 -212 -560 -178
rect -508 -212 -492 -178
rect -398 -212 -382 -178
rect -330 -212 -314 -178
rect -220 -212 -204 -178
rect -152 -212 -136 -178
rect -42 -212 -26 -178
rect 26 -212 42 -178
rect 136 -212 152 -178
rect 204 -212 220 -178
rect 314 -212 330 -178
rect 382 -212 398 -178
rect 492 -212 508 -178
rect 560 -212 576 -178
rect 670 -212 686 -178
rect 738 -212 754 -178
rect 848 -212 864 -178
rect 916 -212 932 -178
rect 1026 -212 1042 -178
rect 1094 -212 1110 -178
rect 1204 -212 1220 -178
rect 1272 -212 1288 -178
rect 1382 -212 1398 -178
rect 1450 -212 1466 -178
rect 1560 -212 1576 -178
rect 1628 -212 1644 -178
rect 1738 -212 1754 -178
rect 1806 -212 1822 -178
rect 1916 -212 1932 -178
rect 1984 -212 2000 -178
rect 2094 -212 2110 -178
rect 2162 -212 2178 -178
rect 2272 -212 2288 -178
rect 2340 -212 2420 -178
<< viali >>
rect -2162 178 -2110 212
rect -1984 178 -1932 212
rect -1806 178 -1754 212
rect -1628 178 -1576 212
rect -1450 178 -1398 212
rect -1272 178 -1220 212
rect -1094 178 -1042 212
rect -916 178 -864 212
rect -738 178 -686 212
rect -560 178 -508 212
rect -382 178 -330 212
rect -204 178 -152 212
rect -26 178 26 212
rect 152 178 204 212
rect 330 178 382 212
rect 508 178 560 212
rect 686 178 738 212
rect 864 178 916 212
rect 1042 178 1094 212
rect 1220 178 1272 212
rect 1398 178 1450 212
rect 1576 178 1628 212
rect 1754 178 1806 212
rect 1932 178 1984 212
rect 2110 178 2162 212
rect -2162 -212 -2110 -178
rect -1984 -212 -1932 -178
rect -1806 -212 -1754 -178
rect -1628 -212 -1576 -178
rect -1450 -212 -1398 -178
rect -1272 -212 -1220 -178
rect -1094 -212 -1042 -178
rect -916 -212 -864 -178
rect -738 -212 -686 -178
rect -560 -212 -508 -178
rect -382 -212 -330 -178
rect -204 -212 -152 -178
rect -26 -212 26 -178
rect 152 -212 204 -178
rect 330 -212 382 -178
rect 508 -212 560 -178
rect 686 -212 738 -178
rect 864 -212 916 -178
rect 1042 -212 1094 -178
rect 1220 -212 1272 -178
rect 1398 -212 1450 -178
rect 1576 -212 1628 -178
rect 1754 -212 1806 -178
rect 1932 -212 1984 -178
rect 2110 -212 2162 -178
<< metal1 >>
rect -2174 212 -2098 218
rect -2174 178 -2162 212
rect -2110 178 -2098 212
rect -2174 172 -2098 178
rect -1996 212 -1920 218
rect -1996 178 -1984 212
rect -1932 178 -1920 212
rect -1996 172 -1920 178
rect -1818 212 -1742 218
rect -1818 178 -1806 212
rect -1754 178 -1742 212
rect -1818 172 -1742 178
rect -1640 212 -1564 218
rect -1640 178 -1628 212
rect -1576 178 -1564 212
rect -1640 172 -1564 178
rect -1462 212 -1386 218
rect -1462 178 -1450 212
rect -1398 178 -1386 212
rect -1462 172 -1386 178
rect -1284 212 -1208 218
rect -1284 178 -1272 212
rect -1220 178 -1208 212
rect -1284 172 -1208 178
rect -1106 212 -1030 218
rect -1106 178 -1094 212
rect -1042 178 -1030 212
rect -1106 172 -1030 178
rect -928 212 -852 218
rect -928 178 -916 212
rect -864 178 -852 212
rect -928 172 -852 178
rect -750 212 -674 218
rect -750 178 -738 212
rect -686 178 -674 212
rect -750 172 -674 178
rect -572 212 -496 218
rect -572 178 -560 212
rect -508 178 -496 212
rect -572 172 -496 178
rect -394 212 -318 218
rect -394 178 -382 212
rect -330 178 -318 212
rect -394 172 -318 178
rect -216 212 -140 218
rect -216 178 -204 212
rect -152 178 -140 212
rect -216 172 -140 178
rect -38 212 38 218
rect -38 178 -26 212
rect 26 178 38 212
rect -38 172 38 178
rect 140 212 216 218
rect 140 178 152 212
rect 204 178 216 212
rect 140 172 216 178
rect 318 212 394 218
rect 318 178 330 212
rect 382 178 394 212
rect 318 172 394 178
rect 496 212 572 218
rect 496 178 508 212
rect 560 178 572 212
rect 496 172 572 178
rect 674 212 750 218
rect 674 178 686 212
rect 738 178 750 212
rect 674 172 750 178
rect 852 212 928 218
rect 852 178 864 212
rect 916 178 928 212
rect 852 172 928 178
rect 1030 212 1106 218
rect 1030 178 1042 212
rect 1094 178 1106 212
rect 1030 172 1106 178
rect 1208 212 1284 218
rect 1208 178 1220 212
rect 1272 178 1284 212
rect 1208 172 1284 178
rect 1386 212 1462 218
rect 1386 178 1398 212
rect 1450 178 1462 212
rect 1386 172 1462 178
rect 1564 212 1640 218
rect 1564 178 1576 212
rect 1628 178 1640 212
rect 1564 172 1640 178
rect 1742 212 1818 218
rect 1742 178 1754 212
rect 1806 178 1818 212
rect 1742 172 1818 178
rect 1920 212 1996 218
rect 1920 178 1932 212
rect 1984 178 1996 212
rect 1920 172 1996 178
rect 2098 212 2174 218
rect 2098 178 2110 212
rect 2162 178 2174 212
rect 2098 172 2174 178
rect -2174 -178 -2098 -172
rect -2174 -212 -2162 -178
rect -2110 -212 -2098 -178
rect -2174 -218 -2098 -212
rect -1996 -178 -1920 -172
rect -1996 -212 -1984 -178
rect -1932 -212 -1920 -178
rect -1996 -218 -1920 -212
rect -1818 -178 -1742 -172
rect -1818 -212 -1806 -178
rect -1754 -212 -1742 -178
rect -1818 -218 -1742 -212
rect -1640 -178 -1564 -172
rect -1640 -212 -1628 -178
rect -1576 -212 -1564 -178
rect -1640 -218 -1564 -212
rect -1462 -178 -1386 -172
rect -1462 -212 -1450 -178
rect -1398 -212 -1386 -178
rect -1462 -218 -1386 -212
rect -1284 -178 -1208 -172
rect -1284 -212 -1272 -178
rect -1220 -212 -1208 -178
rect -1284 -218 -1208 -212
rect -1106 -178 -1030 -172
rect -1106 -212 -1094 -178
rect -1042 -212 -1030 -178
rect -1106 -218 -1030 -212
rect -928 -178 -852 -172
rect -928 -212 -916 -178
rect -864 -212 -852 -178
rect -928 -218 -852 -212
rect -750 -178 -674 -172
rect -750 -212 -738 -178
rect -686 -212 -674 -178
rect -750 -218 -674 -212
rect -572 -178 -496 -172
rect -572 -212 -560 -178
rect -508 -212 -496 -178
rect -572 -218 -496 -212
rect -394 -178 -318 -172
rect -394 -212 -382 -178
rect -330 -212 -318 -178
rect -394 -218 -318 -212
rect -216 -178 -140 -172
rect -216 -212 -204 -178
rect -152 -212 -140 -178
rect -216 -218 -140 -212
rect -38 -178 38 -172
rect -38 -212 -26 -178
rect 26 -212 38 -178
rect -38 -218 38 -212
rect 140 -178 216 -172
rect 140 -212 152 -178
rect 204 -212 216 -178
rect 140 -218 216 -212
rect 318 -178 394 -172
rect 318 -212 330 -178
rect 382 -212 394 -178
rect 318 -218 394 -212
rect 496 -178 572 -172
rect 496 -212 508 -178
rect 560 -212 572 -178
rect 496 -218 572 -212
rect 674 -178 750 -172
rect 674 -212 686 -178
rect 738 -212 750 -178
rect 674 -218 750 -212
rect 852 -178 928 -172
rect 852 -212 864 -178
rect 916 -212 928 -178
rect 852 -218 928 -212
rect 1030 -178 1106 -172
rect 1030 -212 1042 -178
rect 1094 -212 1106 -178
rect 1030 -218 1106 -212
rect 1208 -178 1284 -172
rect 1208 -212 1220 -178
rect 1272 -212 1284 -178
rect 1208 -218 1284 -212
rect 1386 -178 1462 -172
rect 1386 -212 1398 -178
rect 1450 -212 1462 -178
rect 1386 -218 1462 -212
rect 1564 -178 1640 -172
rect 1564 -212 1576 -178
rect 1628 -212 1640 -178
rect 1564 -218 1640 -212
rect 1742 -178 1818 -172
rect 1742 -212 1754 -178
rect 1806 -212 1818 -178
rect 1742 -218 1818 -212
rect 1920 -178 1996 -172
rect 1920 -212 1932 -178
rect 1984 -212 1996 -178
rect 1920 -218 1996 -212
rect 2098 -178 2174 -172
rect 2098 -212 2110 -178
rect 2162 -212 2174 -178
rect 2098 -218 2174 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 27 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
