magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -1469 172 -1411 178
rect -1277 172 -1219 178
rect -1085 172 -1027 178
rect -893 172 -835 178
rect -701 172 -643 178
rect -509 172 -451 178
rect -317 172 -259 178
rect -125 172 -67 178
rect 67 172 125 178
rect 259 172 317 178
rect 451 172 509 178
rect 643 172 701 178
rect 835 172 893 178
rect 1027 172 1085 178
rect 1219 172 1277 178
rect 1411 172 1469 178
rect -1469 138 -1457 172
rect -1277 138 -1265 172
rect -1085 138 -1073 172
rect -893 138 -881 172
rect -701 138 -689 172
rect -509 138 -497 172
rect -317 138 -305 172
rect -125 138 -113 172
rect 67 138 79 172
rect 259 138 271 172
rect 451 138 463 172
rect 643 138 655 172
rect 835 138 847 172
rect 1027 138 1039 172
rect 1219 138 1231 172
rect 1411 138 1423 172
rect -1469 132 -1411 138
rect -1277 132 -1219 138
rect -1085 132 -1027 138
rect -893 132 -835 138
rect -701 132 -643 138
rect -509 132 -451 138
rect -317 132 -259 138
rect -125 132 -67 138
rect 67 132 125 138
rect 259 132 317 138
rect 451 132 509 138
rect 643 132 701 138
rect 835 132 893 138
rect 1027 132 1085 138
rect 1219 132 1277 138
rect 1411 132 1469 138
<< pwell >>
rect -1789 -300 1789 300
<< nmos >>
rect -1599 -100 -1569 100
rect -1503 -100 -1473 100
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
rect 1473 -100 1503 100
rect 1569 -100 1599 100
<< ndiff >>
rect -1661 85 -1599 100
rect -1661 51 -1649 85
rect -1615 51 -1599 85
rect -1661 17 -1599 51
rect -1661 -17 -1649 17
rect -1615 -17 -1599 17
rect -1661 -51 -1599 -17
rect -1661 -85 -1649 -51
rect -1615 -85 -1599 -51
rect -1661 -100 -1599 -85
rect -1569 85 -1503 100
rect -1569 51 -1553 85
rect -1519 51 -1503 85
rect -1569 17 -1503 51
rect -1569 -17 -1553 17
rect -1519 -17 -1503 17
rect -1569 -51 -1503 -17
rect -1569 -85 -1553 -51
rect -1519 -85 -1503 -51
rect -1569 -100 -1503 -85
rect -1473 85 -1407 100
rect -1473 51 -1457 85
rect -1423 51 -1407 85
rect -1473 17 -1407 51
rect -1473 -17 -1457 17
rect -1423 -17 -1407 17
rect -1473 -51 -1407 -17
rect -1473 -85 -1457 -51
rect -1423 -85 -1407 -51
rect -1473 -100 -1407 -85
rect -1377 85 -1311 100
rect -1377 51 -1361 85
rect -1327 51 -1311 85
rect -1377 17 -1311 51
rect -1377 -17 -1361 17
rect -1327 -17 -1311 17
rect -1377 -51 -1311 -17
rect -1377 -85 -1361 -51
rect -1327 -85 -1311 -51
rect -1377 -100 -1311 -85
rect -1281 85 -1215 100
rect -1281 51 -1265 85
rect -1231 51 -1215 85
rect -1281 17 -1215 51
rect -1281 -17 -1265 17
rect -1231 -17 -1215 17
rect -1281 -51 -1215 -17
rect -1281 -85 -1265 -51
rect -1231 -85 -1215 -51
rect -1281 -100 -1215 -85
rect -1185 85 -1119 100
rect -1185 51 -1169 85
rect -1135 51 -1119 85
rect -1185 17 -1119 51
rect -1185 -17 -1169 17
rect -1135 -17 -1119 17
rect -1185 -51 -1119 -17
rect -1185 -85 -1169 -51
rect -1135 -85 -1119 -51
rect -1185 -100 -1119 -85
rect -1089 85 -1023 100
rect -1089 51 -1073 85
rect -1039 51 -1023 85
rect -1089 17 -1023 51
rect -1089 -17 -1073 17
rect -1039 -17 -1023 17
rect -1089 -51 -1023 -17
rect -1089 -85 -1073 -51
rect -1039 -85 -1023 -51
rect -1089 -100 -1023 -85
rect -993 85 -927 100
rect -993 51 -977 85
rect -943 51 -927 85
rect -993 17 -927 51
rect -993 -17 -977 17
rect -943 -17 -927 17
rect -993 -51 -927 -17
rect -993 -85 -977 -51
rect -943 -85 -927 -51
rect -993 -100 -927 -85
rect -897 85 -831 100
rect -897 51 -881 85
rect -847 51 -831 85
rect -897 17 -831 51
rect -897 -17 -881 17
rect -847 -17 -831 17
rect -897 -51 -831 -17
rect -897 -85 -881 -51
rect -847 -85 -831 -51
rect -897 -100 -831 -85
rect -801 85 -735 100
rect -801 51 -785 85
rect -751 51 -735 85
rect -801 17 -735 51
rect -801 -17 -785 17
rect -751 -17 -735 17
rect -801 -51 -735 -17
rect -801 -85 -785 -51
rect -751 -85 -735 -51
rect -801 -100 -735 -85
rect -705 85 -639 100
rect -705 51 -689 85
rect -655 51 -639 85
rect -705 17 -639 51
rect -705 -17 -689 17
rect -655 -17 -639 17
rect -705 -51 -639 -17
rect -705 -85 -689 -51
rect -655 -85 -639 -51
rect -705 -100 -639 -85
rect -609 85 -543 100
rect -609 51 -593 85
rect -559 51 -543 85
rect -609 17 -543 51
rect -609 -17 -593 17
rect -559 -17 -543 17
rect -609 -51 -543 -17
rect -609 -85 -593 -51
rect -559 -85 -543 -51
rect -609 -100 -543 -85
rect -513 85 -447 100
rect -513 51 -497 85
rect -463 51 -447 85
rect -513 17 -447 51
rect -513 -17 -497 17
rect -463 -17 -447 17
rect -513 -51 -447 -17
rect -513 -85 -497 -51
rect -463 -85 -447 -51
rect -513 -100 -447 -85
rect -417 85 -351 100
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -100 -351 -85
rect -321 85 -255 100
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -100 -255 -85
rect -225 85 -159 100
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 225 100
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -100 225 -85
rect 255 85 321 100
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -100 321 -85
rect 351 85 417 100
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -100 417 -85
rect 447 85 513 100
rect 447 51 463 85
rect 497 51 513 85
rect 447 17 513 51
rect 447 -17 463 17
rect 497 -17 513 17
rect 447 -51 513 -17
rect 447 -85 463 -51
rect 497 -85 513 -51
rect 447 -100 513 -85
rect 543 85 609 100
rect 543 51 559 85
rect 593 51 609 85
rect 543 17 609 51
rect 543 -17 559 17
rect 593 -17 609 17
rect 543 -51 609 -17
rect 543 -85 559 -51
rect 593 -85 609 -51
rect 543 -100 609 -85
rect 639 85 705 100
rect 639 51 655 85
rect 689 51 705 85
rect 639 17 705 51
rect 639 -17 655 17
rect 689 -17 705 17
rect 639 -51 705 -17
rect 639 -85 655 -51
rect 689 -85 705 -51
rect 639 -100 705 -85
rect 735 85 801 100
rect 735 51 751 85
rect 785 51 801 85
rect 735 17 801 51
rect 735 -17 751 17
rect 785 -17 801 17
rect 735 -51 801 -17
rect 735 -85 751 -51
rect 785 -85 801 -51
rect 735 -100 801 -85
rect 831 85 897 100
rect 831 51 847 85
rect 881 51 897 85
rect 831 17 897 51
rect 831 -17 847 17
rect 881 -17 897 17
rect 831 -51 897 -17
rect 831 -85 847 -51
rect 881 -85 897 -51
rect 831 -100 897 -85
rect 927 85 993 100
rect 927 51 943 85
rect 977 51 993 85
rect 927 17 993 51
rect 927 -17 943 17
rect 977 -17 993 17
rect 927 -51 993 -17
rect 927 -85 943 -51
rect 977 -85 993 -51
rect 927 -100 993 -85
rect 1023 85 1089 100
rect 1023 51 1039 85
rect 1073 51 1089 85
rect 1023 17 1089 51
rect 1023 -17 1039 17
rect 1073 -17 1089 17
rect 1023 -51 1089 -17
rect 1023 -85 1039 -51
rect 1073 -85 1089 -51
rect 1023 -100 1089 -85
rect 1119 85 1185 100
rect 1119 51 1135 85
rect 1169 51 1185 85
rect 1119 17 1185 51
rect 1119 -17 1135 17
rect 1169 -17 1185 17
rect 1119 -51 1185 -17
rect 1119 -85 1135 -51
rect 1169 -85 1185 -51
rect 1119 -100 1185 -85
rect 1215 85 1281 100
rect 1215 51 1231 85
rect 1265 51 1281 85
rect 1215 17 1281 51
rect 1215 -17 1231 17
rect 1265 -17 1281 17
rect 1215 -51 1281 -17
rect 1215 -85 1231 -51
rect 1265 -85 1281 -51
rect 1215 -100 1281 -85
rect 1311 85 1377 100
rect 1311 51 1327 85
rect 1361 51 1377 85
rect 1311 17 1377 51
rect 1311 -17 1327 17
rect 1361 -17 1377 17
rect 1311 -51 1377 -17
rect 1311 -85 1327 -51
rect 1361 -85 1377 -51
rect 1311 -100 1377 -85
rect 1407 85 1473 100
rect 1407 51 1423 85
rect 1457 51 1473 85
rect 1407 17 1473 51
rect 1407 -17 1423 17
rect 1457 -17 1473 17
rect 1407 -51 1473 -17
rect 1407 -85 1423 -51
rect 1457 -85 1473 -51
rect 1407 -100 1473 -85
rect 1503 85 1569 100
rect 1503 51 1519 85
rect 1553 51 1569 85
rect 1503 17 1569 51
rect 1503 -17 1519 17
rect 1553 -17 1569 17
rect 1503 -51 1569 -17
rect 1503 -85 1519 -51
rect 1553 -85 1569 -51
rect 1503 -100 1569 -85
rect 1599 85 1661 100
rect 1599 51 1615 85
rect 1649 51 1661 85
rect 1599 17 1661 51
rect 1599 -17 1615 17
rect 1649 -17 1661 17
rect 1599 -51 1661 -17
rect 1599 -85 1615 -51
rect 1649 -85 1661 -51
rect 1599 -100 1661 -85
<< ndiffc >>
rect -1649 51 -1615 85
rect -1649 -17 -1615 17
rect -1649 -85 -1615 -51
rect -1553 51 -1519 85
rect -1553 -17 -1519 17
rect -1553 -85 -1519 -51
rect -1457 51 -1423 85
rect -1457 -17 -1423 17
rect -1457 -85 -1423 -51
rect -1361 51 -1327 85
rect -1361 -17 -1327 17
rect -1361 -85 -1327 -51
rect -1265 51 -1231 85
rect -1265 -17 -1231 17
rect -1265 -85 -1231 -51
rect -1169 51 -1135 85
rect -1169 -17 -1135 17
rect -1169 -85 -1135 -51
rect -1073 51 -1039 85
rect -1073 -17 -1039 17
rect -1073 -85 -1039 -51
rect -977 51 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -51
rect -881 51 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -51
rect -785 51 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -51
rect -689 51 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -51
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
rect 655 51 689 85
rect 655 -17 689 17
rect 655 -85 689 -51
rect 751 51 785 85
rect 751 -17 785 17
rect 751 -85 785 -51
rect 847 51 881 85
rect 847 -17 881 17
rect 847 -85 881 -51
rect 943 51 977 85
rect 943 -17 977 17
rect 943 -85 977 -51
rect 1039 51 1073 85
rect 1039 -17 1073 17
rect 1039 -85 1073 -51
rect 1135 51 1169 85
rect 1135 -17 1169 17
rect 1135 -85 1169 -51
rect 1231 51 1265 85
rect 1231 -17 1265 17
rect 1231 -85 1265 -51
rect 1327 51 1361 85
rect 1327 -17 1361 17
rect 1327 -85 1361 -51
rect 1423 51 1457 85
rect 1423 -17 1457 17
rect 1423 -85 1457 -51
rect 1519 51 1553 85
rect 1519 -17 1553 17
rect 1519 -85 1553 -51
rect 1615 51 1649 85
rect 1615 -17 1649 17
rect 1615 -85 1649 -51
<< psubdiff >>
rect -1763 240 -1649 274
rect -1615 240 -1581 274
rect -1547 240 -1513 274
rect -1479 240 -1445 274
rect -1411 240 -1377 274
rect -1343 240 -1309 274
rect -1275 240 -1241 274
rect -1207 240 -1173 274
rect -1139 240 -1105 274
rect -1071 240 -1037 274
rect -1003 240 -969 274
rect -935 240 -901 274
rect -867 240 -833 274
rect -799 240 -765 274
rect -731 240 -697 274
rect -663 240 -629 274
rect -595 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 595 274
rect 629 240 663 274
rect 697 240 731 274
rect 765 240 799 274
rect 833 240 867 274
rect 901 240 935 274
rect 969 240 1003 274
rect 1037 240 1071 274
rect 1105 240 1139 274
rect 1173 240 1207 274
rect 1241 240 1275 274
rect 1309 240 1343 274
rect 1377 240 1411 274
rect 1445 240 1479 274
rect 1513 240 1547 274
rect 1581 240 1615 274
rect 1649 240 1763 274
rect -1763 153 -1729 240
rect -1763 85 -1729 119
rect 1729 153 1763 240
rect -1763 17 -1729 51
rect -1763 -51 -1729 -17
rect -1763 -119 -1729 -85
rect 1729 85 1763 119
rect 1729 17 1763 51
rect 1729 -51 1763 -17
rect -1763 -240 -1729 -153
rect 1729 -119 1763 -85
rect 1729 -240 1763 -153
rect -1763 -274 -1649 -240
rect -1615 -274 -1581 -240
rect -1547 -274 -1513 -240
rect -1479 -274 -1445 -240
rect -1411 -274 -1377 -240
rect -1343 -274 -1309 -240
rect -1275 -274 -1241 -240
rect -1207 -274 -1173 -240
rect -1139 -274 -1105 -240
rect -1071 -274 -1037 -240
rect -1003 -274 -969 -240
rect -935 -274 -901 -240
rect -867 -274 -833 -240
rect -799 -274 -765 -240
rect -731 -274 -697 -240
rect -663 -274 -629 -240
rect -595 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 595 -240
rect 629 -274 663 -240
rect 697 -274 731 -240
rect 765 -274 799 -240
rect 833 -274 867 -240
rect 901 -274 935 -240
rect 969 -274 1003 -240
rect 1037 -274 1071 -240
rect 1105 -274 1139 -240
rect 1173 -274 1207 -240
rect 1241 -274 1275 -240
rect 1309 -274 1343 -240
rect 1377 -274 1411 -240
rect 1445 -274 1479 -240
rect 1513 -274 1547 -240
rect 1581 -274 1615 -240
rect 1649 -274 1763 -240
<< psubdiffcont >>
rect -1649 240 -1615 274
rect -1581 240 -1547 274
rect -1513 240 -1479 274
rect -1445 240 -1411 274
rect -1377 240 -1343 274
rect -1309 240 -1275 274
rect -1241 240 -1207 274
rect -1173 240 -1139 274
rect -1105 240 -1071 274
rect -1037 240 -1003 274
rect -969 240 -935 274
rect -901 240 -867 274
rect -833 240 -799 274
rect -765 240 -731 274
rect -697 240 -663 274
rect -629 240 -595 274
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect 595 240 629 274
rect 663 240 697 274
rect 731 240 765 274
rect 799 240 833 274
rect 867 240 901 274
rect 935 240 969 274
rect 1003 240 1037 274
rect 1071 240 1105 274
rect 1139 240 1173 274
rect 1207 240 1241 274
rect 1275 240 1309 274
rect 1343 240 1377 274
rect 1411 240 1445 274
rect 1479 240 1513 274
rect 1547 240 1581 274
rect 1615 240 1649 274
rect -1763 119 -1729 153
rect 1729 119 1763 153
rect -1763 51 -1729 85
rect -1763 -17 -1729 17
rect -1763 -85 -1729 -51
rect 1729 51 1763 85
rect 1729 -17 1763 17
rect 1729 -85 1763 -51
rect -1763 -153 -1729 -119
rect 1729 -153 1763 -119
rect -1649 -274 -1615 -240
rect -1581 -274 -1547 -240
rect -1513 -274 -1479 -240
rect -1445 -274 -1411 -240
rect -1377 -274 -1343 -240
rect -1309 -274 -1275 -240
rect -1241 -274 -1207 -240
rect -1173 -274 -1139 -240
rect -1105 -274 -1071 -240
rect -1037 -274 -1003 -240
rect -969 -274 -935 -240
rect -901 -274 -867 -240
rect -833 -274 -799 -240
rect -765 -274 -731 -240
rect -697 -274 -663 -240
rect -629 -274 -595 -240
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
rect 595 -274 629 -240
rect 663 -274 697 -240
rect 731 -274 765 -240
rect 799 -274 833 -240
rect 867 -274 901 -240
rect 935 -274 969 -240
rect 1003 -274 1037 -240
rect 1071 -274 1105 -240
rect 1139 -274 1173 -240
rect 1207 -274 1241 -240
rect 1275 -274 1309 -240
rect 1343 -274 1377 -240
rect 1411 -274 1445 -240
rect 1479 -274 1513 -240
rect 1547 -274 1581 -240
rect 1615 -274 1649 -240
<< poly >>
rect -1521 172 1521 188
rect -1521 138 -1457 172
rect -1423 138 -1265 172
rect -1231 138 -1073 172
rect -1039 138 -881 172
rect -847 138 -689 172
rect -655 138 -497 172
rect -463 138 -305 172
rect -271 138 -113 172
rect -79 138 79 172
rect 113 138 271 172
rect 305 138 463 172
rect 497 138 655 172
rect 689 138 847 172
rect 881 138 1039 172
rect 1073 138 1231 172
rect 1265 138 1423 172
rect 1457 138 1521 172
rect -1599 100 -1569 126
rect -1521 122 1521 138
rect -1503 100 -1473 122
rect -1407 100 -1377 122
rect -1311 100 -1281 122
rect -1215 100 -1185 122
rect -1119 100 -1089 122
rect -1023 100 -993 122
rect -927 100 -897 122
rect -831 100 -801 122
rect -735 100 -705 122
rect -639 100 -609 122
rect -543 100 -513 122
rect -447 100 -417 122
rect -351 100 -321 122
rect -255 100 -225 122
rect -159 100 -129 122
rect -63 100 -33 122
rect 33 100 63 122
rect 129 100 159 122
rect 225 100 255 122
rect 321 100 351 122
rect 417 100 447 122
rect 513 100 543 122
rect 609 100 639 122
rect 705 100 735 122
rect 801 100 831 122
rect 897 100 927 122
rect 993 100 1023 122
rect 1089 100 1119 122
rect 1185 100 1215 122
rect 1281 100 1311 122
rect 1377 100 1407 122
rect 1473 100 1503 122
rect 1569 100 1599 126
rect -1599 -122 -1569 -100
rect -1617 -138 -1551 -122
rect -1503 -126 -1473 -100
rect -1407 -126 -1377 -100
rect -1311 -126 -1281 -100
rect -1215 -126 -1185 -100
rect -1119 -126 -1089 -100
rect -1023 -126 -993 -100
rect -927 -126 -897 -100
rect -831 -126 -801 -100
rect -735 -126 -705 -100
rect -639 -126 -609 -100
rect -543 -126 -513 -100
rect -447 -126 -417 -100
rect -351 -126 -321 -100
rect -255 -126 -225 -100
rect -159 -126 -129 -100
rect -63 -126 -33 -100
rect 33 -126 63 -100
rect 129 -126 159 -100
rect 225 -126 255 -100
rect 321 -126 351 -100
rect 417 -126 447 -100
rect 513 -126 543 -100
rect 609 -126 639 -100
rect 705 -126 735 -100
rect 801 -126 831 -100
rect 897 -126 927 -100
rect 993 -126 1023 -100
rect 1089 -126 1119 -100
rect 1185 -126 1215 -100
rect 1281 -126 1311 -100
rect 1377 -126 1407 -100
rect 1473 -126 1503 -100
rect 1569 -126 1599 -100
rect -1617 -172 -1601 -138
rect -1567 -172 -1551 -138
rect -1617 -188 -1551 -172
rect 1551 -142 1617 -126
rect 1551 -176 1567 -142
rect 1601 -176 1617 -142
rect 1551 -192 1617 -176
<< polycont >>
rect -1457 138 -1423 172
rect -1265 138 -1231 172
rect -1073 138 -1039 172
rect -881 138 -847 172
rect -689 138 -655 172
rect -497 138 -463 172
rect -305 138 -271 172
rect -113 138 -79 172
rect 79 138 113 172
rect 271 138 305 172
rect 463 138 497 172
rect 655 138 689 172
rect 847 138 881 172
rect 1039 138 1073 172
rect 1231 138 1265 172
rect 1423 138 1457 172
rect -1601 -172 -1567 -138
rect 1567 -176 1601 -142
<< locali >>
rect -1763 240 -1649 274
rect -1615 240 -1581 274
rect -1547 240 -1513 274
rect -1479 240 -1445 274
rect -1411 240 -1377 274
rect -1343 240 -1309 274
rect -1275 240 -1241 274
rect -1207 240 -1173 274
rect -1139 240 -1105 274
rect -1071 240 -1037 274
rect -1003 240 -969 274
rect -935 240 -901 274
rect -867 240 -833 274
rect -799 240 -765 274
rect -731 240 -697 274
rect -663 240 -629 274
rect -595 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 595 274
rect 629 240 663 274
rect 697 240 731 274
rect 765 240 799 274
rect 833 240 867 274
rect 901 240 935 274
rect 969 240 1003 274
rect 1037 240 1071 274
rect 1105 240 1139 274
rect 1173 240 1207 274
rect 1241 240 1275 274
rect 1309 240 1343 274
rect 1377 240 1411 274
rect 1445 240 1479 274
rect 1513 240 1547 274
rect 1581 240 1615 274
rect 1649 240 1763 274
rect -1763 153 -1729 240
rect -1473 138 -1457 172
rect -1423 138 -1407 172
rect -1281 138 -1265 172
rect -1231 138 -1215 172
rect -1089 138 -1073 172
rect -1039 138 -1023 172
rect -897 138 -881 172
rect -847 138 -831 172
rect -705 138 -689 172
rect -655 138 -639 172
rect -513 138 -497 172
rect -463 138 -447 172
rect -321 138 -305 172
rect -271 138 -255 172
rect -129 138 -113 172
rect -79 138 -63 172
rect 63 138 79 172
rect 113 138 129 172
rect 255 138 271 172
rect 305 138 321 172
rect 447 138 463 172
rect 497 138 513 172
rect 639 138 655 172
rect 689 138 705 172
rect 831 138 847 172
rect 881 138 897 172
rect 1023 138 1039 172
rect 1073 138 1089 172
rect 1215 138 1231 172
rect 1265 138 1281 172
rect 1407 138 1423 172
rect 1457 138 1473 172
rect 1729 153 1763 240
rect -1763 85 -1729 119
rect -1763 17 -1729 51
rect -1763 -51 -1729 -17
rect -1763 -119 -1729 -85
rect -1763 -240 -1729 -153
rect -1649 85 -1615 104
rect -1649 17 -1615 51
rect -1649 -51 -1615 -17
rect -1649 -138 -1615 -85
rect -1553 85 -1519 104
rect -1553 17 -1519 51
rect -1553 -51 -1519 -17
rect -1553 -104 -1519 -85
rect -1457 85 -1423 104
rect -1457 17 -1423 51
rect -1457 -51 -1423 -17
rect -1457 -104 -1423 -85
rect -1361 85 -1327 104
rect -1361 17 -1327 51
rect -1361 -51 -1327 -17
rect -1361 -104 -1327 -85
rect -1265 85 -1231 104
rect -1265 17 -1231 51
rect -1265 -51 -1231 -17
rect -1265 -104 -1231 -85
rect -1169 85 -1135 104
rect -1169 17 -1135 51
rect -1169 -51 -1135 -17
rect -1169 -104 -1135 -85
rect -1073 85 -1039 104
rect -1073 17 -1039 51
rect -1073 -51 -1039 -17
rect -1073 -104 -1039 -85
rect -977 85 -943 104
rect -977 17 -943 51
rect -977 -51 -943 -17
rect -977 -104 -943 -85
rect -881 85 -847 104
rect -881 17 -847 51
rect -881 -51 -847 -17
rect -881 -104 -847 -85
rect -785 85 -751 104
rect -785 17 -751 51
rect -785 -51 -751 -17
rect -785 -104 -751 -85
rect -689 85 -655 104
rect -689 17 -655 51
rect -689 -51 -655 -17
rect -689 -104 -655 -85
rect -593 85 -559 104
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -104 -559 -85
rect -497 85 -463 104
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -104 -463 -85
rect -401 85 -367 104
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -104 -367 -85
rect -305 85 -271 104
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -104 -271 -85
rect -209 85 -175 104
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -104 209 -85
rect 271 85 305 104
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -104 305 -85
rect 367 85 401 104
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -104 401 -85
rect 463 85 497 104
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -104 497 -85
rect 559 85 593 104
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -104 593 -85
rect 655 85 689 104
rect 655 17 689 51
rect 655 -51 689 -17
rect 655 -104 689 -85
rect 751 85 785 104
rect 751 17 785 51
rect 751 -51 785 -17
rect 751 -104 785 -85
rect 847 85 881 104
rect 847 17 881 51
rect 847 -51 881 -17
rect 847 -104 881 -85
rect 943 85 977 104
rect 943 17 977 51
rect 943 -51 977 -17
rect 943 -104 977 -85
rect 1039 85 1073 104
rect 1039 17 1073 51
rect 1039 -51 1073 -17
rect 1039 -104 1073 -85
rect 1135 85 1169 104
rect 1135 17 1169 51
rect 1135 -51 1169 -17
rect 1135 -104 1169 -85
rect 1231 85 1265 104
rect 1231 17 1265 51
rect 1231 -51 1265 -17
rect 1231 -104 1265 -85
rect 1327 85 1361 104
rect 1327 17 1361 51
rect 1327 -51 1361 -17
rect 1327 -104 1361 -85
rect 1423 85 1457 104
rect 1423 17 1457 51
rect 1423 -51 1457 -17
rect 1423 -104 1457 -85
rect 1519 85 1553 104
rect 1519 17 1553 51
rect 1519 -51 1553 -17
rect 1519 -104 1553 -85
rect 1615 85 1649 104
rect 1615 17 1649 51
rect 1615 -51 1649 -17
rect -1649 -172 -1601 -138
rect -1567 -172 -1551 -138
rect 1615 -142 1649 -85
rect -1649 -240 -1615 -172
rect 1551 -176 1567 -142
rect 1601 -176 1649 -142
rect 1615 -240 1649 -176
rect 1729 85 1763 119
rect 1729 17 1763 51
rect 1729 -51 1763 -17
rect 1729 -119 1763 -85
rect 1729 -240 1763 -153
rect -1763 -274 -1649 -240
rect -1615 -274 -1581 -240
rect -1547 -274 -1513 -240
rect -1479 -274 -1445 -240
rect -1411 -274 -1377 -240
rect -1343 -274 -1309 -240
rect -1275 -274 -1241 -240
rect -1207 -274 -1173 -240
rect -1139 -274 -1105 -240
rect -1071 -274 -1037 -240
rect -1003 -274 -969 -240
rect -935 -274 -901 -240
rect -867 -274 -833 -240
rect -799 -274 -765 -240
rect -731 -274 -697 -240
rect -663 -274 -629 -240
rect -595 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 595 -240
rect 629 -274 663 -240
rect 697 -274 731 -240
rect 765 -274 799 -240
rect 833 -274 867 -240
rect 901 -274 935 -240
rect 969 -274 1003 -240
rect 1037 -274 1071 -240
rect 1105 -274 1139 -240
rect 1173 -274 1207 -240
rect 1241 -274 1275 -240
rect 1309 -274 1343 -240
rect 1377 -274 1411 -240
rect 1445 -274 1479 -240
rect 1513 -274 1547 -240
rect 1581 -274 1615 -240
rect 1649 -274 1763 -240
<< viali >>
rect -1457 138 -1423 172
rect -1265 138 -1231 172
rect -1073 138 -1039 172
rect -881 138 -847 172
rect -689 138 -655 172
rect -497 138 -463 172
rect -305 138 -271 172
rect -113 138 -79 172
rect 79 138 113 172
rect 271 138 305 172
rect 463 138 497 172
rect 655 138 689 172
rect 847 138 881 172
rect 1039 138 1073 172
rect 1231 138 1265 172
rect 1423 138 1457 172
<< metal1 >>
rect -1469 172 -1411 178
rect -1469 138 -1457 172
rect -1423 138 -1411 172
rect -1469 132 -1411 138
rect -1277 172 -1219 178
rect -1277 138 -1265 172
rect -1231 138 -1219 172
rect -1277 132 -1219 138
rect -1085 172 -1027 178
rect -1085 138 -1073 172
rect -1039 138 -1027 172
rect -1085 132 -1027 138
rect -893 172 -835 178
rect -893 138 -881 172
rect -847 138 -835 172
rect -893 132 -835 138
rect -701 172 -643 178
rect -701 138 -689 172
rect -655 138 -643 172
rect -701 132 -643 138
rect -509 172 -451 178
rect -509 138 -497 172
rect -463 138 -451 172
rect -509 132 -451 138
rect -317 172 -259 178
rect -317 138 -305 172
rect -271 138 -259 172
rect -317 132 -259 138
rect -125 172 -67 178
rect -125 138 -113 172
rect -79 138 -67 172
rect -125 132 -67 138
rect 67 172 125 178
rect 67 138 79 172
rect 113 138 125 172
rect 67 132 125 138
rect 259 172 317 178
rect 259 138 271 172
rect 305 138 317 172
rect 259 132 317 138
rect 451 172 509 178
rect 451 138 463 172
rect 497 138 509 172
rect 451 132 509 138
rect 643 172 701 178
rect 643 138 655 172
rect 689 138 701 172
rect 643 132 701 138
rect 835 172 893 178
rect 835 138 847 172
rect 881 138 893 172
rect 835 132 893 138
rect 1027 172 1085 178
rect 1027 138 1039 172
rect 1073 138 1085 172
rect 1027 132 1085 138
rect 1219 172 1277 178
rect 1219 138 1231 172
rect 1265 138 1277 172
rect 1219 132 1277 138
rect 1411 172 1469 178
rect 1411 138 1423 172
rect 1457 138 1469 172
rect 1411 132 1469 138
<< properties >>
string FIXED_BBOX -1746 -256 1746 256
<< end >>
