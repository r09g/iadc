magic
tech sky130A
magscale 1 2
timestamp 1654598415
<< pwell >>
rect -646 -262 648 200
<< nmos >>
rect -446 -52 -416 52
rect -350 -52 -320 52
rect -254 -52 -224 52
rect -158 -52 -128 52
rect -62 -52 -32 52
rect 34 -52 64 52
rect 130 -52 160 52
rect 226 -52 256 52
rect 322 -52 352 52
rect 418 -52 448 52
<< ndiff >>
rect -508 40 -446 52
rect -508 -40 -496 40
rect -462 -40 -446 40
rect -508 -52 -446 -40
rect -416 40 -350 52
rect -416 -40 -400 40
rect -366 -40 -350 40
rect -416 -52 -350 -40
rect -320 40 -254 52
rect -320 -40 -304 40
rect -270 -40 -254 40
rect -320 -52 -254 -40
rect -224 40 -158 52
rect -224 -40 -208 40
rect -174 -40 -158 40
rect -224 -52 -158 -40
rect -128 40 -62 52
rect -128 -40 -112 40
rect -78 -40 -62 40
rect -128 -52 -62 -40
rect -32 40 34 52
rect -32 -40 -16 40
rect 18 -40 34 40
rect -32 -52 34 -40
rect 64 40 130 52
rect 64 -40 80 40
rect 114 -40 130 40
rect 64 -52 130 -40
rect 160 40 226 52
rect 160 -40 176 40
rect 210 -40 226 40
rect 160 -52 226 -40
rect 256 40 322 52
rect 256 -40 272 40
rect 306 -40 322 40
rect 256 -52 322 -40
rect 352 40 418 52
rect 352 -40 368 40
rect 402 -40 418 40
rect 352 -52 418 -40
rect 448 40 510 52
rect 448 -40 464 40
rect 498 -40 510 40
rect 448 -52 510 -40
<< ndiffc >>
rect -496 -40 -462 40
rect -400 -40 -366 40
rect -304 -40 -270 40
rect -208 -40 -174 40
rect -112 -40 -78 40
rect -16 -40 18 40
rect 80 -40 114 40
rect 176 -40 210 40
rect 272 -40 306 40
rect 368 -40 402 40
rect 464 -40 498 40
<< psubdiff >>
rect -610 130 -514 164
rect 516 130 612 164
rect -610 68 -576 130
rect 578 68 612 130
rect -610 -192 -576 -130
rect 578 -192 612 -130
rect -610 -226 -514 -192
rect 516 -226 612 -192
<< psubdiffcont >>
rect -514 130 516 164
rect -610 -130 -576 68
rect 578 -130 612 68
rect -514 -226 516 -192
<< poly >>
rect -446 52 -416 78
rect -350 52 -320 78
rect -254 52 -224 78
rect -158 52 -128 78
rect -62 52 -32 78
rect 34 52 64 78
rect 130 52 160 78
rect 226 52 256 78
rect 322 52 352 78
rect 418 52 448 78
rect -446 -83 -416 -52
rect -350 -83 -320 -52
rect -254 -83 -224 -52
rect -158 -83 -128 -52
rect -62 -83 -32 -52
rect 34 -83 64 -52
rect 130 -83 160 -52
rect 226 -83 256 -52
rect 322 -83 352 -52
rect 418 -83 448 -52
rect -512 -99 514 -83
rect -512 -133 -496 -99
rect -462 -133 -304 -99
rect -270 -133 -112 -99
rect -78 -133 80 -99
rect 114 -133 272 -99
rect 306 -133 464 -99
rect 498 -133 514 -99
rect -512 -149 514 -133
<< polycont >>
rect -496 -133 -462 -99
rect -304 -133 -270 -99
rect -112 -133 -78 -99
rect 80 -133 114 -99
rect 272 -133 306 -99
rect 464 -133 498 -99
<< locali >>
rect -610 130 -514 164
rect 516 130 612 164
rect -610 68 -576 130
rect 578 68 612 130
rect -496 40 -462 56
rect -496 -56 -462 -40
rect -400 40 -366 56
rect -400 -56 -366 -40
rect -304 40 -270 56
rect -304 -56 -270 -40
rect -208 40 -174 56
rect -208 -56 -174 -40
rect -112 40 -78 56
rect -112 -56 -78 -40
rect -16 40 18 56
rect -16 -56 18 -40
rect 80 40 114 56
rect 80 -56 114 -40
rect 176 40 210 56
rect 176 -56 210 -40
rect 272 40 306 56
rect 272 -56 306 -40
rect 368 40 402 56
rect 368 -56 402 -40
rect 464 40 498 56
rect 464 -56 498 -40
rect -610 -192 -576 -130
rect -512 -99 514 -91
rect -512 -133 -496 -99
rect -462 -133 -304 -99
rect -270 -133 -112 -99
rect -78 -133 80 -99
rect 114 -133 272 -99
rect 306 -133 464 -99
rect 498 -133 514 -99
rect -512 -141 514 -133
rect 578 -192 612 -130
rect -610 -226 -514 -192
rect 516 -226 612 -192
<< viali >>
rect -496 -40 -462 40
rect -400 -40 -366 40
rect -304 -40 -270 40
rect -208 -40 -174 40
rect -112 -40 -78 40
rect -16 -40 18 40
rect 80 -40 114 40
rect 176 -40 210 40
rect 272 -40 306 40
rect 368 -40 402 40
rect 464 -40 498 40
<< metal1 >>
rect -502 40 -456 52
rect -502 -40 -496 40
rect -462 -40 -456 40
rect -502 -52 -456 -40
rect -406 40 -360 52
rect -406 -40 -400 40
rect -366 -40 -360 40
rect -406 -52 -360 -40
rect -310 40 -264 52
rect -310 -40 -304 40
rect -270 -40 -264 40
rect -310 -52 -264 -40
rect -214 40 -168 52
rect -214 -40 -208 40
rect -174 -40 -168 40
rect -214 -52 -168 -40
rect -118 40 -72 52
rect -118 -40 -112 40
rect -78 -40 -72 40
rect -118 -52 -72 -40
rect -22 40 24 52
rect -22 -40 -16 40
rect 18 -40 24 40
rect -22 -52 24 -40
rect 74 40 120 52
rect 74 -40 80 40
rect 114 -40 120 40
rect 74 -52 120 -40
rect 170 40 216 52
rect 170 -40 176 40
rect 210 -40 216 40
rect 170 -52 216 -40
rect 266 40 312 52
rect 266 -40 272 40
rect 306 -40 312 40
rect 266 -52 312 -40
rect 362 40 408 52
rect 362 -40 368 40
rect 402 -40 408 40
rect 362 -52 408 -40
rect 458 40 504 52
rect 458 -40 464 40
rect 498 -40 504 40
rect 458 -52 504 -40
<< properties >>
string FIXED_BBOX -594 -210 594 210
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.53 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
