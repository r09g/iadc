magic
tech sky130A
magscale 1 2
timestamp 1654899744
<< nwell >>
rect -3152 6932 -2673 8059
rect 1443 8056 2009 8212
rect -3154 6887 -2673 6932
rect 6080 6889 6614 8059
rect -3693 5999 -3238 6015
rect -3788 5636 -3150 5999
rect -3788 5635 -3668 5636
rect -3250 5635 -3150 5636
rect -3291 5573 -3213 5619
rect -3304 3617 -3219 3663
rect 6700 5999 7155 6015
rect 6612 5636 7250 5999
rect 6612 5635 6712 5636
rect 7130 5635 7250 5636
rect 6675 5573 6753 5619
rect 6681 3617 6766 3663
<< pwell >>
rect 1230 9436 1385 10632
rect 1203 9003 1385 9436
rect 1203 8939 1393 9003
rect 1203 8242 1385 8939
rect 2067 8242 2249 10632
rect -2789 -193 6262 6567
<< psubdiff >>
rect -2744 6497 -2648 6531
rect 6130 6497 6226 6531
rect -2744 6435 -2710 6497
rect -2744 4697 -2710 4759
rect 6192 6435 6226 6497
rect 6192 4697 6226 4759
rect -2744 4663 -2648 4697
rect 6130 4663 6226 4697
rect -2744 4242 -2648 4276
rect 6130 4242 6226 4276
rect -2744 4180 -2710 4242
rect -2744 682 -2710 745
rect 6192 4180 6226 4242
rect 6192 682 6226 745
rect -2744 648 -2647 682
rect 6129 648 6226 682
<< psubdiffcont >>
rect -2648 6497 6130 6531
rect -2744 4759 -2710 6435
rect 6192 4759 6226 6435
rect -2648 4663 6130 4697
rect -2648 4242 6130 4276
rect -2744 745 -2710 4180
rect 6192 745 6226 4180
rect -2647 648 6129 682
<< locali >>
rect -2744 6497 -2648 6531
rect 6130 6497 6226 6531
rect -2744 6435 -2710 6497
rect 6192 6435 6226 6497
rect 6076 6395 6192 6429
rect -2710 6085 -2596 6119
rect 6076 5955 6192 5989
rect -2710 5649 -2596 5683
rect 6076 5515 6192 5549
rect -2710 5205 -2596 5239
rect 6076 5075 6192 5109
rect -2710 4765 -2596 4799
rect -2744 4697 -2710 4759
rect 6192 4697 6226 4759
rect -2744 4663 -2648 4697
rect 6130 4663 6226 4697
rect -2744 4242 -2648 4276
rect 6130 4242 6226 4276
rect -2744 4180 -2710 4242
rect 6192 4180 6226 4242
rect 6076 4140 6192 4174
rect -2710 3830 -2596 3864
rect 6076 3700 6192 3734
rect -2324 3458 -2290 3474
rect -2210 3458 -2176 3474
rect -2114 3458 -2080 3474
rect -2000 3458 -1966 3474
rect -1904 3458 -1870 3474
rect -1790 3458 -1756 3474
rect -1694 3458 -1660 3474
rect -1580 3458 -1546 3474
rect -1484 3458 -1450 3474
rect -1370 3458 -1336 3474
rect -1274 3458 -1240 3474
rect -1160 3458 -1126 3474
rect -1064 3458 -1030 3474
rect -950 3458 -916 3474
rect -854 3458 -820 3474
rect -740 3458 -706 3474
rect -644 3458 -610 3474
rect -530 3458 -496 3474
rect -434 3458 -400 3474
rect -320 3458 -286 3474
rect -224 3458 -190 3474
rect -110 3458 -76 3474
rect -14 3458 20 3474
rect 100 3458 134 3474
rect 196 3458 230 3474
rect 310 3458 344 3474
rect 406 3458 440 3474
rect 520 3458 554 3474
rect 616 3458 650 3474
rect 730 3458 764 3474
rect 826 3458 860 3474
rect 940 3458 974 3474
rect 1036 3458 1070 3474
rect 1150 3458 1184 3474
rect 1246 3458 1280 3474
rect 1360 3458 1394 3474
rect 1456 3458 1490 3474
rect 1570 3458 1604 3474
rect 1666 3458 1700 3474
rect 1780 3458 1814 3474
rect 1876 3458 1910 3474
rect 1990 3458 2024 3474
rect 2086 3458 2120 3474
rect 2200 3458 2234 3474
rect 2296 3458 2330 3474
rect 2410 3458 2444 3474
rect 2506 3458 2540 3474
rect 2620 3458 2654 3474
rect 2716 3458 2750 3474
rect 2830 3458 2864 3474
rect 2926 3458 2960 3474
rect 3040 3458 3074 3474
rect 3136 3458 3170 3474
rect 3250 3458 3284 3474
rect 3346 3458 3380 3474
rect 3460 3458 3494 3474
rect 3556 3458 3590 3474
rect 3670 3458 3704 3474
rect 3766 3458 3800 3474
rect 3880 3458 3914 3474
rect 3976 3458 4010 3474
rect 4090 3458 4124 3474
rect 4186 3458 4220 3474
rect 4300 3458 4334 3474
rect 4396 3458 4430 3474
rect 4510 3458 4544 3474
rect 4606 3458 4640 3474
rect 4720 3458 4754 3474
rect 4816 3458 4850 3474
rect 4930 3458 4964 3474
rect 5026 3458 5060 3474
rect 5140 3458 5174 3474
rect 5236 3458 5270 3474
rect 5350 3458 5384 3474
rect 5446 3458 5480 3474
rect 5560 3458 5594 3474
rect 5656 3458 5690 3474
rect 5770 3458 5804 3474
rect 5866 3458 5900 3474
rect -2710 3390 -2595 3424
rect 6076 3260 6192 3294
rect -2324 3018 -2290 3034
rect -2210 3018 -2176 3034
rect -2114 3018 -2080 3034
rect -2000 3018 -1966 3034
rect -1904 3018 -1870 3034
rect -1790 3018 -1756 3034
rect -1694 3018 -1660 3034
rect -1580 3018 -1546 3034
rect -1484 3018 -1450 3034
rect -1370 3018 -1336 3034
rect -1274 3018 -1240 3034
rect -1160 3018 -1126 3034
rect -1064 3018 -1030 3034
rect -950 3018 -916 3034
rect -854 3018 -820 3034
rect -740 3018 -706 3034
rect -644 3018 -610 3034
rect -530 3018 -496 3034
rect -434 3018 -400 3034
rect -320 3018 -286 3034
rect -224 3018 -190 3034
rect -110 3018 -76 3034
rect -14 3018 20 3034
rect 100 3018 134 3034
rect 196 3018 230 3034
rect 310 3018 344 3034
rect 406 3018 440 3034
rect 520 3018 554 3034
rect 616 3018 650 3034
rect 730 3018 764 3034
rect 826 3018 860 3034
rect 940 3018 974 3034
rect 1036 3018 1070 3034
rect 1150 3018 1184 3034
rect 1246 3018 1280 3034
rect 1360 3018 1394 3034
rect 1456 3018 1490 3034
rect 1570 3018 1604 3034
rect 1666 3018 1700 3034
rect 1780 3018 1814 3034
rect 1876 3018 1910 3034
rect 1990 3018 2024 3034
rect 2086 3018 2120 3034
rect 2200 3018 2234 3034
rect 2296 3018 2330 3034
rect 2410 3018 2444 3034
rect 2506 3018 2540 3034
rect 2620 3018 2654 3034
rect 2716 3018 2750 3034
rect 2830 3018 2864 3034
rect 2926 3018 2960 3034
rect 3040 3018 3074 3034
rect 3136 3018 3170 3034
rect 3250 3018 3284 3034
rect 3346 3018 3380 3034
rect 3460 3018 3494 3034
rect 3556 3018 3590 3034
rect 3670 3018 3704 3034
rect 3766 3018 3800 3034
rect 3880 3018 3914 3034
rect 3976 3018 4010 3034
rect 4090 3018 4124 3034
rect 4186 3018 4220 3034
rect 4300 3018 4334 3034
rect 4396 3018 4430 3034
rect 4510 3018 4544 3034
rect 4606 3018 4640 3034
rect 4720 3018 4754 3034
rect 4816 3018 4850 3034
rect 4930 3018 4964 3034
rect 5026 3018 5060 3034
rect 5140 3018 5174 3034
rect 5236 3018 5270 3034
rect 5350 3018 5384 3034
rect 5446 3018 5480 3034
rect 5560 3018 5594 3034
rect 5656 3018 5690 3034
rect 5770 3018 5804 3034
rect 5866 3018 5900 3034
rect -2710 2950 -2596 2984
rect 6076 2820 6192 2854
rect -2324 2578 -2290 2594
rect -2210 2578 -2176 2594
rect -2114 2578 -2080 2594
rect -2000 2578 -1966 2594
rect -1904 2578 -1870 2594
rect -1790 2578 -1756 2594
rect -1694 2578 -1660 2594
rect -1580 2578 -1546 2594
rect -1484 2578 -1450 2594
rect -1370 2578 -1336 2594
rect -1274 2578 -1240 2594
rect -1160 2578 -1126 2594
rect -1064 2578 -1030 2594
rect -950 2578 -916 2594
rect -854 2578 -820 2594
rect -740 2578 -706 2594
rect -644 2578 -610 2594
rect -530 2578 -496 2594
rect -434 2578 -400 2594
rect -320 2578 -286 2594
rect -224 2578 -190 2594
rect -110 2578 -76 2594
rect -14 2578 20 2594
rect 100 2578 134 2594
rect 196 2578 230 2594
rect 310 2578 344 2594
rect 406 2578 440 2594
rect 520 2578 554 2594
rect 616 2578 650 2594
rect 730 2578 764 2594
rect 826 2578 860 2594
rect 940 2578 974 2594
rect 1036 2578 1070 2594
rect 1150 2578 1184 2594
rect 1246 2578 1280 2594
rect 1360 2578 1394 2594
rect 1456 2578 1490 2594
rect 1570 2578 1604 2594
rect 1666 2578 1700 2594
rect 1780 2578 1814 2594
rect 1876 2578 1910 2594
rect 1990 2578 2024 2594
rect 2086 2578 2120 2594
rect 2200 2578 2234 2594
rect 2296 2578 2330 2594
rect 2410 2578 2444 2594
rect 2506 2578 2540 2594
rect 2620 2578 2654 2594
rect 2716 2578 2750 2594
rect 2830 2578 2864 2594
rect 2926 2578 2960 2594
rect 3040 2578 3074 2594
rect 3136 2578 3170 2594
rect 3250 2578 3284 2594
rect 3346 2578 3380 2594
rect 3460 2578 3494 2594
rect 3556 2578 3590 2594
rect 3670 2578 3704 2594
rect 3766 2578 3800 2594
rect 3880 2578 3914 2594
rect 3976 2578 4010 2594
rect 4090 2578 4124 2594
rect 4186 2578 4220 2594
rect 4300 2578 4334 2594
rect 4396 2578 4430 2594
rect 4510 2578 4544 2594
rect 4606 2578 4640 2594
rect 4720 2578 4754 2594
rect 4816 2578 4850 2594
rect 4930 2578 4964 2594
rect 5026 2578 5060 2594
rect 5140 2578 5174 2594
rect 5236 2578 5270 2594
rect 5350 2578 5384 2594
rect 5446 2578 5480 2594
rect 5560 2578 5594 2594
rect 5656 2578 5690 2594
rect 5770 2578 5804 2594
rect 5866 2578 5900 2594
rect -2710 2510 -2596 2544
rect 6076 2380 6192 2414
rect -2324 2138 -2290 2154
rect -2210 2138 -2176 2154
rect -2114 2138 -2080 2154
rect -2000 2138 -1966 2154
rect -1904 2138 -1870 2154
rect -1790 2138 -1756 2154
rect -1694 2138 -1660 2154
rect -1580 2138 -1546 2154
rect -1484 2138 -1450 2154
rect -1370 2138 -1336 2154
rect -1274 2138 -1240 2154
rect -1160 2138 -1126 2154
rect -1064 2138 -1030 2154
rect -950 2138 -916 2154
rect -854 2138 -820 2154
rect -740 2138 -706 2154
rect -644 2138 -610 2154
rect -530 2138 -496 2154
rect -434 2138 -400 2154
rect -320 2138 -286 2154
rect -224 2138 -190 2154
rect -110 2138 -76 2154
rect -14 2138 20 2154
rect 100 2138 134 2154
rect 196 2138 230 2154
rect 310 2138 344 2154
rect 406 2138 440 2154
rect 520 2138 554 2154
rect 616 2138 650 2154
rect 730 2138 764 2154
rect 826 2138 860 2154
rect 940 2138 974 2154
rect 1036 2138 1070 2154
rect 1150 2138 1184 2154
rect 1246 2138 1280 2154
rect 1360 2138 1394 2154
rect 1456 2138 1490 2154
rect 1570 2138 1604 2154
rect 1666 2138 1700 2154
rect 1780 2138 1814 2154
rect 1876 2138 1910 2154
rect 1990 2138 2024 2154
rect 2086 2138 2120 2154
rect 2200 2138 2234 2154
rect 2296 2138 2330 2154
rect 2410 2138 2444 2154
rect 2506 2138 2540 2154
rect 2620 2138 2654 2154
rect 2716 2138 2750 2154
rect 2830 2138 2864 2154
rect 2926 2138 2960 2154
rect 3040 2138 3074 2154
rect 3136 2138 3170 2154
rect 3250 2138 3284 2154
rect 3346 2138 3380 2154
rect 3460 2138 3494 2154
rect 3556 2138 3590 2154
rect 3670 2138 3704 2154
rect 3766 2138 3800 2154
rect 3880 2138 3914 2154
rect 3976 2138 4010 2154
rect 4090 2138 4124 2154
rect 4186 2138 4220 2154
rect 4300 2138 4334 2154
rect 4396 2138 4430 2154
rect 4510 2138 4544 2154
rect 4606 2138 4640 2154
rect 4720 2138 4754 2154
rect 4816 2138 4850 2154
rect 4930 2138 4964 2154
rect 5026 2138 5060 2154
rect 5140 2138 5174 2154
rect 5236 2138 5270 2154
rect 5350 2138 5384 2154
rect 5446 2138 5480 2154
rect 5560 2138 5594 2154
rect 5656 2138 5690 2154
rect 5770 2138 5804 2154
rect 5866 2138 5900 2154
rect -2710 2070 -2596 2104
rect 6076 1940 6192 1974
rect -2324 1698 -2290 1714
rect -2210 1698 -2176 1714
rect -2114 1698 -2080 1714
rect -2000 1698 -1966 1714
rect -1904 1698 -1870 1714
rect -1790 1698 -1756 1714
rect -1694 1698 -1660 1714
rect -1580 1698 -1546 1714
rect -1484 1698 -1450 1714
rect -1370 1698 -1336 1714
rect -1274 1698 -1240 1714
rect -1160 1698 -1126 1714
rect -1064 1698 -1030 1714
rect -950 1698 -916 1714
rect -854 1698 -820 1714
rect -740 1698 -706 1714
rect -644 1698 -610 1714
rect -530 1698 -496 1714
rect -434 1698 -400 1714
rect -320 1698 -286 1714
rect -224 1698 -190 1714
rect -110 1698 -76 1714
rect -14 1698 20 1714
rect 100 1698 134 1714
rect 196 1698 230 1714
rect 310 1698 344 1714
rect 406 1698 440 1714
rect 520 1698 554 1714
rect 616 1698 650 1714
rect 730 1698 764 1714
rect 826 1698 860 1714
rect 940 1698 974 1714
rect 1036 1698 1070 1714
rect 1150 1698 1184 1714
rect 1246 1698 1280 1714
rect 1360 1698 1394 1714
rect 1456 1698 1490 1714
rect 1570 1698 1604 1714
rect 1666 1698 1700 1714
rect 1780 1698 1814 1714
rect 1876 1698 1910 1714
rect 1990 1698 2024 1714
rect 2086 1698 2120 1714
rect 2200 1698 2234 1714
rect 2296 1698 2330 1714
rect 2410 1698 2444 1714
rect 2506 1698 2540 1714
rect 2620 1698 2654 1714
rect 2716 1698 2750 1714
rect 2830 1698 2864 1714
rect 2926 1698 2960 1714
rect 3040 1698 3074 1714
rect 3136 1698 3170 1714
rect 3250 1698 3284 1714
rect 3346 1698 3380 1714
rect 3460 1698 3494 1714
rect 3556 1698 3590 1714
rect 3670 1698 3704 1714
rect 3766 1698 3800 1714
rect 3880 1698 3914 1714
rect 3976 1698 4010 1714
rect 4090 1698 4124 1714
rect 4186 1698 4220 1714
rect 4300 1698 4334 1714
rect 4396 1698 4430 1714
rect 4510 1698 4544 1714
rect 4606 1698 4640 1714
rect 4720 1698 4754 1714
rect 4816 1698 4850 1714
rect 4930 1698 4964 1714
rect 5026 1698 5060 1714
rect 5140 1698 5174 1714
rect 5236 1698 5270 1714
rect 5350 1698 5384 1714
rect 5446 1698 5480 1714
rect 5560 1698 5594 1714
rect 5656 1698 5690 1714
rect 5770 1698 5804 1714
rect 5866 1698 5900 1714
rect -2710 1630 -2596 1664
rect 6076 1500 6192 1534
rect -2324 1258 -2290 1274
rect -2210 1258 -2176 1274
rect -2114 1258 -2080 1274
rect -2000 1258 -1966 1274
rect -1904 1258 -1870 1274
rect -1790 1258 -1756 1274
rect -1694 1258 -1660 1274
rect -1580 1258 -1546 1274
rect -1484 1258 -1450 1274
rect -1370 1258 -1336 1274
rect -1274 1258 -1240 1274
rect -1160 1258 -1126 1274
rect -1064 1258 -1030 1274
rect -950 1258 -916 1274
rect -854 1258 -820 1274
rect -740 1258 -706 1274
rect -644 1258 -610 1274
rect -530 1258 -496 1274
rect -434 1258 -400 1274
rect -320 1258 -286 1274
rect -224 1258 -190 1274
rect -110 1258 -76 1274
rect -14 1258 20 1274
rect 100 1258 134 1274
rect 196 1258 230 1274
rect 310 1258 344 1274
rect 406 1258 440 1274
rect 520 1258 554 1274
rect 616 1258 650 1274
rect 730 1258 764 1274
rect 826 1258 860 1274
rect 940 1258 974 1274
rect 1036 1258 1070 1274
rect 1150 1258 1184 1274
rect 1246 1258 1280 1274
rect 1360 1258 1394 1274
rect 1456 1258 1490 1274
rect 1570 1258 1604 1274
rect 1666 1258 1700 1274
rect 1780 1258 1814 1274
rect 1876 1258 1910 1274
rect 1990 1258 2024 1274
rect 2086 1258 2120 1274
rect 2200 1258 2234 1274
rect 2296 1258 2330 1274
rect 2410 1258 2444 1274
rect 2506 1258 2540 1274
rect 2620 1258 2654 1274
rect 2716 1258 2750 1274
rect 2830 1258 2864 1274
rect 2926 1258 2960 1274
rect 3040 1258 3074 1274
rect 3136 1258 3170 1274
rect 3250 1258 3284 1274
rect 3346 1258 3380 1274
rect 3460 1258 3494 1274
rect 3556 1258 3590 1274
rect 3670 1258 3704 1274
rect 3766 1258 3800 1274
rect 3880 1258 3914 1274
rect 3976 1258 4010 1274
rect 4090 1258 4124 1274
rect 4186 1258 4220 1274
rect 4300 1258 4334 1274
rect 4396 1258 4430 1274
rect 4510 1258 4544 1274
rect 4606 1258 4640 1274
rect 4720 1258 4754 1274
rect 4816 1258 4850 1274
rect 4930 1258 4964 1274
rect 5026 1258 5060 1274
rect 5140 1258 5174 1274
rect 5236 1258 5270 1274
rect 5350 1258 5384 1274
rect 5446 1258 5480 1274
rect 5560 1258 5594 1274
rect 5656 1258 5690 1274
rect 5770 1258 5804 1274
rect 5866 1258 5900 1274
rect -2710 1190 -2593 1224
rect 6076 1059 6192 1093
rect -2324 818 -2290 834
rect -2210 818 -2176 834
rect -2114 818 -2080 834
rect -2000 818 -1966 834
rect -1904 818 -1870 834
rect -1790 818 -1756 834
rect -1694 818 -1660 834
rect -1580 818 -1546 834
rect -1484 818 -1450 834
rect -1370 818 -1336 834
rect -1274 818 -1240 834
rect -1160 818 -1126 834
rect -1064 818 -1030 834
rect -950 818 -916 834
rect -854 818 -820 834
rect -740 818 -706 834
rect -644 818 -610 834
rect -530 818 -496 834
rect -434 818 -400 834
rect -320 818 -286 834
rect -224 818 -190 834
rect -110 818 -76 834
rect -14 818 20 834
rect 100 818 134 834
rect 196 818 230 834
rect 310 818 344 834
rect 406 818 440 834
rect 520 818 554 834
rect 616 818 650 834
rect 730 818 764 834
rect 826 818 860 834
rect 940 818 974 834
rect 1036 818 1070 834
rect 1150 818 1184 834
rect 1246 818 1280 834
rect 1360 818 1394 834
rect 1456 818 1490 834
rect 1570 818 1604 834
rect 1666 818 1700 834
rect 1780 818 1814 834
rect 1876 818 1910 834
rect 1990 818 2024 834
rect 2086 818 2120 834
rect 2200 818 2234 834
rect 2296 818 2330 834
rect 2410 818 2444 834
rect 2506 818 2540 834
rect 2620 818 2654 834
rect 2716 818 2750 834
rect 2830 818 2864 834
rect 2926 818 2960 834
rect 3040 818 3074 834
rect 3136 818 3170 834
rect 3250 818 3284 834
rect 3346 818 3380 834
rect 3460 818 3494 834
rect 3556 818 3590 834
rect 3670 818 3704 834
rect 3766 818 3800 834
rect 3880 818 3914 834
rect 3976 818 4010 834
rect 4090 818 4124 834
rect 4186 818 4220 834
rect 4300 818 4334 834
rect 4396 818 4430 834
rect 4510 818 4544 834
rect 4606 818 4640 834
rect 4720 818 4754 834
rect 4816 818 4850 834
rect 4930 818 4964 834
rect 5026 818 5060 834
rect 5140 818 5174 834
rect 5236 818 5270 834
rect 5350 818 5384 834
rect 5446 818 5480 834
rect 5560 818 5594 834
rect 5656 818 5690 834
rect 5770 818 5804 834
rect 5866 818 5900 834
rect -2710 750 -2596 784
rect -2744 682 -2710 745
rect 6192 682 6226 745
rect -2744 648 -2647 682
rect 6129 648 6226 682
rect 282 -123 316 14
rect 474 -123 508 14
rect 666 -123 700 14
rect 858 -123 892 14
rect 1050 -123 1084 14
rect 1242 -123 1276 14
rect 1434 -123 1468 14
rect 1626 -123 1660 14
rect 1818 -123 1852 14
rect 2010 -123 2044 14
rect 2202 -123 2236 14
rect 2394 -123 2428 14
rect 2586 -123 2620 14
rect 2778 -123 2812 14
rect 2970 -123 3004 14
rect 3162 -123 3196 14
<< viali >>
rect 1404 9322 1438 9356
rect 2016 9330 2050 9364
rect 1404 9231 1438 9265
rect 2015 9224 2049 9258
rect 1317 8955 1351 8989
rect 1403 8955 1437 8989
rect 1497 8948 1531 8982
rect 1599 8948 1633 8982
rect 1820 8948 1854 8982
rect 1921 8948 1955 8982
rect 2016 8955 2050 8989
rect 2102 8955 2136 8989
rect 1404 8746 1438 8780
rect 2012 8745 2046 8779
rect 1404 8660 1438 8694
rect 2012 8659 2046 8693
rect 1306 8463 1341 8498
rect 1518 8463 1552 8497
rect 1898 8462 1932 8496
rect 2109 8462 2144 8497
rect 1397 8278 1431 8312
rect 2022 8279 2056 8313
rect -3656 7989 -3282 8023
rect -2662 7989 6114 8023
rect 6744 7989 7118 8023
rect -3415 7779 -3381 7813
rect -2434 7794 -2400 7828
rect -2224 7794 -2190 7828
rect -2014 7794 -1980 7828
rect -1804 7794 -1770 7828
rect -1594 7794 -1560 7828
rect -1384 7794 -1350 7828
rect -1174 7794 -1140 7828
rect -964 7794 -930 7828
rect -754 7794 -720 7828
rect -544 7794 -510 7828
rect -334 7794 -300 7828
rect -124 7794 -90 7828
rect 86 7794 120 7828
rect 296 7794 330 7828
rect 506 7794 540 7828
rect 716 7794 750 7828
rect 926 7794 960 7828
rect 1136 7794 1170 7828
rect 1346 7794 1380 7828
rect 1556 7794 1590 7828
rect 1766 7794 1800 7828
rect 1976 7794 2010 7828
rect 2186 7794 2220 7828
rect 2396 7794 2430 7828
rect 2606 7794 2640 7828
rect 2816 7794 2850 7828
rect 3026 7794 3060 7828
rect 3236 7794 3270 7828
rect 3446 7794 3480 7828
rect 3656 7794 3690 7828
rect 3866 7794 3900 7828
rect 4076 7794 4110 7828
rect 4286 7794 4320 7828
rect 4496 7794 4530 7828
rect 4706 7794 4740 7828
rect 4916 7794 4950 7828
rect 5126 7794 5160 7828
rect 5336 7794 5370 7828
rect 5546 7794 5580 7828
rect 5756 7794 5790 7828
rect 6843 7779 6877 7813
rect -3557 7683 -3523 7717
rect -2338 7652 -2304 7686
rect -2128 7652 -2094 7686
rect -1918 7652 -1884 7686
rect -1708 7652 -1674 7686
rect -1498 7652 -1464 7686
rect -1288 7652 -1254 7686
rect -1078 7652 -1044 7686
rect -868 7652 -834 7686
rect -658 7652 -624 7686
rect -448 7652 -414 7686
rect -238 7652 -204 7686
rect -28 7652 6 7686
rect 182 7652 216 7686
rect 392 7652 426 7686
rect 602 7652 636 7686
rect 812 7652 846 7686
rect 1022 7652 1056 7686
rect 1232 7652 1266 7686
rect 1442 7652 1476 7686
rect 1652 7652 1686 7686
rect 1862 7652 1896 7686
rect 2072 7652 2106 7686
rect 2282 7652 2316 7686
rect 2492 7652 2526 7686
rect 2702 7652 2736 7686
rect 2912 7652 2946 7686
rect 3122 7652 3156 7686
rect 3332 7652 3366 7686
rect 3542 7652 3576 7686
rect 3752 7652 3786 7686
rect 3962 7652 3996 7686
rect 4172 7652 4206 7686
rect 4382 7652 4416 7686
rect 4592 7652 4626 7686
rect 4802 7652 4836 7686
rect 5012 7652 5046 7686
rect 5222 7652 5256 7686
rect 5432 7652 5466 7686
rect 5642 7652 5676 7686
rect 5852 7652 5886 7686
rect 6985 7683 7019 7717
rect -3415 7587 -3381 7621
rect 6843 7587 6877 7621
rect -3557 7491 -3523 7525
rect 6985 7491 7019 7525
rect -3415 7395 -3381 7429
rect 6843 7395 6877 7429
rect -3557 7299 -3523 7333
rect 6985 7299 7019 7333
rect -2432 7262 -2398 7296
rect -2222 7262 -2188 7296
rect -2012 7262 -1978 7296
rect -1802 7262 -1768 7296
rect -1592 7262 -1558 7296
rect -1382 7262 -1348 7296
rect -1172 7262 -1138 7296
rect -962 7262 -928 7296
rect -752 7262 -718 7296
rect -542 7262 -508 7296
rect -332 7262 -298 7296
rect -122 7262 -88 7296
rect 88 7262 122 7296
rect 298 7262 332 7296
rect 508 7262 542 7296
rect 718 7262 752 7296
rect 928 7262 962 7296
rect 1138 7262 1172 7296
rect 1348 7262 1382 7296
rect 1558 7262 1592 7296
rect 1768 7262 1802 7296
rect 1978 7262 2012 7296
rect 2188 7262 2222 7296
rect 2398 7262 2432 7296
rect 2608 7262 2642 7296
rect 2818 7262 2852 7296
rect 3028 7262 3062 7296
rect 3238 7262 3272 7296
rect 3448 7262 3482 7296
rect 3658 7262 3692 7296
rect 3868 7262 3902 7296
rect 4078 7262 4112 7296
rect 4288 7262 4322 7296
rect 4498 7262 4532 7296
rect 4708 7262 4742 7296
rect 4918 7262 4952 7296
rect 5128 7262 5162 7296
rect 5338 7262 5372 7296
rect 5548 7262 5582 7296
rect 5758 7262 5792 7296
rect -3415 7203 -3381 7237
rect 6843 7203 6877 7237
rect -3557 7107 -3523 7141
rect -2336 7120 -2302 7154
rect -2126 7120 -2092 7154
rect -1916 7120 -1882 7154
rect -1706 7120 -1672 7154
rect -1496 7120 -1462 7154
rect -1286 7120 -1252 7154
rect -1076 7120 -1042 7154
rect -866 7120 -832 7154
rect -656 7120 -622 7154
rect -446 7120 -412 7154
rect -236 7120 -202 7154
rect -26 7120 8 7154
rect 184 7120 218 7154
rect 394 7120 428 7154
rect 604 7120 638 7154
rect 814 7120 848 7154
rect 1024 7120 1058 7154
rect 1234 7120 1268 7154
rect 1444 7120 1478 7154
rect 1654 7120 1688 7154
rect 1864 7120 1898 7154
rect 2074 7120 2108 7154
rect 2284 7120 2318 7154
rect 2494 7120 2528 7154
rect 2704 7120 2738 7154
rect 2914 7120 2948 7154
rect 3124 7120 3158 7154
rect 3334 7120 3368 7154
rect 3544 7120 3578 7154
rect 3754 7120 3788 7154
rect 3964 7120 3998 7154
rect 4174 7120 4208 7154
rect 4384 7120 4418 7154
rect 4594 7120 4628 7154
rect 4804 7120 4838 7154
rect 5014 7120 5048 7154
rect 5224 7120 5258 7154
rect 5434 7120 5468 7154
rect 5644 7120 5678 7154
rect 5854 7120 5888 7154
rect 6985 7107 7019 7141
rect -3415 7011 -3381 7045
rect 6843 7011 6877 7045
rect -3557 6915 -3523 6949
rect 6985 6915 7019 6949
rect -3415 6819 -3381 6853
rect 6843 6819 6877 6853
rect -3557 6723 -3523 6757
rect 6985 6723 7019 6757
rect -3415 6627 -3381 6661
rect 6843 6627 6877 6661
rect -3557 6531 -3523 6565
rect 6985 6531 7019 6565
rect -3415 6435 -3381 6469
rect -3557 6339 -3523 6373
rect -3415 6243 -3381 6277
rect -3656 6033 -3282 6067
rect -3656 5579 -3282 5613
rect -3415 5369 -3381 5403
rect -3557 5273 -3523 5307
rect -3415 5177 -3381 5211
rect -3557 5081 -3523 5115
rect -3415 4985 -3381 5019
rect -3557 4889 -3523 4923
rect -3415 4793 -3381 4827
rect -2744 4759 -2710 6435
rect 6843 6435 6877 6469
rect -3557 4697 -3523 4731
rect 6192 4759 6226 6435
rect 6985 6339 7019 6373
rect 6843 6243 6877 6277
rect 6744 6033 7118 6067
rect 6744 5579 7118 5613
rect 6843 5369 6877 5403
rect 6985 5273 7019 5307
rect 6843 5177 6877 5211
rect 6985 5081 7019 5115
rect 6843 4985 6877 5019
rect 6985 4889 7019 4923
rect 6843 4793 6877 4827
rect 6985 4697 7019 4731
rect -3415 4601 -3381 4635
rect 6843 4601 6877 4635
rect -3557 4505 -3523 4539
rect 6985 4505 7019 4539
rect -3415 4409 -3381 4443
rect 6843 4409 6877 4443
rect -3557 4313 -3523 4347
rect 6985 4313 7019 4347
rect -3415 4217 -3381 4251
rect -3557 4121 -3523 4155
rect -3415 4025 -3381 4059
rect -3557 3929 -3523 3963
rect -3415 3833 -3381 3867
rect -3656 3623 -3282 3657
rect -2744 745 -2710 4180
rect 6843 4217 6877 4251
rect -2420 4056 -2386 4090
rect -2210 4056 -2176 4090
rect -2000 4056 -1966 4090
rect -1790 4056 -1756 4090
rect -1580 4056 -1546 4090
rect -1370 4056 -1336 4090
rect -1160 4056 -1126 4090
rect -950 4056 -916 4090
rect -740 4056 -706 4090
rect -530 4056 -496 4090
rect -320 4056 -286 4090
rect -110 4056 -76 4090
rect 100 4056 134 4090
rect 310 4056 344 4090
rect 520 4056 554 4090
rect 730 4056 764 4090
rect 940 4056 974 4090
rect 1150 4056 1184 4090
rect 1360 4056 1394 4090
rect 1570 4056 1604 4090
rect 1780 4056 1814 4090
rect 1990 4056 2024 4090
rect 2200 4056 2234 4090
rect 2410 4056 2444 4090
rect 2620 4056 2654 4090
rect 2830 4056 2864 4090
rect 3040 4056 3074 4090
rect 3250 4056 3284 4090
rect 3460 4056 3494 4090
rect 3670 4056 3704 4090
rect 3880 4056 3914 4090
rect 4090 4056 4124 4090
rect 4300 4056 4334 4090
rect 4510 4056 4544 4090
rect 4720 4056 4754 4090
rect 4930 4056 4964 4090
rect 5140 4056 5174 4090
rect 5350 4056 5384 4090
rect 5560 4056 5594 4090
rect 5770 4056 5804 4090
rect -2324 3914 -2290 3948
rect -2114 3914 -2080 3948
rect -1904 3914 -1870 3948
rect -1694 3914 -1660 3948
rect -1484 3914 -1450 3948
rect -1274 3914 -1240 3948
rect -1064 3914 -1030 3948
rect -854 3914 -820 3948
rect -644 3914 -610 3948
rect -434 3914 -400 3948
rect -224 3914 -190 3948
rect -14 3914 20 3948
rect 196 3914 230 3948
rect 406 3914 440 3948
rect 616 3914 650 3948
rect 826 3914 860 3948
rect 1036 3914 1070 3948
rect 1246 3914 1280 3948
rect 1456 3914 1490 3948
rect 1666 3914 1700 3948
rect 1876 3914 1910 3948
rect 2086 3914 2120 3948
rect 2296 3914 2330 3948
rect 2506 3914 2540 3948
rect 2716 3914 2750 3948
rect 2926 3914 2960 3948
rect 3136 3914 3170 3948
rect 3346 3914 3380 3948
rect 3556 3914 3590 3948
rect 3766 3914 3800 3948
rect 3976 3914 4010 3948
rect 4186 3914 4220 3948
rect 4396 3914 4430 3948
rect 4606 3914 4640 3948
rect 4816 3914 4850 3948
rect 5026 3914 5060 3948
rect 5236 3914 5270 3948
rect 5446 3914 5480 3948
rect 5656 3914 5690 3948
rect 5866 3914 5900 3948
rect -2420 3616 -2386 3650
rect -2210 3616 -2176 3650
rect -2000 3616 -1966 3650
rect -1790 3616 -1756 3650
rect -1580 3616 -1546 3650
rect -1370 3616 -1336 3650
rect -1160 3616 -1126 3650
rect -950 3616 -916 3650
rect -740 3616 -706 3650
rect -530 3616 -496 3650
rect -320 3616 -286 3650
rect -110 3616 -76 3650
rect 100 3616 134 3650
rect 310 3616 344 3650
rect 520 3616 554 3650
rect 730 3616 764 3650
rect 940 3616 974 3650
rect 1150 3616 1184 3650
rect 1360 3616 1394 3650
rect 1570 3616 1604 3650
rect 1780 3616 1814 3650
rect 1990 3616 2024 3650
rect 2200 3616 2234 3650
rect 2410 3616 2444 3650
rect 2620 3616 2654 3650
rect 2830 3616 2864 3650
rect 3040 3616 3074 3650
rect 3250 3616 3284 3650
rect 3460 3616 3494 3650
rect 3670 3616 3704 3650
rect 3880 3616 3914 3650
rect 4090 3616 4124 3650
rect 4300 3616 4334 3650
rect 4510 3616 4544 3650
rect 4720 3616 4754 3650
rect 4930 3616 4964 3650
rect 5140 3616 5174 3650
rect 5350 3616 5384 3650
rect 5560 3616 5594 3650
rect 5770 3616 5804 3650
rect -2324 3474 -2290 3508
rect -2114 3474 -2080 3508
rect -1904 3474 -1870 3508
rect -1694 3474 -1660 3508
rect -1484 3474 -1450 3508
rect -1274 3474 -1240 3508
rect -1064 3474 -1030 3508
rect -854 3474 -820 3508
rect -644 3474 -610 3508
rect -434 3474 -400 3508
rect -224 3474 -190 3508
rect -14 3474 20 3508
rect 196 3474 230 3508
rect 406 3474 440 3508
rect 616 3474 650 3508
rect 826 3474 860 3508
rect 1036 3474 1070 3508
rect 1246 3474 1280 3508
rect 1456 3474 1490 3508
rect 1666 3474 1700 3508
rect 1876 3474 1910 3508
rect 2086 3474 2120 3508
rect 2296 3474 2330 3508
rect 2506 3474 2540 3508
rect 2716 3474 2750 3508
rect 2926 3474 2960 3508
rect 3136 3474 3170 3508
rect 3346 3474 3380 3508
rect 3556 3474 3590 3508
rect 3766 3474 3800 3508
rect 3976 3474 4010 3508
rect 4186 3474 4220 3508
rect 4396 3474 4430 3508
rect 4606 3474 4640 3508
rect 4816 3474 4850 3508
rect 5026 3474 5060 3508
rect 5236 3474 5270 3508
rect 5446 3474 5480 3508
rect 5656 3474 5690 3508
rect 5866 3474 5900 3508
rect -2420 3176 -2386 3210
rect -2210 3176 -2176 3210
rect -2000 3176 -1966 3210
rect -1790 3176 -1756 3210
rect -1580 3176 -1546 3210
rect -1370 3176 -1336 3210
rect -1160 3176 -1126 3210
rect -950 3176 -916 3210
rect -740 3176 -706 3210
rect -530 3176 -496 3210
rect -320 3176 -286 3210
rect -110 3176 -76 3210
rect 100 3176 134 3210
rect 310 3176 344 3210
rect 520 3176 554 3210
rect 730 3176 764 3210
rect 940 3176 974 3210
rect 1150 3176 1184 3210
rect 1360 3176 1394 3210
rect 1570 3176 1604 3210
rect 1780 3176 1814 3210
rect 1990 3176 2024 3210
rect 2200 3176 2234 3210
rect 2410 3176 2444 3210
rect 2620 3176 2654 3210
rect 2830 3176 2864 3210
rect 3040 3176 3074 3210
rect 3250 3176 3284 3210
rect 3460 3176 3494 3210
rect 3670 3176 3704 3210
rect 3880 3176 3914 3210
rect 4090 3176 4124 3210
rect 4300 3176 4334 3210
rect 4510 3176 4544 3210
rect 4720 3176 4754 3210
rect 4930 3176 4964 3210
rect 5140 3176 5174 3210
rect 5350 3176 5384 3210
rect 5560 3176 5594 3210
rect 5770 3176 5804 3210
rect -2324 3034 -2290 3068
rect -2114 3034 -2080 3068
rect -1904 3034 -1870 3068
rect -1694 3034 -1660 3068
rect -1484 3034 -1450 3068
rect -1274 3034 -1240 3068
rect -1064 3034 -1030 3068
rect -854 3034 -820 3068
rect -644 3034 -610 3068
rect -434 3034 -400 3068
rect -224 3034 -190 3068
rect -14 3034 20 3068
rect 196 3034 230 3068
rect 406 3034 440 3068
rect 616 3034 650 3068
rect 826 3034 860 3068
rect 1036 3034 1070 3068
rect 1246 3034 1280 3068
rect 1456 3034 1490 3068
rect 1666 3034 1700 3068
rect 1876 3034 1910 3068
rect 2086 3034 2120 3068
rect 2296 3034 2330 3068
rect 2506 3034 2540 3068
rect 2716 3034 2750 3068
rect 2926 3034 2960 3068
rect 3136 3034 3170 3068
rect 3346 3034 3380 3068
rect 3556 3034 3590 3068
rect 3766 3034 3800 3068
rect 3976 3034 4010 3068
rect 4186 3034 4220 3068
rect 4396 3034 4430 3068
rect 4606 3034 4640 3068
rect 4816 3034 4850 3068
rect 5026 3034 5060 3068
rect 5236 3034 5270 3068
rect 5446 3034 5480 3068
rect 5656 3034 5690 3068
rect 5866 3034 5900 3068
rect -2420 2736 -2386 2770
rect -2210 2736 -2176 2770
rect -2000 2736 -1966 2770
rect -1790 2736 -1756 2770
rect -1580 2736 -1546 2770
rect -1370 2736 -1336 2770
rect -1160 2736 -1126 2770
rect -950 2736 -916 2770
rect -740 2736 -706 2770
rect -530 2736 -496 2770
rect -320 2736 -286 2770
rect -110 2736 -76 2770
rect 100 2736 134 2770
rect 310 2736 344 2770
rect 520 2736 554 2770
rect 730 2736 764 2770
rect 940 2736 974 2770
rect 1150 2736 1184 2770
rect 1360 2736 1394 2770
rect 1570 2736 1604 2770
rect 1780 2736 1814 2770
rect 1990 2736 2024 2770
rect 2200 2736 2234 2770
rect 2410 2736 2444 2770
rect 2620 2736 2654 2770
rect 2830 2736 2864 2770
rect 3040 2736 3074 2770
rect 3250 2736 3284 2770
rect 3460 2736 3494 2770
rect 3670 2736 3704 2770
rect 3880 2736 3914 2770
rect 4090 2736 4124 2770
rect 4300 2736 4334 2770
rect 4510 2736 4544 2770
rect 4720 2736 4754 2770
rect 4930 2736 4964 2770
rect 5140 2736 5174 2770
rect 5350 2736 5384 2770
rect 5560 2736 5594 2770
rect 5770 2736 5804 2770
rect -2324 2594 -2290 2628
rect -2114 2594 -2080 2628
rect -1904 2594 -1870 2628
rect -1694 2594 -1660 2628
rect -1484 2594 -1450 2628
rect -1274 2594 -1240 2628
rect -1064 2594 -1030 2628
rect -854 2594 -820 2628
rect -644 2594 -610 2628
rect -434 2594 -400 2628
rect -224 2594 -190 2628
rect -14 2594 20 2628
rect 196 2594 230 2628
rect 406 2594 440 2628
rect 616 2594 650 2628
rect 826 2594 860 2628
rect 1036 2594 1070 2628
rect 1246 2594 1280 2628
rect 1456 2594 1490 2628
rect 1666 2594 1700 2628
rect 1876 2594 1910 2628
rect 2086 2594 2120 2628
rect 2296 2594 2330 2628
rect 2506 2594 2540 2628
rect 2716 2594 2750 2628
rect 2926 2594 2960 2628
rect 3136 2594 3170 2628
rect 3346 2594 3380 2628
rect 3556 2594 3590 2628
rect 3766 2594 3800 2628
rect 3976 2594 4010 2628
rect 4186 2594 4220 2628
rect 4396 2594 4430 2628
rect 4606 2594 4640 2628
rect 4816 2594 4850 2628
rect 5026 2594 5060 2628
rect 5236 2594 5270 2628
rect 5446 2594 5480 2628
rect 5656 2594 5690 2628
rect 5866 2594 5900 2628
rect -2420 2296 -2386 2330
rect -2210 2296 -2176 2330
rect -2000 2296 -1966 2330
rect -1790 2296 -1756 2330
rect -1580 2296 -1546 2330
rect -1370 2296 -1336 2330
rect -1160 2296 -1126 2330
rect -950 2296 -916 2330
rect -740 2296 -706 2330
rect -530 2296 -496 2330
rect -320 2296 -286 2330
rect -110 2296 -76 2330
rect 100 2296 134 2330
rect 310 2296 344 2330
rect 520 2296 554 2330
rect 730 2296 764 2330
rect 940 2296 974 2330
rect 1150 2296 1184 2330
rect 1360 2296 1394 2330
rect 1570 2296 1604 2330
rect 1780 2296 1814 2330
rect 1990 2296 2024 2330
rect 2200 2296 2234 2330
rect 2410 2296 2444 2330
rect 2620 2296 2654 2330
rect 2830 2296 2864 2330
rect 3040 2296 3074 2330
rect 3250 2296 3284 2330
rect 3460 2296 3494 2330
rect 3670 2296 3704 2330
rect 3880 2296 3914 2330
rect 4090 2296 4124 2330
rect 4300 2296 4334 2330
rect 4510 2296 4544 2330
rect 4720 2296 4754 2330
rect 4930 2296 4964 2330
rect 5140 2296 5174 2330
rect 5350 2296 5384 2330
rect 5560 2296 5594 2330
rect 5770 2296 5804 2330
rect -2324 2154 -2290 2188
rect -2114 2154 -2080 2188
rect -1904 2154 -1870 2188
rect -1694 2154 -1660 2188
rect -1484 2154 -1450 2188
rect -1274 2154 -1240 2188
rect -1064 2154 -1030 2188
rect -854 2154 -820 2188
rect -644 2154 -610 2188
rect -434 2154 -400 2188
rect -224 2154 -190 2188
rect -14 2154 20 2188
rect 196 2154 230 2188
rect 406 2154 440 2188
rect 616 2154 650 2188
rect 826 2154 860 2188
rect 1036 2154 1070 2188
rect 1246 2154 1280 2188
rect 1456 2154 1490 2188
rect 1666 2154 1700 2188
rect 1876 2154 1910 2188
rect 2086 2154 2120 2188
rect 2296 2154 2330 2188
rect 2506 2154 2540 2188
rect 2716 2154 2750 2188
rect 2926 2154 2960 2188
rect 3136 2154 3170 2188
rect 3346 2154 3380 2188
rect 3556 2154 3590 2188
rect 3766 2154 3800 2188
rect 3976 2154 4010 2188
rect 4186 2154 4220 2188
rect 4396 2154 4430 2188
rect 4606 2154 4640 2188
rect 4816 2154 4850 2188
rect 5026 2154 5060 2188
rect 5236 2154 5270 2188
rect 5446 2154 5480 2188
rect 5656 2154 5690 2188
rect 5866 2154 5900 2188
rect -2420 1856 -2386 1890
rect -2210 1856 -2176 1890
rect -2000 1856 -1966 1890
rect -1790 1856 -1756 1890
rect -1580 1856 -1546 1890
rect -1370 1856 -1336 1890
rect -1160 1856 -1126 1890
rect -950 1856 -916 1890
rect -740 1856 -706 1890
rect -530 1856 -496 1890
rect -320 1856 -286 1890
rect -110 1856 -76 1890
rect 100 1856 134 1890
rect 310 1856 344 1890
rect 520 1856 554 1890
rect 730 1856 764 1890
rect 940 1856 974 1890
rect 1150 1856 1184 1890
rect 1360 1856 1394 1890
rect 1570 1856 1604 1890
rect 1780 1856 1814 1890
rect 1990 1856 2024 1890
rect 2200 1856 2234 1890
rect 2410 1856 2444 1890
rect 2620 1856 2654 1890
rect 2830 1856 2864 1890
rect 3040 1856 3074 1890
rect 3250 1856 3284 1890
rect 3460 1856 3494 1890
rect 3670 1856 3704 1890
rect 3880 1856 3914 1890
rect 4090 1856 4124 1890
rect 4300 1856 4334 1890
rect 4510 1856 4544 1890
rect 4720 1856 4754 1890
rect 4930 1856 4964 1890
rect 5140 1856 5174 1890
rect 5350 1856 5384 1890
rect 5560 1856 5594 1890
rect 5770 1856 5804 1890
rect -2324 1714 -2290 1748
rect -2114 1714 -2080 1748
rect -1904 1714 -1870 1748
rect -1694 1714 -1660 1748
rect -1484 1714 -1450 1748
rect -1274 1714 -1240 1748
rect -1064 1714 -1030 1748
rect -854 1714 -820 1748
rect -644 1714 -610 1748
rect -434 1714 -400 1748
rect -224 1714 -190 1748
rect -14 1714 20 1748
rect 196 1714 230 1748
rect 406 1714 440 1748
rect 616 1714 650 1748
rect 826 1714 860 1748
rect 1036 1714 1070 1748
rect 1246 1714 1280 1748
rect 1456 1714 1490 1748
rect 1666 1714 1700 1748
rect 1876 1714 1910 1748
rect 2086 1714 2120 1748
rect 2296 1714 2330 1748
rect 2506 1714 2540 1748
rect 2716 1714 2750 1748
rect 2926 1714 2960 1748
rect 3136 1714 3170 1748
rect 3346 1714 3380 1748
rect 3556 1714 3590 1748
rect 3766 1714 3800 1748
rect 3976 1714 4010 1748
rect 4186 1714 4220 1748
rect 4396 1714 4430 1748
rect 4606 1714 4640 1748
rect 4816 1714 4850 1748
rect 5026 1714 5060 1748
rect 5236 1714 5270 1748
rect 5446 1714 5480 1748
rect 5656 1714 5690 1748
rect 5866 1714 5900 1748
rect -2420 1416 -2386 1450
rect -2210 1416 -2176 1450
rect -2000 1416 -1966 1450
rect -1790 1416 -1756 1450
rect -1580 1416 -1546 1450
rect -1370 1416 -1336 1450
rect -1160 1416 -1126 1450
rect -950 1416 -916 1450
rect -740 1416 -706 1450
rect -530 1416 -496 1450
rect -320 1416 -286 1450
rect -110 1416 -76 1450
rect 100 1416 134 1450
rect 310 1416 344 1450
rect 520 1416 554 1450
rect 730 1416 764 1450
rect 940 1416 974 1450
rect 1150 1416 1184 1450
rect 1360 1416 1394 1450
rect 1570 1416 1604 1450
rect 1780 1416 1814 1450
rect 1990 1416 2024 1450
rect 2200 1416 2234 1450
rect 2410 1416 2444 1450
rect 2620 1416 2654 1450
rect 2830 1416 2864 1450
rect 3040 1416 3074 1450
rect 3250 1416 3284 1450
rect 3460 1416 3494 1450
rect 3670 1416 3704 1450
rect 3880 1416 3914 1450
rect 4090 1416 4124 1450
rect 4300 1416 4334 1450
rect 4510 1416 4544 1450
rect 4720 1416 4754 1450
rect 4930 1416 4964 1450
rect 5140 1416 5174 1450
rect 5350 1416 5384 1450
rect 5560 1416 5594 1450
rect 5770 1416 5804 1450
rect -2324 1274 -2290 1308
rect -2114 1274 -2080 1308
rect -1904 1274 -1870 1308
rect -1694 1274 -1660 1308
rect -1484 1274 -1450 1308
rect -1274 1274 -1240 1308
rect -1064 1274 -1030 1308
rect -854 1274 -820 1308
rect -644 1274 -610 1308
rect -434 1274 -400 1308
rect -224 1274 -190 1308
rect -14 1274 20 1308
rect 196 1274 230 1308
rect 406 1274 440 1308
rect 616 1274 650 1308
rect 826 1274 860 1308
rect 1036 1274 1070 1308
rect 1246 1274 1280 1308
rect 1456 1274 1490 1308
rect 1666 1274 1700 1308
rect 1876 1274 1910 1308
rect 2086 1274 2120 1308
rect 2296 1274 2330 1308
rect 2506 1274 2540 1308
rect 2716 1274 2750 1308
rect 2926 1274 2960 1308
rect 3136 1274 3170 1308
rect 3346 1274 3380 1308
rect 3556 1274 3590 1308
rect 3766 1274 3800 1308
rect 3976 1274 4010 1308
rect 4186 1274 4220 1308
rect 4396 1274 4430 1308
rect 4606 1274 4640 1308
rect 4816 1274 4850 1308
rect 5026 1274 5060 1308
rect 5236 1274 5270 1308
rect 5446 1274 5480 1308
rect 5656 1274 5690 1308
rect 5866 1274 5900 1308
rect -2420 976 -2386 1010
rect -2210 976 -2176 1010
rect -2000 976 -1966 1010
rect -1790 976 -1756 1010
rect -1580 976 -1546 1010
rect -1370 976 -1336 1010
rect -1160 976 -1126 1010
rect -950 976 -916 1010
rect -740 976 -706 1010
rect -530 976 -496 1010
rect -320 976 -286 1010
rect -110 976 -76 1010
rect 100 976 134 1010
rect 310 976 344 1010
rect 520 976 554 1010
rect 730 976 764 1010
rect 940 976 974 1010
rect 1150 976 1184 1010
rect 1360 976 1394 1010
rect 1570 976 1604 1010
rect 1780 976 1814 1010
rect 1990 976 2024 1010
rect 2200 976 2234 1010
rect 2410 976 2444 1010
rect 2620 976 2654 1010
rect 2830 976 2864 1010
rect 3040 976 3074 1010
rect 3250 976 3284 1010
rect 3460 976 3494 1010
rect 3670 976 3704 1010
rect 3880 976 3914 1010
rect 4090 976 4124 1010
rect 4300 976 4334 1010
rect 4510 976 4544 1010
rect 4720 976 4754 1010
rect 4930 976 4964 1010
rect 5140 976 5174 1010
rect 5350 976 5384 1010
rect 5560 976 5594 1010
rect 5770 976 5804 1010
rect -2324 834 -2290 868
rect -2114 834 -2080 868
rect -1904 834 -1870 868
rect -1694 834 -1660 868
rect -1484 834 -1450 868
rect -1274 834 -1240 868
rect -1064 834 -1030 868
rect -854 834 -820 868
rect -644 834 -610 868
rect -434 834 -400 868
rect -224 834 -190 868
rect -14 834 20 868
rect 196 834 230 868
rect 406 834 440 868
rect 616 834 650 868
rect 826 834 860 868
rect 1036 834 1070 868
rect 1246 834 1280 868
rect 1456 834 1490 868
rect 1666 834 1700 868
rect 1876 834 1910 868
rect 2086 834 2120 868
rect 2296 834 2330 868
rect 2506 834 2540 868
rect 2716 834 2750 868
rect 2926 834 2960 868
rect 3136 834 3170 868
rect 3346 834 3380 868
rect 3556 834 3590 868
rect 3766 834 3800 868
rect 3976 834 4010 868
rect 4186 834 4220 868
rect 4396 834 4430 868
rect 4606 834 4640 868
rect 4816 834 4850 868
rect 5026 834 5060 868
rect 5236 834 5270 868
rect 5446 834 5480 868
rect 5656 834 5690 868
rect 5866 834 5900 868
rect 6192 745 6226 4180
rect 6985 4121 7019 4155
rect 6843 4025 6877 4059
rect 6985 3929 7019 3963
rect 6843 3833 6877 3867
rect 6744 3623 7118 3657
rect 186 171 220 205
rect 378 171 412 205
rect 570 171 604 205
rect 762 171 796 205
rect 954 171 988 205
rect 1146 171 1180 205
rect 1338 171 1372 205
rect 1530 171 1564 205
rect 1722 171 1756 205
rect 1914 171 1948 205
rect 2106 171 2140 205
rect 2298 171 2332 205
rect 2490 171 2524 205
rect 2682 171 2716 205
rect 2874 171 2908 205
rect 3066 171 3100 205
rect 3258 171 3292 205
rect 282 29 316 63
rect 474 29 508 63
rect 666 29 700 63
rect 858 29 892 63
rect 1050 29 1084 63
rect 1242 29 1276 63
rect 1434 29 1468 63
rect 1626 29 1660 63
rect 1818 29 1852 63
rect 2010 29 2044 63
rect 2202 29 2236 63
rect 2394 29 2428 63
rect 2586 29 2620 63
rect 2778 29 2812 63
rect 2970 29 3004 63
rect 3162 29 3196 63
rect 72 -157 3406 -123
<< metal1 >>
rect 1134 9790 1230 10729
rect 1134 9738 1156 9790
rect 1208 9738 1230 9790
rect 1134 9649 1230 9738
rect 1134 9597 1156 9649
rect 1208 9597 1230 9649
rect 1134 9508 1230 9597
rect 1134 9456 1156 9508
rect 1208 9456 1230 9508
rect 1134 9367 1230 9456
rect 1134 9315 1156 9367
rect 1208 9315 1230 9367
rect 1134 9226 1230 9315
rect 1134 9174 1156 9226
rect 1208 9174 1230 9226
rect 1134 8241 1230 9174
rect 1317 8995 1351 10729
rect 1397 9362 1449 9374
rect 1392 9356 1450 9362
rect 1392 9322 1404 9356
rect 1438 9322 1450 9356
rect 1392 9316 1450 9322
rect 1397 9271 1449 9316
rect 1392 9265 1450 9271
rect 1566 9268 1576 9320
rect 1628 9268 1638 9320
rect 1392 9231 1404 9265
rect 1438 9231 1450 9265
rect 1392 9225 1450 9231
rect 1397 9154 1449 9225
rect 1387 9102 1397 9154
rect 1449 9102 1459 9154
rect 1305 8989 1363 8995
rect 1391 8989 1449 8995
rect 1576 8991 1628 9268
rect 1305 8955 1317 8989
rect 1351 8955 1403 8989
rect 1437 8955 1449 8989
rect 1305 8949 1363 8955
rect 1391 8949 1449 8955
rect 1477 8939 1487 8991
rect 1539 8939 1576 8991
rect 1628 8988 1638 8991
rect 1628 8982 1645 8988
rect 1633 8948 1645 8982
rect 1628 8942 1645 8948
rect 1628 8939 1638 8942
rect 1392 8780 1450 8786
rect 1392 8746 1404 8780
rect 1438 8746 1450 8780
rect 1392 8740 1450 8746
rect 1403 8700 1438 8740
rect 1392 8694 1450 8700
rect 1392 8660 1404 8694
rect 1438 8660 1450 8694
rect 1392 8654 1450 8660
rect 1403 8505 1438 8654
rect 1294 8498 1564 8505
rect 1294 8463 1306 8498
rect 1341 8497 1564 8498
rect 1341 8470 1518 8497
rect 1341 8463 1353 8470
rect 1294 8457 1353 8463
rect 1506 8463 1518 8470
rect 1552 8463 1564 8497
rect 1506 8457 1564 8463
rect 1379 8270 1389 8322
rect 1441 8270 1451 8322
rect 1678 8131 1774 10729
rect 1993 9320 2003 9372
rect 2055 9320 2065 9372
rect 2003 9268 2055 9320
rect 1993 9216 2003 9268
rect 2055 9216 2065 9268
rect 1813 9102 1823 9154
rect 1875 9102 1885 9154
rect 1823 8991 1875 9102
rect 2102 8995 2136 10729
rect 2222 9792 2318 10729
rect 2222 9740 2244 9792
rect 2296 9740 2318 9792
rect 2222 9651 2318 9740
rect 2222 9599 2244 9651
rect 2296 9599 2318 9651
rect 2222 9510 2318 9599
rect 2222 9458 2244 9510
rect 2296 9458 2318 9510
rect 2222 9369 2318 9458
rect 2222 9317 2244 9369
rect 2296 9317 2318 9369
rect 2222 9228 2318 9317
rect 2222 9176 2244 9228
rect 2296 9176 2318 9228
rect 1813 8988 1823 8991
rect 1808 8982 1823 8988
rect 1808 8948 1820 8982
rect 1808 8942 1823 8948
rect 1813 8939 1823 8942
rect 1875 8939 1912 8991
rect 1964 8939 1974 8991
rect 2004 8989 2148 8995
rect 2004 8955 2016 8989
rect 2050 8955 2102 8989
rect 2136 8955 2148 8989
rect 2004 8949 2148 8955
rect 2000 8779 2058 8785
rect 2000 8745 2012 8779
rect 2046 8745 2058 8779
rect 2000 8739 2058 8745
rect 2012 8699 2047 8739
rect 2000 8693 2058 8699
rect 2000 8659 2012 8693
rect 2046 8659 2058 8693
rect 2000 8653 2058 8659
rect 2012 8504 2047 8653
rect 2222 8611 2318 9176
rect 2271 8578 2318 8611
rect 2230 8530 2254 8543
rect 2313 8530 2318 8578
rect 2230 8525 2318 8530
rect 1886 8497 2156 8504
rect 1886 8496 2109 8497
rect 1886 8462 1898 8496
rect 1932 8469 2109 8496
rect 1932 8462 1944 8469
rect 1886 8456 1944 8462
rect 2097 8462 2109 8469
rect 2144 8462 2156 8497
rect 2097 8456 2156 8462
rect 2003 8271 2013 8323
rect 2065 8271 2075 8323
rect 2222 8241 2318 8525
rect -3788 8041 7250 8131
rect -3788 8023 -1286 8041
rect -1234 8023 287 8041
rect 339 8023 3230 8041
rect 3282 8023 4699 8041
rect 4751 8023 7250 8041
rect -3788 7989 -3656 8023
rect -3282 7989 -2662 8023
rect 6114 7989 6744 8023
rect 7118 7989 7250 8023
rect -3788 7983 7250 7989
rect -3557 7723 -3523 7983
rect -3427 7813 -3369 7819
rect -3427 7779 -3415 7813
rect -3381 7779 -3369 7813
rect -3427 7773 -3369 7779
rect -3569 7717 -3511 7723
rect -3650 7581 -3616 7685
rect -3569 7683 -3557 7717
rect -3523 7683 -3511 7717
rect -3569 7677 -3511 7683
rect -3672 7529 -3662 7581
rect -3610 7529 -3600 7581
rect -3557 7531 -3523 7677
rect -3415 7627 -3381 7773
rect -3427 7621 -3369 7627
rect -3427 7587 -3415 7621
rect -3381 7587 -3369 7621
rect -3427 7581 -3369 7587
rect -3322 7581 -3288 7781
rect -3650 6431 -3616 7529
rect -3569 7525 -3511 7531
rect -3569 7491 -3557 7525
rect -3523 7491 -3511 7525
rect -3569 7485 -3511 7491
rect -3557 7339 -3523 7485
rect -3415 7435 -3381 7581
rect -3341 7529 -3331 7581
rect -3279 7529 -3269 7581
rect -3427 7429 -3369 7435
rect -3427 7395 -3415 7429
rect -3381 7395 -3369 7429
rect -3427 7389 -3369 7395
rect -3569 7333 -3511 7339
rect -3569 7299 -3557 7333
rect -3523 7299 -3511 7333
rect -3569 7293 -3511 7299
rect -3557 7147 -3523 7293
rect -3415 7243 -3381 7389
rect -3427 7237 -3369 7243
rect -3427 7203 -3415 7237
rect -3381 7203 -3369 7237
rect -3427 7197 -3369 7203
rect -3569 7141 -3511 7147
rect -3569 7107 -3557 7141
rect -3523 7107 -3511 7141
rect -3569 7101 -3511 7107
rect -3557 6955 -3523 7101
rect -3415 7051 -3381 7197
rect -3427 7045 -3369 7051
rect -3427 7011 -3415 7045
rect -3381 7011 -3369 7045
rect -3427 7005 -3369 7011
rect -3569 6949 -3511 6955
rect -3569 6915 -3557 6949
rect -3523 6915 -3511 6949
rect -3569 6909 -3511 6915
rect -3557 6763 -3523 6909
rect -3415 6859 -3381 7005
rect -3427 6853 -3369 6859
rect -3427 6819 -3415 6853
rect -3381 6819 -3369 6853
rect -3427 6813 -3369 6819
rect -3569 6757 -3511 6763
rect -3569 6723 -3557 6757
rect -3523 6723 -3511 6757
rect -3569 6717 -3511 6723
rect -3415 6720 -3381 6813
rect -3557 6571 -3523 6717
rect -3433 6668 -3423 6720
rect -3371 6668 -3361 6720
rect -3427 6661 -3369 6668
rect -3427 6627 -3415 6661
rect -3381 6627 -3369 6661
rect -3427 6621 -3369 6627
rect -3569 6565 -3511 6571
rect -3569 6531 -3557 6565
rect -3523 6531 -3511 6565
rect -3569 6525 -3511 6531
rect -3670 6379 -3660 6431
rect -3608 6379 -3598 6431
rect -3557 6379 -3523 6525
rect -3415 6475 -3381 6621
rect -3427 6469 -3369 6475
rect -3427 6435 -3415 6469
rect -3381 6435 -3369 6469
rect -3427 6429 -3369 6435
rect -3322 6431 -3288 7529
rect -3650 6275 -3616 6379
rect -3569 6373 -3511 6379
rect -3569 6339 -3557 6373
rect -3523 6339 -3511 6373
rect -3569 6333 -3511 6339
rect -3557 6073 -3523 6333
rect -3415 6283 -3381 6429
rect -3341 6379 -3331 6431
rect -3279 6379 -3269 6431
rect -3322 6371 -3288 6379
rect -3427 6277 -3369 6283
rect -3427 6243 -3415 6277
rect -3381 6243 -3369 6277
rect -3427 6237 -3369 6243
rect -3220 6073 -3150 7983
rect 1960 7921 1970 7930
rect -2446 7887 1970 7921
rect 1960 7878 1970 7887
rect 2022 7921 2032 7930
rect 2022 7887 5898 7921
rect 2022 7878 2032 7887
rect -2446 7828 -2388 7834
rect -2236 7828 -2178 7834
rect -2026 7828 -1968 7834
rect -1816 7828 -1758 7834
rect -1606 7828 -1548 7834
rect -1396 7828 -1338 7834
rect -1186 7828 -1128 7834
rect -976 7828 -918 7834
rect -766 7828 -708 7834
rect -556 7828 -498 7834
rect -346 7828 -288 7834
rect -136 7828 -78 7834
rect 74 7828 132 7834
rect 284 7828 342 7834
rect 494 7828 552 7834
rect 704 7828 762 7834
rect 914 7828 972 7834
rect 1124 7828 1182 7834
rect 1334 7828 1392 7834
rect 1544 7828 1602 7834
rect 1754 7828 1812 7834
rect 1964 7828 2022 7834
rect 2174 7828 2232 7834
rect 2384 7828 2442 7834
rect 2594 7828 2652 7834
rect 2804 7828 2862 7834
rect 3014 7828 3072 7834
rect 3224 7828 3282 7834
rect 3434 7828 3492 7834
rect 3644 7828 3702 7834
rect 3854 7828 3912 7834
rect 4064 7828 4122 7834
rect 4274 7828 4332 7834
rect 4484 7828 4542 7834
rect 4694 7828 4752 7834
rect 4904 7828 4962 7834
rect 5114 7828 5172 7834
rect 5324 7828 5382 7834
rect 5534 7828 5592 7834
rect 5744 7828 5802 7834
rect -2446 7794 -2434 7828
rect -2400 7794 -2224 7828
rect -2190 7794 -2014 7828
rect -1980 7794 -1804 7828
rect -1770 7794 -1594 7828
rect -1560 7794 -1384 7828
rect -1350 7794 -1286 7828
rect -2446 7788 -2388 7794
rect -2236 7788 -2178 7794
rect -2026 7788 -1968 7794
rect -1816 7788 -1758 7794
rect -1606 7788 -1548 7794
rect -1396 7788 -1338 7794
rect -1296 7776 -1286 7794
rect -1234 7794 -1174 7828
rect -1140 7794 -964 7828
rect -930 7794 -754 7828
rect -720 7794 -544 7828
rect -510 7794 -334 7828
rect -300 7794 -124 7828
rect -90 7794 86 7828
rect 120 7794 287 7828
rect 339 7794 506 7828
rect 540 7794 716 7828
rect 750 7794 926 7828
rect 960 7794 1136 7828
rect 1170 7794 1346 7828
rect 1380 7794 1556 7828
rect 1590 7794 1766 7828
rect 1800 7794 1976 7828
rect 2010 7794 2186 7828
rect 2220 7794 2396 7828
rect 2430 7794 2606 7828
rect 2640 7794 2816 7828
rect 2850 7794 3026 7828
rect 3060 7794 3230 7828
rect 3282 7794 3446 7828
rect 3480 7794 3656 7828
rect 3690 7794 3866 7828
rect 3900 7794 4076 7828
rect 4110 7794 4286 7828
rect 4320 7794 4496 7828
rect 4530 7794 4699 7828
rect 4751 7794 4916 7828
rect 4950 7794 5126 7828
rect 5160 7794 5336 7828
rect 5370 7794 5546 7828
rect 5580 7794 5756 7828
rect 5790 7794 5898 7828
rect -1234 7776 -1224 7794
rect -1186 7788 -1128 7794
rect -976 7788 -918 7794
rect -766 7788 -708 7794
rect -556 7788 -498 7794
rect -346 7788 -288 7794
rect -136 7788 -78 7794
rect 74 7788 132 7794
rect 277 7776 287 7794
rect 339 7776 349 7794
rect 494 7788 552 7794
rect 704 7788 762 7794
rect 914 7788 972 7794
rect 1124 7788 1182 7794
rect 1334 7788 1392 7794
rect 1544 7788 1602 7794
rect 1749 7776 1821 7794
rect 1964 7788 2022 7794
rect 2174 7788 2232 7794
rect 2384 7788 2442 7794
rect 2594 7788 2652 7794
rect 2804 7788 2862 7794
rect 3014 7788 3072 7794
rect 3220 7776 3230 7794
rect 3282 7776 3292 7794
rect 3434 7788 3492 7794
rect 3644 7788 3702 7794
rect 3854 7788 3912 7794
rect 4064 7788 4122 7794
rect 4274 7788 4332 7794
rect 4484 7788 4542 7794
rect 4689 7776 4699 7794
rect 4751 7776 4761 7794
rect 4904 7788 4962 7794
rect 5114 7788 5172 7794
rect 5324 7788 5382 7794
rect 5534 7788 5592 7794
rect 5744 7788 5802 7794
rect -2350 7686 -2292 7692
rect -2140 7686 -2082 7692
rect -1930 7686 -1872 7692
rect -1720 7686 -1662 7692
rect -1510 7686 -1452 7692
rect -1300 7686 -1242 7692
rect -1090 7686 -1032 7692
rect -880 7686 -822 7692
rect -670 7686 -612 7692
rect -460 7686 -402 7692
rect -250 7686 -192 7692
rect -40 7686 18 7692
rect 170 7686 228 7692
rect 380 7686 438 7692
rect 590 7686 648 7692
rect 800 7686 858 7692
rect 1010 7686 1068 7692
rect 1220 7686 1278 7692
rect 1430 7686 1488 7692
rect 1640 7686 1698 7692
rect 1850 7686 1908 7692
rect 2060 7686 2118 7692
rect 2270 7686 2328 7692
rect 2391 7686 2401 7704
rect -2446 7652 -2338 7686
rect -2304 7652 -2128 7686
rect -2094 7652 -1918 7686
rect -1884 7652 -1708 7686
rect -1674 7652 -1498 7686
rect -1464 7652 -1288 7686
rect -1254 7652 -1078 7686
rect -1044 7652 -868 7686
rect -834 7652 -658 7686
rect -624 7652 -448 7686
rect -414 7652 -238 7686
rect -204 7652 -28 7686
rect 6 7652 182 7686
rect 216 7652 392 7686
rect 426 7652 602 7686
rect 636 7652 812 7686
rect 846 7652 1022 7686
rect 1056 7652 1232 7686
rect 1266 7652 1442 7686
rect 1476 7652 1652 7686
rect 1686 7652 1862 7686
rect 1896 7652 2072 7686
rect 2106 7652 2282 7686
rect 2316 7652 2401 7686
rect 2453 7692 2463 7704
rect 2453 7686 2538 7692
rect 2690 7686 2748 7692
rect 2900 7686 2958 7692
rect 3110 7686 3168 7692
rect 3320 7686 3378 7692
rect 3530 7686 3588 7692
rect 3740 7686 3798 7692
rect 3861 7686 3871 7704
rect 2453 7652 2492 7686
rect 2526 7652 2702 7686
rect 2736 7652 2912 7686
rect 2946 7652 3122 7686
rect 3156 7652 3332 7686
rect 3366 7652 3542 7686
rect 3576 7652 3752 7686
rect 3786 7652 3871 7686
rect 3923 7692 3933 7704
rect 3923 7686 4008 7692
rect 4160 7686 4218 7692
rect 4370 7686 4428 7692
rect 4580 7686 4638 7692
rect 4790 7686 4848 7692
rect 5000 7686 5058 7692
rect 5210 7686 5268 7692
rect 5330 7686 5340 7704
rect 3923 7652 3962 7686
rect 3996 7652 4172 7686
rect 4206 7652 4382 7686
rect 4416 7652 4592 7686
rect 4626 7652 4802 7686
rect 4836 7652 5012 7686
rect 5046 7652 5222 7686
rect 5256 7652 5340 7686
rect 5392 7692 5402 7704
rect 5392 7686 5478 7692
rect 5630 7686 5688 7692
rect 5840 7686 5898 7692
rect 5392 7652 5432 7686
rect 5466 7652 5642 7686
rect 5676 7652 5852 7686
rect 5886 7652 5898 7686
rect -2350 7646 -2292 7652
rect -2140 7646 -2082 7652
rect -1930 7646 -1872 7652
rect -1720 7646 -1662 7652
rect -1510 7646 -1452 7652
rect -1300 7646 -1242 7652
rect -1090 7646 -1032 7652
rect -880 7646 -822 7652
rect -670 7646 -612 7652
rect -460 7646 -402 7652
rect -250 7646 -192 7652
rect -40 7646 18 7652
rect 170 7646 228 7652
rect 380 7646 438 7652
rect 590 7646 648 7652
rect 800 7646 858 7652
rect 1010 7646 1068 7652
rect 1220 7646 1278 7652
rect 1430 7646 1488 7652
rect 1640 7646 1698 7652
rect 1850 7646 1908 7652
rect 2060 7646 2118 7652
rect 2270 7646 2328 7652
rect 2480 7646 2538 7652
rect 2690 7646 2748 7652
rect 2900 7646 2958 7652
rect 3110 7646 3168 7652
rect 3320 7646 3378 7652
rect 3530 7646 3588 7652
rect 3740 7646 3798 7652
rect 3950 7646 4008 7652
rect 4160 7646 4218 7652
rect 4370 7646 4428 7652
rect 4580 7646 4638 7652
rect 4790 7646 4848 7652
rect 5000 7646 5058 7652
rect 5210 7646 5268 7652
rect 5420 7646 5478 7652
rect 5630 7646 5688 7652
rect 5840 7646 5898 7652
rect 1960 7593 1970 7602
rect -2444 7559 1970 7593
rect 1960 7550 1970 7559
rect 2022 7593 2032 7602
rect 2022 7559 5898 7593
rect 2022 7550 2032 7559
rect 1436 7389 1458 7400
rect -2444 7355 1458 7389
rect 1436 7349 1458 7355
rect 1448 7348 1458 7349
rect 1510 7389 1520 7400
rect 1510 7355 5900 7389
rect 1510 7348 1520 7355
rect -2444 7296 -2386 7302
rect -2234 7296 -2176 7302
rect -2024 7296 -1966 7302
rect -1814 7296 -1756 7302
rect -1604 7296 -1546 7302
rect -1394 7296 -1336 7302
rect -1184 7296 -1126 7302
rect -974 7296 -916 7302
rect -764 7296 -706 7302
rect -554 7296 -496 7302
rect -344 7296 -286 7302
rect -134 7296 -76 7302
rect 76 7296 134 7302
rect 286 7296 344 7302
rect 496 7296 554 7302
rect 706 7296 764 7302
rect 916 7296 974 7302
rect 1126 7296 1184 7302
rect 1336 7296 1394 7302
rect 1546 7296 1604 7302
rect 1756 7296 1814 7302
rect 1966 7296 2024 7302
rect 2176 7296 2234 7302
rect 2386 7296 2444 7302
rect 2596 7296 2654 7302
rect 2806 7296 2864 7302
rect 3016 7296 3074 7302
rect 3226 7296 3284 7302
rect 3436 7296 3494 7302
rect 3646 7296 3704 7302
rect 3856 7296 3914 7302
rect 4066 7296 4124 7302
rect 4276 7296 4334 7302
rect 4486 7296 4544 7302
rect 4696 7296 4754 7302
rect 4906 7296 4964 7302
rect 5116 7296 5174 7302
rect 5326 7296 5384 7302
rect 5536 7296 5594 7302
rect 5746 7296 5804 7302
rect -2444 7262 -2432 7296
rect -2398 7262 -2222 7296
rect -2188 7262 -2012 7296
rect -1978 7262 -1802 7296
rect -1768 7262 -1592 7296
rect -1558 7262 -1382 7296
rect -1348 7262 -1286 7296
rect -2444 7256 -2386 7262
rect -2234 7256 -2176 7262
rect -2024 7256 -1966 7262
rect -1814 7256 -1756 7262
rect -1604 7256 -1546 7262
rect -1394 7256 -1336 7262
rect -1296 7244 -1286 7262
rect -1234 7262 -1172 7296
rect -1138 7262 -962 7296
rect -928 7262 -752 7296
rect -718 7262 -542 7296
rect -508 7262 -332 7296
rect -298 7262 -122 7296
rect -88 7262 88 7296
rect 122 7262 287 7296
rect 339 7262 508 7296
rect 542 7262 718 7296
rect 752 7262 928 7296
rect 962 7262 1138 7296
rect 1172 7262 1348 7296
rect 1382 7262 1558 7296
rect 1592 7262 1768 7296
rect 1802 7262 1978 7296
rect 2012 7262 2188 7296
rect 2222 7262 2398 7296
rect 2432 7262 2608 7296
rect 2642 7262 2818 7296
rect 2852 7262 3028 7296
rect 3062 7262 3230 7296
rect 3282 7262 3448 7296
rect 3482 7262 3658 7296
rect 3692 7262 3868 7296
rect 3902 7262 4078 7296
rect 4112 7262 4288 7296
rect 4322 7262 4498 7296
rect 4532 7262 4699 7296
rect 4751 7262 4918 7296
rect 4952 7262 5128 7296
rect 5162 7262 5338 7296
rect 5372 7262 5548 7296
rect 5582 7262 5758 7296
rect 5792 7262 5900 7296
rect -1234 7244 -1224 7262
rect -1184 7256 -1126 7262
rect -974 7256 -916 7262
rect -764 7256 -706 7262
rect -554 7256 -496 7262
rect -344 7256 -286 7262
rect -134 7256 -76 7262
rect 76 7256 134 7262
rect 277 7244 287 7262
rect 339 7244 349 7262
rect 496 7256 554 7262
rect 706 7256 764 7262
rect 916 7256 974 7262
rect 1126 7256 1184 7262
rect 1336 7256 1394 7262
rect 1546 7256 1604 7262
rect 1749 7244 1821 7262
rect 1966 7256 2024 7262
rect 2176 7256 2234 7262
rect 2386 7256 2444 7262
rect 2596 7256 2654 7262
rect 2806 7256 2864 7262
rect 3016 7256 3074 7262
rect 3220 7244 3230 7262
rect 3282 7244 3292 7262
rect 3436 7256 3494 7262
rect 3646 7256 3704 7262
rect 3856 7256 3914 7262
rect 4066 7256 4124 7262
rect 4276 7256 4334 7262
rect 4486 7256 4544 7262
rect 4689 7244 4699 7262
rect 4751 7244 4761 7262
rect 4906 7256 4964 7262
rect 5116 7256 5174 7262
rect 5326 7256 5384 7262
rect 5536 7256 5594 7262
rect 5746 7256 5804 7262
rect -2348 7154 -2290 7160
rect -2138 7154 -2080 7160
rect -2019 7154 -2009 7172
rect -2444 7120 -2336 7154
rect -2302 7120 -2126 7154
rect -2092 7120 -2009 7154
rect -1957 7160 -1947 7172
rect -1957 7154 -1870 7160
rect -1718 7154 -1660 7160
rect -1508 7154 -1450 7160
rect -1298 7154 -1240 7160
rect -1088 7154 -1030 7160
rect -878 7154 -820 7160
rect -668 7154 -610 7160
rect -549 7154 -539 7172
rect -1957 7120 -1916 7154
rect -1882 7120 -1706 7154
rect -1672 7120 -1496 7154
rect -1462 7120 -1286 7154
rect -1252 7120 -1076 7154
rect -1042 7120 -866 7154
rect -832 7120 -656 7154
rect -622 7120 -539 7154
rect -487 7160 -477 7172
rect -487 7154 -400 7160
rect -248 7154 -190 7160
rect -38 7154 20 7160
rect 172 7154 230 7160
rect 382 7154 440 7160
rect 592 7154 650 7160
rect 802 7154 860 7160
rect 921 7154 931 7172
rect -487 7120 -446 7154
rect -412 7120 -236 7154
rect -202 7120 -26 7154
rect 8 7120 184 7154
rect 218 7120 394 7154
rect 428 7120 604 7154
rect 638 7120 814 7154
rect 848 7120 931 7154
rect 983 7160 993 7172
rect 983 7154 1070 7160
rect 1222 7154 1280 7160
rect 1432 7154 1490 7160
rect 1642 7154 1700 7160
rect 1852 7154 1910 7160
rect 2062 7154 2120 7160
rect 2272 7154 2330 7160
rect 2482 7154 2540 7160
rect 2692 7154 2750 7160
rect 2902 7154 2960 7160
rect 3112 7154 3170 7160
rect 3322 7154 3380 7160
rect 3532 7154 3590 7160
rect 3742 7154 3800 7160
rect 3952 7154 4010 7160
rect 4162 7154 4220 7160
rect 4372 7154 4430 7160
rect 4582 7154 4640 7160
rect 4792 7154 4850 7160
rect 5002 7154 5060 7160
rect 5212 7154 5270 7160
rect 5422 7154 5480 7160
rect 5632 7154 5690 7160
rect 5842 7154 5900 7160
rect 983 7120 1024 7154
rect 1058 7120 1234 7154
rect 1268 7120 1444 7154
rect 1478 7120 1654 7154
rect 1688 7120 1864 7154
rect 1898 7120 2074 7154
rect 2108 7120 2284 7154
rect 2318 7120 2494 7154
rect 2528 7120 2704 7154
rect 2738 7120 2914 7154
rect 2948 7120 3124 7154
rect 3158 7120 3334 7154
rect 3368 7120 3544 7154
rect 3578 7120 3754 7154
rect 3788 7120 3964 7154
rect 3998 7120 4174 7154
rect 4208 7120 4384 7154
rect 4418 7120 4594 7154
rect 4628 7120 4804 7154
rect 4838 7120 5014 7154
rect 5048 7120 5224 7154
rect 5258 7120 5434 7154
rect 5468 7120 5644 7154
rect 5678 7120 5854 7154
rect 5888 7120 5900 7154
rect -2348 7114 -2290 7120
rect -2138 7114 -2080 7120
rect -1928 7114 -1870 7120
rect -1718 7114 -1660 7120
rect -1508 7114 -1450 7120
rect -1298 7114 -1240 7120
rect -1088 7114 -1030 7120
rect -878 7114 -820 7120
rect -668 7114 -610 7120
rect -458 7114 -400 7120
rect -248 7114 -190 7120
rect -38 7114 20 7120
rect 172 7114 230 7120
rect 382 7114 440 7120
rect 592 7114 650 7120
rect 802 7114 860 7120
rect 1012 7114 1070 7120
rect 1222 7114 1280 7120
rect 1432 7114 1490 7120
rect 1642 7114 1700 7120
rect 1852 7114 1910 7120
rect 2062 7114 2120 7120
rect 2272 7114 2330 7120
rect 2482 7114 2540 7120
rect 2692 7114 2750 7120
rect 2902 7114 2960 7120
rect 3112 7114 3170 7120
rect 3322 7114 3380 7120
rect 3532 7114 3590 7120
rect 3742 7114 3800 7120
rect 3952 7114 4010 7120
rect 4162 7114 4220 7120
rect 4372 7114 4430 7120
rect 4582 7114 4640 7120
rect 4792 7114 4850 7120
rect 5002 7114 5060 7120
rect 5212 7114 5270 7120
rect 5422 7114 5480 7120
rect 5632 7114 5690 7120
rect 5842 7114 5900 7120
rect 1448 7061 1458 7070
rect -2432 7027 1458 7061
rect 1448 7018 1458 7027
rect 1510 7061 1520 7070
rect 1510 7027 5912 7061
rect 1510 7018 1520 7027
rect 921 6793 931 6845
rect 983 6793 1970 6845
rect 2022 6793 2032 6845
rect -3082 6668 -3072 6720
rect -3020 6668 -2009 6720
rect -1957 6668 -1379 6720
rect -1327 6668 -539 6720
rect -487 6668 301 6720
rect 353 6668 931 6720
rect 983 6668 994 6720
rect 2390 6668 2401 6720
rect 2453 6668 3031 6720
rect 3083 6668 3871 6720
rect 3923 6668 4711 6720
rect 4763 6668 5340 6720
rect 5392 6668 6482 6720
rect 6534 6668 6544 6720
rect 1448 6536 1458 6588
rect 1510 6536 2401 6588
rect 2453 6536 2463 6588
rect -3668 6067 -3150 6073
rect -3668 6033 -3656 6067
rect -3282 6033 -3150 6067
rect -3668 6027 -3150 6033
rect -3220 5619 -3150 6027
rect -3668 5613 -3150 5619
rect -3668 5579 -3656 5613
rect -3282 5579 -3150 5613
rect -3668 5573 -3150 5579
rect -3557 5313 -3523 5573
rect -3427 5403 -3369 5409
rect -3427 5369 -3415 5403
rect -3381 5369 -3369 5403
rect -3427 5363 -3369 5369
rect -3569 5307 -3511 5313
rect -3650 5173 -3616 5275
rect -3569 5273 -3557 5307
rect -3523 5273 -3511 5307
rect -3569 5267 -3511 5273
rect -3670 5121 -3660 5173
rect -3608 5121 -3598 5173
rect -3557 5121 -3523 5267
rect -3415 5217 -3381 5363
rect -3427 5211 -3369 5217
rect -3427 5177 -3415 5211
rect -3381 5177 -3369 5211
rect -3427 5171 -3369 5177
rect -3322 5173 -3288 5371
rect -3650 4021 -3616 5121
rect -3569 5115 -3511 5121
rect -3569 5081 -3557 5115
rect -3523 5081 -3511 5115
rect -3569 5075 -3511 5081
rect -3557 4929 -3523 5075
rect -3415 5025 -3381 5171
rect -3339 5121 -3329 5173
rect -3277 5121 -3267 5173
rect -3427 5019 -3369 5025
rect -3427 4985 -3415 5019
rect -3381 4985 -3369 5019
rect -3427 4979 -3369 4985
rect -3569 4923 -3511 4929
rect -3569 4889 -3557 4923
rect -3523 4889 -3511 4923
rect -3569 4883 -3511 4889
rect -3557 4737 -3523 4883
rect -3415 4833 -3381 4979
rect -3427 4827 -3369 4833
rect -3427 4793 -3415 4827
rect -3381 4793 -3369 4827
rect -3427 4787 -3369 4793
rect -3569 4731 -3511 4737
rect -3569 4697 -3557 4731
rect -3523 4697 -3511 4731
rect -3569 4691 -3511 4697
rect -3557 4545 -3523 4691
rect -3415 4641 -3381 4787
rect -3427 4635 -3369 4641
rect -3427 4601 -3415 4635
rect -3381 4601 -3369 4635
rect -3427 4595 -3369 4601
rect -3569 4539 -3511 4545
rect -3569 4505 -3557 4539
rect -3523 4505 -3511 4539
rect -3569 4499 -3511 4505
rect -3557 4353 -3523 4499
rect -3415 4497 -3381 4595
rect -3435 4445 -3425 4497
rect -3373 4445 -3363 4497
rect -3427 4443 -3369 4445
rect -3427 4409 -3415 4443
rect -3381 4409 -3369 4443
rect -3427 4403 -3369 4409
rect -3569 4347 -3511 4353
rect -3569 4313 -3557 4347
rect -3523 4313 -3511 4347
rect -3569 4307 -3511 4313
rect -3557 4161 -3523 4307
rect -3415 4257 -3381 4403
rect -3427 4251 -3369 4257
rect -3427 4217 -3415 4251
rect -3381 4217 -3369 4251
rect -3427 4211 -3369 4217
rect -3569 4155 -3511 4161
rect -3569 4121 -3557 4155
rect -3523 4121 -3511 4155
rect -3569 4115 -3511 4121
rect -3670 3969 -3660 4021
rect -3608 3969 -3598 4021
rect -3557 3969 -3523 4115
rect -3415 4065 -3381 4211
rect -3427 4059 -3369 4065
rect -3427 4025 -3415 4059
rect -3381 4025 -3369 4059
rect -3427 4019 -3369 4025
rect -3322 4021 -3288 5121
rect -3650 3865 -3616 3969
rect -3569 3963 -3511 3969
rect -3569 3929 -3557 3963
rect -3523 3929 -3511 3963
rect -3569 3923 -3511 3929
rect -3415 3873 -3381 4019
rect -3341 3969 -3331 4021
rect -3279 3969 -3269 4021
rect -3322 3961 -3288 3969
rect -3427 3867 -3369 3873
rect -3427 3833 -3415 3867
rect -3381 3833 -3369 3867
rect -3427 3827 -3369 3833
rect -3220 3663 -3150 5573
rect -2845 6435 -2704 6447
rect -2845 6412 -2744 6435
rect -2845 6360 -2798 6412
rect -2746 6360 -2744 6412
rect -2845 6271 -2744 6360
rect -2845 6219 -2798 6271
rect -2746 6219 -2744 6271
rect -2845 6130 -2744 6219
rect -2845 6078 -2798 6130
rect -2746 6078 -2744 6130
rect -2845 5989 -2744 6078
rect -2845 5937 -2798 5989
rect -2746 5937 -2744 5989
rect -2845 5848 -2744 5937
rect -2845 5796 -2798 5848
rect -2746 5796 -2744 5848
rect -2845 5707 -2744 5796
rect -2845 5655 -2798 5707
rect -2746 5655 -2744 5707
rect -2845 5566 -2744 5655
rect -2845 5514 -2798 5566
rect -2746 5514 -2744 5566
rect -2845 5425 -2744 5514
rect -2845 5373 -2798 5425
rect -2746 5373 -2744 5425
rect -2845 5284 -2744 5373
rect -2845 5232 -2798 5284
rect -2746 5232 -2744 5284
rect -2845 5143 -2744 5232
rect -2845 5091 -2798 5143
rect -2746 5091 -2744 5143
rect -2845 5002 -2744 5091
rect -2845 4950 -2798 5002
rect -2746 4950 -2744 5002
rect -2845 4861 -2744 4950
rect -2845 4809 -2798 4861
rect -2746 4809 -2744 4861
rect -2845 4759 -2744 4809
rect -2710 4759 -2704 6435
rect 1960 6429 1970 6438
rect -2432 6395 1970 6429
rect 1960 6386 1970 6395
rect 2022 6429 2032 6438
rect 6186 6435 6322 6447
rect 2022 6395 5900 6429
rect 2022 6386 2032 6395
rect 3021 6293 3031 6345
rect 3083 6293 3093 6345
rect 4701 6293 4711 6345
rect 4763 6293 4773 6345
rect 2391 6169 2401 6221
rect 2453 6169 2463 6221
rect 3861 6169 3871 6221
rect 3923 6169 3933 6221
rect 5330 6169 5340 6221
rect 5392 6169 5402 6221
rect 1960 6119 1970 6128
rect -2432 6085 1970 6119
rect 1960 6076 1970 6085
rect 2022 6119 2032 6128
rect 2022 6085 5900 6119
rect 2022 6076 2032 6085
rect 1448 5989 1458 5998
rect -2432 5955 1458 5989
rect 1448 5946 1458 5955
rect 1510 5989 1520 5998
rect 1510 5955 5900 5989
rect 1510 5946 1520 5955
rect -1389 5853 -1379 5905
rect -1327 5853 -1317 5905
rect 291 5853 301 5905
rect 353 5853 363 5905
rect -2019 5729 -2009 5781
rect -1957 5729 -1947 5781
rect -549 5729 -539 5781
rect -487 5729 -477 5781
rect 921 5729 931 5781
rect 983 5729 993 5781
rect 1448 5679 1458 5686
rect -2432 5645 1458 5679
rect 1448 5634 1458 5645
rect 1510 5679 1520 5686
rect 1510 5645 5900 5679
rect 1510 5634 1520 5645
rect 1448 5549 1458 5558
rect -2432 5515 1458 5549
rect 1448 5506 1458 5515
rect 1510 5549 1520 5558
rect 1510 5515 5900 5549
rect 1510 5506 1520 5515
rect -1389 5413 -1379 5465
rect -1327 5413 -1317 5465
rect 291 5413 301 5465
rect 353 5413 363 5465
rect -2019 5289 -2009 5341
rect -1957 5289 -1947 5341
rect -549 5289 -539 5341
rect -487 5289 -477 5341
rect 921 5289 931 5341
rect 983 5289 993 5341
rect 1448 5239 1458 5245
rect -2432 5205 1458 5239
rect 1448 5193 1458 5205
rect 1510 5239 1520 5245
rect 1510 5205 5900 5239
rect 1510 5193 1520 5205
rect 1960 5109 1970 5119
rect -2432 5075 1970 5109
rect 1960 5067 1970 5075
rect 2022 5109 2032 5119
rect 2022 5075 5900 5109
rect 2022 5067 2032 5075
rect 3021 4973 3031 5025
rect 3083 4973 3093 5025
rect 4701 4973 4711 5025
rect 4763 4973 4773 5025
rect 2391 4849 2401 4901
rect 2453 4849 2463 4901
rect 3861 4849 3871 4901
rect 3923 4849 3933 4901
rect 5330 4849 5340 4901
rect 5392 4849 5402 4901
rect 1960 4799 1970 4808
rect -2432 4765 1970 4799
rect -2845 4747 -2704 4759
rect 1960 4756 1970 4765
rect 2022 4799 2032 4808
rect 2022 4765 5900 4799
rect 2022 4756 2032 4765
rect 6186 4759 6192 6435
rect 6226 6412 6322 6435
rect 6226 6360 6229 6412
rect 6281 6360 6322 6412
rect 6226 6271 6322 6360
rect 6226 6219 6229 6271
rect 6281 6219 6322 6271
rect 6226 6130 6322 6219
rect 6226 6078 6229 6130
rect 6281 6078 6322 6130
rect 6226 5989 6322 6078
rect 6226 5937 6229 5989
rect 6281 5937 6322 5989
rect 6226 5848 6322 5937
rect 6226 5796 6229 5848
rect 6281 5796 6322 5848
rect 6226 5707 6322 5796
rect 6226 5655 6229 5707
rect 6281 5655 6322 5707
rect 6226 5566 6322 5655
rect 6226 5514 6229 5566
rect 6281 5514 6322 5566
rect 6226 5425 6322 5514
rect 6226 5373 6229 5425
rect 6281 5373 6322 5425
rect 6226 5284 6322 5373
rect 6226 5232 6229 5284
rect 6281 5232 6322 5284
rect 6226 5143 6322 5232
rect 6226 5091 6229 5143
rect 6281 5091 6322 5143
rect 6226 5002 6322 5091
rect 6226 4950 6229 5002
rect 6281 4950 6322 5002
rect 6226 4861 6322 4950
rect 6226 4809 6229 4861
rect 6281 4809 6322 4861
rect 6226 4759 6322 4809
rect 6186 4747 6322 4759
rect 6612 6073 6682 7983
rect 6831 7813 6889 7819
rect 6750 7581 6784 7781
rect 6831 7779 6843 7813
rect 6877 7779 6889 7813
rect 6831 7773 6889 7779
rect 6843 7627 6877 7773
rect 6985 7723 7019 7983
rect 6973 7717 7031 7723
rect 6973 7683 6985 7717
rect 7019 7683 7031 7717
rect 6973 7677 7031 7683
rect 6831 7621 6889 7627
rect 6831 7587 6843 7621
rect 6877 7587 6889 7621
rect 6831 7581 6889 7587
rect 6731 7529 6741 7581
rect 6793 7529 6803 7581
rect 6750 6431 6784 7529
rect 6843 7435 6877 7581
rect 6985 7531 7019 7677
rect 7078 7581 7112 7685
rect 6973 7525 7031 7531
rect 7062 7529 7072 7581
rect 7124 7529 7134 7581
rect 6973 7491 6985 7525
rect 7019 7491 7031 7525
rect 6973 7485 7031 7491
rect 6831 7429 6889 7435
rect 6831 7395 6843 7429
rect 6877 7395 6889 7429
rect 6831 7389 6889 7395
rect 6843 7243 6877 7389
rect 6985 7339 7019 7485
rect 6973 7333 7031 7339
rect 6973 7299 6985 7333
rect 7019 7299 7031 7333
rect 6973 7293 7031 7299
rect 6831 7237 6889 7243
rect 6831 7203 6843 7237
rect 6877 7203 6889 7237
rect 6831 7197 6889 7203
rect 6843 7051 6877 7197
rect 6985 7147 7019 7293
rect 6973 7141 7031 7147
rect 6973 7107 6985 7141
rect 7019 7107 7031 7141
rect 6973 7101 7031 7107
rect 6831 7045 6889 7051
rect 6831 7011 6843 7045
rect 6877 7011 6889 7045
rect 6831 7005 6889 7011
rect 6843 6859 6877 7005
rect 6985 6955 7019 7101
rect 6973 6949 7031 6955
rect 6973 6915 6985 6949
rect 7019 6915 7031 6949
rect 6973 6909 7031 6915
rect 6831 6853 6889 6859
rect 6831 6819 6843 6853
rect 6877 6819 6889 6853
rect 6831 6813 6889 6819
rect 6843 6720 6877 6813
rect 6985 6763 7019 6909
rect 6973 6757 7031 6763
rect 6973 6723 6985 6757
rect 7019 6723 7031 6757
rect 6823 6668 6833 6720
rect 6885 6668 6895 6720
rect 6973 6717 7031 6723
rect 6831 6661 6889 6668
rect 6831 6627 6843 6661
rect 6877 6627 6889 6661
rect 6831 6621 6889 6627
rect 6843 6475 6877 6621
rect 6985 6571 7019 6717
rect 6973 6565 7031 6571
rect 6973 6531 6985 6565
rect 7019 6531 7031 6565
rect 6973 6525 7031 6531
rect 6831 6469 6889 6475
rect 6831 6435 6843 6469
rect 6877 6435 6889 6469
rect 6731 6379 6741 6431
rect 6793 6379 6803 6431
rect 6831 6429 6889 6435
rect 6750 6371 6784 6379
rect 6843 6283 6877 6429
rect 6985 6379 7019 6525
rect 7078 6431 7112 7529
rect 7060 6379 7070 6431
rect 7122 6379 7132 6431
rect 6973 6373 7031 6379
rect 6973 6339 6985 6373
rect 7019 6339 7031 6373
rect 6973 6333 7031 6339
rect 6831 6277 6889 6283
rect 6831 6243 6843 6277
rect 6877 6243 6889 6277
rect 6831 6237 6889 6243
rect 6985 6073 7019 6333
rect 7078 6275 7112 6379
rect 6612 6067 7130 6073
rect 6612 6033 6744 6067
rect 7118 6033 7130 6067
rect 6612 6027 7130 6033
rect 6612 5619 6682 6027
rect 6612 5613 7130 5619
rect 6612 5579 6744 5613
rect 7118 5579 7130 5613
rect 6612 5573 7130 5579
rect -3082 4445 -3072 4497
rect -3020 4445 -2009 4497
rect -1957 4445 -539 4497
rect -487 4445 931 4497
rect 983 4445 999 4497
rect 2391 4445 2401 4497
rect 2453 4445 3871 4497
rect 3923 4445 5340 4497
rect 5392 4445 6482 4497
rect 6534 4445 6544 4497
rect -3668 3657 -3150 3663
rect -3668 3623 -3656 3657
rect -3282 3623 -3150 3657
rect -3668 3617 -3150 3623
rect -3220 3587 -3150 3617
rect -2845 4180 -2704 4192
rect -2845 4144 -2744 4180
rect -2845 4092 -2798 4144
rect -2746 4092 -2744 4144
rect -2845 4003 -2744 4092
rect -2845 3951 -2798 4003
rect -2746 3951 -2744 4003
rect -2845 3862 -2744 3951
rect -2845 3810 -2798 3862
rect -2746 3810 -2744 3862
rect -2845 3721 -2744 3810
rect -2845 3669 -2798 3721
rect -2746 3669 -2744 3721
rect -2845 3580 -2744 3669
rect -2845 3528 -2798 3580
rect -2746 3528 -2744 3580
rect -2845 3439 -2744 3528
rect -2845 3387 -2798 3439
rect -2746 3387 -2744 3439
rect -2845 3298 -2744 3387
rect -2845 3246 -2798 3298
rect -2746 3246 -2744 3298
rect -2845 3157 -2744 3246
rect -2845 3105 -2798 3157
rect -2746 3105 -2744 3157
rect -2845 3016 -2744 3105
rect -2845 2964 -2798 3016
rect -2746 2964 -2744 3016
rect -2845 2875 -2744 2964
rect -2845 2823 -2798 2875
rect -2746 2823 -2744 2875
rect -2845 2734 -2744 2823
rect -2845 2682 -2798 2734
rect -2746 2682 -2744 2734
rect -2845 1549 -2744 2682
rect -2845 1497 -2798 1549
rect -2746 1497 -2744 1549
rect -2845 1408 -2744 1497
rect -2845 1356 -2798 1408
rect -2746 1356 -2744 1408
rect -2845 1267 -2744 1356
rect -2845 1215 -2798 1267
rect -2746 1215 -2744 1267
rect -2845 1126 -2744 1215
rect -2845 1074 -2798 1126
rect -2746 1074 -2744 1126
rect -2845 985 -2744 1074
rect -2845 933 -2798 985
rect -2746 933 -2744 985
rect -2845 844 -2744 933
rect -2845 792 -2798 844
rect -2746 792 -2744 844
rect -2845 745 -2744 792
rect -2710 745 -2704 4180
rect -2598 4131 -2588 4183
rect -2536 4174 -2526 4183
rect -2391 4174 -2319 4183
rect -1551 4174 -1479 4183
rect -711 4174 -639 4183
rect 129 4174 201 4183
rect 969 4174 1041 4183
rect 6186 4180 6322 4192
rect -2536 4140 5912 4174
rect -2536 4131 -2526 4140
rect -2391 4131 -2319 4140
rect -1551 4131 -1479 4140
rect -711 4131 -639 4140
rect 129 4131 201 4140
rect 969 4131 1041 4140
rect -2432 4090 -2374 4096
rect -2229 4090 -2157 4096
rect -2012 4090 -1954 4096
rect -1802 4090 -1744 4096
rect -1592 4090 -1534 4096
rect -1382 4090 -1324 4096
rect -1172 4090 -1114 4096
rect -962 4090 -904 4096
rect -752 4090 -694 4096
rect -549 4090 -539 4096
rect -487 4090 -477 4096
rect -332 4090 -274 4096
rect -122 4090 -64 4096
rect 88 4090 146 4096
rect 298 4090 356 4096
rect 508 4090 566 4096
rect 718 4090 776 4096
rect 928 4090 986 4096
rect 1138 4090 1196 4096
rect 1348 4090 1406 4096
rect 1558 4090 1616 4096
rect 1768 4090 1826 4096
rect 1978 4090 2036 4096
rect 2188 4090 2246 4096
rect 2398 4090 2456 4096
rect 2608 4090 2666 4096
rect 2818 4090 2876 4096
rect 3028 4090 3086 4096
rect 3238 4090 3296 4096
rect 3448 4090 3506 4096
rect 3658 4090 3716 4096
rect 3868 4090 3926 4096
rect 4078 4090 4136 4096
rect 4288 4090 4346 4096
rect 4498 4090 4556 4096
rect 4708 4090 4766 4096
rect 4918 4090 4976 4096
rect 5128 4090 5186 4096
rect 5338 4090 5396 4096
rect 5548 4090 5606 4096
rect 5758 4090 5816 4096
rect -2432 4056 -2420 4090
rect -2386 4056 -2210 4090
rect -2176 4056 -2009 4090
rect -1957 4056 -1790 4090
rect -1756 4056 -1580 4090
rect -1546 4056 -1370 4090
rect -1336 4056 -1160 4090
rect -1126 4056 -950 4090
rect -916 4056 -740 4090
rect -706 4056 -539 4090
rect -487 4056 -320 4090
rect -286 4056 -110 4090
rect -76 4056 100 4090
rect 134 4056 310 4090
rect 344 4056 520 4090
rect 554 4056 730 4090
rect 764 4056 931 4090
rect 983 4056 1150 4090
rect 1184 4056 1360 4090
rect 1394 4056 1570 4090
rect 1604 4056 1780 4090
rect 1814 4056 1990 4090
rect 2024 4056 2200 4090
rect 2234 4056 2410 4090
rect 2444 4056 2620 4090
rect 2654 4056 2830 4090
rect 2864 4056 3040 4090
rect 3074 4056 3250 4090
rect 3284 4056 3460 4090
rect 3494 4056 3670 4090
rect 3704 4056 3880 4090
rect 3914 4056 4090 4090
rect 4124 4056 4300 4090
rect 4334 4056 4510 4090
rect 4544 4056 4720 4090
rect 4754 4056 4930 4090
rect 4964 4056 5140 4090
rect 5174 4056 5350 4090
rect 5384 4056 5560 4090
rect 5594 4056 5770 4090
rect 5804 4056 5816 4090
rect -2432 4050 -2374 4056
rect -2229 4044 -2157 4056
rect -2019 4038 -2009 4056
rect -1957 4038 -1947 4056
rect -1802 4050 -1744 4056
rect -1592 4050 -1534 4056
rect -1382 4050 -1324 4056
rect -1172 4050 -1114 4056
rect -962 4050 -904 4056
rect -752 4050 -694 4056
rect -549 4044 -539 4056
rect -487 4044 -477 4056
rect -332 4050 -274 4056
rect -122 4050 -64 4056
rect 88 4050 146 4056
rect 298 4050 356 4056
rect 508 4050 566 4056
rect 718 4050 776 4056
rect 921 4038 931 4056
rect 983 4038 993 4056
rect 1138 4050 1196 4056
rect 1348 4050 1406 4056
rect 1558 4050 1616 4056
rect 1768 4050 1826 4056
rect 1978 4050 2036 4056
rect 2188 4050 2246 4056
rect 2398 4050 2456 4056
rect 2608 4050 2666 4056
rect 2818 4050 2876 4056
rect 3028 4050 3086 4056
rect 3238 4050 3296 4056
rect 3448 4050 3506 4056
rect 3658 4050 3716 4056
rect 3868 4050 3926 4056
rect 4078 4050 4136 4056
rect 4288 4050 4346 4056
rect 4498 4050 4556 4056
rect 4708 4050 4766 4056
rect 4918 4050 4976 4056
rect 5128 4050 5186 4056
rect 5338 4050 5396 4056
rect 5548 4050 5606 4056
rect 5758 4050 5816 4056
rect -2336 3948 -2278 3954
rect -2126 3948 -2068 3954
rect -1916 3948 -1858 3954
rect -1706 3948 -1648 3954
rect -1496 3948 -1438 3954
rect -1293 3948 -1283 3960
rect -1231 3948 -1221 3960
rect -1076 3948 -1018 3954
rect -866 3948 -808 3954
rect -656 3948 -598 3954
rect -446 3948 -388 3954
rect -236 3948 -178 3954
rect -26 3948 32 3954
rect 184 3948 242 3954
rect 292 3948 302 3960
rect -2336 3914 -2324 3948
rect -2290 3914 -2114 3948
rect -2080 3914 -1904 3948
rect -1870 3914 -1694 3948
rect -1660 3914 -1484 3948
rect -1450 3914 -1283 3948
rect -1231 3914 -1064 3948
rect -1030 3914 -854 3948
rect -820 3914 -644 3948
rect -610 3914 -434 3948
rect -400 3914 -224 3948
rect -190 3914 -14 3948
rect 20 3914 196 3948
rect 230 3914 302 3948
rect -2336 3908 -2278 3914
rect -2126 3908 -2068 3914
rect -1916 3908 -1858 3914
rect -1706 3908 -1648 3914
rect -1496 3908 -1438 3914
rect -1293 3908 -1283 3914
rect -1231 3908 -1221 3914
rect -1076 3908 -1018 3914
rect -866 3908 -808 3914
rect -656 3908 -598 3914
rect -446 3908 -388 3914
rect -236 3908 -178 3914
rect -26 3908 32 3914
rect 184 3908 242 3914
rect 292 3908 302 3914
rect 354 3948 364 3960
rect 394 3948 452 3954
rect 604 3948 662 3954
rect 814 3948 872 3954
rect 1024 3948 1082 3954
rect 1234 3948 1292 3954
rect 1444 3948 1502 3954
rect 1647 3948 1657 3960
rect 1709 3948 1719 3960
rect 1864 3948 1922 3954
rect 2074 3948 2132 3954
rect 2284 3948 2342 3954
rect 2494 3948 2552 3954
rect 2704 3948 2762 3954
rect 2907 3948 2917 3960
rect 2969 3948 2979 3960
rect 3124 3948 3182 3954
rect 3334 3948 3392 3954
rect 3544 3948 3602 3954
rect 3754 3948 3812 3954
rect 3964 3948 4022 3954
rect 4174 3948 4232 3954
rect 4384 3948 4442 3954
rect 4594 3948 4652 3954
rect 4804 3948 4862 3954
rect 4911 3948 4921 3960
rect 354 3914 406 3948
rect 440 3914 616 3948
rect 650 3914 826 3948
rect 860 3914 1036 3948
rect 1070 3914 1246 3948
rect 1280 3914 1456 3948
rect 1490 3914 1657 3948
rect 1709 3914 1876 3948
rect 1910 3914 2086 3948
rect 2120 3914 2296 3948
rect 2330 3914 2506 3948
rect 2540 3914 2716 3948
rect 2750 3914 2917 3948
rect 2969 3914 3136 3948
rect 3170 3914 3346 3948
rect 3380 3914 3556 3948
rect 3590 3914 3766 3948
rect 3800 3914 3976 3948
rect 4010 3914 4186 3948
rect 4220 3914 4396 3948
rect 4430 3914 4606 3948
rect 4640 3914 4816 3948
rect 4850 3914 4921 3948
rect 354 3908 364 3914
rect 394 3908 452 3914
rect 604 3908 662 3914
rect 814 3908 872 3914
rect 1024 3908 1082 3914
rect 1234 3908 1292 3914
rect 1444 3908 1502 3914
rect 1647 3908 1657 3914
rect 1709 3908 1719 3914
rect 1864 3908 1922 3914
rect 2074 3908 2132 3914
rect 2284 3908 2342 3914
rect 2494 3908 2552 3914
rect 2704 3908 2762 3914
rect 2907 3908 2917 3914
rect 2969 3908 2979 3914
rect 3124 3908 3182 3914
rect 3334 3908 3392 3914
rect 3544 3908 3602 3914
rect 3754 3908 3812 3914
rect 3964 3908 4022 3914
rect 4174 3908 4232 3914
rect 4384 3908 4442 3914
rect 4594 3908 4652 3914
rect 4804 3908 4862 3914
rect 4911 3908 4921 3914
rect 4973 3948 4983 3960
rect 5014 3948 5072 3954
rect 5224 3948 5282 3954
rect 5434 3948 5492 3954
rect 5644 3948 5702 3954
rect 5854 3948 5912 3954
rect 4973 3914 5026 3948
rect 5060 3914 5236 3948
rect 5270 3914 5446 3948
rect 5480 3914 5656 3948
rect 5690 3914 5866 3948
rect 5900 3914 5912 3948
rect 4973 3908 4983 3914
rect 5014 3908 5072 3914
rect 5224 3908 5282 3914
rect 5434 3908 5492 3914
rect 5644 3908 5702 3914
rect 5854 3908 5912 3914
rect -2598 3821 -2588 3873
rect -2536 3864 -2526 3873
rect -2181 3864 -2109 3873
rect -1341 3864 -1269 3873
rect -501 3864 -429 3873
rect 339 3864 411 3873
rect 1179 3864 1251 3873
rect -2536 3830 5912 3864
rect -2536 3821 -2526 3830
rect -2181 3821 -2109 3830
rect -1341 3821 -1269 3830
rect -501 3821 -429 3830
rect 339 3821 411 3830
rect 1179 3821 1251 3830
rect -1971 3734 -1899 3743
rect -291 3734 -219 3743
rect 1389 3734 1461 3743
rect 6010 3734 6020 3743
rect -2432 3700 6020 3734
rect -1971 3691 -1899 3700
rect -291 3691 -219 3700
rect 1389 3691 1461 3700
rect 6010 3691 6020 3700
rect 6072 3691 6082 3743
rect -2432 3650 -2374 3656
rect -2222 3650 -2164 3656
rect -2012 3650 -1954 3656
rect -1802 3650 -1744 3656
rect -1592 3650 -1534 3656
rect -1382 3650 -1324 3656
rect -1172 3650 -1114 3656
rect -962 3650 -904 3656
rect -752 3650 -694 3656
rect -542 3650 -484 3656
rect -332 3650 -274 3656
rect -122 3650 -64 3656
rect 88 3650 146 3656
rect 298 3650 356 3656
rect 508 3650 566 3656
rect 718 3650 776 3656
rect 928 3650 986 3656
rect 1138 3650 1196 3656
rect 1348 3650 1406 3656
rect 1558 3650 1616 3656
rect 1768 3650 1826 3656
rect 1978 3650 2036 3656
rect 2188 3650 2246 3656
rect 2398 3650 2456 3656
rect 2608 3650 2666 3656
rect 2818 3650 2876 3656
rect 3028 3650 3086 3656
rect 3238 3650 3296 3656
rect 3448 3650 3506 3656
rect 3658 3650 3716 3656
rect 3868 3650 3926 3656
rect 4078 3650 4136 3656
rect 4288 3650 4346 3656
rect 4498 3650 4556 3656
rect 4708 3650 4766 3656
rect 4918 3650 4976 3656
rect 5128 3650 5186 3656
rect 5338 3650 5396 3656
rect 5548 3650 5606 3656
rect 5758 3650 5816 3656
rect -2432 3616 -2420 3650
rect -2386 3616 -2210 3650
rect -2176 3616 -2000 3650
rect -1966 3616 -1790 3650
rect -1756 3616 -1580 3650
rect -1546 3616 -1370 3650
rect -1336 3616 -1160 3650
rect -1126 3616 -950 3650
rect -916 3616 -740 3650
rect -706 3616 -530 3650
rect -496 3616 -320 3650
rect -286 3616 -110 3650
rect -76 3616 100 3650
rect 134 3616 310 3650
rect 344 3616 520 3650
rect 554 3616 730 3650
rect 764 3616 940 3650
rect 974 3616 1150 3650
rect 1184 3616 1360 3650
rect 1394 3616 1570 3650
rect 1604 3616 1780 3650
rect 1814 3616 1990 3650
rect 2024 3616 2200 3650
rect 2234 3616 2401 3650
rect 2453 3616 2620 3650
rect 2654 3616 2830 3650
rect 2864 3616 3040 3650
rect 3074 3616 3250 3650
rect 3284 3616 3460 3650
rect 3494 3616 3670 3650
rect 3704 3616 3871 3650
rect 3923 3616 4090 3650
rect 4124 3616 4300 3650
rect 4334 3616 4510 3650
rect 4544 3616 4720 3650
rect 4754 3616 4930 3650
rect 4964 3616 5140 3650
rect 5174 3616 5340 3650
rect 5392 3616 5560 3650
rect 5594 3616 5770 3650
rect 5804 3616 5816 3650
rect -2432 3610 -2374 3616
rect -2222 3610 -2164 3616
rect -2012 3610 -1954 3616
rect -1802 3610 -1744 3616
rect -1592 3610 -1534 3616
rect -1382 3610 -1324 3616
rect -1172 3610 -1114 3616
rect -962 3610 -904 3616
rect -752 3610 -694 3616
rect -542 3610 -484 3616
rect -332 3610 -274 3616
rect -122 3610 -64 3616
rect 88 3610 146 3616
rect 298 3610 356 3616
rect 508 3610 566 3616
rect 718 3610 776 3616
rect 928 3610 986 3616
rect 1138 3610 1196 3616
rect 1348 3610 1406 3616
rect 1558 3610 1616 3616
rect 1768 3610 1826 3616
rect 1978 3610 2036 3616
rect 2188 3610 2246 3616
rect 2391 3598 2401 3616
rect 2453 3598 2463 3616
rect 2608 3610 2666 3616
rect 2818 3610 2876 3616
rect 3028 3610 3086 3616
rect 3238 3610 3296 3616
rect 3448 3610 3506 3616
rect 3658 3610 3716 3616
rect 3861 3598 3871 3616
rect 3923 3598 3933 3616
rect 4078 3610 4136 3616
rect 4288 3610 4346 3616
rect 4498 3610 4556 3616
rect 4708 3610 4766 3616
rect 4918 3610 4976 3616
rect 5128 3610 5186 3616
rect 5330 3598 5340 3616
rect 5392 3598 5402 3616
rect 5548 3610 5606 3616
rect 5758 3610 5816 3616
rect -2336 3508 -2278 3514
rect -2126 3508 -2068 3514
rect -1916 3508 -1858 3514
rect -1706 3508 -1648 3514
rect -1496 3508 -1438 3514
rect -1293 3508 -1283 3520
rect -1231 3508 -1221 3520
rect -1076 3508 -1018 3514
rect -866 3508 -808 3514
rect -656 3508 -598 3514
rect -446 3508 -388 3514
rect -236 3508 -178 3514
rect -26 3508 32 3514
rect 184 3508 242 3514
rect 292 3508 302 3520
rect -2336 3474 -2324 3508
rect -2290 3474 -2114 3508
rect -2080 3474 -1904 3508
rect -1870 3474 -1694 3508
rect -1660 3474 -1484 3508
rect -1450 3474 -1283 3508
rect -1231 3474 -1064 3508
rect -1030 3474 -854 3508
rect -820 3474 -644 3508
rect -610 3474 -434 3508
rect -400 3474 -224 3508
rect -190 3474 -14 3508
rect 20 3474 196 3508
rect 230 3474 302 3508
rect -2336 3468 -2278 3474
rect -2126 3468 -2068 3474
rect -1916 3468 -1858 3474
rect -1706 3468 -1648 3474
rect -1496 3468 -1438 3474
rect -1293 3468 -1283 3474
rect -1231 3468 -1221 3474
rect -1076 3468 -1018 3474
rect -866 3468 -808 3474
rect -656 3468 -598 3474
rect -446 3468 -388 3474
rect -236 3468 -178 3474
rect -26 3468 32 3474
rect 184 3468 242 3474
rect 292 3468 302 3474
rect 354 3508 364 3520
rect 394 3508 452 3514
rect 604 3508 662 3514
rect 814 3508 872 3514
rect 1024 3508 1082 3514
rect 1234 3508 1292 3514
rect 1444 3508 1502 3514
rect 1647 3508 1657 3520
rect 1709 3508 1719 3520
rect 1864 3508 1922 3514
rect 2074 3508 2132 3514
rect 2284 3508 2342 3514
rect 2494 3508 2552 3514
rect 2704 3508 2762 3514
rect 2907 3508 2917 3520
rect 2969 3508 2979 3520
rect 3124 3508 3182 3514
rect 3334 3508 3392 3514
rect 3544 3508 3602 3514
rect 3754 3508 3812 3514
rect 3964 3508 4022 3514
rect 4174 3508 4232 3514
rect 4384 3508 4442 3514
rect 4594 3508 4652 3514
rect 4804 3508 4862 3514
rect 4911 3508 4921 3520
rect 354 3474 406 3508
rect 440 3474 616 3508
rect 650 3474 826 3508
rect 860 3474 1036 3508
rect 1070 3474 1246 3508
rect 1280 3474 1456 3508
rect 1490 3474 1657 3508
rect 1709 3474 1876 3508
rect 1910 3474 2086 3508
rect 2120 3474 2296 3508
rect 2330 3474 2506 3508
rect 2540 3474 2716 3508
rect 2750 3474 2917 3508
rect 2969 3474 3136 3508
rect 3170 3474 3346 3508
rect 3380 3474 3556 3508
rect 3590 3474 3766 3508
rect 3800 3474 3976 3508
rect 4010 3474 4186 3508
rect 4220 3474 4396 3508
rect 4430 3474 4606 3508
rect 4640 3474 4816 3508
rect 4850 3474 4921 3508
rect 354 3468 364 3474
rect 394 3468 452 3474
rect 604 3468 662 3474
rect 814 3468 872 3474
rect 1024 3468 1082 3474
rect 1234 3468 1292 3474
rect 1444 3468 1502 3474
rect 1647 3468 1657 3474
rect 1709 3468 1719 3474
rect 1864 3468 1922 3474
rect 2074 3468 2132 3474
rect 2284 3468 2342 3474
rect 2494 3468 2552 3474
rect 2704 3468 2762 3474
rect 2907 3468 2917 3474
rect 2969 3468 2979 3474
rect 3124 3468 3182 3474
rect 3334 3468 3392 3474
rect 3544 3468 3602 3474
rect 3754 3468 3812 3474
rect 3964 3468 4022 3474
rect 4174 3468 4232 3474
rect 4384 3468 4442 3474
rect 4594 3468 4652 3474
rect 4804 3468 4862 3474
rect 4911 3468 4921 3474
rect 4973 3508 4983 3520
rect 5014 3508 5072 3514
rect 5224 3508 5282 3514
rect 5434 3508 5492 3514
rect 5644 3508 5702 3514
rect 5854 3508 5912 3514
rect 4973 3474 5026 3508
rect 5060 3474 5236 3508
rect 5270 3474 5446 3508
rect 5480 3474 5656 3508
rect 5690 3474 5866 3508
rect 5900 3474 5912 3508
rect 4973 3468 4983 3474
rect 5014 3468 5072 3474
rect 5224 3468 5282 3474
rect 5434 3468 5492 3474
rect 5644 3468 5702 3474
rect 5854 3468 5912 3474
rect -1761 3424 -1689 3433
rect -81 3424 -9 3433
rect 1599 3424 1671 3433
rect 6010 3424 6020 3433
rect -2432 3390 6020 3424
rect -1761 3381 -1689 3390
rect -81 3381 -9 3390
rect 1599 3381 1671 3390
rect 6010 3381 6020 3390
rect 6072 3381 6082 3433
rect -2391 3294 -2319 3303
rect -1551 3294 -1479 3303
rect -711 3294 -639 3303
rect 129 3294 201 3303
rect 969 3294 1041 3303
rect 6010 3294 6020 3305
rect -2432 3260 6020 3294
rect -2391 3251 -2319 3260
rect -1551 3251 -1479 3260
rect -711 3251 -639 3260
rect 129 3251 201 3260
rect 969 3251 1041 3260
rect 6010 3253 6020 3260
rect 6072 3253 6082 3305
rect -2432 3210 -2374 3216
rect -2222 3210 -2164 3216
rect -2012 3210 -1954 3216
rect -1802 3210 -1744 3216
rect -1592 3210 -1534 3216
rect -1382 3210 -1324 3216
rect -1172 3210 -1114 3216
rect -962 3210 -904 3216
rect -752 3210 -694 3216
rect -542 3210 -484 3216
rect -332 3210 -274 3216
rect -122 3210 -64 3216
rect 88 3210 146 3216
rect 298 3210 356 3216
rect 508 3210 566 3216
rect 718 3210 776 3216
rect 928 3210 986 3216
rect 1138 3210 1196 3216
rect 1348 3210 1406 3216
rect 1558 3210 1616 3216
rect 1768 3210 1826 3216
rect 1978 3210 2036 3216
rect 2188 3210 2246 3216
rect 2398 3210 2456 3216
rect 2608 3210 2666 3216
rect 2818 3210 2876 3216
rect 3028 3210 3086 3216
rect 3238 3210 3296 3216
rect 3448 3210 3506 3216
rect 3658 3210 3716 3216
rect 3868 3210 3926 3216
rect 4078 3210 4136 3216
rect 4288 3210 4346 3216
rect 4498 3210 4556 3216
rect 4708 3210 4766 3216
rect 4918 3210 4976 3216
rect 5128 3210 5186 3216
rect 5338 3210 5396 3216
rect 5548 3210 5606 3216
rect 5758 3210 5816 3216
rect -2432 3176 -2420 3210
rect -2386 3176 -2210 3210
rect -2176 3176 -2000 3210
rect -1966 3176 -1790 3210
rect -1756 3176 -1580 3210
rect -1546 3176 -1370 3210
rect -1336 3176 -1160 3210
rect -1126 3176 -950 3210
rect -916 3176 -740 3210
rect -706 3176 -530 3210
rect -496 3176 -320 3210
rect -286 3176 -110 3210
rect -76 3176 100 3210
rect 134 3176 310 3210
rect 344 3176 520 3210
rect 554 3176 730 3210
rect 764 3176 940 3210
rect 974 3176 1150 3210
rect 1184 3176 1360 3210
rect 1394 3176 1570 3210
rect 1604 3176 1780 3210
rect 1814 3176 1990 3210
rect 2024 3176 2200 3210
rect 2234 3176 2401 3210
rect 2453 3176 2620 3210
rect 2654 3176 2830 3210
rect 2864 3176 3040 3210
rect 3074 3176 3250 3210
rect 3284 3176 3460 3210
rect 3494 3176 3670 3210
rect 3704 3176 3871 3210
rect 3923 3176 4090 3210
rect 4124 3176 4300 3210
rect 4334 3176 4510 3210
rect 4544 3176 4720 3210
rect 4754 3176 4930 3210
rect 4964 3176 5140 3210
rect 5174 3176 5340 3210
rect 5392 3176 5560 3210
rect 5594 3176 5770 3210
rect 5804 3176 5816 3210
rect -2432 3170 -2374 3176
rect -2222 3170 -2164 3176
rect -2012 3170 -1954 3176
rect -1802 3170 -1744 3176
rect -1592 3170 -1534 3176
rect -1382 3170 -1324 3176
rect -1172 3170 -1114 3176
rect -962 3170 -904 3176
rect -752 3170 -694 3176
rect -542 3170 -484 3176
rect -332 3170 -274 3176
rect -122 3170 -64 3176
rect 88 3170 146 3176
rect 298 3170 356 3176
rect 508 3170 566 3176
rect 718 3170 776 3176
rect 928 3170 986 3176
rect 1138 3170 1196 3176
rect 1348 3170 1406 3176
rect 1558 3170 1616 3176
rect 1768 3170 1826 3176
rect 1978 3170 2036 3176
rect 2188 3170 2246 3176
rect 2391 3158 2401 3176
rect 2453 3158 2463 3176
rect 2608 3170 2666 3176
rect 2818 3170 2876 3176
rect 3028 3170 3086 3176
rect 3238 3170 3296 3176
rect 3448 3170 3506 3176
rect 3658 3170 3716 3176
rect 3861 3158 3871 3176
rect 3923 3158 3933 3176
rect 4078 3170 4136 3176
rect 4288 3170 4346 3176
rect 4498 3170 4556 3176
rect 4708 3170 4766 3176
rect 4918 3170 4976 3176
rect 5128 3170 5186 3176
rect 5330 3158 5340 3176
rect 5392 3158 5402 3176
rect 5548 3170 5606 3176
rect 5758 3170 5816 3176
rect -2336 3068 -2278 3074
rect -2126 3068 -2068 3074
rect -1916 3068 -1858 3074
rect -1706 3068 -1648 3074
rect -1496 3068 -1438 3074
rect -1293 3068 -1283 3080
rect -1231 3068 -1221 3080
rect -1076 3068 -1018 3074
rect -866 3068 -808 3074
rect -656 3068 -598 3074
rect -446 3068 -388 3074
rect -236 3068 -178 3074
rect -26 3068 32 3074
rect 184 3068 242 3074
rect 292 3068 302 3080
rect -2336 3034 -2324 3068
rect -2290 3034 -2114 3068
rect -2080 3034 -1904 3068
rect -1870 3034 -1694 3068
rect -1660 3034 -1484 3068
rect -1450 3034 -1283 3068
rect -1231 3034 -1064 3068
rect -1030 3034 -854 3068
rect -820 3034 -644 3068
rect -610 3034 -434 3068
rect -400 3034 -224 3068
rect -190 3034 -14 3068
rect 20 3034 196 3068
rect 230 3034 302 3068
rect -2336 3028 -2278 3034
rect -2126 3028 -2068 3034
rect -1916 3028 -1858 3034
rect -1706 3028 -1648 3034
rect -1496 3028 -1438 3034
rect -1293 3028 -1283 3034
rect -1231 3028 -1221 3034
rect -1076 3028 -1018 3034
rect -866 3028 -808 3034
rect -656 3028 -598 3034
rect -446 3028 -388 3034
rect -236 3028 -178 3034
rect -26 3028 32 3034
rect 184 3028 242 3034
rect 292 3028 302 3034
rect 354 3068 364 3080
rect 394 3068 452 3074
rect 604 3068 662 3074
rect 814 3068 872 3074
rect 1024 3068 1082 3074
rect 1234 3068 1292 3074
rect 1444 3068 1502 3074
rect 1647 3068 1657 3080
rect 1709 3068 1719 3080
rect 1864 3068 1922 3074
rect 2074 3068 2132 3074
rect 2284 3068 2342 3074
rect 2494 3068 2552 3074
rect 2704 3068 2762 3074
rect 2907 3068 2917 3080
rect 2969 3068 2979 3080
rect 3124 3068 3182 3074
rect 3334 3068 3392 3074
rect 3544 3068 3602 3074
rect 3754 3068 3812 3074
rect 3964 3068 4022 3074
rect 4174 3068 4232 3074
rect 4384 3068 4442 3074
rect 4594 3068 4652 3074
rect 4804 3068 4862 3074
rect 4911 3068 4921 3080
rect 354 3034 406 3068
rect 440 3034 616 3068
rect 650 3034 826 3068
rect 860 3034 1036 3068
rect 1070 3034 1246 3068
rect 1280 3034 1456 3068
rect 1490 3034 1657 3068
rect 1709 3034 1876 3068
rect 1910 3034 2086 3068
rect 2120 3034 2296 3068
rect 2330 3034 2506 3068
rect 2540 3034 2716 3068
rect 2750 3034 2917 3068
rect 2969 3034 3136 3068
rect 3170 3034 3346 3068
rect 3380 3034 3556 3068
rect 3590 3034 3766 3068
rect 3800 3034 3976 3068
rect 4010 3034 4186 3068
rect 4220 3034 4396 3068
rect 4430 3034 4606 3068
rect 4640 3034 4816 3068
rect 4850 3034 4921 3068
rect 354 3028 364 3034
rect 394 3028 452 3034
rect 604 3028 662 3034
rect 814 3028 872 3034
rect 1024 3028 1082 3034
rect 1234 3028 1292 3034
rect 1444 3028 1502 3034
rect 1647 3028 1657 3034
rect 1709 3028 1719 3034
rect 1864 3028 1922 3034
rect 2074 3028 2132 3034
rect 2284 3028 2342 3034
rect 2494 3028 2552 3034
rect 2704 3028 2762 3034
rect 2907 3028 2917 3034
rect 2969 3028 2979 3034
rect 3124 3028 3182 3034
rect 3334 3028 3392 3034
rect 3544 3028 3602 3034
rect 3754 3028 3812 3034
rect 3964 3028 4022 3034
rect 4174 3028 4232 3034
rect 4384 3028 4442 3034
rect 4594 3028 4652 3034
rect 4804 3028 4862 3034
rect 4911 3028 4921 3034
rect 4973 3068 4983 3080
rect 5014 3068 5072 3074
rect 5224 3068 5282 3074
rect 5434 3068 5492 3074
rect 5644 3068 5702 3074
rect 5854 3068 5912 3074
rect 4973 3034 5026 3068
rect 5060 3034 5236 3068
rect 5270 3034 5446 3068
rect 5480 3034 5656 3068
rect 5690 3034 5866 3068
rect 5900 3034 5912 3068
rect 4973 3028 4983 3034
rect 5014 3028 5072 3034
rect 5224 3028 5282 3034
rect 5434 3028 5492 3034
rect 5644 3028 5702 3034
rect 5854 3028 5912 3034
rect -2181 2984 -2109 2993
rect -1341 2984 -1269 2993
rect -501 2984 -429 2993
rect 339 2984 411 2993
rect 1179 2984 1251 2993
rect 6010 2984 6020 2991
rect -2432 2950 6020 2984
rect -2181 2941 -2109 2950
rect -1341 2941 -1269 2950
rect -501 2941 -429 2950
rect 339 2941 411 2950
rect 1179 2941 1251 2950
rect 6010 2939 6020 2950
rect 6072 2939 6082 2991
rect -2598 2811 -2588 2863
rect -2536 2854 -2526 2863
rect -1971 2854 -1899 2863
rect -291 2854 -219 2863
rect 1389 2854 1461 2863
rect -2536 2820 5912 2854
rect -2536 2811 -2526 2820
rect -1971 2811 -1899 2820
rect -291 2811 -219 2820
rect 1389 2811 1461 2820
rect -2432 2770 -2374 2776
rect -2229 2770 -2157 2776
rect -2012 2770 -1954 2776
rect -1802 2770 -1744 2776
rect -1592 2770 -1534 2776
rect -1382 2770 -1324 2776
rect -1172 2770 -1114 2776
rect -962 2770 -904 2776
rect -752 2770 -694 2776
rect -549 2770 -539 2776
rect -487 2770 -477 2776
rect -332 2770 -274 2776
rect -122 2770 -64 2776
rect 88 2770 146 2776
rect 298 2770 356 2776
rect 508 2770 566 2776
rect 718 2770 776 2776
rect 928 2770 986 2776
rect 1138 2770 1196 2776
rect 1348 2770 1406 2776
rect 1558 2770 1616 2776
rect 1768 2770 1826 2776
rect 1978 2770 2036 2776
rect 2188 2770 2246 2776
rect 2398 2770 2456 2776
rect 2608 2770 2666 2776
rect 2818 2770 2876 2776
rect 3028 2770 3086 2776
rect 3238 2770 3296 2776
rect 3448 2770 3506 2776
rect 3658 2770 3716 2776
rect 3868 2770 3926 2776
rect 4078 2770 4136 2776
rect 4288 2770 4346 2776
rect 4498 2770 4556 2776
rect 4708 2770 4766 2776
rect 4918 2770 4976 2776
rect 5128 2770 5186 2776
rect 5338 2770 5396 2776
rect 5548 2770 5606 2776
rect 5758 2770 5816 2776
rect -2432 2736 -2420 2770
rect -2386 2736 -2210 2770
rect -2176 2736 -2009 2770
rect -1957 2736 -1790 2770
rect -1756 2736 -1580 2770
rect -1546 2736 -1370 2770
rect -1336 2736 -1160 2770
rect -1126 2736 -950 2770
rect -916 2736 -740 2770
rect -706 2736 -539 2770
rect -487 2736 -320 2770
rect -286 2736 -110 2770
rect -76 2736 100 2770
rect 134 2736 310 2770
rect 344 2736 520 2770
rect 554 2736 730 2770
rect 764 2736 931 2770
rect 983 2736 1150 2770
rect 1184 2736 1360 2770
rect 1394 2736 1570 2770
rect 1604 2736 1780 2770
rect 1814 2736 1990 2770
rect 2024 2736 2200 2770
rect 2234 2736 2410 2770
rect 2444 2736 2620 2770
rect 2654 2736 2830 2770
rect 2864 2736 3040 2770
rect 3074 2736 3250 2770
rect 3284 2736 3460 2770
rect 3494 2736 3670 2770
rect 3704 2736 3880 2770
rect 3914 2736 4090 2770
rect 4124 2736 4300 2770
rect 4334 2736 4510 2770
rect 4544 2736 4720 2770
rect 4754 2736 4930 2770
rect 4964 2736 5140 2770
rect 5174 2736 5350 2770
rect 5384 2736 5560 2770
rect 5594 2736 5770 2770
rect 5804 2736 5816 2770
rect -2432 2730 -2374 2736
rect -2229 2724 -2157 2736
rect -2019 2718 -2009 2736
rect -1957 2718 -1947 2736
rect -1802 2730 -1744 2736
rect -1592 2730 -1534 2736
rect -1382 2730 -1324 2736
rect -1172 2730 -1114 2736
rect -962 2730 -904 2736
rect -752 2730 -694 2736
rect -549 2724 -539 2736
rect -487 2724 -477 2736
rect -332 2730 -274 2736
rect -122 2730 -64 2736
rect 88 2730 146 2736
rect 298 2730 356 2736
rect 508 2730 566 2736
rect 718 2730 776 2736
rect 921 2718 931 2736
rect 983 2718 993 2736
rect 1138 2730 1196 2736
rect 1348 2730 1406 2736
rect 1558 2730 1616 2736
rect 1768 2730 1826 2736
rect 1978 2730 2036 2736
rect 2188 2730 2246 2736
rect 2398 2730 2456 2736
rect 2608 2730 2666 2736
rect 2818 2730 2876 2736
rect 3028 2730 3086 2736
rect 3238 2730 3296 2736
rect 3448 2730 3506 2736
rect 3658 2730 3716 2736
rect 3868 2730 3926 2736
rect 4078 2730 4136 2736
rect 4288 2730 4346 2736
rect 4498 2730 4556 2736
rect 4708 2730 4766 2736
rect 4918 2730 4976 2736
rect 5128 2730 5186 2736
rect 5338 2730 5396 2736
rect 5548 2730 5606 2736
rect 5758 2730 5816 2736
rect -2336 2628 -2278 2634
rect -2126 2628 -2068 2634
rect -1916 2628 -1858 2634
rect -1706 2628 -1648 2634
rect -1496 2628 -1438 2634
rect -1293 2628 -1283 2640
rect -1231 2628 -1221 2640
rect -1076 2628 -1018 2634
rect -866 2628 -808 2634
rect -656 2628 -598 2634
rect -446 2628 -388 2634
rect -236 2628 -178 2634
rect -26 2628 32 2634
rect 184 2628 242 2634
rect 292 2628 302 2640
rect -2336 2594 -2324 2628
rect -2290 2594 -2114 2628
rect -2080 2594 -1904 2628
rect -1870 2594 -1694 2628
rect -1660 2594 -1484 2628
rect -1450 2594 -1283 2628
rect -1231 2594 -1064 2628
rect -1030 2594 -854 2628
rect -820 2594 -644 2628
rect -610 2594 -434 2628
rect -400 2594 -224 2628
rect -190 2594 -14 2628
rect 20 2594 196 2628
rect 230 2594 302 2628
rect -2336 2588 -2278 2594
rect -2126 2588 -2068 2594
rect -1916 2588 -1858 2594
rect -1706 2588 -1648 2594
rect -1496 2588 -1438 2594
rect -1293 2588 -1283 2594
rect -1231 2588 -1221 2594
rect -1076 2588 -1018 2594
rect -866 2588 -808 2594
rect -656 2588 -598 2594
rect -446 2588 -388 2594
rect -236 2588 -178 2594
rect -26 2588 32 2594
rect 184 2588 242 2594
rect 292 2588 302 2594
rect 354 2628 364 2640
rect 394 2628 452 2634
rect 604 2628 662 2634
rect 814 2628 872 2634
rect 1024 2628 1082 2634
rect 1234 2628 1292 2634
rect 1444 2628 1502 2634
rect 1647 2628 1657 2640
rect 1709 2628 1719 2640
rect 1864 2628 1922 2634
rect 2074 2628 2132 2634
rect 2284 2628 2342 2634
rect 2494 2628 2552 2634
rect 2704 2628 2762 2634
rect 2907 2628 2917 2640
rect 2969 2628 2979 2640
rect 3124 2628 3182 2634
rect 3334 2628 3392 2634
rect 3544 2628 3602 2634
rect 3754 2628 3812 2634
rect 3964 2628 4022 2634
rect 4174 2628 4232 2634
rect 4384 2628 4442 2634
rect 4594 2628 4652 2634
rect 4804 2628 4862 2634
rect 4911 2628 4921 2640
rect 354 2594 406 2628
rect 440 2594 616 2628
rect 650 2594 826 2628
rect 860 2594 1036 2628
rect 1070 2594 1246 2628
rect 1280 2594 1456 2628
rect 1490 2594 1657 2628
rect 1709 2594 1876 2628
rect 1910 2594 2086 2628
rect 2120 2594 2296 2628
rect 2330 2594 2506 2628
rect 2540 2594 2716 2628
rect 2750 2594 2917 2628
rect 2969 2594 3136 2628
rect 3170 2594 3346 2628
rect 3380 2594 3556 2628
rect 3590 2594 3766 2628
rect 3800 2594 3976 2628
rect 4010 2594 4186 2628
rect 4220 2594 4396 2628
rect 4430 2594 4606 2628
rect 4640 2594 4816 2628
rect 4850 2594 4921 2628
rect 354 2588 364 2594
rect 394 2588 452 2594
rect 604 2588 662 2594
rect 814 2588 872 2594
rect 1024 2588 1082 2594
rect 1234 2588 1292 2594
rect 1444 2588 1502 2594
rect 1647 2588 1657 2594
rect 1709 2588 1719 2594
rect 1864 2588 1922 2594
rect 2074 2588 2132 2594
rect 2284 2588 2342 2594
rect 2494 2588 2552 2594
rect 2704 2588 2762 2594
rect 2907 2588 2917 2594
rect 2969 2588 2979 2594
rect 3124 2588 3182 2594
rect 3334 2588 3392 2594
rect 3544 2588 3602 2594
rect 3754 2588 3812 2594
rect 3964 2588 4022 2594
rect 4174 2588 4232 2594
rect 4384 2588 4442 2594
rect 4594 2588 4652 2594
rect 4804 2588 4862 2594
rect 4911 2588 4921 2594
rect 4973 2628 4983 2640
rect 5014 2628 5072 2634
rect 5224 2628 5282 2634
rect 5434 2628 5492 2634
rect 5644 2628 5702 2634
rect 5854 2628 5912 2634
rect 4973 2594 5026 2628
rect 5060 2594 5236 2628
rect 5270 2594 5446 2628
rect 5480 2594 5656 2628
rect 5690 2594 5866 2628
rect 5900 2594 5912 2628
rect 4973 2588 4983 2594
rect 5014 2588 5072 2594
rect 5224 2588 5282 2594
rect 5434 2588 5492 2594
rect 5644 2588 5702 2594
rect 5854 2588 5912 2594
rect -2598 2501 -2588 2553
rect -2536 2544 -2526 2553
rect -1761 2544 -1689 2553
rect -81 2544 -9 2553
rect 1599 2544 1671 2553
rect -2536 2510 5912 2544
rect -2536 2501 -2526 2510
rect -1761 2501 -1689 2510
rect -81 2501 -9 2510
rect 1599 2501 1671 2510
rect -2598 2424 -2546 2501
rect -2598 2372 -2588 2424
rect -2536 2414 -2526 2424
rect -2391 2414 -2319 2423
rect -1551 2414 -1479 2423
rect -711 2414 -639 2423
rect 129 2414 201 2423
rect 969 2414 1041 2423
rect -2536 2380 5912 2414
rect -2536 2372 -2526 2380
rect -2391 2371 -2319 2380
rect -1551 2371 -1479 2380
rect -711 2371 -639 2380
rect 129 2371 201 2380
rect 969 2371 1041 2380
rect -2432 2330 -2374 2336
rect -2229 2330 -2157 2336
rect -2012 2330 -1954 2336
rect -1802 2330 -1744 2336
rect -1592 2330 -1534 2336
rect -1382 2330 -1324 2336
rect -1172 2330 -1114 2336
rect -962 2330 -904 2336
rect -752 2330 -694 2336
rect -549 2330 -539 2336
rect -487 2330 -477 2336
rect -332 2330 -274 2336
rect -122 2330 -64 2336
rect 88 2330 146 2336
rect 298 2330 356 2336
rect 508 2330 566 2336
rect 718 2330 776 2336
rect 928 2330 986 2336
rect 1138 2330 1196 2336
rect 1348 2330 1406 2336
rect 1558 2330 1616 2336
rect 1768 2330 1826 2336
rect 1978 2330 2036 2336
rect 2188 2330 2246 2336
rect 2398 2330 2456 2336
rect 2608 2330 2666 2336
rect 2818 2330 2876 2336
rect 3028 2330 3086 2336
rect 3238 2330 3296 2336
rect 3448 2330 3506 2336
rect 3658 2330 3716 2336
rect 3868 2330 3926 2336
rect 4078 2330 4136 2336
rect 4288 2330 4346 2336
rect 4498 2330 4556 2336
rect 4708 2330 4766 2336
rect 4918 2330 4976 2336
rect 5128 2330 5186 2336
rect 5338 2330 5396 2336
rect 5548 2330 5606 2336
rect 5758 2330 5816 2336
rect -2432 2296 -2420 2330
rect -2386 2296 -2210 2330
rect -2176 2296 -2009 2330
rect -1957 2296 -1790 2330
rect -1756 2296 -1580 2330
rect -1546 2296 -1370 2330
rect -1336 2296 -1160 2330
rect -1126 2296 -950 2330
rect -916 2296 -740 2330
rect -706 2296 -539 2330
rect -487 2296 -320 2330
rect -286 2296 -110 2330
rect -76 2296 100 2330
rect 134 2296 310 2330
rect 344 2296 520 2330
rect 554 2296 730 2330
rect 764 2296 931 2330
rect 983 2296 1150 2330
rect 1184 2296 1360 2330
rect 1394 2296 1570 2330
rect 1604 2296 1780 2330
rect 1814 2296 1990 2330
rect 2024 2296 2200 2330
rect 2234 2296 2410 2330
rect 2444 2296 2620 2330
rect 2654 2296 2830 2330
rect 2864 2296 3040 2330
rect 3074 2296 3250 2330
rect 3284 2296 3460 2330
rect 3494 2296 3670 2330
rect 3704 2296 3880 2330
rect 3914 2296 4090 2330
rect 4124 2296 4300 2330
rect 4334 2296 4510 2330
rect 4544 2296 4720 2330
rect 4754 2296 4930 2330
rect 4964 2296 5140 2330
rect 5174 2296 5350 2330
rect 5384 2296 5560 2330
rect 5594 2296 5770 2330
rect 5804 2296 5816 2330
rect -2432 2290 -2374 2296
rect -2229 2284 -2157 2296
rect -2019 2278 -2009 2296
rect -1957 2278 -1947 2296
rect -1802 2290 -1744 2296
rect -1592 2290 -1534 2296
rect -1382 2290 -1324 2296
rect -1172 2290 -1114 2296
rect -962 2290 -904 2296
rect -752 2290 -694 2296
rect -549 2284 -539 2296
rect -487 2284 -477 2296
rect -332 2290 -274 2296
rect -122 2290 -64 2296
rect 88 2290 146 2296
rect 298 2290 356 2296
rect 508 2290 566 2296
rect 718 2290 776 2296
rect 921 2278 931 2296
rect 983 2278 993 2296
rect 1138 2290 1196 2296
rect 1348 2290 1406 2296
rect 1558 2290 1616 2296
rect 1768 2290 1826 2296
rect 1978 2290 2036 2296
rect 2188 2290 2246 2296
rect 2398 2290 2456 2296
rect 2608 2290 2666 2296
rect 2818 2290 2876 2296
rect 3028 2290 3086 2296
rect 3238 2290 3296 2296
rect 3448 2290 3506 2296
rect 3658 2290 3716 2296
rect 3868 2290 3926 2296
rect 4078 2290 4136 2296
rect 4288 2290 4346 2296
rect 4498 2290 4556 2296
rect 4708 2290 4766 2296
rect 4918 2290 4976 2296
rect 5128 2290 5186 2296
rect 5338 2290 5396 2296
rect 5548 2290 5606 2296
rect 5758 2290 5816 2296
rect -2336 2188 -2278 2194
rect -2126 2188 -2068 2194
rect -1916 2188 -1858 2194
rect -1706 2188 -1648 2194
rect -1496 2188 -1438 2194
rect -1293 2188 -1283 2200
rect -1231 2188 -1221 2200
rect -1076 2188 -1018 2194
rect -866 2188 -808 2194
rect -656 2188 -598 2194
rect -446 2188 -388 2194
rect -236 2188 -178 2194
rect -26 2188 32 2194
rect 184 2188 242 2194
rect 292 2188 302 2200
rect -2336 2154 -2324 2188
rect -2290 2154 -2114 2188
rect -2080 2154 -1904 2188
rect -1870 2154 -1694 2188
rect -1660 2154 -1484 2188
rect -1450 2154 -1283 2188
rect -1231 2154 -1064 2188
rect -1030 2154 -854 2188
rect -820 2154 -644 2188
rect -610 2154 -434 2188
rect -400 2154 -224 2188
rect -190 2154 -14 2188
rect 20 2154 196 2188
rect 230 2154 302 2188
rect -2336 2148 -2278 2154
rect -2126 2148 -2068 2154
rect -1916 2148 -1858 2154
rect -1706 2148 -1648 2154
rect -1496 2148 -1438 2154
rect -1293 2148 -1283 2154
rect -1231 2148 -1221 2154
rect -1076 2148 -1018 2154
rect -866 2148 -808 2154
rect -656 2148 -598 2154
rect -446 2148 -388 2154
rect -236 2148 -178 2154
rect -26 2148 32 2154
rect 184 2148 242 2154
rect 292 2148 302 2154
rect 354 2188 364 2200
rect 394 2188 452 2194
rect 604 2188 662 2194
rect 814 2188 872 2194
rect 1024 2188 1082 2194
rect 1234 2188 1292 2194
rect 1444 2188 1502 2194
rect 1647 2188 1657 2200
rect 1709 2188 1719 2200
rect 1864 2188 1922 2194
rect 2074 2188 2132 2194
rect 2284 2188 2342 2194
rect 2494 2188 2552 2194
rect 2704 2188 2762 2194
rect 2907 2188 2917 2200
rect 2969 2188 2979 2200
rect 3124 2188 3182 2194
rect 3334 2188 3392 2194
rect 3544 2188 3602 2194
rect 3754 2188 3812 2194
rect 3964 2188 4022 2194
rect 4174 2188 4232 2194
rect 4384 2188 4442 2194
rect 4594 2188 4652 2194
rect 4804 2188 4862 2194
rect 4911 2188 4921 2200
rect 354 2154 406 2188
rect 440 2154 616 2188
rect 650 2154 826 2188
rect 860 2154 1036 2188
rect 1070 2154 1246 2188
rect 1280 2154 1456 2188
rect 1490 2154 1657 2188
rect 1709 2154 1876 2188
rect 1910 2154 2086 2188
rect 2120 2154 2296 2188
rect 2330 2154 2506 2188
rect 2540 2154 2716 2188
rect 2750 2154 2917 2188
rect 2969 2154 3136 2188
rect 3170 2154 3346 2188
rect 3380 2154 3556 2188
rect 3590 2154 3766 2188
rect 3800 2154 3976 2188
rect 4010 2154 4186 2188
rect 4220 2154 4396 2188
rect 4430 2154 4606 2188
rect 4640 2154 4816 2188
rect 4850 2154 4921 2188
rect 354 2148 364 2154
rect 394 2148 452 2154
rect 604 2148 662 2154
rect 814 2148 872 2154
rect 1024 2148 1082 2154
rect 1234 2148 1292 2154
rect 1444 2148 1502 2154
rect 1647 2148 1657 2154
rect 1709 2148 1719 2154
rect 1864 2148 1922 2154
rect 2074 2148 2132 2154
rect 2284 2148 2342 2154
rect 2494 2148 2552 2154
rect 2704 2148 2762 2154
rect 2907 2148 2917 2154
rect 2969 2148 2979 2154
rect 3124 2148 3182 2154
rect 3334 2148 3392 2154
rect 3544 2148 3602 2154
rect 3754 2148 3812 2154
rect 3964 2148 4022 2154
rect 4174 2148 4232 2154
rect 4384 2148 4442 2154
rect 4594 2148 4652 2154
rect 4804 2148 4862 2154
rect 4911 2148 4921 2154
rect 4973 2188 4983 2200
rect 5014 2188 5072 2194
rect 5224 2188 5282 2194
rect 5434 2188 5492 2194
rect 5644 2188 5702 2194
rect 5854 2188 5912 2194
rect 4973 2154 5026 2188
rect 5060 2154 5236 2188
rect 5270 2154 5446 2188
rect 5480 2154 5656 2188
rect 5690 2154 5866 2188
rect 5900 2154 5912 2188
rect 4973 2148 4983 2154
rect 5014 2148 5072 2154
rect 5224 2148 5282 2154
rect 5434 2148 5492 2154
rect 5644 2148 5702 2154
rect 5854 2148 5912 2154
rect -2598 2061 -2588 2113
rect -2536 2104 -2526 2113
rect -2181 2104 -2109 2113
rect -1341 2104 -1269 2113
rect -501 2104 -429 2113
rect 339 2104 411 2113
rect 1179 2104 1251 2113
rect -2536 2070 5912 2104
rect -2536 2061 -2526 2070
rect -2181 2061 -2109 2070
rect -1341 2061 -1269 2070
rect -501 2061 -429 2070
rect 339 2061 411 2070
rect 1179 2061 1251 2070
rect -1971 1974 -1899 1983
rect -291 1974 -219 1983
rect 1389 1974 1461 1983
rect 6010 1974 6020 1985
rect -2432 1940 6020 1974
rect -1971 1931 -1899 1940
rect -291 1931 -219 1940
rect 1389 1931 1461 1940
rect 6010 1933 6020 1940
rect 6072 1974 6082 1985
rect 6072 1940 6088 1974
rect 6072 1933 6082 1940
rect -2432 1890 -2374 1896
rect -2222 1890 -2164 1896
rect -2012 1890 -1954 1896
rect -1802 1890 -1744 1896
rect -1592 1890 -1534 1896
rect -1382 1890 -1324 1896
rect -1172 1890 -1114 1896
rect -962 1890 -904 1896
rect -752 1890 -694 1896
rect -542 1890 -484 1896
rect -332 1890 -274 1896
rect -122 1890 -64 1896
rect 88 1890 146 1896
rect 298 1890 356 1896
rect 508 1890 566 1896
rect 718 1890 776 1896
rect 928 1890 986 1896
rect 1138 1890 1196 1896
rect 1348 1890 1406 1896
rect 1558 1890 1616 1896
rect 1768 1890 1826 1896
rect 1978 1890 2036 1896
rect 2188 1890 2246 1896
rect 2398 1890 2456 1896
rect 2608 1890 2666 1896
rect 2818 1890 2876 1896
rect 3028 1890 3086 1896
rect 3238 1890 3296 1896
rect 3448 1890 3506 1896
rect 3658 1890 3716 1896
rect 3868 1890 3926 1896
rect 4078 1890 4136 1896
rect 4288 1890 4346 1896
rect 4498 1890 4556 1896
rect 4708 1890 4766 1896
rect 4918 1890 4976 1896
rect 5128 1890 5186 1896
rect 5338 1890 5396 1896
rect 5548 1890 5606 1896
rect 5758 1890 5816 1896
rect -2432 1856 -2420 1890
rect -2386 1856 -2210 1890
rect -2176 1856 -2000 1890
rect -1966 1856 -1790 1890
rect -1756 1856 -1580 1890
rect -1546 1856 -1370 1890
rect -1336 1856 -1160 1890
rect -1126 1856 -950 1890
rect -916 1856 -740 1890
rect -706 1856 -530 1890
rect -496 1856 -320 1890
rect -286 1856 -110 1890
rect -76 1856 100 1890
rect 134 1856 310 1890
rect 344 1856 520 1890
rect 554 1856 730 1890
rect 764 1856 940 1890
rect 974 1856 1150 1890
rect 1184 1856 1360 1890
rect 1394 1856 1570 1890
rect 1604 1856 1780 1890
rect 1814 1856 1990 1890
rect 2024 1856 2200 1890
rect 2234 1856 2401 1890
rect 2453 1856 2620 1890
rect 2654 1856 2830 1890
rect 2864 1856 3040 1890
rect 3074 1856 3250 1890
rect 3284 1856 3460 1890
rect 3494 1856 3670 1890
rect 3704 1856 3871 1890
rect 3923 1856 4090 1890
rect 4124 1856 4300 1890
rect 4334 1856 4510 1890
rect 4544 1856 4720 1890
rect 4754 1856 4930 1890
rect 4964 1856 5140 1890
rect 5174 1856 5340 1890
rect 5392 1856 5560 1890
rect 5594 1856 5770 1890
rect 5804 1856 5816 1890
rect -2432 1850 -2374 1856
rect -2222 1850 -2164 1856
rect -2012 1850 -1954 1856
rect -1802 1850 -1744 1856
rect -1592 1850 -1534 1856
rect -1382 1850 -1324 1856
rect -1172 1850 -1114 1856
rect -962 1850 -904 1856
rect -752 1850 -694 1856
rect -542 1850 -484 1856
rect -332 1850 -274 1856
rect -122 1850 -64 1856
rect 88 1850 146 1856
rect 298 1850 356 1856
rect 508 1850 566 1856
rect 718 1850 776 1856
rect 928 1850 986 1856
rect 1138 1850 1196 1856
rect 1348 1850 1406 1856
rect 1558 1850 1616 1856
rect 1768 1850 1826 1856
rect 1978 1850 2036 1856
rect 2188 1850 2246 1856
rect 2391 1838 2401 1856
rect 2453 1838 2463 1856
rect 2608 1850 2666 1856
rect 2818 1850 2876 1856
rect 3028 1850 3086 1856
rect 3238 1850 3296 1856
rect 3448 1850 3506 1856
rect 3658 1850 3716 1856
rect 3861 1838 3871 1856
rect 3923 1838 3933 1856
rect 4078 1850 4136 1856
rect 4288 1850 4346 1856
rect 4498 1850 4556 1856
rect 4708 1850 4766 1856
rect 4918 1850 4976 1856
rect 5128 1850 5186 1856
rect 5330 1838 5340 1856
rect 5392 1838 5402 1856
rect 5548 1850 5606 1856
rect 5758 1850 5816 1856
rect -2336 1748 -2278 1754
rect -2126 1748 -2068 1754
rect -1916 1748 -1858 1754
rect -1706 1748 -1648 1754
rect -1496 1748 -1438 1754
rect -1293 1748 -1283 1760
rect -1231 1748 -1221 1760
rect -1076 1748 -1018 1754
rect -866 1748 -808 1754
rect -656 1748 -598 1754
rect -446 1748 -388 1754
rect -236 1748 -178 1754
rect -26 1748 32 1754
rect 184 1748 242 1754
rect 292 1748 302 1760
rect -2336 1714 -2324 1748
rect -2290 1714 -2114 1748
rect -2080 1714 -1904 1748
rect -1870 1714 -1694 1748
rect -1660 1714 -1484 1748
rect -1450 1714 -1283 1748
rect -1231 1714 -1064 1748
rect -1030 1714 -854 1748
rect -820 1714 -644 1748
rect -610 1714 -434 1748
rect -400 1714 -224 1748
rect -190 1714 -14 1748
rect 20 1714 196 1748
rect 230 1714 302 1748
rect -2336 1708 -2278 1714
rect -2126 1708 -2068 1714
rect -1916 1708 -1858 1714
rect -1706 1708 -1648 1714
rect -1496 1708 -1438 1714
rect -1293 1708 -1283 1714
rect -1231 1708 -1221 1714
rect -1076 1708 -1018 1714
rect -866 1708 -808 1714
rect -656 1708 -598 1714
rect -446 1708 -388 1714
rect -236 1708 -178 1714
rect -26 1708 32 1714
rect 184 1708 242 1714
rect 292 1708 302 1714
rect 354 1748 364 1760
rect 394 1748 452 1754
rect 604 1748 662 1754
rect 814 1748 872 1754
rect 1024 1748 1082 1754
rect 1234 1748 1292 1754
rect 1444 1748 1502 1754
rect 1647 1748 1657 1760
rect 1709 1748 1719 1760
rect 1864 1748 1922 1754
rect 2074 1748 2132 1754
rect 2284 1748 2342 1754
rect 2494 1748 2552 1754
rect 2704 1748 2762 1754
rect 2907 1748 2917 1760
rect 2969 1748 2979 1760
rect 3124 1748 3182 1754
rect 3334 1748 3392 1754
rect 3544 1748 3602 1754
rect 3754 1748 3812 1754
rect 3964 1748 4022 1754
rect 4174 1748 4232 1754
rect 4384 1748 4442 1754
rect 4594 1748 4652 1754
rect 4804 1748 4862 1754
rect 4911 1748 4921 1760
rect 354 1714 406 1748
rect 440 1714 616 1748
rect 650 1714 826 1748
rect 860 1714 1036 1748
rect 1070 1714 1246 1748
rect 1280 1714 1456 1748
rect 1490 1714 1657 1748
rect 1709 1714 1876 1748
rect 1910 1714 2086 1748
rect 2120 1714 2296 1748
rect 2330 1714 2506 1748
rect 2540 1714 2716 1748
rect 2750 1714 2917 1748
rect 2969 1714 3136 1748
rect 3170 1714 3346 1748
rect 3380 1714 3556 1748
rect 3590 1714 3766 1748
rect 3800 1714 3976 1748
rect 4010 1714 4186 1748
rect 4220 1714 4396 1748
rect 4430 1714 4606 1748
rect 4640 1714 4816 1748
rect 4850 1714 4921 1748
rect 354 1708 364 1714
rect 394 1708 452 1714
rect 604 1708 662 1714
rect 814 1708 872 1714
rect 1024 1708 1082 1714
rect 1234 1708 1292 1714
rect 1444 1708 1502 1714
rect 1647 1708 1657 1714
rect 1709 1708 1719 1714
rect 1864 1708 1922 1714
rect 2074 1708 2132 1714
rect 2284 1708 2342 1714
rect 2494 1708 2552 1714
rect 2704 1708 2762 1714
rect 2907 1708 2917 1714
rect 2969 1708 2979 1714
rect 3124 1708 3182 1714
rect 3334 1708 3392 1714
rect 3544 1708 3602 1714
rect 3754 1708 3812 1714
rect 3964 1708 4022 1714
rect 4174 1708 4232 1714
rect 4384 1708 4442 1714
rect 4594 1708 4652 1714
rect 4804 1708 4862 1714
rect 4911 1708 4921 1714
rect 4973 1748 4983 1760
rect 5014 1748 5072 1754
rect 5224 1748 5282 1754
rect 5434 1748 5492 1754
rect 5644 1748 5702 1754
rect 5854 1748 5912 1754
rect 4973 1714 5026 1748
rect 5060 1714 5236 1748
rect 5270 1714 5446 1748
rect 5480 1714 5656 1748
rect 5690 1714 5866 1748
rect 5900 1714 5912 1748
rect 4973 1708 4983 1714
rect 5014 1708 5072 1714
rect 5224 1708 5282 1714
rect 5434 1708 5492 1714
rect 5644 1708 5702 1714
rect 5854 1708 5912 1714
rect -1761 1664 -1689 1673
rect -81 1664 -9 1673
rect 1599 1664 1671 1673
rect 6010 1664 6020 1671
rect -2432 1630 6020 1664
rect -1761 1621 -1689 1630
rect -81 1621 -9 1630
rect 1599 1621 1671 1630
rect 6010 1619 6020 1630
rect 6072 1664 6082 1671
rect 6072 1630 6083 1664
rect 6072 1619 6082 1630
rect -2391 1534 -2319 1543
rect -1551 1534 -1479 1543
rect -711 1534 -639 1543
rect 129 1534 201 1543
rect 969 1534 1041 1543
rect 6010 1534 6020 1544
rect -2432 1500 6020 1534
rect -2391 1491 -2319 1500
rect -1551 1491 -1479 1500
rect -711 1491 -639 1500
rect 129 1491 201 1500
rect 969 1491 1041 1500
rect 6010 1492 6020 1500
rect 6072 1492 6082 1544
rect -2432 1450 -2374 1456
rect -2222 1450 -2164 1456
rect -2012 1450 -1954 1456
rect -1802 1450 -1744 1456
rect -1592 1450 -1534 1456
rect -1382 1450 -1324 1456
rect -1172 1450 -1114 1456
rect -962 1450 -904 1456
rect -752 1450 -694 1456
rect -542 1450 -484 1456
rect -332 1450 -274 1456
rect -122 1450 -64 1456
rect 88 1450 146 1456
rect 298 1450 356 1456
rect 508 1450 566 1456
rect 718 1450 776 1456
rect 928 1450 986 1456
rect 1138 1450 1196 1456
rect 1348 1450 1406 1456
rect 1558 1450 1616 1456
rect 1768 1450 1826 1456
rect 1978 1450 2036 1456
rect 2188 1450 2246 1456
rect 2398 1450 2456 1456
rect 2608 1450 2666 1456
rect 2818 1450 2876 1456
rect 3028 1450 3086 1456
rect 3238 1450 3296 1456
rect 3448 1450 3506 1456
rect 3658 1450 3716 1456
rect 3868 1450 3926 1456
rect 4078 1450 4136 1456
rect 4288 1450 4346 1456
rect 4498 1450 4556 1456
rect 4708 1450 4766 1456
rect 4918 1450 4976 1456
rect 5128 1450 5186 1456
rect 5338 1450 5396 1456
rect 5548 1450 5606 1456
rect 5758 1450 5816 1456
rect -2432 1416 -2420 1450
rect -2386 1416 -2210 1450
rect -2176 1416 -2000 1450
rect -1966 1416 -1790 1450
rect -1756 1416 -1580 1450
rect -1546 1416 -1370 1450
rect -1336 1416 -1160 1450
rect -1126 1416 -950 1450
rect -916 1416 -740 1450
rect -706 1416 -530 1450
rect -496 1416 -320 1450
rect -286 1416 -110 1450
rect -76 1416 100 1450
rect 134 1416 310 1450
rect 344 1416 520 1450
rect 554 1416 730 1450
rect 764 1416 940 1450
rect 974 1416 1150 1450
rect 1184 1416 1360 1450
rect 1394 1416 1570 1450
rect 1604 1416 1780 1450
rect 1814 1416 1990 1450
rect 2024 1416 2200 1450
rect 2234 1416 2401 1450
rect 2453 1416 2620 1450
rect 2654 1416 2830 1450
rect 2864 1416 3040 1450
rect 3074 1416 3250 1450
rect 3284 1416 3460 1450
rect 3494 1416 3670 1450
rect 3704 1416 3871 1450
rect 3923 1416 4090 1450
rect 4124 1416 4300 1450
rect 4334 1416 4510 1450
rect 4544 1416 4720 1450
rect 4754 1416 4930 1450
rect 4964 1416 5140 1450
rect 5174 1416 5340 1450
rect 5392 1416 5560 1450
rect 5594 1416 5770 1450
rect 5804 1416 5816 1450
rect -2432 1410 -2374 1416
rect -2222 1410 -2164 1416
rect -2012 1410 -1954 1416
rect -1802 1410 -1744 1416
rect -1592 1410 -1534 1416
rect -1382 1410 -1324 1416
rect -1172 1410 -1114 1416
rect -962 1410 -904 1416
rect -752 1410 -694 1416
rect -542 1410 -484 1416
rect -332 1410 -274 1416
rect -122 1410 -64 1416
rect 88 1410 146 1416
rect 298 1410 356 1416
rect 508 1410 566 1416
rect 718 1410 776 1416
rect 928 1410 986 1416
rect 1138 1410 1196 1416
rect 1348 1410 1406 1416
rect 1558 1410 1616 1416
rect 1768 1410 1826 1416
rect 1978 1410 2036 1416
rect 2188 1410 2246 1416
rect 2391 1398 2401 1416
rect 2453 1398 2463 1416
rect 2608 1410 2666 1416
rect 2818 1410 2876 1416
rect 3028 1410 3086 1416
rect 3238 1410 3296 1416
rect 3448 1410 3506 1416
rect 3658 1410 3716 1416
rect 3861 1398 3871 1416
rect 3923 1398 3933 1416
rect 4078 1410 4136 1416
rect 4288 1410 4346 1416
rect 4498 1410 4556 1416
rect 4708 1410 4766 1416
rect 4918 1410 4976 1416
rect 5128 1410 5186 1416
rect 5330 1398 5340 1416
rect 5392 1398 5402 1416
rect 5548 1410 5606 1416
rect 5758 1410 5816 1416
rect -2336 1308 -2278 1314
rect -2126 1308 -2068 1314
rect -1916 1308 -1858 1314
rect -1706 1308 -1648 1314
rect -1496 1308 -1438 1314
rect -1293 1308 -1283 1320
rect -1231 1308 -1221 1320
rect -1076 1308 -1018 1314
rect -866 1308 -808 1314
rect -656 1308 -598 1314
rect -446 1308 -388 1314
rect -236 1308 -178 1314
rect -26 1308 32 1314
rect 184 1308 242 1314
rect 292 1308 302 1320
rect -2336 1274 -2324 1308
rect -2290 1274 -2114 1308
rect -2080 1274 -1904 1308
rect -1870 1274 -1694 1308
rect -1660 1274 -1484 1308
rect -1450 1274 -1283 1308
rect -1231 1274 -1064 1308
rect -1030 1274 -854 1308
rect -820 1274 -644 1308
rect -610 1274 -434 1308
rect -400 1274 -224 1308
rect -190 1274 -14 1308
rect 20 1274 196 1308
rect 230 1274 302 1308
rect -2336 1268 -2278 1274
rect -2126 1268 -2068 1274
rect -1916 1268 -1858 1274
rect -1706 1268 -1648 1274
rect -1496 1268 -1438 1274
rect -1293 1268 -1283 1274
rect -1231 1268 -1221 1274
rect -1076 1268 -1018 1274
rect -866 1268 -808 1274
rect -656 1268 -598 1274
rect -446 1268 -388 1274
rect -236 1268 -178 1274
rect -26 1268 32 1274
rect 184 1268 242 1274
rect 292 1268 302 1274
rect 354 1308 364 1320
rect 394 1308 452 1314
rect 604 1308 662 1314
rect 814 1308 872 1314
rect 1024 1308 1082 1314
rect 1234 1308 1292 1314
rect 1444 1308 1502 1314
rect 1647 1308 1657 1320
rect 1709 1308 1719 1320
rect 1864 1308 1922 1314
rect 2074 1308 2132 1314
rect 2284 1308 2342 1314
rect 2494 1308 2552 1314
rect 2704 1308 2762 1314
rect 2907 1308 2917 1320
rect 2969 1308 2979 1320
rect 3124 1308 3182 1314
rect 3334 1308 3392 1314
rect 3544 1308 3602 1314
rect 3754 1308 3812 1314
rect 3964 1308 4022 1314
rect 4174 1308 4232 1314
rect 4384 1308 4442 1314
rect 4594 1308 4652 1314
rect 4804 1308 4862 1314
rect 4911 1308 4921 1320
rect 354 1274 406 1308
rect 440 1274 616 1308
rect 650 1274 826 1308
rect 860 1274 1036 1308
rect 1070 1274 1246 1308
rect 1280 1274 1456 1308
rect 1490 1274 1657 1308
rect 1709 1274 1876 1308
rect 1910 1274 2086 1308
rect 2120 1274 2296 1308
rect 2330 1274 2506 1308
rect 2540 1274 2716 1308
rect 2750 1274 2917 1308
rect 2969 1274 3136 1308
rect 3170 1274 3346 1308
rect 3380 1274 3556 1308
rect 3590 1274 3766 1308
rect 3800 1274 3976 1308
rect 4010 1274 4186 1308
rect 4220 1274 4396 1308
rect 4430 1274 4606 1308
rect 4640 1274 4816 1308
rect 4850 1274 4921 1308
rect 354 1268 364 1274
rect 394 1268 452 1274
rect 604 1268 662 1274
rect 814 1268 872 1274
rect 1024 1268 1082 1274
rect 1234 1268 1292 1274
rect 1444 1268 1502 1274
rect 1647 1268 1657 1274
rect 1709 1268 1719 1274
rect 1864 1268 1922 1274
rect 2074 1268 2132 1274
rect 2284 1268 2342 1274
rect 2494 1268 2552 1274
rect 2704 1268 2762 1274
rect 2907 1268 2917 1274
rect 2969 1268 2979 1274
rect 3124 1268 3182 1274
rect 3334 1268 3392 1274
rect 3544 1268 3602 1274
rect 3754 1268 3812 1274
rect 3964 1268 4022 1274
rect 4174 1268 4232 1274
rect 4384 1268 4442 1274
rect 4594 1268 4652 1274
rect 4804 1268 4862 1274
rect 4911 1268 4921 1274
rect 4973 1308 4983 1320
rect 5014 1308 5072 1314
rect 5224 1308 5282 1314
rect 5434 1308 5492 1314
rect 5644 1308 5702 1314
rect 5854 1308 5912 1314
rect 4973 1274 5026 1308
rect 5060 1274 5236 1308
rect 5270 1274 5446 1308
rect 5480 1274 5656 1308
rect 5690 1274 5866 1308
rect 5900 1274 5912 1308
rect 4973 1268 4983 1274
rect 5014 1268 5072 1274
rect 5224 1268 5282 1274
rect 5434 1268 5492 1274
rect 5644 1268 5702 1274
rect 5854 1268 5912 1274
rect -2181 1224 -2109 1233
rect -1341 1224 -1269 1233
rect -501 1224 -429 1233
rect 339 1224 411 1233
rect 1179 1224 1251 1233
rect 6010 1224 6020 1233
rect -2432 1190 6020 1224
rect -2181 1181 -2109 1190
rect -1341 1181 -1269 1190
rect -501 1181 -429 1190
rect 339 1181 411 1190
rect 1179 1181 1251 1190
rect 6010 1181 6020 1190
rect 6072 1181 6082 1233
rect -2598 1051 -2588 1103
rect -2536 1094 -2526 1103
rect -1971 1094 -1899 1103
rect -291 1094 -219 1103
rect 1389 1094 1461 1103
rect -2536 1060 5912 1094
rect -2536 1051 -2526 1060
rect -1971 1051 -1899 1060
rect -291 1051 -219 1060
rect 1389 1051 1461 1060
rect -2432 1010 -2374 1016
rect -2229 1010 -2157 1016
rect -2012 1010 -1954 1016
rect -1802 1010 -1744 1016
rect -1592 1010 -1534 1016
rect -1382 1010 -1324 1016
rect -1172 1010 -1114 1016
rect -962 1010 -904 1016
rect -752 1010 -694 1016
rect -549 1010 -539 1016
rect -487 1010 -477 1016
rect -332 1010 -274 1016
rect -122 1010 -64 1016
rect 88 1010 146 1016
rect 298 1010 356 1016
rect 508 1010 566 1016
rect 718 1010 776 1016
rect 928 1010 986 1016
rect 1138 1010 1196 1016
rect 1348 1010 1406 1016
rect 1558 1010 1616 1016
rect 1768 1010 1826 1016
rect 1978 1010 2036 1016
rect 2188 1010 2246 1016
rect 2398 1010 2456 1016
rect 2608 1010 2666 1016
rect 2818 1010 2876 1016
rect 3028 1010 3086 1016
rect 3238 1010 3296 1016
rect 3448 1010 3506 1016
rect 3658 1010 3716 1016
rect 3868 1010 3926 1016
rect 4078 1010 4136 1016
rect 4288 1010 4346 1016
rect 4498 1010 4556 1016
rect 4708 1010 4766 1016
rect 4918 1010 4976 1016
rect 5128 1010 5186 1016
rect 5338 1010 5396 1016
rect 5548 1010 5606 1016
rect 5758 1010 5816 1016
rect -2432 976 -2420 1010
rect -2386 976 -2210 1010
rect -2176 976 -2009 1010
rect -1957 976 -1790 1010
rect -1756 976 -1580 1010
rect -1546 976 -1370 1010
rect -1336 976 -1160 1010
rect -1126 976 -950 1010
rect -916 976 -740 1010
rect -706 976 -539 1010
rect -487 976 -320 1010
rect -286 976 -110 1010
rect -76 976 100 1010
rect 134 976 310 1010
rect 344 976 520 1010
rect 554 976 730 1010
rect 764 976 931 1010
rect 983 976 1150 1010
rect 1184 976 1360 1010
rect 1394 976 1570 1010
rect 1604 976 1780 1010
rect 1814 976 1990 1010
rect 2024 976 2200 1010
rect 2234 976 2410 1010
rect 2444 976 2620 1010
rect 2654 976 2830 1010
rect 2864 976 3040 1010
rect 3074 976 3250 1010
rect 3284 976 3460 1010
rect 3494 976 3670 1010
rect 3704 976 3880 1010
rect 3914 976 4090 1010
rect 4124 976 4300 1010
rect 4334 976 4510 1010
rect 4544 976 4720 1010
rect 4754 976 4930 1010
rect 4964 976 5140 1010
rect 5174 976 5350 1010
rect 5384 976 5560 1010
rect 5594 976 5770 1010
rect 5804 976 5816 1010
rect -2432 970 -2374 976
rect -2229 964 -2157 976
rect -2019 958 -2009 976
rect -1957 958 -1947 976
rect -1802 970 -1744 976
rect -1592 970 -1534 976
rect -1382 970 -1324 976
rect -1172 970 -1114 976
rect -962 970 -904 976
rect -752 970 -694 976
rect -549 964 -539 976
rect -487 964 -477 976
rect -332 970 -274 976
rect -122 970 -64 976
rect 88 970 146 976
rect 298 970 356 976
rect 508 970 566 976
rect 718 970 776 976
rect 921 958 931 976
rect 983 958 993 976
rect 1138 970 1196 976
rect 1348 970 1406 976
rect 1558 970 1616 976
rect 1768 970 1826 976
rect 1978 970 2036 976
rect 2188 970 2246 976
rect 2398 970 2456 976
rect 2608 970 2666 976
rect 2818 970 2876 976
rect 3028 970 3086 976
rect 3238 970 3296 976
rect 3448 970 3506 976
rect 3658 970 3716 976
rect 3868 970 3926 976
rect 4078 970 4136 976
rect 4288 970 4346 976
rect 4498 970 4556 976
rect 4708 970 4766 976
rect 4918 970 4976 976
rect 5128 970 5186 976
rect 5338 970 5396 976
rect 5548 970 5606 976
rect 5758 970 5816 976
rect -2336 868 -2278 874
rect -2126 868 -2068 874
rect -1916 868 -1858 874
rect -1706 868 -1648 874
rect -1496 868 -1438 874
rect -1293 868 -1283 880
rect -1231 868 -1221 880
rect -1076 868 -1018 874
rect -866 868 -808 874
rect -656 868 -598 874
rect -446 868 -388 874
rect -236 868 -178 874
rect -26 868 32 874
rect 184 868 242 874
rect 292 868 302 880
rect -2336 834 -2324 868
rect -2290 834 -2114 868
rect -2080 834 -1904 868
rect -1870 834 -1694 868
rect -1660 834 -1484 868
rect -1450 834 -1283 868
rect -1231 834 -1064 868
rect -1030 834 -854 868
rect -820 834 -644 868
rect -610 834 -434 868
rect -400 834 -224 868
rect -190 834 -14 868
rect 20 834 196 868
rect 230 834 302 868
rect -2336 828 -2278 834
rect -2126 828 -2068 834
rect -1916 828 -1858 834
rect -1706 828 -1648 834
rect -1496 828 -1438 834
rect -1293 828 -1283 834
rect -1231 828 -1221 834
rect -1076 828 -1018 834
rect -866 828 -808 834
rect -656 828 -598 834
rect -446 828 -388 834
rect -236 828 -178 834
rect -26 828 32 834
rect 184 828 242 834
rect 292 828 302 834
rect 354 868 364 880
rect 394 868 452 874
rect 604 868 662 874
rect 814 868 872 874
rect 1024 868 1082 874
rect 1234 868 1292 874
rect 1444 868 1502 874
rect 1647 868 1657 880
rect 1709 868 1719 880
rect 1864 868 1922 874
rect 2074 868 2132 874
rect 2284 868 2342 874
rect 2494 868 2552 874
rect 2704 868 2762 874
rect 2907 868 2917 880
rect 2969 868 2979 880
rect 3124 868 3182 874
rect 3334 868 3392 874
rect 3544 868 3602 874
rect 3754 868 3812 874
rect 3964 868 4022 874
rect 4174 868 4232 874
rect 4384 868 4442 874
rect 4594 868 4652 874
rect 4804 868 4862 874
rect 4911 868 4921 880
rect 354 834 406 868
rect 440 834 616 868
rect 650 834 826 868
rect 860 834 1036 868
rect 1070 834 1246 868
rect 1280 834 1456 868
rect 1490 834 1657 868
rect 1709 834 1876 868
rect 1910 834 2086 868
rect 2120 834 2296 868
rect 2330 834 2506 868
rect 2540 834 2716 868
rect 2750 834 2917 868
rect 2969 834 3136 868
rect 3170 834 3346 868
rect 3380 834 3556 868
rect 3590 834 3766 868
rect 3800 834 3976 868
rect 4010 834 4186 868
rect 4220 834 4396 868
rect 4430 834 4606 868
rect 4640 834 4816 868
rect 4850 834 4921 868
rect 354 828 364 834
rect 394 828 452 834
rect 604 828 662 834
rect 814 828 872 834
rect 1024 828 1082 834
rect 1234 828 1292 834
rect 1444 828 1502 834
rect 1647 828 1657 834
rect 1709 828 1719 834
rect 1864 828 1922 834
rect 2074 828 2132 834
rect 2284 828 2342 834
rect 2494 828 2552 834
rect 2704 828 2762 834
rect 2907 828 2917 834
rect 2969 828 2979 834
rect 3124 828 3182 834
rect 3334 828 3392 834
rect 3544 828 3602 834
rect 3754 828 3812 834
rect 3964 828 4022 834
rect 4174 828 4232 834
rect 4384 828 4442 834
rect 4594 828 4652 834
rect 4804 828 4862 834
rect 4911 828 4921 834
rect 4973 868 4983 880
rect 5014 868 5072 874
rect 5224 868 5282 874
rect 5434 868 5492 874
rect 5644 868 5702 874
rect 5854 868 5912 874
rect 4973 834 5026 868
rect 5060 834 5236 868
rect 5270 834 5446 868
rect 5480 834 5656 868
rect 5690 834 5866 868
rect 5900 834 5912 868
rect 4973 828 4983 834
rect 5014 828 5072 834
rect 5224 828 5282 834
rect 5434 828 5492 834
rect 5644 828 5702 834
rect 5854 828 5912 834
rect -2845 733 -2704 745
rect -2598 741 -2588 793
rect -2536 784 -2526 793
rect -1761 784 -1689 793
rect -81 784 -9 793
rect 1599 784 1671 793
rect -2536 750 5912 784
rect -2536 741 -2526 750
rect -1761 741 -1689 750
rect -81 741 -9 750
rect 1599 741 1671 750
rect 6186 745 6192 4180
rect 6226 4144 6322 4180
rect 6226 4092 6229 4144
rect 6281 4092 6322 4144
rect 6226 4003 6322 4092
rect 6226 3951 6229 4003
rect 6281 3951 6322 4003
rect 6226 3862 6322 3951
rect 6226 3810 6229 3862
rect 6281 3810 6322 3862
rect 6226 3721 6322 3810
rect 6226 3669 6229 3721
rect 6281 3669 6322 3721
rect 6226 3580 6322 3669
rect 6612 3663 6682 5573
rect 6831 5403 6889 5409
rect 6750 5173 6784 5371
rect 6831 5369 6843 5403
rect 6877 5369 6889 5403
rect 6831 5363 6889 5369
rect 6843 5217 6877 5363
rect 6985 5313 7019 5573
rect 6973 5307 7031 5313
rect 6973 5273 6985 5307
rect 7019 5273 7031 5307
rect 6973 5267 7031 5273
rect 6831 5211 6889 5217
rect 6831 5177 6843 5211
rect 6877 5177 6889 5211
rect 6729 5121 6739 5173
rect 6791 5121 6801 5173
rect 6831 5171 6889 5177
rect 6750 4021 6784 5121
rect 6843 5025 6877 5171
rect 6985 5121 7019 5267
rect 7078 5173 7112 5275
rect 7060 5121 7070 5173
rect 7122 5121 7132 5173
rect 6973 5115 7031 5121
rect 6973 5081 6985 5115
rect 7019 5081 7031 5115
rect 6973 5075 7031 5081
rect 6831 5019 6889 5025
rect 6831 4985 6843 5019
rect 6877 4985 6889 5019
rect 6831 4979 6889 4985
rect 6843 4833 6877 4979
rect 6985 4929 7019 5075
rect 6973 4923 7031 4929
rect 6973 4889 6985 4923
rect 7019 4889 7031 4923
rect 6973 4883 7031 4889
rect 6831 4827 6889 4833
rect 6831 4793 6843 4827
rect 6877 4793 6889 4827
rect 6831 4787 6889 4793
rect 6843 4641 6877 4787
rect 6985 4737 7019 4883
rect 6973 4731 7031 4737
rect 6973 4697 6985 4731
rect 7019 4697 7031 4731
rect 6973 4691 7031 4697
rect 6831 4635 6889 4641
rect 6831 4601 6843 4635
rect 6877 4601 6889 4635
rect 6831 4595 6889 4601
rect 6843 4497 6877 4595
rect 6985 4545 7019 4691
rect 6973 4539 7031 4545
rect 6973 4505 6985 4539
rect 7019 4505 7031 4539
rect 6973 4499 7031 4505
rect 6825 4445 6835 4497
rect 6887 4445 6897 4497
rect 6831 4443 6889 4445
rect 6831 4409 6843 4443
rect 6877 4409 6889 4443
rect 6831 4403 6889 4409
rect 6843 4257 6877 4403
rect 6985 4353 7019 4499
rect 6973 4347 7031 4353
rect 6973 4313 6985 4347
rect 7019 4313 7031 4347
rect 6973 4307 7031 4313
rect 6831 4251 6889 4257
rect 6831 4217 6843 4251
rect 6877 4217 6889 4251
rect 6831 4211 6889 4217
rect 6843 4065 6877 4211
rect 6985 4161 7019 4307
rect 6973 4155 7031 4161
rect 6973 4121 6985 4155
rect 7019 4121 7031 4155
rect 6973 4115 7031 4121
rect 6831 4059 6889 4065
rect 6831 4025 6843 4059
rect 6877 4025 6889 4059
rect 6731 3969 6741 4021
rect 6793 3969 6803 4021
rect 6831 4019 6889 4025
rect 6750 3961 6784 3969
rect 6843 3873 6877 4019
rect 6985 3969 7019 4115
rect 7078 4021 7112 5121
rect 7060 3969 7070 4021
rect 7122 3969 7132 4021
rect 6973 3963 7031 3969
rect 6973 3929 6985 3963
rect 7019 3929 7031 3963
rect 6973 3923 7031 3929
rect 6831 3867 6889 3873
rect 6831 3833 6843 3867
rect 6877 3833 6889 3867
rect 7078 3865 7112 3969
rect 6831 3827 6889 3833
rect 6612 3657 7130 3663
rect 6612 3623 6744 3657
rect 7118 3623 7130 3657
rect 6612 3617 7130 3623
rect 6612 3587 6682 3617
rect 6226 3528 6229 3580
rect 6281 3528 6322 3580
rect 6226 3439 6322 3528
rect 6226 3387 6229 3439
rect 6281 3387 6322 3439
rect 6226 3298 6322 3387
rect 6226 3246 6229 3298
rect 6281 3246 6322 3298
rect 6226 3157 6322 3246
rect 6226 3105 6229 3157
rect 6281 3105 6322 3157
rect 6226 3016 6322 3105
rect 6226 2964 6229 3016
rect 6281 2964 6322 3016
rect 6226 2875 6322 2964
rect 6226 2823 6229 2875
rect 6281 2823 6322 2875
rect 6226 2734 6322 2823
rect 6226 2682 6229 2734
rect 6281 2682 6322 2734
rect 6226 1549 6322 2682
rect 6226 1497 6229 1549
rect 6281 1497 6322 1549
rect 6226 1408 6322 1497
rect 6226 1356 6229 1408
rect 6281 1356 6322 1408
rect 6226 1267 6322 1356
rect 6226 1215 6229 1267
rect 6281 1215 6322 1267
rect 6226 1126 6322 1215
rect 6226 1074 6229 1126
rect 6281 1074 6322 1126
rect 6226 985 6322 1074
rect 6226 933 6229 985
rect 6281 933 6322 985
rect 6226 844 6322 933
rect 6226 792 6229 844
rect 6281 792 6322 844
rect 6226 745 6322 792
rect 6186 733 6322 745
rect -1297 463 -1283 567
rect -1231 463 302 567
rect 354 463 1657 567
rect 1709 463 2917 567
rect 2969 463 4921 567
rect 4973 463 4983 567
rect -1297 462 4983 463
rect 1032 289 1042 303
rect 218 255 1042 289
rect 1032 251 1042 255
rect 1094 289 1104 303
rect 2375 289 2385 303
rect 1094 255 2385 289
rect 1094 251 1104 255
rect 2375 251 2385 255
rect 2437 289 2447 303
rect 2437 255 3208 289
rect 2437 251 2447 255
rect 174 205 232 211
rect 292 205 302 211
rect 174 171 186 205
rect 220 171 302 205
rect 174 165 232 171
rect 292 159 302 171
rect 354 205 424 211
rect 558 205 616 211
rect 750 205 808 211
rect 942 205 1000 211
rect 1134 205 1192 211
rect 1326 205 1384 211
rect 1518 205 1576 211
rect 1647 205 1657 211
rect 354 171 378 205
rect 412 171 570 205
rect 604 171 762 205
rect 796 171 954 205
rect 988 171 1146 205
rect 1180 171 1338 205
rect 1372 171 1530 205
rect 1564 171 1657 205
rect 354 165 424 171
rect 558 165 616 171
rect 750 165 808 171
rect 942 165 1000 171
rect 1134 165 1192 171
rect 1326 165 1384 171
rect 1518 165 1576 171
rect 354 159 364 165
rect 1647 159 1657 171
rect 1709 205 1768 211
rect 1902 205 1960 211
rect 2094 205 2152 211
rect 2286 205 2344 211
rect 2478 205 2536 211
rect 2670 205 2728 211
rect 2862 205 2917 211
rect 1709 171 1722 205
rect 1756 171 1914 205
rect 1948 171 2106 205
rect 2140 171 2298 205
rect 2332 171 2490 205
rect 2524 171 2682 205
rect 2716 171 2874 205
rect 2908 171 2917 205
rect 1709 165 1768 171
rect 1902 165 1960 171
rect 2094 165 2152 171
rect 2286 165 2344 171
rect 2478 165 2536 171
rect 2670 165 2728 171
rect 2862 165 2917 171
rect 1709 159 1719 165
rect 2907 159 2917 165
rect 2969 205 2979 211
rect 3054 205 3112 211
rect 3246 205 3304 211
rect 2969 171 3066 205
rect 3100 171 3258 205
rect 3292 171 3304 205
rect 2969 159 2979 171
rect 3054 165 3112 171
rect 3246 165 3304 171
rect 270 63 328 69
rect 462 63 520 69
rect 654 63 712 69
rect 846 63 904 69
rect 1038 63 1096 69
rect 1230 63 1288 69
rect 1422 63 1480 69
rect 1614 63 1672 69
rect 1806 63 1864 69
rect 1998 63 2056 69
rect 2190 63 2248 69
rect 2382 63 2440 69
rect 2574 63 2632 69
rect 2766 63 2824 69
rect 2958 63 3016 69
rect 3150 63 3208 69
rect 270 29 282 63
rect 316 29 474 63
rect 508 29 666 63
rect 700 29 858 63
rect 892 29 1050 63
rect 1084 29 1242 63
rect 1276 29 1434 63
rect 1468 29 1626 63
rect 1660 29 1818 63
rect 1852 29 2010 63
rect 2044 29 2202 63
rect 2236 29 2394 63
rect 2428 29 2586 63
rect 2620 29 2778 63
rect 2812 29 2970 63
rect 3004 29 3162 63
rect 3196 29 3208 63
rect 270 23 328 29
rect 462 23 520 29
rect 654 23 712 29
rect 846 23 904 29
rect 1038 23 1096 29
rect 1230 23 1288 29
rect 1422 23 1480 29
rect 1614 23 1672 29
rect 1806 23 1864 29
rect 1998 23 2056 29
rect 2190 23 2248 29
rect 2382 23 2440 29
rect 2574 23 2632 29
rect 2766 23 2824 29
rect 2958 23 3016 29
rect 3150 23 3208 29
rect -3246 -114 6607 -82
rect -3246 -115 5523 -114
rect -3246 -167 -2798 -115
rect -2746 -167 -2657 -115
rect -2605 -167 -2516 -115
rect -2464 -167 -2375 -115
rect -2323 -167 -2234 -115
rect -2182 -167 -2093 -115
rect -2041 -123 5523 -115
rect -2041 -157 72 -123
rect 3406 -157 5523 -123
rect -2041 -166 5523 -157
rect 5575 -166 5664 -114
rect 5716 -166 5805 -114
rect 5857 -166 5946 -114
rect 5998 -166 6087 -114
rect 6139 -166 6228 -114
rect 6280 -166 6607 -114
rect -2041 -167 6607 -166
rect -3246 -193 6607 -167
<< via1 >>
rect 1156 9738 1208 9790
rect 1156 9597 1208 9649
rect 1156 9456 1208 9508
rect 1156 9315 1208 9367
rect 1156 9174 1208 9226
rect 1576 9268 1628 9320
rect 1397 9102 1449 9154
rect 1487 8982 1539 8991
rect 1487 8948 1497 8982
rect 1497 8948 1531 8982
rect 1531 8948 1539 8982
rect 1487 8939 1539 8948
rect 1576 8982 1628 8991
rect 1576 8948 1599 8982
rect 1599 8948 1628 8982
rect 1576 8939 1628 8948
rect 1389 8312 1441 8322
rect 1389 8278 1397 8312
rect 1397 8278 1431 8312
rect 1431 8278 1441 8312
rect 1389 8270 1441 8278
rect 2003 9364 2055 9372
rect 2003 9330 2016 9364
rect 2016 9330 2050 9364
rect 2050 9330 2055 9364
rect 2003 9320 2055 9330
rect 2003 9258 2055 9268
rect 2003 9224 2015 9258
rect 2015 9224 2049 9258
rect 2049 9224 2055 9258
rect 2003 9216 2055 9224
rect 1823 9102 1875 9154
rect 2244 9740 2296 9792
rect 2244 9599 2296 9651
rect 2244 9458 2296 9510
rect 2244 9317 2296 9369
rect 2244 9176 2296 9228
rect 1823 8982 1875 8991
rect 1823 8948 1854 8982
rect 1854 8948 1875 8982
rect 1823 8939 1875 8948
rect 1912 8982 1964 8991
rect 1912 8948 1921 8982
rect 1921 8948 1955 8982
rect 1955 8948 1964 8982
rect 1912 8939 1964 8948
rect 2013 8313 2065 8323
rect 2013 8279 2022 8313
rect 2022 8279 2056 8313
rect 2056 8279 2065 8313
rect 2013 8271 2065 8279
rect -1286 8023 -1234 8041
rect 287 8023 339 8041
rect 3230 8023 3282 8041
rect 4699 8023 4751 8041
rect -1286 7989 -1234 8023
rect 287 7989 339 8023
rect 3230 7989 3282 8023
rect 4699 7989 4751 8023
rect -3662 7529 -3610 7581
rect -3331 7529 -3279 7581
rect -3423 6668 -3371 6720
rect -3660 6379 -3608 6431
rect -3331 6379 -3279 6431
rect 1970 7878 2022 7930
rect -1286 7776 -1234 7828
rect 287 7794 296 7828
rect 296 7794 330 7828
rect 330 7794 339 7828
rect 3230 7794 3236 7828
rect 3236 7794 3270 7828
rect 3270 7794 3282 7828
rect 4699 7794 4706 7828
rect 4706 7794 4740 7828
rect 4740 7794 4751 7828
rect 287 7776 339 7794
rect 3230 7776 3282 7794
rect 4699 7776 4751 7794
rect 2401 7652 2453 7704
rect 3871 7652 3923 7704
rect 5340 7652 5392 7704
rect 1970 7550 2022 7602
rect 1458 7348 1510 7400
rect -1286 7244 -1234 7296
rect 287 7262 298 7296
rect 298 7262 332 7296
rect 332 7262 339 7296
rect 3230 7262 3238 7296
rect 3238 7262 3272 7296
rect 3272 7262 3282 7296
rect 4699 7262 4708 7296
rect 4708 7262 4742 7296
rect 4742 7262 4751 7296
rect 287 7244 339 7262
rect 3230 7244 3282 7262
rect 4699 7244 4751 7262
rect -2009 7120 -1957 7172
rect -539 7120 -487 7172
rect 931 7120 983 7172
rect 1458 7018 1510 7070
rect 931 6793 983 6845
rect 1970 6793 2022 6845
rect -3072 6668 -3020 6720
rect -2009 6668 -1957 6720
rect -1379 6668 -1327 6720
rect -539 6668 -487 6720
rect 301 6668 353 6720
rect 931 6668 983 6720
rect 2401 6668 2453 6720
rect 3031 6668 3083 6720
rect 3871 6668 3923 6720
rect 4711 6668 4763 6720
rect 5340 6668 5392 6720
rect 6482 6668 6534 6720
rect 1458 6536 1510 6588
rect 2401 6536 2453 6588
rect -3660 5121 -3608 5173
rect -3329 5121 -3277 5173
rect -3425 4445 -3373 4497
rect -3660 3969 -3608 4021
rect -3331 3969 -3279 4021
rect -2798 6360 -2746 6412
rect -2798 6219 -2746 6271
rect -2798 6078 -2746 6130
rect -2798 5937 -2746 5989
rect -2798 5796 -2746 5848
rect -2798 5655 -2746 5707
rect -2798 5514 -2746 5566
rect -2798 5373 -2746 5425
rect -2798 5232 -2746 5284
rect -2798 5091 -2746 5143
rect -2798 4950 -2746 5002
rect -2798 4809 -2746 4861
rect 1970 6386 2022 6438
rect 3031 6293 3083 6345
rect 4711 6293 4763 6345
rect 2401 6169 2453 6221
rect 3871 6169 3923 6221
rect 5340 6169 5392 6221
rect 1970 6076 2022 6128
rect 1458 5946 1510 5998
rect -1379 5853 -1327 5905
rect 301 5853 353 5905
rect -2009 5729 -1957 5781
rect -539 5729 -487 5781
rect 931 5729 983 5781
rect 1458 5634 1510 5686
rect 1458 5506 1510 5558
rect -1379 5413 -1327 5465
rect 301 5413 353 5465
rect -2009 5289 -1957 5341
rect -539 5289 -487 5341
rect 931 5289 983 5341
rect 1458 5193 1510 5245
rect 1970 5067 2022 5119
rect 3031 4973 3083 5025
rect 4711 4973 4763 5025
rect 2401 4849 2453 4901
rect 3871 4849 3923 4901
rect 5340 4849 5392 4901
rect 1970 4756 2022 4808
rect 6229 6360 6281 6412
rect 6229 6219 6281 6271
rect 6229 6078 6281 6130
rect 6229 5937 6281 5989
rect 6229 5796 6281 5848
rect 6229 5655 6281 5707
rect 6229 5514 6281 5566
rect 6229 5373 6281 5425
rect 6229 5232 6281 5284
rect 6229 5091 6281 5143
rect 6229 4950 6281 5002
rect 6229 4809 6281 4861
rect 6741 7529 6793 7581
rect 7072 7529 7124 7581
rect 6833 6668 6885 6720
rect 6741 6379 6793 6431
rect 7070 6379 7122 6431
rect -3072 4445 -3020 4497
rect -2009 4445 -1957 4497
rect -539 4445 -487 4497
rect 931 4445 983 4497
rect 2401 4445 2453 4497
rect 3871 4445 3923 4497
rect 5340 4445 5392 4497
rect 6482 4445 6534 4497
rect -2798 4092 -2746 4144
rect -2798 3951 -2746 4003
rect -2798 3810 -2746 3862
rect -2798 3669 -2746 3721
rect -2798 3528 -2746 3580
rect -2798 3387 -2746 3439
rect -2798 3246 -2746 3298
rect -2798 3105 -2746 3157
rect -2798 2964 -2746 3016
rect -2798 2823 -2746 2875
rect -2798 2682 -2746 2734
rect -2798 1497 -2746 1549
rect -2798 1356 -2746 1408
rect -2798 1215 -2746 1267
rect -2798 1074 -2746 1126
rect -2798 933 -2746 985
rect -2798 792 -2746 844
rect -2588 4131 -2536 4183
rect -539 4090 -487 4096
rect -2009 4056 -2000 4090
rect -2000 4056 -1966 4090
rect -1966 4056 -1957 4090
rect -539 4056 -530 4090
rect -530 4056 -496 4090
rect -496 4056 -487 4090
rect 931 4056 940 4090
rect 940 4056 974 4090
rect 974 4056 983 4090
rect -2009 4038 -1957 4056
rect -539 4044 -487 4056
rect 931 4038 983 4056
rect -1283 3948 -1231 3960
rect -1283 3914 -1274 3948
rect -1274 3914 -1240 3948
rect -1240 3914 -1231 3948
rect -1283 3908 -1231 3914
rect 302 3908 354 3960
rect 1657 3948 1709 3960
rect 2917 3948 2969 3960
rect 1657 3914 1666 3948
rect 1666 3914 1700 3948
rect 1700 3914 1709 3948
rect 2917 3914 2926 3948
rect 2926 3914 2960 3948
rect 2960 3914 2969 3948
rect 1657 3908 1709 3914
rect 2917 3908 2969 3914
rect 4921 3908 4973 3960
rect -2588 3821 -2536 3873
rect 6020 3691 6072 3743
rect 2401 3616 2410 3650
rect 2410 3616 2444 3650
rect 2444 3616 2453 3650
rect 3871 3616 3880 3650
rect 3880 3616 3914 3650
rect 3914 3616 3923 3650
rect 5340 3616 5350 3650
rect 5350 3616 5384 3650
rect 5384 3616 5392 3650
rect 2401 3598 2453 3616
rect 3871 3598 3923 3616
rect 5340 3598 5392 3616
rect -1283 3508 -1231 3520
rect -1283 3474 -1274 3508
rect -1274 3474 -1240 3508
rect -1240 3474 -1231 3508
rect -1283 3468 -1231 3474
rect 302 3468 354 3520
rect 1657 3508 1709 3520
rect 2917 3508 2969 3520
rect 1657 3474 1666 3508
rect 1666 3474 1700 3508
rect 1700 3474 1709 3508
rect 2917 3474 2926 3508
rect 2926 3474 2960 3508
rect 2960 3474 2969 3508
rect 1657 3468 1709 3474
rect 2917 3468 2969 3474
rect 4921 3468 4973 3520
rect 6020 3381 6072 3433
rect 6020 3253 6072 3305
rect 2401 3176 2410 3210
rect 2410 3176 2444 3210
rect 2444 3176 2453 3210
rect 3871 3176 3880 3210
rect 3880 3176 3914 3210
rect 3914 3176 3923 3210
rect 5340 3176 5350 3210
rect 5350 3176 5384 3210
rect 5384 3176 5392 3210
rect 2401 3158 2453 3176
rect 3871 3158 3923 3176
rect 5340 3158 5392 3176
rect -1283 3068 -1231 3080
rect -1283 3034 -1274 3068
rect -1274 3034 -1240 3068
rect -1240 3034 -1231 3068
rect -1283 3028 -1231 3034
rect 302 3028 354 3080
rect 1657 3068 1709 3080
rect 2917 3068 2969 3080
rect 1657 3034 1666 3068
rect 1666 3034 1700 3068
rect 1700 3034 1709 3068
rect 2917 3034 2926 3068
rect 2926 3034 2960 3068
rect 2960 3034 2969 3068
rect 1657 3028 1709 3034
rect 2917 3028 2969 3034
rect 4921 3028 4973 3080
rect 6020 2939 6072 2991
rect -2588 2811 -2536 2863
rect -539 2770 -487 2776
rect -2009 2736 -2000 2770
rect -2000 2736 -1966 2770
rect -1966 2736 -1957 2770
rect -539 2736 -530 2770
rect -530 2736 -496 2770
rect -496 2736 -487 2770
rect 931 2736 940 2770
rect 940 2736 974 2770
rect 974 2736 983 2770
rect -2009 2718 -1957 2736
rect -539 2724 -487 2736
rect 931 2718 983 2736
rect -1283 2628 -1231 2640
rect -1283 2594 -1274 2628
rect -1274 2594 -1240 2628
rect -1240 2594 -1231 2628
rect -1283 2588 -1231 2594
rect 302 2588 354 2640
rect 1657 2628 1709 2640
rect 2917 2628 2969 2640
rect 1657 2594 1666 2628
rect 1666 2594 1700 2628
rect 1700 2594 1709 2628
rect 2917 2594 2926 2628
rect 2926 2594 2960 2628
rect 2960 2594 2969 2628
rect 1657 2588 1709 2594
rect 2917 2588 2969 2594
rect 4921 2588 4973 2640
rect -2588 2501 -2536 2553
rect -2588 2372 -2536 2424
rect -539 2330 -487 2336
rect -2009 2296 -2000 2330
rect -2000 2296 -1966 2330
rect -1966 2296 -1957 2330
rect -539 2296 -530 2330
rect -530 2296 -496 2330
rect -496 2296 -487 2330
rect 931 2296 940 2330
rect 940 2296 974 2330
rect 974 2296 983 2330
rect -2009 2278 -1957 2296
rect -539 2284 -487 2296
rect 931 2278 983 2296
rect -1283 2188 -1231 2200
rect -1283 2154 -1274 2188
rect -1274 2154 -1240 2188
rect -1240 2154 -1231 2188
rect -1283 2148 -1231 2154
rect 302 2148 354 2200
rect 1657 2188 1709 2200
rect 2917 2188 2969 2200
rect 1657 2154 1666 2188
rect 1666 2154 1700 2188
rect 1700 2154 1709 2188
rect 2917 2154 2926 2188
rect 2926 2154 2960 2188
rect 2960 2154 2969 2188
rect 1657 2148 1709 2154
rect 2917 2148 2969 2154
rect 4921 2148 4973 2200
rect -2588 2061 -2536 2113
rect 6020 1933 6072 1985
rect 2401 1856 2410 1890
rect 2410 1856 2444 1890
rect 2444 1856 2453 1890
rect 3871 1856 3880 1890
rect 3880 1856 3914 1890
rect 3914 1856 3923 1890
rect 5340 1856 5350 1890
rect 5350 1856 5384 1890
rect 5384 1856 5392 1890
rect 2401 1838 2453 1856
rect 3871 1838 3923 1856
rect 5340 1838 5392 1856
rect -1283 1748 -1231 1760
rect -1283 1714 -1274 1748
rect -1274 1714 -1240 1748
rect -1240 1714 -1231 1748
rect -1283 1708 -1231 1714
rect 302 1708 354 1760
rect 1657 1748 1709 1760
rect 2917 1748 2969 1760
rect 1657 1714 1666 1748
rect 1666 1714 1700 1748
rect 1700 1714 1709 1748
rect 2917 1714 2926 1748
rect 2926 1714 2960 1748
rect 2960 1714 2969 1748
rect 1657 1708 1709 1714
rect 2917 1708 2969 1714
rect 4921 1708 4973 1760
rect 6020 1619 6072 1671
rect 6020 1492 6072 1544
rect 2401 1416 2410 1450
rect 2410 1416 2444 1450
rect 2444 1416 2453 1450
rect 3871 1416 3880 1450
rect 3880 1416 3914 1450
rect 3914 1416 3923 1450
rect 5340 1416 5350 1450
rect 5350 1416 5384 1450
rect 5384 1416 5392 1450
rect 2401 1398 2453 1416
rect 3871 1398 3923 1416
rect 5340 1398 5392 1416
rect -1283 1308 -1231 1320
rect -1283 1274 -1274 1308
rect -1274 1274 -1240 1308
rect -1240 1274 -1231 1308
rect -1283 1268 -1231 1274
rect 302 1268 354 1320
rect 1657 1308 1709 1320
rect 2917 1308 2969 1320
rect 1657 1274 1666 1308
rect 1666 1274 1700 1308
rect 1700 1274 1709 1308
rect 2917 1274 2926 1308
rect 2926 1274 2960 1308
rect 2960 1274 2969 1308
rect 1657 1268 1709 1274
rect 2917 1268 2969 1274
rect 4921 1268 4973 1320
rect 6020 1181 6072 1233
rect -2588 1051 -2536 1103
rect -539 1010 -487 1016
rect -2009 976 -2000 1010
rect -2000 976 -1966 1010
rect -1966 976 -1957 1010
rect -539 976 -530 1010
rect -530 976 -496 1010
rect -496 976 -487 1010
rect 931 976 940 1010
rect 940 976 974 1010
rect 974 976 983 1010
rect -2009 958 -1957 976
rect -539 964 -487 976
rect 931 958 983 976
rect -1283 868 -1231 880
rect -1283 834 -1274 868
rect -1274 834 -1240 868
rect -1240 834 -1231 868
rect -1283 828 -1231 834
rect 302 828 354 880
rect 1657 868 1709 880
rect 2917 868 2969 880
rect 1657 834 1666 868
rect 1666 834 1700 868
rect 1700 834 1709 868
rect 2917 834 2926 868
rect 2926 834 2960 868
rect 2960 834 2969 868
rect 1657 828 1709 834
rect 2917 828 2969 834
rect 4921 828 4973 880
rect -2588 741 -2536 793
rect 6229 4092 6281 4144
rect 6229 3951 6281 4003
rect 6229 3810 6281 3862
rect 6229 3669 6281 3721
rect 6739 5121 6791 5173
rect 7070 5121 7122 5173
rect 6835 4445 6887 4497
rect 6741 3969 6793 4021
rect 7070 3969 7122 4021
rect 6229 3528 6281 3580
rect 6229 3387 6281 3439
rect 6229 3246 6281 3298
rect 6229 3105 6281 3157
rect 6229 2964 6281 3016
rect 6229 2823 6281 2875
rect 6229 2682 6281 2734
rect 6229 1497 6281 1549
rect 6229 1356 6281 1408
rect 6229 1215 6281 1267
rect 6229 1074 6281 1126
rect 6229 933 6281 985
rect 6229 792 6281 844
rect -1283 463 -1231 567
rect 302 463 354 567
rect 1657 463 1709 567
rect 2917 463 2969 567
rect 4921 463 4973 567
rect 1042 251 1094 303
rect 2385 251 2437 303
rect 302 159 354 211
rect 1657 159 1709 211
rect 2917 159 2969 211
rect -2798 -167 -2746 -115
rect -2657 -167 -2605 -115
rect -2516 -167 -2464 -115
rect -2375 -167 -2323 -115
rect -2234 -167 -2182 -115
rect -2093 -167 -2041 -115
rect 5523 -166 5575 -114
rect 5664 -166 5716 -114
rect 5805 -166 5857 -114
rect 5946 -166 5998 -114
rect 6087 -166 6139 -114
rect 6228 -166 6280 -114
<< metal2 >>
rect 1134 9790 1230 9800
rect 1134 9738 1156 9790
rect 1208 9738 1230 9790
rect 1134 9649 1230 9738
rect 1134 9597 1156 9649
rect 1208 9597 1230 9649
rect 1134 9553 1230 9597
rect -2845 9508 1230 9553
rect -2845 9456 1156 9508
rect 1208 9456 1230 9508
rect -2845 9412 1230 9456
rect -3662 7581 -3610 7591
rect -3331 7581 -3279 7591
rect -3610 7529 -3331 7581
rect -3662 7519 -3608 7529
rect -3331 7519 -3279 7529
rect -3660 6431 -3608 7519
rect -3423 6720 -3371 6730
rect -3072 6720 -3020 6730
rect -3427 6668 -3423 6720
rect -3371 6668 -3072 6720
rect -3020 6668 -3010 6720
rect -3423 6658 -3371 6668
rect -3072 6658 -3020 6668
rect -3331 6431 -3279 6441
rect -3608 6379 -3331 6431
rect -3660 5871 -3608 6379
rect -3331 6369 -3279 6379
rect -2845 6412 -2704 9412
rect 1134 9367 1230 9412
rect 2222 9792 2318 9802
rect 2222 9740 2244 9792
rect 2296 9740 2318 9792
rect 2222 9651 2318 9740
rect 2222 9599 2244 9651
rect 2296 9599 2318 9651
rect 2222 9552 2318 9599
rect 2222 9510 6322 9552
rect 2222 9458 2244 9510
rect 2296 9458 6322 9510
rect 2222 9416 6322 9458
rect 1134 9315 1156 9367
rect 1208 9315 1230 9367
rect 2003 9372 2055 9382
rect 1134 9226 1230 9315
rect 1576 9320 1628 9330
rect 1628 9268 2055 9320
rect 1576 9258 1628 9268
rect 1134 9174 1156 9226
rect 1208 9174 1230 9226
rect 2003 9206 2055 9216
rect 2222 9369 2318 9416
rect 2222 9317 2244 9369
rect 2296 9317 2318 9369
rect 2222 9228 2318 9317
rect 1134 9164 1230 9174
rect 2222 9176 2244 9228
rect 2296 9176 2318 9228
rect 2222 9166 2318 9176
rect 1397 9154 1449 9164
rect 1823 9154 1875 9164
rect 1449 9102 1823 9154
rect 1397 9092 1449 9102
rect 1823 9092 1875 9102
rect 1487 8991 1628 9001
rect 1539 8939 1576 8991
rect 1487 8929 1539 8939
rect 1576 8929 1628 8939
rect 1823 8991 1875 9001
rect 1912 8991 1964 9001
rect 1875 8939 1912 8991
rect 1823 8929 1875 8939
rect 1912 8929 1964 8939
rect 1389 8322 1441 8332
rect 2013 8323 2065 8333
rect 1379 8270 1389 8322
rect 1441 8270 1510 8322
rect 1389 8260 1510 8270
rect -1286 8041 -1234 8051
rect -1286 7828 -1234 7989
rect -1286 7296 -1234 7776
rect -1286 7234 -1234 7244
rect 287 8041 339 8051
rect 287 7828 339 7989
rect 287 7296 339 7776
rect 287 7234 339 7244
rect 1458 7400 1510 8260
rect -2009 7172 -1957 7182
rect -2009 6720 -1957 7120
rect -539 7172 -487 7182
rect -2009 6652 -1957 6668
rect -1379 6720 -1327 6727
rect -2845 6360 -2798 6412
rect -2746 6360 -2704 6412
rect -2845 6271 -2704 6360
rect -2845 6219 -2798 6271
rect -2746 6219 -2704 6271
rect -2845 6130 -2704 6219
rect -2845 6078 -2798 6130
rect -2746 6078 -2704 6130
rect -2845 5989 -2704 6078
rect -2845 5937 -2798 5989
rect -2746 5937 -2704 5989
rect -3667 5861 -3603 5871
rect -3667 5787 -3603 5797
rect -2845 5848 -2704 5937
rect -2845 5796 -2798 5848
rect -2746 5796 -2704 5848
rect -1379 5905 -1327 6668
rect -539 6720 -487 7120
rect 931 7172 983 7182
rect 931 6845 983 7120
rect -539 6652 -487 6668
rect 301 6720 353 6730
rect -3660 5173 -3608 5787
rect -2845 5707 -2704 5796
rect -2845 5655 -2798 5707
rect -2746 5655 -2704 5707
rect -2845 5566 -2704 5655
rect -2845 5514 -2798 5566
rect -2746 5514 -2704 5566
rect -2845 5425 -2704 5514
rect -2845 5373 -2798 5425
rect -2746 5373 -2704 5425
rect -2845 5284 -2704 5373
rect -2845 5232 -2798 5284
rect -2746 5232 -2704 5284
rect -3329 5173 -3277 5183
rect -3608 5121 -3329 5173
rect -3660 4021 -3608 5121
rect -3329 5111 -3277 5121
rect -2845 5143 -2704 5232
rect -2845 5091 -2798 5143
rect -2746 5091 -2704 5143
rect -2845 5002 -2704 5091
rect -2845 4950 -2798 5002
rect -2746 4950 -2704 5002
rect -2845 4861 -2704 4950
rect -2845 4809 -2798 4861
rect -2746 4809 -2704 4861
rect -3425 4497 -3373 4507
rect -3072 4497 -3020 4507
rect -3427 4445 -3425 4497
rect -3373 4445 -3072 4497
rect -3020 4445 -3010 4497
rect -3425 4435 -3373 4445
rect -3072 4435 -3020 4445
rect -2845 4144 -2704 4809
rect -2009 5781 -1957 5796
rect -2009 5341 -1957 5729
rect -1379 5465 -1327 5853
rect 301 5905 353 6668
rect 931 6720 983 6793
rect 931 6652 983 6668
rect 1458 7070 1510 7348
rect -1379 5403 -1327 5413
rect -539 5781 -487 5791
rect -2009 4497 -1957 5289
rect -2845 4092 -2798 4144
rect -2746 4092 -2704 4144
rect -3331 4021 -3279 4031
rect -3608 3969 -3331 4021
rect -3660 3959 -3608 3969
rect -3331 3959 -3279 3969
rect -2845 4003 -2704 4092
rect -2845 3951 -2798 4003
rect -2746 3951 -2704 4003
rect -2845 3862 -2704 3951
rect -2845 3810 -2798 3862
rect -2746 3810 -2704 3862
rect -2845 3721 -2704 3810
rect -2845 3669 -2798 3721
rect -2746 3669 -2704 3721
rect -2845 3580 -2704 3669
rect -2845 3528 -2798 3580
rect -2746 3528 -2704 3580
rect -2845 3439 -2704 3528
rect -2845 3387 -2798 3439
rect -2746 3387 -2704 3439
rect -2845 3298 -2704 3387
rect -2845 3246 -2798 3298
rect -2746 3246 -2704 3298
rect -2845 3157 -2704 3246
rect -2845 3105 -2798 3157
rect -2746 3105 -2704 3157
rect -2845 3016 -2704 3105
rect -2845 2964 -2798 3016
rect -2746 2964 -2704 3016
rect -2845 2875 -2704 2964
rect -2845 2823 -2798 2875
rect -2746 2823 -2704 2875
rect -2845 2734 -2704 2823
rect -2845 2682 -2798 2734
rect -2746 2682 -2704 2734
rect -2845 2672 -2704 2682
rect -2588 4183 -2536 4193
rect -2588 3873 -2536 4131
rect -2588 2863 -2536 3821
rect -2588 2553 -2536 2811
rect -2588 2424 -2536 2501
rect -2588 2113 -2536 2372
rect -2845 1549 -2704 1559
rect -2845 1497 -2798 1549
rect -2746 1497 -2704 1549
rect -2845 1408 -2704 1497
rect -2845 1356 -2798 1408
rect -2746 1356 -2704 1408
rect -2845 1267 -2704 1356
rect -2845 1215 -2798 1267
rect -2746 1215 -2704 1267
rect -2845 1126 -2704 1215
rect -2845 1074 -2798 1126
rect -2746 1074 -2704 1126
rect -2845 985 -2704 1074
rect -2845 933 -2798 985
rect -2746 933 -2704 985
rect -2845 844 -2704 933
rect -2845 792 -2798 844
rect -2746 792 -2704 844
rect -2845 -52 -2704 792
rect -2588 1103 -2536 2061
rect -2588 793 -2536 1051
rect -2009 4090 -1957 4445
rect -2009 2770 -1957 4038
rect -539 5341 -487 5729
rect 301 5465 353 5853
rect 1458 6588 1510 7018
rect 1458 5998 1510 6536
rect 301 5403 353 5413
rect 931 5781 983 5794
rect -539 4497 -487 5289
rect -539 4096 -487 4445
rect -2009 2330 -1957 2718
rect -2009 1010 -1957 2278
rect -2009 948 -1957 958
rect -1283 3960 -1231 3970
rect -1283 3520 -1231 3908
rect -1283 3080 -1231 3468
rect -1283 2640 -1231 3028
rect -1283 2200 -1231 2588
rect -1283 1760 -1231 2148
rect -1283 1320 -1231 1708
rect -2588 731 -2536 741
rect -1283 880 -1231 1268
rect -539 2776 -487 4044
rect 931 5341 983 5729
rect 931 4497 983 5289
rect 1458 5686 1510 5946
rect 1458 5558 1510 5634
rect 1458 5245 1510 5506
rect 1458 5183 1510 5193
rect 1970 8271 2013 8323
rect 2065 8271 2071 8323
rect 1970 8261 2065 8271
rect 1970 7930 2022 8261
rect 1970 7602 2022 7878
rect 3230 8041 3282 8051
rect 3230 7828 3282 7989
rect 1970 6845 2022 7550
rect 1970 6438 2022 6793
rect 2401 7704 2453 7711
rect 2401 6720 2453 7652
rect 3230 7296 3282 7776
rect 4699 8041 4751 8051
rect 4699 7828 4751 7989
rect 3230 7234 3282 7244
rect 3871 7704 3923 7714
rect 2401 6588 2453 6668
rect 2401 6526 2453 6536
rect 3031 6720 3083 6730
rect 1970 6128 2022 6386
rect 3031 6345 3083 6668
rect 3871 6720 3923 7652
rect 4699 7296 4751 7776
rect 4699 7234 4751 7244
rect 5340 7704 5392 7714
rect 3871 6657 3923 6668
rect 4711 6720 4763 6730
rect 1970 5119 2022 6076
rect 1970 4808 2022 5067
rect 1970 4746 2022 4756
rect 2401 6221 2453 6240
rect 2401 4901 2453 6169
rect 3031 5025 3083 6293
rect 4711 6345 4763 6668
rect 5340 6720 5392 7652
rect 5340 6657 5392 6668
rect 3031 4963 3083 4973
rect 3871 6221 3923 6236
rect 931 4090 983 4445
rect -539 2336 -487 2724
rect -539 1016 -487 2284
rect -539 954 -487 964
rect 302 3960 354 3970
rect 302 3520 354 3908
rect 302 3080 354 3468
rect 302 2640 354 3028
rect 302 2200 354 2588
rect 302 1760 354 2148
rect 302 1320 354 1708
rect -1283 567 -1231 828
rect -1283 457 -1231 463
rect 302 880 354 1268
rect 931 2770 983 4038
rect 2401 4497 2453 4849
rect 931 2330 983 2718
rect 931 1010 983 2278
rect 931 948 983 958
rect 1657 3960 1709 3975
rect 1657 3520 1709 3908
rect 1657 3080 1709 3468
rect 1657 2640 1709 3028
rect 1657 2200 1709 2588
rect 1657 1760 1709 2148
rect 1657 1320 1709 1708
rect 2401 3650 2453 4445
rect 3871 4901 3923 6169
rect 4711 5025 4763 6293
rect 6186 6412 6322 9416
rect 6741 7581 6793 7591
rect 7072 7581 7124 7591
rect 6793 7529 7072 7581
rect 6741 7519 6793 7529
rect 7070 7519 7124 7529
rect 6482 6720 6534 6730
rect 6833 6720 6885 6730
rect 6462 6668 6482 6720
rect 6534 6668 6833 6720
rect 6885 6668 6889 6720
rect 6482 6658 6534 6668
rect 6833 6658 6885 6668
rect 6186 6360 6229 6412
rect 6281 6360 6322 6412
rect 6741 6431 6793 6441
rect 7070 6431 7122 7519
rect 6793 6379 7070 6431
rect 6741 6369 6793 6379
rect 6186 6271 6322 6360
rect 4711 4963 4763 4973
rect 5340 6221 5392 6237
rect 3871 4497 3923 4849
rect 2401 3210 2453 3598
rect 2401 1890 2453 3158
rect 2401 1450 2453 1838
rect 2401 1388 2453 1398
rect 2917 3960 2969 3974
rect 2917 3520 2969 3908
rect 2917 3080 2969 3468
rect 2917 2640 2969 3028
rect 2917 2200 2969 2588
rect 2917 1760 2969 2148
rect 302 567 354 828
rect 302 211 354 463
rect 1657 880 1709 1268
rect 1657 567 1709 828
rect 1036 313 1100 323
rect 1036 239 1100 249
rect 302 149 354 159
rect 1657 211 1709 463
rect 2917 1320 2969 1708
rect 3871 3650 3923 4445
rect 5340 4901 5392 6169
rect 5340 4497 5392 4849
rect 3871 3210 3923 3598
rect 3871 1890 3923 3158
rect 3871 1450 3923 1838
rect 3871 1388 3923 1398
rect 4921 3960 4973 3970
rect 4921 3520 4973 3908
rect 4921 3080 4973 3468
rect 4921 2640 4973 3028
rect 4921 2200 4973 2588
rect 4921 1760 4973 2148
rect 2917 880 2969 1268
rect 2917 567 2969 828
rect 2380 313 2444 323
rect 2380 239 2444 249
rect 1657 149 1709 159
rect 2917 211 2969 463
rect 4921 1320 4973 1708
rect 5340 3650 5392 4445
rect 6186 6219 6229 6271
rect 6281 6219 6322 6271
rect 6186 6130 6322 6219
rect 6186 6078 6229 6130
rect 6281 6078 6322 6130
rect 6186 5989 6322 6078
rect 6186 5937 6229 5989
rect 6281 5937 6322 5989
rect 6186 5848 6322 5937
rect 7070 5871 7122 6379
rect 6186 5796 6229 5848
rect 6281 5796 6322 5848
rect 6186 5707 6322 5796
rect 7064 5861 7128 5871
rect 7064 5787 7128 5797
rect 6186 5655 6229 5707
rect 6281 5655 6322 5707
rect 6186 5566 6322 5655
rect 6186 5514 6229 5566
rect 6281 5514 6322 5566
rect 6186 5425 6322 5514
rect 6186 5373 6229 5425
rect 6281 5373 6322 5425
rect 6186 5284 6322 5373
rect 6186 5232 6229 5284
rect 6281 5232 6322 5284
rect 6186 5143 6322 5232
rect 6186 5091 6229 5143
rect 6281 5091 6322 5143
rect 6739 5173 6791 5183
rect 7070 5173 7122 5787
rect 6791 5121 7070 5173
rect 6739 5111 6791 5121
rect 6186 5002 6322 5091
rect 6186 4950 6229 5002
rect 6281 4950 6322 5002
rect 6186 4861 6322 4950
rect 6186 4809 6229 4861
rect 6281 4809 6322 4861
rect 6186 4144 6322 4809
rect 6482 4497 6534 4507
rect 6835 4497 6887 4507
rect 6462 4445 6482 4497
rect 6534 4445 6835 4497
rect 6887 4445 6889 4497
rect 6482 4435 6534 4445
rect 6835 4435 6887 4445
rect 6186 4092 6229 4144
rect 6281 4092 6322 4144
rect 6186 4003 6322 4092
rect 6186 3951 6229 4003
rect 6281 3951 6322 4003
rect 6741 4021 6793 4031
rect 7070 4021 7122 5121
rect 6793 3969 7070 4021
rect 6741 3959 6793 3969
rect 7070 3959 7122 3969
rect 6186 3862 6322 3951
rect 6186 3810 6229 3862
rect 6281 3810 6322 3862
rect 5340 3210 5392 3598
rect 5340 1890 5392 3158
rect 5340 1450 5392 1838
rect 5340 1388 5392 1398
rect 6020 3743 6072 3753
rect 6020 3433 6072 3691
rect 6020 3305 6072 3381
rect 6020 2991 6072 3253
rect 6020 1985 6072 2939
rect 6186 3721 6322 3810
rect 6186 3669 6229 3721
rect 6281 3669 6322 3721
rect 6186 3580 6322 3669
rect 6186 3528 6229 3580
rect 6281 3528 6322 3580
rect 6186 3439 6322 3528
rect 6186 3387 6229 3439
rect 6281 3387 6322 3439
rect 6186 3298 6322 3387
rect 6186 3246 6229 3298
rect 6281 3246 6322 3298
rect 6186 3157 6322 3246
rect 6186 3105 6229 3157
rect 6281 3105 6322 3157
rect 6186 3016 6322 3105
rect 6186 2964 6229 3016
rect 6281 2964 6322 3016
rect 6186 2875 6322 2964
rect 6186 2823 6229 2875
rect 6281 2823 6322 2875
rect 6186 2734 6322 2823
rect 6186 2682 6229 2734
rect 6281 2682 6322 2734
rect 6186 2672 6322 2682
rect 6020 1671 6072 1933
rect 6020 1544 6072 1619
rect 4921 880 4973 1268
rect 6020 1233 6072 1492
rect 6020 1168 6072 1181
rect 6186 1549 6322 1559
rect 6186 1497 6229 1549
rect 6281 1497 6322 1549
rect 6186 1408 6322 1497
rect 6186 1356 6229 1408
rect 6281 1356 6322 1408
rect 6186 1267 6322 1356
rect 6186 1215 6229 1267
rect 6281 1215 6322 1267
rect 4921 567 4973 828
rect 4921 453 4973 463
rect 6186 1126 6322 1215
rect 6186 1074 6229 1126
rect 6281 1074 6322 1126
rect 6186 985 6322 1074
rect 6186 933 6229 985
rect 6281 933 6322 985
rect 6186 844 6322 933
rect 6186 792 6229 844
rect 6281 792 6322 844
rect 2917 149 2969 159
rect -2845 -115 -2004 -52
rect 6186 -57 6322 792
rect -2845 -167 -2798 -115
rect -2746 -167 -2657 -115
rect -2605 -167 -2516 -115
rect -2464 -167 -2375 -115
rect -2323 -167 -2234 -115
rect -2182 -167 -2093 -115
rect -2041 -167 -2004 -115
rect -2845 -193 -2004 -167
rect 5496 -114 6322 -57
rect 5496 -166 5523 -114
rect 5575 -166 5664 -114
rect 5716 -166 5805 -114
rect 5857 -166 5946 -114
rect 5998 -166 6087 -114
rect 6139 -166 6228 -114
rect 6280 -166 6322 -114
rect 5496 -193 6322 -166
<< via2 >>
rect -3667 5797 -3603 5861
rect 1036 303 1100 313
rect 1036 251 1042 303
rect 1042 251 1094 303
rect 1094 251 1100 303
rect 1036 249 1100 251
rect 2380 303 2444 313
rect 2380 251 2385 303
rect 2385 251 2437 303
rect 2437 251 2444 303
rect 2380 249 2444 251
rect 7064 5797 7128 5861
<< metal3 >>
rect -3677 5861 -3593 5866
rect 7054 5861 7138 5866
rect -3677 5797 -3667 5861
rect -3603 5797 7064 5861
rect 7128 5797 7138 5861
rect -3677 5792 -3593 5797
rect 1698 492 1762 5797
rect 7054 5792 7138 5797
rect 1036 428 2444 492
rect 1036 318 1100 428
rect 2380 318 2444 428
rect 1026 313 1110 318
rect 1026 249 1036 313
rect 1100 249 1110 313
rect 1026 244 1110 249
rect 2370 313 2454 318
rect 2370 249 2380 313
rect 2444 249 2454 313
rect 2370 244 2454 249
rect 2380 242 2444 244
use current_tail  current_tail_0
timestamp 1654898484
transform 1 0 1739 0 1 118
box -1799 -310 1799 310
use input_diff_pair  input_diff_pair_0
timestamp 1654898484
transform 1 0 -2641 0 1 3815
box -1 -3081 8763 375
use latch_nmos_pair  latch_nmos_pair_0
timestamp 1654898484
transform 1 0 -2642 0 1 6069
box 0 -1320 8764 376
use latch_pmos_pair  latch_pmos_pair_0
timestamp 1654898484
transform 1 0 -2735 0 1 7455
box -59 -567 8981 604
use precharge_pmos  precharge_pmos_0
timestamp 1654898484
transform 0 1 -3736 -1 0 8008
box -52 -52 2010 586
use precharge_pmos  precharge_pmos_1
timestamp 1654898484
transform 0 1 -3734 -1 0 5598
box -52 -52 2010 586
use sky130_fd_pr__pfet_01v8_VCG74W  sky130_fd_pr__pfet_01v8_VCG74W_0
timestamp 1654898484
transform 0 -1 6931 -1 0 7029
box -1031 -319 1031 319
use sky130_fd_pr__pfet_01v8_VCG74W  sky130_fd_pr__pfet_01v8_VCG74W_1
timestamp 1654898484
transform 0 -1 6931 -1 0 4619
box -1031 -319 1031 319
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654629081
transform 0 -1 2270 1 0 8241
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1654629081
transform 0 1 1182 1 0 8241
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654629081
transform 0 1 1182 -1 0 10633
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1654629081
transform 0 -1 2270 1 0 9529
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654629081
transform 0 1 1182 -1 0 9437
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_1
timestamp 1654629081
transform 0 -1 2270 -1 0 9437
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654629081
transform 0 1 1182 -1 0 9529
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654629081
transform 0 -1 2270 1 0 9437
box -38 -48 130 592
<< labels >>
flabel metal1 1334 10724 1334 10724 5 FreeSans 400 0 0 0 outn
port 5 s
flabel metal1 2119 10721 2119 10721 1 FreeSans 400 0 0 0 outp
port 4 n
flabel metal3 1730 4459 1730 4459 1 FreeSans 400 0 0 0 clk
port 1 n
flabel metal1 -3776 8059 -3776 8059 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 -3228 -136 -3228 -136 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal2 6063 2476 6063 2476 1 FreeSans 400 0 0 0 in
port 3 n
flabel metal2 -2580 2466 -2580 2466 1 FreeSans 400 0 0 0 ip
port 2 n
<< end >>
