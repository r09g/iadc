magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -4124 172 -4066 178
rect -3704 172 -3646 178
rect -3284 172 -3226 178
rect -2864 172 -2806 178
rect -2444 172 -2386 178
rect -2024 172 -1966 178
rect -1604 172 -1546 178
rect -1184 172 -1126 178
rect -764 172 -706 178
rect -344 172 -286 178
rect 76 172 134 178
rect 496 172 554 178
rect 916 172 974 178
rect 1336 172 1394 178
rect 1756 172 1814 178
rect 2176 172 2234 178
rect 2596 172 2654 178
rect 3016 172 3074 178
rect 3436 172 3494 178
rect 3856 172 3914 178
rect -4124 138 -4112 172
rect -3704 138 -3692 172
rect -3284 138 -3272 172
rect -2864 138 -2852 172
rect -2444 138 -2432 172
rect -2024 138 -2012 172
rect -1604 138 -1592 172
rect -1184 138 -1172 172
rect -764 138 -752 172
rect -344 138 -332 172
rect 76 138 88 172
rect 496 138 508 172
rect 916 138 928 172
rect 1336 138 1348 172
rect 1756 138 1768 172
rect 2176 138 2188 172
rect 2596 138 2608 172
rect 3016 138 3028 172
rect 3436 138 3448 172
rect 3856 138 3868 172
rect -4124 132 -4066 138
rect -3704 132 -3646 138
rect -3284 132 -3226 138
rect -2864 132 -2806 138
rect -2444 132 -2386 138
rect -2024 132 -1966 138
rect -1604 132 -1546 138
rect -1184 132 -1126 138
rect -764 132 -706 138
rect -344 132 -286 138
rect 76 132 134 138
rect 496 132 554 138
rect 916 132 974 138
rect 1336 132 1394 138
rect 1756 132 1814 138
rect 2176 132 2234 138
rect 2596 132 2654 138
rect 3016 132 3074 138
rect 3436 132 3494 138
rect 3856 132 3914 138
rect -3914 -138 -3856 -132
rect -3494 -138 -3436 -132
rect -3074 -138 -3016 -132
rect -2654 -138 -2596 -132
rect -2234 -138 -2176 -132
rect -1814 -138 -1756 -132
rect -1394 -138 -1336 -132
rect -974 -138 -916 -132
rect -554 -138 -496 -132
rect -134 -138 -76 -132
rect 286 -138 344 -132
rect 706 -138 764 -132
rect 1126 -138 1184 -132
rect 1546 -138 1604 -132
rect 1966 -138 2024 -132
rect 2386 -138 2444 -132
rect 2806 -138 2864 -132
rect 3226 -138 3284 -132
rect 3646 -138 3704 -132
rect 4066 -138 4124 -132
rect -3914 -172 -3902 -138
rect -3494 -172 -3482 -138
rect -3074 -172 -3062 -138
rect -2654 -172 -2642 -138
rect -2234 -172 -2222 -138
rect -1814 -172 -1802 -138
rect -1394 -172 -1382 -138
rect -974 -172 -962 -138
rect -554 -172 -542 -138
rect -134 -172 -122 -138
rect 286 -172 298 -138
rect 706 -172 718 -138
rect 1126 -172 1138 -138
rect 1546 -172 1558 -138
rect 1966 -172 1978 -138
rect 2386 -172 2398 -138
rect 2806 -172 2818 -138
rect 3226 -172 3238 -138
rect 3646 -172 3658 -138
rect 4066 -172 4078 -138
rect -3914 -178 -3856 -172
rect -3494 -178 -3436 -172
rect -3074 -178 -3016 -172
rect -2654 -178 -2596 -172
rect -2234 -178 -2176 -172
rect -1814 -178 -1756 -172
rect -1394 -178 -1336 -172
rect -974 -178 -916 -172
rect -554 -178 -496 -172
rect -134 -178 -76 -172
rect 286 -178 344 -172
rect 706 -178 764 -172
rect 1126 -178 1184 -172
rect 1546 -178 1604 -172
rect 1966 -178 2024 -172
rect 2386 -178 2444 -172
rect 2806 -178 2864 -172
rect 3226 -178 3284 -172
rect 3646 -178 3704 -172
rect 4066 -178 4124 -172
<< pwell >>
rect -4408 -126 4408 126
<< nmos >>
rect -4320 -100 -4290 100
rect -4110 -100 -4080 100
rect -3900 -100 -3870 100
rect -3690 -100 -3660 100
rect -3480 -100 -3450 100
rect -3270 -100 -3240 100
rect -3060 -100 -3030 100
rect -2850 -100 -2820 100
rect -2640 -100 -2610 100
rect -2430 -100 -2400 100
rect -2220 -100 -2190 100
rect -2010 -100 -1980 100
rect -1800 -100 -1770 100
rect -1590 -100 -1560 100
rect -1380 -100 -1350 100
rect -1170 -100 -1140 100
rect -960 -100 -930 100
rect -750 -100 -720 100
rect -540 -100 -510 100
rect -330 -100 -300 100
rect -120 -100 -90 100
rect 90 -100 120 100
rect 300 -100 330 100
rect 510 -100 540 100
rect 720 -100 750 100
rect 930 -100 960 100
rect 1140 -100 1170 100
rect 1350 -100 1380 100
rect 1560 -100 1590 100
rect 1770 -100 1800 100
rect 1980 -100 2010 100
rect 2190 -100 2220 100
rect 2400 -100 2430 100
rect 2610 -100 2640 100
rect 2820 -100 2850 100
rect 3030 -100 3060 100
rect 3240 -100 3270 100
rect 3450 -100 3480 100
rect 3660 -100 3690 100
rect 3870 -100 3900 100
rect 4080 -100 4110 100
rect 4290 -100 4320 100
<< ndiff >>
rect -4382 85 -4320 100
rect -4382 51 -4370 85
rect -4336 51 -4320 85
rect -4382 17 -4320 51
rect -4382 -17 -4370 17
rect -4336 -17 -4320 17
rect -4382 -51 -4320 -17
rect -4382 -85 -4370 -51
rect -4336 -85 -4320 -51
rect -4382 -100 -4320 -85
rect -4290 85 -4228 100
rect -4290 51 -4274 85
rect -4240 51 -4228 85
rect -4290 17 -4228 51
rect -4290 -17 -4274 17
rect -4240 -17 -4228 17
rect -4290 -51 -4228 -17
rect -4290 -85 -4274 -51
rect -4240 -85 -4228 -51
rect -4290 -100 -4228 -85
rect -4172 85 -4110 100
rect -4172 51 -4160 85
rect -4126 51 -4110 85
rect -4172 17 -4110 51
rect -4172 -17 -4160 17
rect -4126 -17 -4110 17
rect -4172 -51 -4110 -17
rect -4172 -85 -4160 -51
rect -4126 -85 -4110 -51
rect -4172 -100 -4110 -85
rect -4080 85 -4018 100
rect -4080 51 -4064 85
rect -4030 51 -4018 85
rect -4080 17 -4018 51
rect -4080 -17 -4064 17
rect -4030 -17 -4018 17
rect -4080 -51 -4018 -17
rect -4080 -85 -4064 -51
rect -4030 -85 -4018 -51
rect -4080 -100 -4018 -85
rect -3962 85 -3900 100
rect -3962 51 -3950 85
rect -3916 51 -3900 85
rect -3962 17 -3900 51
rect -3962 -17 -3950 17
rect -3916 -17 -3900 17
rect -3962 -51 -3900 -17
rect -3962 -85 -3950 -51
rect -3916 -85 -3900 -51
rect -3962 -100 -3900 -85
rect -3870 85 -3808 100
rect -3870 51 -3854 85
rect -3820 51 -3808 85
rect -3870 17 -3808 51
rect -3870 -17 -3854 17
rect -3820 -17 -3808 17
rect -3870 -51 -3808 -17
rect -3870 -85 -3854 -51
rect -3820 -85 -3808 -51
rect -3870 -100 -3808 -85
rect -3752 85 -3690 100
rect -3752 51 -3740 85
rect -3706 51 -3690 85
rect -3752 17 -3690 51
rect -3752 -17 -3740 17
rect -3706 -17 -3690 17
rect -3752 -51 -3690 -17
rect -3752 -85 -3740 -51
rect -3706 -85 -3690 -51
rect -3752 -100 -3690 -85
rect -3660 85 -3598 100
rect -3660 51 -3644 85
rect -3610 51 -3598 85
rect -3660 17 -3598 51
rect -3660 -17 -3644 17
rect -3610 -17 -3598 17
rect -3660 -51 -3598 -17
rect -3660 -85 -3644 -51
rect -3610 -85 -3598 -51
rect -3660 -100 -3598 -85
rect -3542 85 -3480 100
rect -3542 51 -3530 85
rect -3496 51 -3480 85
rect -3542 17 -3480 51
rect -3542 -17 -3530 17
rect -3496 -17 -3480 17
rect -3542 -51 -3480 -17
rect -3542 -85 -3530 -51
rect -3496 -85 -3480 -51
rect -3542 -100 -3480 -85
rect -3450 85 -3388 100
rect -3450 51 -3434 85
rect -3400 51 -3388 85
rect -3450 17 -3388 51
rect -3450 -17 -3434 17
rect -3400 -17 -3388 17
rect -3450 -51 -3388 -17
rect -3450 -85 -3434 -51
rect -3400 -85 -3388 -51
rect -3450 -100 -3388 -85
rect -3332 85 -3270 100
rect -3332 51 -3320 85
rect -3286 51 -3270 85
rect -3332 17 -3270 51
rect -3332 -17 -3320 17
rect -3286 -17 -3270 17
rect -3332 -51 -3270 -17
rect -3332 -85 -3320 -51
rect -3286 -85 -3270 -51
rect -3332 -100 -3270 -85
rect -3240 85 -3178 100
rect -3240 51 -3224 85
rect -3190 51 -3178 85
rect -3240 17 -3178 51
rect -3240 -17 -3224 17
rect -3190 -17 -3178 17
rect -3240 -51 -3178 -17
rect -3240 -85 -3224 -51
rect -3190 -85 -3178 -51
rect -3240 -100 -3178 -85
rect -3122 85 -3060 100
rect -3122 51 -3110 85
rect -3076 51 -3060 85
rect -3122 17 -3060 51
rect -3122 -17 -3110 17
rect -3076 -17 -3060 17
rect -3122 -51 -3060 -17
rect -3122 -85 -3110 -51
rect -3076 -85 -3060 -51
rect -3122 -100 -3060 -85
rect -3030 85 -2968 100
rect -3030 51 -3014 85
rect -2980 51 -2968 85
rect -3030 17 -2968 51
rect -3030 -17 -3014 17
rect -2980 -17 -2968 17
rect -3030 -51 -2968 -17
rect -3030 -85 -3014 -51
rect -2980 -85 -2968 -51
rect -3030 -100 -2968 -85
rect -2912 85 -2850 100
rect -2912 51 -2900 85
rect -2866 51 -2850 85
rect -2912 17 -2850 51
rect -2912 -17 -2900 17
rect -2866 -17 -2850 17
rect -2912 -51 -2850 -17
rect -2912 -85 -2900 -51
rect -2866 -85 -2850 -51
rect -2912 -100 -2850 -85
rect -2820 85 -2758 100
rect -2820 51 -2804 85
rect -2770 51 -2758 85
rect -2820 17 -2758 51
rect -2820 -17 -2804 17
rect -2770 -17 -2758 17
rect -2820 -51 -2758 -17
rect -2820 -85 -2804 -51
rect -2770 -85 -2758 -51
rect -2820 -100 -2758 -85
rect -2702 85 -2640 100
rect -2702 51 -2690 85
rect -2656 51 -2640 85
rect -2702 17 -2640 51
rect -2702 -17 -2690 17
rect -2656 -17 -2640 17
rect -2702 -51 -2640 -17
rect -2702 -85 -2690 -51
rect -2656 -85 -2640 -51
rect -2702 -100 -2640 -85
rect -2610 85 -2548 100
rect -2610 51 -2594 85
rect -2560 51 -2548 85
rect -2610 17 -2548 51
rect -2610 -17 -2594 17
rect -2560 -17 -2548 17
rect -2610 -51 -2548 -17
rect -2610 -85 -2594 -51
rect -2560 -85 -2548 -51
rect -2610 -100 -2548 -85
rect -2492 85 -2430 100
rect -2492 51 -2480 85
rect -2446 51 -2430 85
rect -2492 17 -2430 51
rect -2492 -17 -2480 17
rect -2446 -17 -2430 17
rect -2492 -51 -2430 -17
rect -2492 -85 -2480 -51
rect -2446 -85 -2430 -51
rect -2492 -100 -2430 -85
rect -2400 85 -2338 100
rect -2400 51 -2384 85
rect -2350 51 -2338 85
rect -2400 17 -2338 51
rect -2400 -17 -2384 17
rect -2350 -17 -2338 17
rect -2400 -51 -2338 -17
rect -2400 -85 -2384 -51
rect -2350 -85 -2338 -51
rect -2400 -100 -2338 -85
rect -2282 85 -2220 100
rect -2282 51 -2270 85
rect -2236 51 -2220 85
rect -2282 17 -2220 51
rect -2282 -17 -2270 17
rect -2236 -17 -2220 17
rect -2282 -51 -2220 -17
rect -2282 -85 -2270 -51
rect -2236 -85 -2220 -51
rect -2282 -100 -2220 -85
rect -2190 85 -2128 100
rect -2190 51 -2174 85
rect -2140 51 -2128 85
rect -2190 17 -2128 51
rect -2190 -17 -2174 17
rect -2140 -17 -2128 17
rect -2190 -51 -2128 -17
rect -2190 -85 -2174 -51
rect -2140 -85 -2128 -51
rect -2190 -100 -2128 -85
rect -2072 85 -2010 100
rect -2072 51 -2060 85
rect -2026 51 -2010 85
rect -2072 17 -2010 51
rect -2072 -17 -2060 17
rect -2026 -17 -2010 17
rect -2072 -51 -2010 -17
rect -2072 -85 -2060 -51
rect -2026 -85 -2010 -51
rect -2072 -100 -2010 -85
rect -1980 85 -1918 100
rect -1980 51 -1964 85
rect -1930 51 -1918 85
rect -1980 17 -1918 51
rect -1980 -17 -1964 17
rect -1930 -17 -1918 17
rect -1980 -51 -1918 -17
rect -1980 -85 -1964 -51
rect -1930 -85 -1918 -51
rect -1980 -100 -1918 -85
rect -1862 85 -1800 100
rect -1862 51 -1850 85
rect -1816 51 -1800 85
rect -1862 17 -1800 51
rect -1862 -17 -1850 17
rect -1816 -17 -1800 17
rect -1862 -51 -1800 -17
rect -1862 -85 -1850 -51
rect -1816 -85 -1800 -51
rect -1862 -100 -1800 -85
rect -1770 85 -1708 100
rect -1770 51 -1754 85
rect -1720 51 -1708 85
rect -1770 17 -1708 51
rect -1770 -17 -1754 17
rect -1720 -17 -1708 17
rect -1770 -51 -1708 -17
rect -1770 -85 -1754 -51
rect -1720 -85 -1708 -51
rect -1770 -100 -1708 -85
rect -1652 85 -1590 100
rect -1652 51 -1640 85
rect -1606 51 -1590 85
rect -1652 17 -1590 51
rect -1652 -17 -1640 17
rect -1606 -17 -1590 17
rect -1652 -51 -1590 -17
rect -1652 -85 -1640 -51
rect -1606 -85 -1590 -51
rect -1652 -100 -1590 -85
rect -1560 85 -1498 100
rect -1560 51 -1544 85
rect -1510 51 -1498 85
rect -1560 17 -1498 51
rect -1560 -17 -1544 17
rect -1510 -17 -1498 17
rect -1560 -51 -1498 -17
rect -1560 -85 -1544 -51
rect -1510 -85 -1498 -51
rect -1560 -100 -1498 -85
rect -1442 85 -1380 100
rect -1442 51 -1430 85
rect -1396 51 -1380 85
rect -1442 17 -1380 51
rect -1442 -17 -1430 17
rect -1396 -17 -1380 17
rect -1442 -51 -1380 -17
rect -1442 -85 -1430 -51
rect -1396 -85 -1380 -51
rect -1442 -100 -1380 -85
rect -1350 85 -1288 100
rect -1350 51 -1334 85
rect -1300 51 -1288 85
rect -1350 17 -1288 51
rect -1350 -17 -1334 17
rect -1300 -17 -1288 17
rect -1350 -51 -1288 -17
rect -1350 -85 -1334 -51
rect -1300 -85 -1288 -51
rect -1350 -100 -1288 -85
rect -1232 85 -1170 100
rect -1232 51 -1220 85
rect -1186 51 -1170 85
rect -1232 17 -1170 51
rect -1232 -17 -1220 17
rect -1186 -17 -1170 17
rect -1232 -51 -1170 -17
rect -1232 -85 -1220 -51
rect -1186 -85 -1170 -51
rect -1232 -100 -1170 -85
rect -1140 85 -1078 100
rect -1140 51 -1124 85
rect -1090 51 -1078 85
rect -1140 17 -1078 51
rect -1140 -17 -1124 17
rect -1090 -17 -1078 17
rect -1140 -51 -1078 -17
rect -1140 -85 -1124 -51
rect -1090 -85 -1078 -51
rect -1140 -100 -1078 -85
rect -1022 85 -960 100
rect -1022 51 -1010 85
rect -976 51 -960 85
rect -1022 17 -960 51
rect -1022 -17 -1010 17
rect -976 -17 -960 17
rect -1022 -51 -960 -17
rect -1022 -85 -1010 -51
rect -976 -85 -960 -51
rect -1022 -100 -960 -85
rect -930 85 -868 100
rect -930 51 -914 85
rect -880 51 -868 85
rect -930 17 -868 51
rect -930 -17 -914 17
rect -880 -17 -868 17
rect -930 -51 -868 -17
rect -930 -85 -914 -51
rect -880 -85 -868 -51
rect -930 -100 -868 -85
rect -812 85 -750 100
rect -812 51 -800 85
rect -766 51 -750 85
rect -812 17 -750 51
rect -812 -17 -800 17
rect -766 -17 -750 17
rect -812 -51 -750 -17
rect -812 -85 -800 -51
rect -766 -85 -750 -51
rect -812 -100 -750 -85
rect -720 85 -658 100
rect -720 51 -704 85
rect -670 51 -658 85
rect -720 17 -658 51
rect -720 -17 -704 17
rect -670 -17 -658 17
rect -720 -51 -658 -17
rect -720 -85 -704 -51
rect -670 -85 -658 -51
rect -720 -100 -658 -85
rect -602 85 -540 100
rect -602 51 -590 85
rect -556 51 -540 85
rect -602 17 -540 51
rect -602 -17 -590 17
rect -556 -17 -540 17
rect -602 -51 -540 -17
rect -602 -85 -590 -51
rect -556 -85 -540 -51
rect -602 -100 -540 -85
rect -510 85 -448 100
rect -510 51 -494 85
rect -460 51 -448 85
rect -510 17 -448 51
rect -510 -17 -494 17
rect -460 -17 -448 17
rect -510 -51 -448 -17
rect -510 -85 -494 -51
rect -460 -85 -448 -51
rect -510 -100 -448 -85
rect -392 85 -330 100
rect -392 51 -380 85
rect -346 51 -330 85
rect -392 17 -330 51
rect -392 -17 -380 17
rect -346 -17 -330 17
rect -392 -51 -330 -17
rect -392 -85 -380 -51
rect -346 -85 -330 -51
rect -392 -100 -330 -85
rect -300 85 -238 100
rect -300 51 -284 85
rect -250 51 -238 85
rect -300 17 -238 51
rect -300 -17 -284 17
rect -250 -17 -238 17
rect -300 -51 -238 -17
rect -300 -85 -284 -51
rect -250 -85 -238 -51
rect -300 -100 -238 -85
rect -182 85 -120 100
rect -182 51 -170 85
rect -136 51 -120 85
rect -182 17 -120 51
rect -182 -17 -170 17
rect -136 -17 -120 17
rect -182 -51 -120 -17
rect -182 -85 -170 -51
rect -136 -85 -120 -51
rect -182 -100 -120 -85
rect -90 85 -28 100
rect -90 51 -74 85
rect -40 51 -28 85
rect -90 17 -28 51
rect -90 -17 -74 17
rect -40 -17 -28 17
rect -90 -51 -28 -17
rect -90 -85 -74 -51
rect -40 -85 -28 -51
rect -90 -100 -28 -85
rect 28 85 90 100
rect 28 51 40 85
rect 74 51 90 85
rect 28 17 90 51
rect 28 -17 40 17
rect 74 -17 90 17
rect 28 -51 90 -17
rect 28 -85 40 -51
rect 74 -85 90 -51
rect 28 -100 90 -85
rect 120 85 182 100
rect 120 51 136 85
rect 170 51 182 85
rect 120 17 182 51
rect 120 -17 136 17
rect 170 -17 182 17
rect 120 -51 182 -17
rect 120 -85 136 -51
rect 170 -85 182 -51
rect 120 -100 182 -85
rect 238 85 300 100
rect 238 51 250 85
rect 284 51 300 85
rect 238 17 300 51
rect 238 -17 250 17
rect 284 -17 300 17
rect 238 -51 300 -17
rect 238 -85 250 -51
rect 284 -85 300 -51
rect 238 -100 300 -85
rect 330 85 392 100
rect 330 51 346 85
rect 380 51 392 85
rect 330 17 392 51
rect 330 -17 346 17
rect 380 -17 392 17
rect 330 -51 392 -17
rect 330 -85 346 -51
rect 380 -85 392 -51
rect 330 -100 392 -85
rect 448 85 510 100
rect 448 51 460 85
rect 494 51 510 85
rect 448 17 510 51
rect 448 -17 460 17
rect 494 -17 510 17
rect 448 -51 510 -17
rect 448 -85 460 -51
rect 494 -85 510 -51
rect 448 -100 510 -85
rect 540 85 602 100
rect 540 51 556 85
rect 590 51 602 85
rect 540 17 602 51
rect 540 -17 556 17
rect 590 -17 602 17
rect 540 -51 602 -17
rect 540 -85 556 -51
rect 590 -85 602 -51
rect 540 -100 602 -85
rect 658 85 720 100
rect 658 51 670 85
rect 704 51 720 85
rect 658 17 720 51
rect 658 -17 670 17
rect 704 -17 720 17
rect 658 -51 720 -17
rect 658 -85 670 -51
rect 704 -85 720 -51
rect 658 -100 720 -85
rect 750 85 812 100
rect 750 51 766 85
rect 800 51 812 85
rect 750 17 812 51
rect 750 -17 766 17
rect 800 -17 812 17
rect 750 -51 812 -17
rect 750 -85 766 -51
rect 800 -85 812 -51
rect 750 -100 812 -85
rect 868 85 930 100
rect 868 51 880 85
rect 914 51 930 85
rect 868 17 930 51
rect 868 -17 880 17
rect 914 -17 930 17
rect 868 -51 930 -17
rect 868 -85 880 -51
rect 914 -85 930 -51
rect 868 -100 930 -85
rect 960 85 1022 100
rect 960 51 976 85
rect 1010 51 1022 85
rect 960 17 1022 51
rect 960 -17 976 17
rect 1010 -17 1022 17
rect 960 -51 1022 -17
rect 960 -85 976 -51
rect 1010 -85 1022 -51
rect 960 -100 1022 -85
rect 1078 85 1140 100
rect 1078 51 1090 85
rect 1124 51 1140 85
rect 1078 17 1140 51
rect 1078 -17 1090 17
rect 1124 -17 1140 17
rect 1078 -51 1140 -17
rect 1078 -85 1090 -51
rect 1124 -85 1140 -51
rect 1078 -100 1140 -85
rect 1170 85 1232 100
rect 1170 51 1186 85
rect 1220 51 1232 85
rect 1170 17 1232 51
rect 1170 -17 1186 17
rect 1220 -17 1232 17
rect 1170 -51 1232 -17
rect 1170 -85 1186 -51
rect 1220 -85 1232 -51
rect 1170 -100 1232 -85
rect 1288 85 1350 100
rect 1288 51 1300 85
rect 1334 51 1350 85
rect 1288 17 1350 51
rect 1288 -17 1300 17
rect 1334 -17 1350 17
rect 1288 -51 1350 -17
rect 1288 -85 1300 -51
rect 1334 -85 1350 -51
rect 1288 -100 1350 -85
rect 1380 85 1442 100
rect 1380 51 1396 85
rect 1430 51 1442 85
rect 1380 17 1442 51
rect 1380 -17 1396 17
rect 1430 -17 1442 17
rect 1380 -51 1442 -17
rect 1380 -85 1396 -51
rect 1430 -85 1442 -51
rect 1380 -100 1442 -85
rect 1498 85 1560 100
rect 1498 51 1510 85
rect 1544 51 1560 85
rect 1498 17 1560 51
rect 1498 -17 1510 17
rect 1544 -17 1560 17
rect 1498 -51 1560 -17
rect 1498 -85 1510 -51
rect 1544 -85 1560 -51
rect 1498 -100 1560 -85
rect 1590 85 1652 100
rect 1590 51 1606 85
rect 1640 51 1652 85
rect 1590 17 1652 51
rect 1590 -17 1606 17
rect 1640 -17 1652 17
rect 1590 -51 1652 -17
rect 1590 -85 1606 -51
rect 1640 -85 1652 -51
rect 1590 -100 1652 -85
rect 1708 85 1770 100
rect 1708 51 1720 85
rect 1754 51 1770 85
rect 1708 17 1770 51
rect 1708 -17 1720 17
rect 1754 -17 1770 17
rect 1708 -51 1770 -17
rect 1708 -85 1720 -51
rect 1754 -85 1770 -51
rect 1708 -100 1770 -85
rect 1800 85 1862 100
rect 1800 51 1816 85
rect 1850 51 1862 85
rect 1800 17 1862 51
rect 1800 -17 1816 17
rect 1850 -17 1862 17
rect 1800 -51 1862 -17
rect 1800 -85 1816 -51
rect 1850 -85 1862 -51
rect 1800 -100 1862 -85
rect 1918 85 1980 100
rect 1918 51 1930 85
rect 1964 51 1980 85
rect 1918 17 1980 51
rect 1918 -17 1930 17
rect 1964 -17 1980 17
rect 1918 -51 1980 -17
rect 1918 -85 1930 -51
rect 1964 -85 1980 -51
rect 1918 -100 1980 -85
rect 2010 85 2072 100
rect 2010 51 2026 85
rect 2060 51 2072 85
rect 2010 17 2072 51
rect 2010 -17 2026 17
rect 2060 -17 2072 17
rect 2010 -51 2072 -17
rect 2010 -85 2026 -51
rect 2060 -85 2072 -51
rect 2010 -100 2072 -85
rect 2128 85 2190 100
rect 2128 51 2140 85
rect 2174 51 2190 85
rect 2128 17 2190 51
rect 2128 -17 2140 17
rect 2174 -17 2190 17
rect 2128 -51 2190 -17
rect 2128 -85 2140 -51
rect 2174 -85 2190 -51
rect 2128 -100 2190 -85
rect 2220 85 2282 100
rect 2220 51 2236 85
rect 2270 51 2282 85
rect 2220 17 2282 51
rect 2220 -17 2236 17
rect 2270 -17 2282 17
rect 2220 -51 2282 -17
rect 2220 -85 2236 -51
rect 2270 -85 2282 -51
rect 2220 -100 2282 -85
rect 2338 85 2400 100
rect 2338 51 2350 85
rect 2384 51 2400 85
rect 2338 17 2400 51
rect 2338 -17 2350 17
rect 2384 -17 2400 17
rect 2338 -51 2400 -17
rect 2338 -85 2350 -51
rect 2384 -85 2400 -51
rect 2338 -100 2400 -85
rect 2430 85 2492 100
rect 2430 51 2446 85
rect 2480 51 2492 85
rect 2430 17 2492 51
rect 2430 -17 2446 17
rect 2480 -17 2492 17
rect 2430 -51 2492 -17
rect 2430 -85 2446 -51
rect 2480 -85 2492 -51
rect 2430 -100 2492 -85
rect 2548 85 2610 100
rect 2548 51 2560 85
rect 2594 51 2610 85
rect 2548 17 2610 51
rect 2548 -17 2560 17
rect 2594 -17 2610 17
rect 2548 -51 2610 -17
rect 2548 -85 2560 -51
rect 2594 -85 2610 -51
rect 2548 -100 2610 -85
rect 2640 85 2702 100
rect 2640 51 2656 85
rect 2690 51 2702 85
rect 2640 17 2702 51
rect 2640 -17 2656 17
rect 2690 -17 2702 17
rect 2640 -51 2702 -17
rect 2640 -85 2656 -51
rect 2690 -85 2702 -51
rect 2640 -100 2702 -85
rect 2758 85 2820 100
rect 2758 51 2770 85
rect 2804 51 2820 85
rect 2758 17 2820 51
rect 2758 -17 2770 17
rect 2804 -17 2820 17
rect 2758 -51 2820 -17
rect 2758 -85 2770 -51
rect 2804 -85 2820 -51
rect 2758 -100 2820 -85
rect 2850 85 2912 100
rect 2850 51 2866 85
rect 2900 51 2912 85
rect 2850 17 2912 51
rect 2850 -17 2866 17
rect 2900 -17 2912 17
rect 2850 -51 2912 -17
rect 2850 -85 2866 -51
rect 2900 -85 2912 -51
rect 2850 -100 2912 -85
rect 2968 85 3030 100
rect 2968 51 2980 85
rect 3014 51 3030 85
rect 2968 17 3030 51
rect 2968 -17 2980 17
rect 3014 -17 3030 17
rect 2968 -51 3030 -17
rect 2968 -85 2980 -51
rect 3014 -85 3030 -51
rect 2968 -100 3030 -85
rect 3060 85 3122 100
rect 3060 51 3076 85
rect 3110 51 3122 85
rect 3060 17 3122 51
rect 3060 -17 3076 17
rect 3110 -17 3122 17
rect 3060 -51 3122 -17
rect 3060 -85 3076 -51
rect 3110 -85 3122 -51
rect 3060 -100 3122 -85
rect 3178 85 3240 100
rect 3178 51 3190 85
rect 3224 51 3240 85
rect 3178 17 3240 51
rect 3178 -17 3190 17
rect 3224 -17 3240 17
rect 3178 -51 3240 -17
rect 3178 -85 3190 -51
rect 3224 -85 3240 -51
rect 3178 -100 3240 -85
rect 3270 85 3332 100
rect 3270 51 3286 85
rect 3320 51 3332 85
rect 3270 17 3332 51
rect 3270 -17 3286 17
rect 3320 -17 3332 17
rect 3270 -51 3332 -17
rect 3270 -85 3286 -51
rect 3320 -85 3332 -51
rect 3270 -100 3332 -85
rect 3388 85 3450 100
rect 3388 51 3400 85
rect 3434 51 3450 85
rect 3388 17 3450 51
rect 3388 -17 3400 17
rect 3434 -17 3450 17
rect 3388 -51 3450 -17
rect 3388 -85 3400 -51
rect 3434 -85 3450 -51
rect 3388 -100 3450 -85
rect 3480 85 3542 100
rect 3480 51 3496 85
rect 3530 51 3542 85
rect 3480 17 3542 51
rect 3480 -17 3496 17
rect 3530 -17 3542 17
rect 3480 -51 3542 -17
rect 3480 -85 3496 -51
rect 3530 -85 3542 -51
rect 3480 -100 3542 -85
rect 3598 85 3660 100
rect 3598 51 3610 85
rect 3644 51 3660 85
rect 3598 17 3660 51
rect 3598 -17 3610 17
rect 3644 -17 3660 17
rect 3598 -51 3660 -17
rect 3598 -85 3610 -51
rect 3644 -85 3660 -51
rect 3598 -100 3660 -85
rect 3690 85 3752 100
rect 3690 51 3706 85
rect 3740 51 3752 85
rect 3690 17 3752 51
rect 3690 -17 3706 17
rect 3740 -17 3752 17
rect 3690 -51 3752 -17
rect 3690 -85 3706 -51
rect 3740 -85 3752 -51
rect 3690 -100 3752 -85
rect 3808 85 3870 100
rect 3808 51 3820 85
rect 3854 51 3870 85
rect 3808 17 3870 51
rect 3808 -17 3820 17
rect 3854 -17 3870 17
rect 3808 -51 3870 -17
rect 3808 -85 3820 -51
rect 3854 -85 3870 -51
rect 3808 -100 3870 -85
rect 3900 85 3962 100
rect 3900 51 3916 85
rect 3950 51 3962 85
rect 3900 17 3962 51
rect 3900 -17 3916 17
rect 3950 -17 3962 17
rect 3900 -51 3962 -17
rect 3900 -85 3916 -51
rect 3950 -85 3962 -51
rect 3900 -100 3962 -85
rect 4018 85 4080 100
rect 4018 51 4030 85
rect 4064 51 4080 85
rect 4018 17 4080 51
rect 4018 -17 4030 17
rect 4064 -17 4080 17
rect 4018 -51 4080 -17
rect 4018 -85 4030 -51
rect 4064 -85 4080 -51
rect 4018 -100 4080 -85
rect 4110 85 4172 100
rect 4110 51 4126 85
rect 4160 51 4172 85
rect 4110 17 4172 51
rect 4110 -17 4126 17
rect 4160 -17 4172 17
rect 4110 -51 4172 -17
rect 4110 -85 4126 -51
rect 4160 -85 4172 -51
rect 4110 -100 4172 -85
rect 4228 85 4290 100
rect 4228 51 4240 85
rect 4274 51 4290 85
rect 4228 17 4290 51
rect 4228 -17 4240 17
rect 4274 -17 4290 17
rect 4228 -51 4290 -17
rect 4228 -85 4240 -51
rect 4274 -85 4290 -51
rect 4228 -100 4290 -85
rect 4320 85 4382 100
rect 4320 51 4336 85
rect 4370 51 4382 85
rect 4320 17 4382 51
rect 4320 -17 4336 17
rect 4370 -17 4382 17
rect 4320 -51 4382 -17
rect 4320 -85 4336 -51
rect 4370 -85 4382 -51
rect 4320 -100 4382 -85
<< ndiffc >>
rect -4370 51 -4336 85
rect -4370 -17 -4336 17
rect -4370 -85 -4336 -51
rect -4274 51 -4240 85
rect -4274 -17 -4240 17
rect -4274 -85 -4240 -51
rect -4160 51 -4126 85
rect -4160 -17 -4126 17
rect -4160 -85 -4126 -51
rect -4064 51 -4030 85
rect -4064 -17 -4030 17
rect -4064 -85 -4030 -51
rect -3950 51 -3916 85
rect -3950 -17 -3916 17
rect -3950 -85 -3916 -51
rect -3854 51 -3820 85
rect -3854 -17 -3820 17
rect -3854 -85 -3820 -51
rect -3740 51 -3706 85
rect -3740 -17 -3706 17
rect -3740 -85 -3706 -51
rect -3644 51 -3610 85
rect -3644 -17 -3610 17
rect -3644 -85 -3610 -51
rect -3530 51 -3496 85
rect -3530 -17 -3496 17
rect -3530 -85 -3496 -51
rect -3434 51 -3400 85
rect -3434 -17 -3400 17
rect -3434 -85 -3400 -51
rect -3320 51 -3286 85
rect -3320 -17 -3286 17
rect -3320 -85 -3286 -51
rect -3224 51 -3190 85
rect -3224 -17 -3190 17
rect -3224 -85 -3190 -51
rect -3110 51 -3076 85
rect -3110 -17 -3076 17
rect -3110 -85 -3076 -51
rect -3014 51 -2980 85
rect -3014 -17 -2980 17
rect -3014 -85 -2980 -51
rect -2900 51 -2866 85
rect -2900 -17 -2866 17
rect -2900 -85 -2866 -51
rect -2804 51 -2770 85
rect -2804 -17 -2770 17
rect -2804 -85 -2770 -51
rect -2690 51 -2656 85
rect -2690 -17 -2656 17
rect -2690 -85 -2656 -51
rect -2594 51 -2560 85
rect -2594 -17 -2560 17
rect -2594 -85 -2560 -51
rect -2480 51 -2446 85
rect -2480 -17 -2446 17
rect -2480 -85 -2446 -51
rect -2384 51 -2350 85
rect -2384 -17 -2350 17
rect -2384 -85 -2350 -51
rect -2270 51 -2236 85
rect -2270 -17 -2236 17
rect -2270 -85 -2236 -51
rect -2174 51 -2140 85
rect -2174 -17 -2140 17
rect -2174 -85 -2140 -51
rect -2060 51 -2026 85
rect -2060 -17 -2026 17
rect -2060 -85 -2026 -51
rect -1964 51 -1930 85
rect -1964 -17 -1930 17
rect -1964 -85 -1930 -51
rect -1850 51 -1816 85
rect -1850 -17 -1816 17
rect -1850 -85 -1816 -51
rect -1754 51 -1720 85
rect -1754 -17 -1720 17
rect -1754 -85 -1720 -51
rect -1640 51 -1606 85
rect -1640 -17 -1606 17
rect -1640 -85 -1606 -51
rect -1544 51 -1510 85
rect -1544 -17 -1510 17
rect -1544 -85 -1510 -51
rect -1430 51 -1396 85
rect -1430 -17 -1396 17
rect -1430 -85 -1396 -51
rect -1334 51 -1300 85
rect -1334 -17 -1300 17
rect -1334 -85 -1300 -51
rect -1220 51 -1186 85
rect -1220 -17 -1186 17
rect -1220 -85 -1186 -51
rect -1124 51 -1090 85
rect -1124 -17 -1090 17
rect -1124 -85 -1090 -51
rect -1010 51 -976 85
rect -1010 -17 -976 17
rect -1010 -85 -976 -51
rect -914 51 -880 85
rect -914 -17 -880 17
rect -914 -85 -880 -51
rect -800 51 -766 85
rect -800 -17 -766 17
rect -800 -85 -766 -51
rect -704 51 -670 85
rect -704 -17 -670 17
rect -704 -85 -670 -51
rect -590 51 -556 85
rect -590 -17 -556 17
rect -590 -85 -556 -51
rect -494 51 -460 85
rect -494 -17 -460 17
rect -494 -85 -460 -51
rect -380 51 -346 85
rect -380 -17 -346 17
rect -380 -85 -346 -51
rect -284 51 -250 85
rect -284 -17 -250 17
rect -284 -85 -250 -51
rect -170 51 -136 85
rect -170 -17 -136 17
rect -170 -85 -136 -51
rect -74 51 -40 85
rect -74 -17 -40 17
rect -74 -85 -40 -51
rect 40 51 74 85
rect 40 -17 74 17
rect 40 -85 74 -51
rect 136 51 170 85
rect 136 -17 170 17
rect 136 -85 170 -51
rect 250 51 284 85
rect 250 -17 284 17
rect 250 -85 284 -51
rect 346 51 380 85
rect 346 -17 380 17
rect 346 -85 380 -51
rect 460 51 494 85
rect 460 -17 494 17
rect 460 -85 494 -51
rect 556 51 590 85
rect 556 -17 590 17
rect 556 -85 590 -51
rect 670 51 704 85
rect 670 -17 704 17
rect 670 -85 704 -51
rect 766 51 800 85
rect 766 -17 800 17
rect 766 -85 800 -51
rect 880 51 914 85
rect 880 -17 914 17
rect 880 -85 914 -51
rect 976 51 1010 85
rect 976 -17 1010 17
rect 976 -85 1010 -51
rect 1090 51 1124 85
rect 1090 -17 1124 17
rect 1090 -85 1124 -51
rect 1186 51 1220 85
rect 1186 -17 1220 17
rect 1186 -85 1220 -51
rect 1300 51 1334 85
rect 1300 -17 1334 17
rect 1300 -85 1334 -51
rect 1396 51 1430 85
rect 1396 -17 1430 17
rect 1396 -85 1430 -51
rect 1510 51 1544 85
rect 1510 -17 1544 17
rect 1510 -85 1544 -51
rect 1606 51 1640 85
rect 1606 -17 1640 17
rect 1606 -85 1640 -51
rect 1720 51 1754 85
rect 1720 -17 1754 17
rect 1720 -85 1754 -51
rect 1816 51 1850 85
rect 1816 -17 1850 17
rect 1816 -85 1850 -51
rect 1930 51 1964 85
rect 1930 -17 1964 17
rect 1930 -85 1964 -51
rect 2026 51 2060 85
rect 2026 -17 2060 17
rect 2026 -85 2060 -51
rect 2140 51 2174 85
rect 2140 -17 2174 17
rect 2140 -85 2174 -51
rect 2236 51 2270 85
rect 2236 -17 2270 17
rect 2236 -85 2270 -51
rect 2350 51 2384 85
rect 2350 -17 2384 17
rect 2350 -85 2384 -51
rect 2446 51 2480 85
rect 2446 -17 2480 17
rect 2446 -85 2480 -51
rect 2560 51 2594 85
rect 2560 -17 2594 17
rect 2560 -85 2594 -51
rect 2656 51 2690 85
rect 2656 -17 2690 17
rect 2656 -85 2690 -51
rect 2770 51 2804 85
rect 2770 -17 2804 17
rect 2770 -85 2804 -51
rect 2866 51 2900 85
rect 2866 -17 2900 17
rect 2866 -85 2900 -51
rect 2980 51 3014 85
rect 2980 -17 3014 17
rect 2980 -85 3014 -51
rect 3076 51 3110 85
rect 3076 -17 3110 17
rect 3076 -85 3110 -51
rect 3190 51 3224 85
rect 3190 -17 3224 17
rect 3190 -85 3224 -51
rect 3286 51 3320 85
rect 3286 -17 3320 17
rect 3286 -85 3320 -51
rect 3400 51 3434 85
rect 3400 -17 3434 17
rect 3400 -85 3434 -51
rect 3496 51 3530 85
rect 3496 -17 3530 17
rect 3496 -85 3530 -51
rect 3610 51 3644 85
rect 3610 -17 3644 17
rect 3610 -85 3644 -51
rect 3706 51 3740 85
rect 3706 -17 3740 17
rect 3706 -85 3740 -51
rect 3820 51 3854 85
rect 3820 -17 3854 17
rect 3820 -85 3854 -51
rect 3916 51 3950 85
rect 3916 -17 3950 17
rect 3916 -85 3950 -51
rect 4030 51 4064 85
rect 4030 -17 4064 17
rect 4030 -85 4064 -51
rect 4126 51 4160 85
rect 4126 -17 4160 17
rect 4126 -85 4160 -51
rect 4240 51 4274 85
rect 4240 -17 4274 17
rect 4240 -85 4274 -51
rect 4336 51 4370 85
rect 4336 -17 4370 17
rect 4336 -85 4370 -51
<< poly >>
rect -4128 172 -4062 188
rect -4128 138 -4112 172
rect -4078 138 -4062 172
rect -4320 100 -4290 126
rect -4128 122 -4062 138
rect -3708 172 -3642 188
rect -3708 138 -3692 172
rect -3658 138 -3642 172
rect -4110 100 -4080 122
rect -3900 100 -3870 126
rect -3708 122 -3642 138
rect -3288 172 -3222 188
rect -3288 138 -3272 172
rect -3238 138 -3222 172
rect -3690 100 -3660 122
rect -3480 100 -3450 126
rect -3288 122 -3222 138
rect -2868 172 -2802 188
rect -2868 138 -2852 172
rect -2818 138 -2802 172
rect -3270 100 -3240 122
rect -3060 100 -3030 126
rect -2868 122 -2802 138
rect -2448 172 -2382 188
rect -2448 138 -2432 172
rect -2398 138 -2382 172
rect -2850 100 -2820 122
rect -2640 100 -2610 126
rect -2448 122 -2382 138
rect -2028 172 -1962 188
rect -2028 138 -2012 172
rect -1978 138 -1962 172
rect -2430 100 -2400 122
rect -2220 100 -2190 126
rect -2028 122 -1962 138
rect -1608 172 -1542 188
rect -1608 138 -1592 172
rect -1558 138 -1542 172
rect -2010 100 -1980 122
rect -1800 100 -1770 126
rect -1608 122 -1542 138
rect -1188 172 -1122 188
rect -1188 138 -1172 172
rect -1138 138 -1122 172
rect -1590 100 -1560 122
rect -1380 100 -1350 126
rect -1188 122 -1122 138
rect -768 172 -702 188
rect -768 138 -752 172
rect -718 138 -702 172
rect -1170 100 -1140 122
rect -960 100 -930 126
rect -768 122 -702 138
rect -348 172 -282 188
rect -348 138 -332 172
rect -298 138 -282 172
rect -750 100 -720 122
rect -540 100 -510 126
rect -348 122 -282 138
rect 72 172 138 188
rect 72 138 88 172
rect 122 138 138 172
rect -330 100 -300 122
rect -120 100 -90 126
rect 72 122 138 138
rect 492 172 558 188
rect 492 138 508 172
rect 542 138 558 172
rect 90 100 120 122
rect 300 100 330 126
rect 492 122 558 138
rect 912 172 978 188
rect 912 138 928 172
rect 962 138 978 172
rect 510 100 540 122
rect 720 100 750 126
rect 912 122 978 138
rect 1332 172 1398 188
rect 1332 138 1348 172
rect 1382 138 1398 172
rect 930 100 960 122
rect 1140 100 1170 126
rect 1332 122 1398 138
rect 1752 172 1818 188
rect 1752 138 1768 172
rect 1802 138 1818 172
rect 1350 100 1380 122
rect 1560 100 1590 126
rect 1752 122 1818 138
rect 2172 172 2238 188
rect 2172 138 2188 172
rect 2222 138 2238 172
rect 1770 100 1800 122
rect 1980 100 2010 126
rect 2172 122 2238 138
rect 2592 172 2658 188
rect 2592 138 2608 172
rect 2642 138 2658 172
rect 2190 100 2220 122
rect 2400 100 2430 126
rect 2592 122 2658 138
rect 3012 172 3078 188
rect 3012 138 3028 172
rect 3062 138 3078 172
rect 2610 100 2640 122
rect 2820 100 2850 126
rect 3012 122 3078 138
rect 3432 172 3498 188
rect 3432 138 3448 172
rect 3482 138 3498 172
rect 3030 100 3060 122
rect 3240 100 3270 126
rect 3432 122 3498 138
rect 3852 172 3918 188
rect 3852 138 3868 172
rect 3902 138 3918 172
rect 3450 100 3480 122
rect 3660 100 3690 126
rect 3852 122 3918 138
rect 4272 172 4338 188
rect 4272 138 4288 172
rect 4322 138 4338 172
rect 3870 100 3900 122
rect 4080 100 4110 126
rect 4272 122 4338 138
rect 4290 100 4320 122
rect -4320 -122 -4290 -100
rect -4338 -138 -4272 -122
rect -4110 -126 -4080 -100
rect -3900 -122 -3870 -100
rect -4338 -172 -4322 -138
rect -4288 -172 -4272 -138
rect -4338 -188 -4272 -172
rect -3918 -138 -3852 -122
rect -3690 -126 -3660 -100
rect -3480 -122 -3450 -100
rect -3918 -172 -3902 -138
rect -3868 -172 -3852 -138
rect -3918 -188 -3852 -172
rect -3498 -138 -3432 -122
rect -3270 -126 -3240 -100
rect -3060 -122 -3030 -100
rect -3498 -172 -3482 -138
rect -3448 -172 -3432 -138
rect -3498 -188 -3432 -172
rect -3078 -138 -3012 -122
rect -2850 -126 -2820 -100
rect -2640 -122 -2610 -100
rect -3078 -172 -3062 -138
rect -3028 -172 -3012 -138
rect -3078 -188 -3012 -172
rect -2658 -138 -2592 -122
rect -2430 -126 -2400 -100
rect -2220 -122 -2190 -100
rect -2658 -172 -2642 -138
rect -2608 -172 -2592 -138
rect -2658 -188 -2592 -172
rect -2238 -138 -2172 -122
rect -2010 -126 -1980 -100
rect -1800 -122 -1770 -100
rect -2238 -172 -2222 -138
rect -2188 -172 -2172 -138
rect -2238 -188 -2172 -172
rect -1818 -138 -1752 -122
rect -1590 -126 -1560 -100
rect -1380 -122 -1350 -100
rect -1818 -172 -1802 -138
rect -1768 -172 -1752 -138
rect -1818 -188 -1752 -172
rect -1398 -138 -1332 -122
rect -1170 -126 -1140 -100
rect -960 -122 -930 -100
rect -1398 -172 -1382 -138
rect -1348 -172 -1332 -138
rect -1398 -188 -1332 -172
rect -978 -138 -912 -122
rect -750 -126 -720 -100
rect -540 -122 -510 -100
rect -978 -172 -962 -138
rect -928 -172 -912 -138
rect -978 -188 -912 -172
rect -558 -138 -492 -122
rect -330 -126 -300 -100
rect -120 -122 -90 -100
rect -558 -172 -542 -138
rect -508 -172 -492 -138
rect -558 -188 -492 -172
rect -138 -138 -72 -122
rect 90 -126 120 -100
rect 300 -122 330 -100
rect -138 -172 -122 -138
rect -88 -172 -72 -138
rect -138 -188 -72 -172
rect 282 -138 348 -122
rect 510 -126 540 -100
rect 720 -122 750 -100
rect 282 -172 298 -138
rect 332 -172 348 -138
rect 282 -188 348 -172
rect 702 -138 768 -122
rect 930 -126 960 -100
rect 1140 -122 1170 -100
rect 702 -172 718 -138
rect 752 -172 768 -138
rect 702 -188 768 -172
rect 1122 -138 1188 -122
rect 1350 -126 1380 -100
rect 1560 -122 1590 -100
rect 1122 -172 1138 -138
rect 1172 -172 1188 -138
rect 1122 -188 1188 -172
rect 1542 -138 1608 -122
rect 1770 -126 1800 -100
rect 1980 -122 2010 -100
rect 1542 -172 1558 -138
rect 1592 -172 1608 -138
rect 1542 -188 1608 -172
rect 1962 -138 2028 -122
rect 2190 -126 2220 -100
rect 2400 -122 2430 -100
rect 1962 -172 1978 -138
rect 2012 -172 2028 -138
rect 1962 -188 2028 -172
rect 2382 -138 2448 -122
rect 2610 -126 2640 -100
rect 2820 -122 2850 -100
rect 2382 -172 2398 -138
rect 2432 -172 2448 -138
rect 2382 -188 2448 -172
rect 2802 -138 2868 -122
rect 3030 -126 3060 -100
rect 3240 -122 3270 -100
rect 2802 -172 2818 -138
rect 2852 -172 2868 -138
rect 2802 -188 2868 -172
rect 3222 -138 3288 -122
rect 3450 -126 3480 -100
rect 3660 -122 3690 -100
rect 3222 -172 3238 -138
rect 3272 -172 3288 -138
rect 3222 -188 3288 -172
rect 3642 -138 3708 -122
rect 3870 -126 3900 -100
rect 4080 -122 4110 -100
rect 3642 -172 3658 -138
rect 3692 -172 3708 -138
rect 3642 -188 3708 -172
rect 4062 -138 4128 -122
rect 4290 -126 4320 -100
rect 4062 -172 4078 -138
rect 4112 -172 4128 -138
rect 4062 -188 4128 -172
<< polycont >>
rect -4112 138 -4078 172
rect -3692 138 -3658 172
rect -3272 138 -3238 172
rect -2852 138 -2818 172
rect -2432 138 -2398 172
rect -2012 138 -1978 172
rect -1592 138 -1558 172
rect -1172 138 -1138 172
rect -752 138 -718 172
rect -332 138 -298 172
rect 88 138 122 172
rect 508 138 542 172
rect 928 138 962 172
rect 1348 138 1382 172
rect 1768 138 1802 172
rect 2188 138 2222 172
rect 2608 138 2642 172
rect 3028 138 3062 172
rect 3448 138 3482 172
rect 3868 138 3902 172
rect 4288 138 4322 172
rect -4322 -172 -4288 -138
rect -3902 -172 -3868 -138
rect -3482 -172 -3448 -138
rect -3062 -172 -3028 -138
rect -2642 -172 -2608 -138
rect -2222 -172 -2188 -138
rect -1802 -172 -1768 -138
rect -1382 -172 -1348 -138
rect -962 -172 -928 -138
rect -542 -172 -508 -138
rect -122 -172 -88 -138
rect 298 -172 332 -138
rect 718 -172 752 -138
rect 1138 -172 1172 -138
rect 1558 -172 1592 -138
rect 1978 -172 2012 -138
rect 2398 -172 2432 -138
rect 2818 -172 2852 -138
rect 3238 -172 3272 -138
rect 3658 -172 3692 -138
rect 4078 -172 4112 -138
<< locali >>
rect -4128 138 -4112 172
rect -4078 138 -4062 172
rect -3708 138 -3692 172
rect -3658 138 -3642 172
rect -3288 138 -3272 172
rect -3238 138 -3222 172
rect -2868 138 -2852 172
rect -2818 138 -2802 172
rect -2448 138 -2432 172
rect -2398 138 -2382 172
rect -2028 138 -2012 172
rect -1978 138 -1962 172
rect -1608 138 -1592 172
rect -1558 138 -1542 172
rect -1188 138 -1172 172
rect -1138 138 -1122 172
rect -768 138 -752 172
rect -718 138 -702 172
rect -348 138 -332 172
rect -298 138 -282 172
rect 72 138 88 172
rect 122 138 138 172
rect 492 138 508 172
rect 542 138 558 172
rect 912 138 928 172
rect 962 138 978 172
rect 1332 138 1348 172
rect 1382 138 1398 172
rect 1752 138 1768 172
rect 1802 138 1818 172
rect 2172 138 2188 172
rect 2222 138 2238 172
rect 2592 138 2608 172
rect 2642 138 2658 172
rect 3012 138 3028 172
rect 3062 138 3078 172
rect 3432 138 3448 172
rect 3482 138 3498 172
rect 3852 138 3868 172
rect 3902 138 3918 172
rect 4240 138 4288 172
rect 4322 138 4370 172
rect -4370 85 -4336 104
rect -4370 17 -4336 51
rect -4370 -51 -4336 -17
rect -4370 -138 -4336 -85
rect -4274 85 -4240 104
rect -4274 17 -4240 51
rect -4274 -51 -4240 -17
rect -4274 -138 -4240 -85
rect -4160 88 -4126 104
rect -4160 17 -4126 51
rect -4160 -51 -4126 -17
rect -4160 -104 -4126 -85
rect -4064 85 -4030 104
rect -4064 17 -4030 51
rect -4064 -51 -4030 -17
rect -4064 -104 -4030 -88
rect -3950 88 -3916 104
rect -3950 17 -3916 51
rect -3950 -51 -3916 -17
rect -3950 -104 -3916 -85
rect -3854 85 -3820 104
rect -3854 17 -3820 51
rect -3854 -51 -3820 -17
rect -3854 -104 -3820 -88
rect -3740 88 -3706 104
rect -3740 17 -3706 51
rect -3740 -51 -3706 -17
rect -3740 -104 -3706 -85
rect -3644 85 -3610 104
rect -3644 17 -3610 51
rect -3644 -51 -3610 -17
rect -3644 -104 -3610 -88
rect -3530 88 -3496 104
rect -3530 17 -3496 51
rect -3530 -51 -3496 -17
rect -3530 -104 -3496 -85
rect -3434 85 -3400 104
rect -3434 17 -3400 51
rect -3434 -51 -3400 -17
rect -3434 -104 -3400 -88
rect -3320 88 -3286 104
rect -3320 17 -3286 51
rect -3320 -51 -3286 -17
rect -3320 -104 -3286 -85
rect -3224 85 -3190 104
rect -3224 17 -3190 51
rect -3224 -51 -3190 -17
rect -3224 -104 -3190 -88
rect -3110 88 -3076 104
rect -3110 17 -3076 51
rect -3110 -51 -3076 -17
rect -3110 -104 -3076 -85
rect -3014 85 -2980 104
rect -3014 17 -2980 51
rect -3014 -51 -2980 -17
rect -3014 -104 -2980 -88
rect -2900 88 -2866 104
rect -2900 17 -2866 51
rect -2900 -51 -2866 -17
rect -2900 -104 -2866 -85
rect -2804 85 -2770 104
rect -2804 17 -2770 51
rect -2804 -51 -2770 -17
rect -2804 -104 -2770 -88
rect -2690 88 -2656 104
rect -2690 17 -2656 51
rect -2690 -51 -2656 -17
rect -2690 -104 -2656 -85
rect -2594 85 -2560 104
rect -2594 17 -2560 51
rect -2594 -51 -2560 -17
rect -2594 -104 -2560 -88
rect -2480 88 -2446 104
rect -2480 17 -2446 51
rect -2480 -51 -2446 -17
rect -2480 -104 -2446 -85
rect -2384 85 -2350 104
rect -2384 17 -2350 51
rect -2384 -51 -2350 -17
rect -2384 -104 -2350 -88
rect -2270 88 -2236 104
rect -2270 17 -2236 51
rect -2270 -51 -2236 -17
rect -2270 -104 -2236 -85
rect -2174 85 -2140 104
rect -2174 17 -2140 51
rect -2174 -51 -2140 -17
rect -2174 -104 -2140 -88
rect -2060 88 -2026 104
rect -2060 17 -2026 51
rect -2060 -51 -2026 -17
rect -2060 -104 -2026 -85
rect -1964 85 -1930 104
rect -1964 17 -1930 51
rect -1964 -51 -1930 -17
rect -1964 -104 -1930 -88
rect -1850 88 -1816 104
rect -1850 17 -1816 51
rect -1850 -51 -1816 -17
rect -1850 -104 -1816 -85
rect -1754 85 -1720 104
rect -1754 17 -1720 51
rect -1754 -51 -1720 -17
rect -1754 -104 -1720 -88
rect -1640 88 -1606 104
rect -1640 17 -1606 51
rect -1640 -51 -1606 -17
rect -1640 -104 -1606 -85
rect -1544 85 -1510 104
rect -1544 17 -1510 51
rect -1544 -51 -1510 -17
rect -1544 -104 -1510 -88
rect -1430 88 -1396 104
rect -1430 17 -1396 51
rect -1430 -51 -1396 -17
rect -1430 -104 -1396 -85
rect -1334 85 -1300 104
rect -1334 17 -1300 51
rect -1334 -51 -1300 -17
rect -1334 -104 -1300 -88
rect -1220 88 -1186 104
rect -1220 17 -1186 51
rect -1220 -51 -1186 -17
rect -1220 -104 -1186 -85
rect -1124 85 -1090 104
rect -1124 17 -1090 51
rect -1124 -51 -1090 -17
rect -1124 -104 -1090 -88
rect -1010 88 -976 104
rect -1010 17 -976 51
rect -1010 -51 -976 -17
rect -1010 -104 -976 -85
rect -914 85 -880 104
rect -914 17 -880 51
rect -914 -51 -880 -17
rect -914 -104 -880 -88
rect -800 88 -766 104
rect -800 17 -766 51
rect -800 -51 -766 -17
rect -800 -104 -766 -85
rect -704 85 -670 104
rect -704 17 -670 51
rect -704 -51 -670 -17
rect -704 -104 -670 -88
rect -590 88 -556 104
rect -590 17 -556 51
rect -590 -51 -556 -17
rect -590 -104 -556 -85
rect -494 85 -460 104
rect -494 17 -460 51
rect -494 -51 -460 -17
rect -494 -104 -460 -88
rect -380 88 -346 104
rect -380 17 -346 51
rect -380 -51 -346 -17
rect -380 -104 -346 -85
rect -284 85 -250 104
rect -284 17 -250 51
rect -284 -51 -250 -17
rect -284 -104 -250 -88
rect -170 88 -136 104
rect -170 17 -136 51
rect -170 -51 -136 -17
rect -170 -104 -136 -85
rect -74 85 -40 104
rect -74 17 -40 51
rect -74 -51 -40 -17
rect -74 -104 -40 -88
rect 40 88 74 104
rect 40 17 74 51
rect 40 -51 74 -17
rect 40 -104 74 -85
rect 136 85 170 104
rect 136 17 170 51
rect 136 -51 170 -17
rect 136 -104 170 -88
rect 250 88 284 104
rect 250 17 284 51
rect 250 -51 284 -17
rect 250 -104 284 -85
rect 346 85 380 104
rect 346 17 380 51
rect 346 -51 380 -17
rect 346 -104 380 -88
rect 460 88 494 104
rect 460 17 494 51
rect 460 -51 494 -17
rect 460 -104 494 -85
rect 556 85 590 104
rect 556 17 590 51
rect 556 -51 590 -17
rect 556 -104 590 -88
rect 670 88 704 104
rect 670 17 704 51
rect 670 -51 704 -17
rect 670 -104 704 -85
rect 766 85 800 104
rect 766 17 800 51
rect 766 -51 800 -17
rect 766 -104 800 -88
rect 880 88 914 104
rect 880 17 914 51
rect 880 -51 914 -17
rect 880 -104 914 -85
rect 976 85 1010 104
rect 976 17 1010 51
rect 976 -51 1010 -17
rect 976 -104 1010 -88
rect 1090 88 1124 104
rect 1090 17 1124 51
rect 1090 -51 1124 -17
rect 1090 -104 1124 -85
rect 1186 85 1220 104
rect 1186 17 1220 51
rect 1186 -51 1220 -17
rect 1186 -104 1220 -88
rect 1300 88 1334 104
rect 1300 17 1334 51
rect 1300 -51 1334 -17
rect 1300 -104 1334 -85
rect 1396 85 1430 104
rect 1396 17 1430 51
rect 1396 -51 1430 -17
rect 1396 -104 1430 -88
rect 1510 88 1544 104
rect 1510 17 1544 51
rect 1510 -51 1544 -17
rect 1510 -104 1544 -85
rect 1606 85 1640 104
rect 1606 17 1640 51
rect 1606 -51 1640 -17
rect 1606 -104 1640 -88
rect 1720 88 1754 104
rect 1720 17 1754 51
rect 1720 -51 1754 -17
rect 1720 -104 1754 -85
rect 1816 85 1850 104
rect 1816 17 1850 51
rect 1816 -51 1850 -17
rect 1816 -104 1850 -88
rect 1930 88 1964 104
rect 1930 17 1964 51
rect 1930 -51 1964 -17
rect 1930 -104 1964 -85
rect 2026 85 2060 104
rect 2026 17 2060 51
rect 2026 -51 2060 -17
rect 2026 -104 2060 -88
rect 2140 88 2174 104
rect 2140 17 2174 51
rect 2140 -51 2174 -17
rect 2140 -104 2174 -85
rect 2236 85 2270 104
rect 2236 17 2270 51
rect 2236 -51 2270 -17
rect 2236 -104 2270 -88
rect 2350 88 2384 104
rect 2350 17 2384 51
rect 2350 -51 2384 -17
rect 2350 -104 2384 -85
rect 2446 85 2480 104
rect 2446 17 2480 51
rect 2446 -51 2480 -17
rect 2446 -104 2480 -88
rect 2560 88 2594 104
rect 2560 17 2594 51
rect 2560 -51 2594 -17
rect 2560 -104 2594 -85
rect 2656 85 2690 104
rect 2656 17 2690 51
rect 2656 -51 2690 -17
rect 2656 -104 2690 -88
rect 2770 88 2804 104
rect 2770 17 2804 51
rect 2770 -51 2804 -17
rect 2770 -104 2804 -85
rect 2866 85 2900 104
rect 2866 17 2900 51
rect 2866 -51 2900 -17
rect 2866 -104 2900 -88
rect 2980 88 3014 104
rect 2980 17 3014 51
rect 2980 -51 3014 -17
rect 2980 -104 3014 -85
rect 3076 85 3110 104
rect 3076 17 3110 51
rect 3076 -51 3110 -17
rect 3076 -104 3110 -88
rect 3190 88 3224 104
rect 3190 17 3224 51
rect 3190 -51 3224 -17
rect 3190 -104 3224 -85
rect 3286 85 3320 104
rect 3286 17 3320 51
rect 3286 -51 3320 -17
rect 3286 -104 3320 -88
rect 3400 88 3434 104
rect 3400 17 3434 51
rect 3400 -51 3434 -17
rect 3400 -104 3434 -85
rect 3496 85 3530 104
rect 3496 17 3530 51
rect 3496 -51 3530 -17
rect 3496 -104 3530 -88
rect 3610 88 3644 104
rect 3610 17 3644 51
rect 3610 -51 3644 -17
rect 3610 -104 3644 -85
rect 3706 85 3740 104
rect 3706 17 3740 51
rect 3706 -51 3740 -17
rect 3706 -104 3740 -88
rect 3820 88 3854 104
rect 3820 17 3854 51
rect 3820 -51 3854 -17
rect 3820 -104 3854 -85
rect 3916 85 3950 104
rect 3916 17 3950 51
rect 3916 -51 3950 -17
rect 3916 -104 3950 -88
rect 4030 88 4064 104
rect 4030 17 4064 51
rect 4030 -51 4064 -17
rect 4030 -104 4064 -85
rect 4126 85 4160 104
rect 4126 17 4160 51
rect 4126 -51 4160 -17
rect 4126 -104 4160 -88
rect 4240 85 4274 138
rect 4240 17 4274 51
rect 4240 -51 4274 -17
rect 4240 -104 4274 -85
rect 4336 85 4370 138
rect 4336 17 4370 51
rect 4336 -51 4370 -17
rect 4336 -104 4370 -85
rect -4370 -172 -4322 -138
rect -4288 -172 -4240 -138
rect -3918 -172 -3902 -138
rect -3868 -172 -3852 -138
rect -3498 -172 -3482 -138
rect -3448 -172 -3432 -138
rect -3078 -172 -3062 -138
rect -3028 -172 -3012 -138
rect -2658 -172 -2642 -138
rect -2608 -172 -2592 -138
rect -2238 -172 -2222 -138
rect -2188 -172 -2172 -138
rect -1818 -172 -1802 -138
rect -1768 -172 -1752 -138
rect -1398 -172 -1382 -138
rect -1348 -172 -1332 -138
rect -978 -172 -962 -138
rect -928 -172 -912 -138
rect -558 -172 -542 -138
rect -508 -172 -492 -138
rect -138 -172 -122 -138
rect -88 -172 -72 -138
rect 282 -172 298 -138
rect 332 -172 348 -138
rect 702 -172 718 -138
rect 752 -172 768 -138
rect 1122 -172 1138 -138
rect 1172 -172 1188 -138
rect 1542 -172 1558 -138
rect 1592 -172 1608 -138
rect 1962 -172 1978 -138
rect 2012 -172 2028 -138
rect 2382 -172 2398 -138
rect 2432 -172 2448 -138
rect 2802 -172 2818 -138
rect 2852 -172 2868 -138
rect 3222 -172 3238 -138
rect 3272 -172 3288 -138
rect 3642 -172 3658 -138
rect 3692 -172 3708 -138
rect 4062 -172 4078 -138
rect 4112 -172 4128 -138
<< viali >>
rect -4112 138 -4078 172
rect -3692 138 -3658 172
rect -3272 138 -3238 172
rect -2852 138 -2818 172
rect -2432 138 -2398 172
rect -2012 138 -1978 172
rect -1592 138 -1558 172
rect -1172 138 -1138 172
rect -752 138 -718 172
rect -332 138 -298 172
rect 88 138 122 172
rect 508 138 542 172
rect 928 138 962 172
rect 1348 138 1382 172
rect 1768 138 1802 172
rect 2188 138 2222 172
rect 2608 138 2642 172
rect 3028 138 3062 172
rect 3448 138 3482 172
rect 3868 138 3902 172
rect -4160 85 -4126 88
rect -4160 54 -4126 85
rect -4064 -85 -4030 -54
rect -4064 -88 -4030 -85
rect -3950 85 -3916 88
rect -3950 54 -3916 85
rect -3854 -85 -3820 -54
rect -3854 -88 -3820 -85
rect -3740 85 -3706 88
rect -3740 54 -3706 85
rect -3644 -85 -3610 -54
rect -3644 -88 -3610 -85
rect -3530 85 -3496 88
rect -3530 54 -3496 85
rect -3434 -85 -3400 -54
rect -3434 -88 -3400 -85
rect -3320 85 -3286 88
rect -3320 54 -3286 85
rect -3224 -85 -3190 -54
rect -3224 -88 -3190 -85
rect -3110 85 -3076 88
rect -3110 54 -3076 85
rect -3014 -85 -2980 -54
rect -3014 -88 -2980 -85
rect -2900 85 -2866 88
rect -2900 54 -2866 85
rect -2804 -85 -2770 -54
rect -2804 -88 -2770 -85
rect -2690 85 -2656 88
rect -2690 54 -2656 85
rect -2594 -85 -2560 -54
rect -2594 -88 -2560 -85
rect -2480 85 -2446 88
rect -2480 54 -2446 85
rect -2384 -85 -2350 -54
rect -2384 -88 -2350 -85
rect -2270 85 -2236 88
rect -2270 54 -2236 85
rect -2174 -85 -2140 -54
rect -2174 -88 -2140 -85
rect -2060 85 -2026 88
rect -2060 54 -2026 85
rect -1964 -85 -1930 -54
rect -1964 -88 -1930 -85
rect -1850 85 -1816 88
rect -1850 54 -1816 85
rect -1754 -85 -1720 -54
rect -1754 -88 -1720 -85
rect -1640 85 -1606 88
rect -1640 54 -1606 85
rect -1544 -85 -1510 -54
rect -1544 -88 -1510 -85
rect -1430 85 -1396 88
rect -1430 54 -1396 85
rect -1334 -85 -1300 -54
rect -1334 -88 -1300 -85
rect -1220 85 -1186 88
rect -1220 54 -1186 85
rect -1124 -85 -1090 -54
rect -1124 -88 -1090 -85
rect -1010 85 -976 88
rect -1010 54 -976 85
rect -914 -85 -880 -54
rect -914 -88 -880 -85
rect -800 85 -766 88
rect -800 54 -766 85
rect -704 -85 -670 -54
rect -704 -88 -670 -85
rect -590 85 -556 88
rect -590 54 -556 85
rect -494 -85 -460 -54
rect -494 -88 -460 -85
rect -380 85 -346 88
rect -380 54 -346 85
rect -284 -85 -250 -54
rect -284 -88 -250 -85
rect -170 85 -136 88
rect -170 54 -136 85
rect -74 -85 -40 -54
rect -74 -88 -40 -85
rect 40 85 74 88
rect 40 54 74 85
rect 136 -85 170 -54
rect 136 -88 170 -85
rect 250 85 284 88
rect 250 54 284 85
rect 346 -85 380 -54
rect 346 -88 380 -85
rect 460 85 494 88
rect 460 54 494 85
rect 556 -85 590 -54
rect 556 -88 590 -85
rect 670 85 704 88
rect 670 54 704 85
rect 766 -85 800 -54
rect 766 -88 800 -85
rect 880 85 914 88
rect 880 54 914 85
rect 976 -85 1010 -54
rect 976 -88 1010 -85
rect 1090 85 1124 88
rect 1090 54 1124 85
rect 1186 -85 1220 -54
rect 1186 -88 1220 -85
rect 1300 85 1334 88
rect 1300 54 1334 85
rect 1396 -85 1430 -54
rect 1396 -88 1430 -85
rect 1510 85 1544 88
rect 1510 54 1544 85
rect 1606 -85 1640 -54
rect 1606 -88 1640 -85
rect 1720 85 1754 88
rect 1720 54 1754 85
rect 1816 -85 1850 -54
rect 1816 -88 1850 -85
rect 1930 85 1964 88
rect 1930 54 1964 85
rect 2026 -85 2060 -54
rect 2026 -88 2060 -85
rect 2140 85 2174 88
rect 2140 54 2174 85
rect 2236 -85 2270 -54
rect 2236 -88 2270 -85
rect 2350 85 2384 88
rect 2350 54 2384 85
rect 2446 -85 2480 -54
rect 2446 -88 2480 -85
rect 2560 85 2594 88
rect 2560 54 2594 85
rect 2656 -85 2690 -54
rect 2656 -88 2690 -85
rect 2770 85 2804 88
rect 2770 54 2804 85
rect 2866 -85 2900 -54
rect 2866 -88 2900 -85
rect 2980 85 3014 88
rect 2980 54 3014 85
rect 3076 -85 3110 -54
rect 3076 -88 3110 -85
rect 3190 85 3224 88
rect 3190 54 3224 85
rect 3286 -85 3320 -54
rect 3286 -88 3320 -85
rect 3400 85 3434 88
rect 3400 54 3434 85
rect 3496 -85 3530 -54
rect 3496 -88 3530 -85
rect 3610 85 3644 88
rect 3610 54 3644 85
rect 3706 -85 3740 -54
rect 3706 -88 3740 -85
rect 3820 85 3854 88
rect 3820 54 3854 85
rect 3916 -85 3950 -54
rect 3916 -88 3950 -85
rect 4030 85 4064 88
rect 4030 54 4064 85
rect 4126 -85 4160 -54
rect 4126 -88 4160 -85
rect -3902 -172 -3868 -138
rect -3482 -172 -3448 -138
rect -3062 -172 -3028 -138
rect -2642 -172 -2608 -138
rect -2222 -172 -2188 -138
rect -1802 -172 -1768 -138
rect -1382 -172 -1348 -138
rect -962 -172 -928 -138
rect -542 -172 -508 -138
rect -122 -172 -88 -138
rect 298 -172 332 -138
rect 718 -172 752 -138
rect 1138 -172 1172 -138
rect 1558 -172 1592 -138
rect 1978 -172 2012 -138
rect 2398 -172 2432 -138
rect 2818 -172 2852 -138
rect 3238 -172 3272 -138
rect 3658 -172 3692 -138
rect 4078 -172 4112 -138
<< metal1 >>
rect -4124 172 -4066 178
rect -4124 138 -4112 172
rect -4078 138 -4066 172
rect -4124 132 -4066 138
rect -3704 172 -3646 178
rect -3704 138 -3692 172
rect -3658 138 -3646 172
rect -3704 132 -3646 138
rect -3284 172 -3226 178
rect -3284 138 -3272 172
rect -3238 138 -3226 172
rect -3284 132 -3226 138
rect -2864 172 -2806 178
rect -2864 138 -2852 172
rect -2818 138 -2806 172
rect -2864 132 -2806 138
rect -2444 172 -2386 178
rect -2444 138 -2432 172
rect -2398 138 -2386 172
rect -2444 132 -2386 138
rect -2024 172 -1966 178
rect -2024 138 -2012 172
rect -1978 138 -1966 172
rect -2024 132 -1966 138
rect -1604 172 -1546 178
rect -1604 138 -1592 172
rect -1558 138 -1546 172
rect -1604 132 -1546 138
rect -1184 172 -1126 178
rect -1184 138 -1172 172
rect -1138 138 -1126 172
rect -1184 132 -1126 138
rect -764 172 -706 178
rect -764 138 -752 172
rect -718 138 -706 172
rect -764 132 -706 138
rect -344 172 -286 178
rect -344 138 -332 172
rect -298 138 -286 172
rect -344 132 -286 138
rect 76 172 134 178
rect 76 138 88 172
rect 122 138 134 172
rect 76 132 134 138
rect 496 172 554 178
rect 496 138 508 172
rect 542 138 554 172
rect 496 132 554 138
rect 916 172 974 178
rect 916 138 928 172
rect 962 138 974 172
rect 916 132 974 138
rect 1336 172 1394 178
rect 1336 138 1348 172
rect 1382 138 1394 172
rect 1336 132 1394 138
rect 1756 172 1814 178
rect 1756 138 1768 172
rect 1802 138 1814 172
rect 1756 132 1814 138
rect 2176 172 2234 178
rect 2176 138 2188 172
rect 2222 138 2234 172
rect 2176 132 2234 138
rect 2596 172 2654 178
rect 2596 138 2608 172
rect 2642 138 2654 172
rect 2596 132 2654 138
rect 3016 172 3074 178
rect 3016 138 3028 172
rect 3062 138 3074 172
rect 3016 132 3074 138
rect 3436 172 3494 178
rect 3436 138 3448 172
rect 3482 138 3494 172
rect 3436 132 3494 138
rect 3856 172 3914 178
rect 3856 138 3868 172
rect 3902 138 3914 172
rect 3856 132 3914 138
rect -4172 88 -4114 94
rect -3962 88 -3904 94
rect -3752 88 -3694 94
rect -3542 88 -3484 94
rect -3332 88 -3274 94
rect -3122 88 -3064 94
rect -2912 88 -2854 94
rect -2702 88 -2644 94
rect -2492 88 -2434 94
rect -2282 88 -2224 94
rect -2072 88 -2014 94
rect -1862 88 -1804 94
rect -1652 88 -1594 94
rect -1442 88 -1384 94
rect -1232 88 -1174 94
rect -1022 88 -964 94
rect -812 88 -754 94
rect -602 88 -544 94
rect -392 88 -334 94
rect -182 88 -124 94
rect 28 88 86 94
rect 238 88 296 94
rect 448 88 506 94
rect 658 88 716 94
rect 868 88 926 94
rect 1078 88 1136 94
rect 1288 88 1346 94
rect 1498 88 1556 94
rect 1708 88 1766 94
rect 1918 88 1976 94
rect 2128 88 2186 94
rect 2338 88 2396 94
rect 2548 88 2606 94
rect 2758 88 2816 94
rect 2968 88 3026 94
rect 3178 88 3236 94
rect 3388 88 3446 94
rect 3598 88 3656 94
rect 3808 88 3866 94
rect 4018 88 4076 94
rect -4172 54 -4160 88
rect -4126 54 -3950 88
rect -3916 54 -3740 88
rect -3706 54 -3530 88
rect -3496 54 -3320 88
rect -3286 54 -3110 88
rect -3076 54 -2900 88
rect -2866 54 -2690 88
rect -2656 54 -2480 88
rect -2446 54 -2270 88
rect -2236 54 -2060 88
rect -2026 54 -1850 88
rect -1816 54 -1640 88
rect -1606 54 -1430 88
rect -1396 54 -1220 88
rect -1186 54 -1010 88
rect -976 54 -800 88
rect -766 54 -590 88
rect -556 54 -380 88
rect -346 54 -170 88
rect -136 54 40 88
rect 74 54 250 88
rect 284 54 460 88
rect 494 54 670 88
rect 704 54 880 88
rect 914 54 1090 88
rect 1124 54 1300 88
rect 1334 54 1510 88
rect 1544 54 1720 88
rect 1754 54 1930 88
rect 1964 54 2140 88
rect 2174 54 2350 88
rect 2384 54 2560 88
rect 2594 54 2770 88
rect 2804 54 2980 88
rect 3014 54 3190 88
rect 3224 54 3400 88
rect 3434 54 3610 88
rect 3644 54 3820 88
rect 3854 54 4030 88
rect 4064 54 4172 88
rect -4172 48 -4114 54
rect -3962 48 -3904 54
rect -3752 48 -3694 54
rect -3542 48 -3484 54
rect -3332 48 -3274 54
rect -3122 48 -3064 54
rect -2912 48 -2854 54
rect -2702 48 -2644 54
rect -2492 48 -2434 54
rect -2282 48 -2224 54
rect -2072 48 -2014 54
rect -1862 48 -1804 54
rect -1652 48 -1594 54
rect -1442 48 -1384 54
rect -1232 48 -1174 54
rect -1022 48 -964 54
rect -812 48 -754 54
rect -602 48 -544 54
rect -392 48 -334 54
rect -182 48 -124 54
rect 28 48 86 54
rect 238 48 296 54
rect 448 48 506 54
rect 658 48 716 54
rect 868 48 926 54
rect 1078 48 1136 54
rect 1288 48 1346 54
rect 1498 48 1556 54
rect 1708 48 1766 54
rect 1918 48 1976 54
rect 2128 48 2186 54
rect 2338 48 2396 54
rect 2548 48 2606 54
rect 2758 48 2816 54
rect 2968 48 3026 54
rect 3178 48 3236 54
rect 3388 48 3446 54
rect 3598 48 3656 54
rect 3808 48 3866 54
rect 4018 48 4076 54
rect -4076 -54 -4018 -48
rect -3866 -54 -3808 -48
rect -3656 -54 -3598 -48
rect -3446 -54 -3388 -48
rect -3236 -54 -3178 -48
rect -3026 -54 -2968 -48
rect -2816 -54 -2758 -48
rect -2606 -54 -2548 -48
rect -2396 -54 -2338 -48
rect -2186 -54 -2128 -48
rect -1976 -54 -1918 -48
rect -1766 -54 -1708 -48
rect -1556 -54 -1498 -48
rect -1346 -54 -1288 -48
rect -1136 -54 -1078 -48
rect -926 -54 -868 -48
rect -716 -54 -658 -48
rect -506 -54 -448 -48
rect -296 -54 -238 -48
rect -86 -54 -28 -48
rect 124 -54 182 -48
rect 334 -54 392 -48
rect 544 -54 602 -48
rect 754 -54 812 -48
rect 964 -54 1022 -48
rect 1174 -54 1232 -48
rect 1384 -54 1442 -48
rect 1594 -54 1652 -48
rect 1804 -54 1862 -48
rect 2014 -54 2072 -48
rect 2224 -54 2282 -48
rect 2434 -54 2492 -48
rect 2644 -54 2702 -48
rect 2854 -54 2912 -48
rect 3064 -54 3122 -48
rect 3274 -54 3332 -48
rect 3484 -54 3542 -48
rect 3694 -54 3752 -48
rect 3904 -54 3962 -48
rect 4114 -54 4172 -48
rect -4172 -88 -4064 -54
rect -4030 -88 -3854 -54
rect -3820 -88 -3644 -54
rect -3610 -88 -3434 -54
rect -3400 -88 -3224 -54
rect -3190 -88 -3014 -54
rect -2980 -88 -2804 -54
rect -2770 -88 -2594 -54
rect -2560 -88 -2384 -54
rect -2350 -88 -2174 -54
rect -2140 -88 -1964 -54
rect -1930 -88 -1754 -54
rect -1720 -88 -1544 -54
rect -1510 -88 -1334 -54
rect -1300 -88 -1124 -54
rect -1090 -88 -914 -54
rect -880 -88 -704 -54
rect -670 -88 -494 -54
rect -460 -88 -284 -54
rect -250 -88 -74 -54
rect -40 -88 136 -54
rect 170 -88 346 -54
rect 380 -88 556 -54
rect 590 -88 766 -54
rect 800 -88 976 -54
rect 1010 -88 1186 -54
rect 1220 -88 1396 -54
rect 1430 -88 1606 -54
rect 1640 -88 1816 -54
rect 1850 -88 2026 -54
rect 2060 -88 2236 -54
rect 2270 -88 2446 -54
rect 2480 -88 2656 -54
rect 2690 -88 2866 -54
rect 2900 -88 3076 -54
rect 3110 -88 3286 -54
rect 3320 -88 3496 -54
rect 3530 -88 3706 -54
rect 3740 -88 3916 -54
rect 3950 -88 4126 -54
rect 4160 -88 4172 -54
rect -4076 -94 -4018 -88
rect -3866 -94 -3808 -88
rect -3656 -94 -3598 -88
rect -3446 -94 -3388 -88
rect -3236 -94 -3178 -88
rect -3026 -94 -2968 -88
rect -2816 -94 -2758 -88
rect -2606 -94 -2548 -88
rect -2396 -94 -2338 -88
rect -2186 -94 -2128 -88
rect -1976 -94 -1918 -88
rect -1766 -94 -1708 -88
rect -1556 -94 -1498 -88
rect -1346 -94 -1288 -88
rect -1136 -94 -1078 -88
rect -926 -94 -868 -88
rect -716 -94 -658 -88
rect -506 -94 -448 -88
rect -296 -94 -238 -88
rect -86 -94 -28 -88
rect 124 -94 182 -88
rect 334 -94 392 -88
rect 544 -94 602 -88
rect 754 -94 812 -88
rect 964 -94 1022 -88
rect 1174 -94 1232 -88
rect 1384 -94 1442 -88
rect 1594 -94 1652 -88
rect 1804 -94 1862 -88
rect 2014 -94 2072 -88
rect 2224 -94 2282 -88
rect 2434 -94 2492 -88
rect 2644 -94 2702 -88
rect 2854 -94 2912 -88
rect 3064 -94 3122 -88
rect 3274 -94 3332 -88
rect 3484 -94 3542 -88
rect 3694 -94 3752 -88
rect 3904 -94 3962 -88
rect 4114 -94 4172 -88
rect -3914 -138 -3856 -132
rect -3914 -172 -3902 -138
rect -3868 -172 -3856 -138
rect -3914 -178 -3856 -172
rect -3494 -138 -3436 -132
rect -3494 -172 -3482 -138
rect -3448 -172 -3436 -138
rect -3494 -178 -3436 -172
rect -3074 -138 -3016 -132
rect -3074 -172 -3062 -138
rect -3028 -172 -3016 -138
rect -3074 -178 -3016 -172
rect -2654 -138 -2596 -132
rect -2654 -172 -2642 -138
rect -2608 -172 -2596 -138
rect -2654 -178 -2596 -172
rect -2234 -138 -2176 -132
rect -2234 -172 -2222 -138
rect -2188 -172 -2176 -138
rect -2234 -178 -2176 -172
rect -1814 -138 -1756 -132
rect -1814 -172 -1802 -138
rect -1768 -172 -1756 -138
rect -1814 -178 -1756 -172
rect -1394 -138 -1336 -132
rect -1394 -172 -1382 -138
rect -1348 -172 -1336 -138
rect -1394 -178 -1336 -172
rect -974 -138 -916 -132
rect -974 -172 -962 -138
rect -928 -172 -916 -138
rect -974 -178 -916 -172
rect -554 -138 -496 -132
rect -554 -172 -542 -138
rect -508 -172 -496 -138
rect -554 -178 -496 -172
rect -134 -138 -76 -132
rect -134 -172 -122 -138
rect -88 -172 -76 -138
rect -134 -178 -76 -172
rect 286 -138 344 -132
rect 286 -172 298 -138
rect 332 -172 344 -138
rect 286 -178 344 -172
rect 706 -138 764 -132
rect 706 -172 718 -138
rect 752 -172 764 -138
rect 706 -178 764 -172
rect 1126 -138 1184 -132
rect 1126 -172 1138 -138
rect 1172 -172 1184 -138
rect 1126 -178 1184 -172
rect 1546 -138 1604 -132
rect 1546 -172 1558 -138
rect 1592 -172 1604 -138
rect 1546 -178 1604 -172
rect 1966 -138 2024 -132
rect 1966 -172 1978 -138
rect 2012 -172 2024 -138
rect 1966 -178 2024 -172
rect 2386 -138 2444 -132
rect 2386 -172 2398 -138
rect 2432 -172 2444 -138
rect 2386 -178 2444 -172
rect 2806 -138 2864 -132
rect 2806 -172 2818 -138
rect 2852 -172 2864 -138
rect 2806 -178 2864 -172
rect 3226 -138 3284 -132
rect 3226 -172 3238 -138
rect 3272 -172 3284 -138
rect 3226 -178 3284 -172
rect 3646 -138 3704 -132
rect 3646 -172 3658 -138
rect 3692 -172 3704 -138
rect 3646 -178 3704 -172
rect 4066 -138 4124 -132
rect 4066 -172 4078 -138
rect 4112 -172 4124 -138
rect 4066 -178 4124 -172
<< end >>
