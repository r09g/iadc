magic
tech sky130A
magscale 1 2
timestamp 1654585951
<< metal3 >>
rect 79999 131172 80009 131408
rect 80245 131172 80255 131408
rect 40081 109395 40317 114465
rect 68084 109367 68320 114465
rect 80009 113632 80245 131172
rect 114815 99999 120001 100235
rect 93224 92601 120001 92837
rect 114890 85163 120001 85399
rect 109850 79125 120001 79361
rect -51382 77232 -45234 77292
rect -27446 77232 -22586 77292
rect 112280 74910 120001 75146
rect -12556 74178 1476 74179
rect -22849 74060 -22586 74120
rect -12654 73942 -12644 74178
rect -12408 73943 1476 74178
rect -12408 73942 -12398 73943
rect -51382 73816 -48635 73876
rect 114815 71171 120001 71407
rect -28366 71010 -22586 71070
rect -51382 70400 -44682 70460
rect -33334 67960 -22586 68020
rect 103602 67576 120001 67812
rect -51382 66984 -42474 67044
rect -22744 65074 -16420 65076
rect -22744 64840 -16650 65074
rect -16660 64838 -16650 64840
rect -16414 64838 -16404 65074
rect 114823 64190 120001 64426
rect -51382 63446 -51119 63506
rect -27354 61860 -22586 61920
rect -9268 61572 9074 61593
rect -9268 61357 -9256 61572
rect -9266 61336 -9256 61357
rect -9020 61357 9074 61572
rect -9020 61336 -9010 61357
rect 112240 60882 120001 61118
rect -51382 60030 -45510 60090
rect -33702 58810 -22586 58870
rect 109895 57420 120001 57656
rect -51382 56614 -39990 56674
rect -22724 55612 -9260 55848
rect -9024 55612 -9014 55848
rect 107700 54257 120001 54493
rect -51382 53198 -34099 53258
rect -26802 52710 -22586 52770
rect -51382 49660 -35850 49720
rect -22778 49560 -12644 49796
rect -12408 49560 -12398 49796
rect 0 48959 16511 49195
rect 104876 46522 120001 46758
rect 0 41418 16508 41654
rect 104793 29588 120001 29824
rect 104809 22648 120001 22884
rect 55973 2 56209 5159
<< via3 >>
rect 80009 131172 80245 131408
rect -12644 73942 -12408 74178
rect -16650 64838 -16414 65074
rect -9256 61336 -9020 61572
rect -9260 55612 -9024 55848
rect -12644 49560 -12408 49796
<< metal4 >>
rect 80008 131408 80246 131409
rect -16662 131172 80009 131408
rect 80245 131172 80246 131408
rect -16652 65075 -16416 131172
rect 80008 131171 80246 131172
rect -3940 75048 6128 75112
rect -12645 74178 -12407 74179
rect -12645 73942 -12644 74178
rect -12408 73942 -12407 74178
rect -12645 73941 -12407 73942
rect -16652 65074 -16413 65075
rect -16652 64838 -16650 65074
rect -16414 64838 -16413 65074
rect -16652 64837 -16413 64838
rect -16652 64812 -16416 64837
rect -12644 49797 -12408 73941
rect -3940 73276 -3876 75048
rect -2040 73340 6128 75048
rect -2040 73276 7880 73340
rect -9257 61572 -9019 61573
rect -9257 61336 -9256 61572
rect -9020 61336 -9019 61572
rect -9257 61335 -9019 61336
rect -9256 55849 -9020 61335
rect -9261 55848 -9020 55849
rect -9261 55612 -9260 55848
rect -9024 55782 -9020 55848
rect -9024 55612 -9023 55782
rect -9261 55611 -9023 55612
rect -12645 49796 -12407 49797
rect -12645 49560 -12644 49796
rect -12408 49560 -12407 49796
rect -12645 49559 -12407 49560
rect 1 6003 2083 8003
rect 1 2003 6083 4003
<< via4 >>
rect -3876 73212 -2040 75048
rect 6128 73340 7964 75176
<< metal5 >>
rect 6104 75176 7988 75200
rect -3900 75048 -2016 75072
rect -3900 74984 -3876 75048
rect -24928 73212 -3876 74984
rect -2040 73212 -2016 75048
rect 6104 73340 6128 75176
rect 7964 73340 7988 75176
rect 6104 73316 7988 73340
rect -24928 73188 -2016 73212
rect -24928 73148 -2830 73188
rect -24850 54782 4001 56782
use analog_top  analog_top_0
timestamp 1654583406
transform 1 0 57094 0 1 24024
box -57094 -24022 62907 90442
use digital_top  digital_top_0
timestamp 1654583406
transform -1 0 -22586 0 1 49556
box 0 0 28796 27744
<< labels >>
flabel metal3 -51336 77260 -51336 77260 1 FreeSans 3200 0 0 0 data_out_6
flabel metal3 -51322 73844 -51322 73844 1 FreeSans 3200 0 0 0 data_out_5
flabel metal3 -51310 70428 -51310 70428 1 FreeSans 3200 0 0 0 data_out_4
flabel metal3 -51310 67008 -51310 67008 1 FreeSans 3200 0 0 0 data_out_3
flabel metal3 -51302 63474 -51302 63474 1 FreeSans 3200 0 0 0 data_out_2
flabel metal5 -22622 74092 -22622 74092 1 FreeSans 3200 0 0 0 data_out_8
flabel metal3 -22664 71038 -22664 71038 1 FreeSans 3200 0 0 0 data_out_9
flabel metal3 -22672 77272 -22672 77272 1 FreeSans 3200 0 0 0 data_out_7
flabel metal3 -22676 67992 -22676 67992 1 FreeSans 3200 0 0 0 data_out_10
flabel metal3 -22642 64986 -22642 64986 1 FreeSans 3200 0 0 0 clk
flabel metal3 -22672 61894 -22672 61894 1 FreeSans 3200 0 0 0 sclk
flabel metal3 -22658 58842 -22658 58842 1 FreeSans 3200 0 0 0 data_out_11
flabel metal5 -16090 55724 -16090 55724 1 FreeSans 3200 0 0 0 mod_op
flabel metal3 -22666 52736 -22666 52736 1 FreeSans 3200 0 0 0 cs_n
flabel metal3 -22420 49676 -22420 49686 1 FreeSans 3200 0 0 0 rst_n
flabel metal3 -51304 49692 -51304 49692 1 FreeSans 3200 0 0 0 serial_data_out
flabel metal3 -51322 56646 -51322 56646 1 FreeSans 3200 0 0 0 data_out_0
flabel metal3 -51312 60056 -51312 60056 1 FreeSans 3200 0 0 0 data_out_1
flabel metal3 -51296 53228 -51296 53228 1 FreeSans 3200 0 0 0 new_data
flabel metal3 1562 49086 1562 49086 1 FreeSans 3200 0 0 0 ip
flabel metal3 2148 41534 2148 41534 1 FreeSans 3200 0 0 0 in
flabel metal4 672 6976 672 6976 1 FreeSans 3200 0 0 0 VDD
flabel metal4 542 2938 542 2938 1 FreeSans 3200 0 0 0 VSS
flabel metal3 56082 670 56082 670 1 FreeSans 3200 0 0 0 i_bias_1
flabel metal3 118940 29730 118940 29730 1 FreeSans 3200 0 0 0 a_probe_2
flabel metal3 118762 22744 118762 22744 1 FreeSans 3200 0 0 0 a_probe_3
flabel metal3 118950 46648 118950 46648 1 FreeSans 3200 0 0 0 a_probe_0
flabel metal3 118798 54340 118798 54340 1 FreeSans 3200 0 0 0 d_probe_3
flabel metal3 118798 57566 118798 57566 1 FreeSans 3200 0 0 0 d_probe_2
flabel metal3 118742 60962 118742 60962 1 FreeSans 3200 0 0 0 d_clk_grp_2_ctrl_1
flabel metal3 118598 64324 118598 64324 1 FreeSans 3200 0 0 0 d_clk_grp_2_ctrl_0
flabel metal3 119018 67684 119018 67684 1 FreeSans 3200 0 0 0 d_probe_1
flabel metal3 118846 71310 118846 71310 1 FreeSans 3200 0 0 0 d_probe_0
flabel metal3 118904 75034 118904 75034 1 FreeSans 3200 0 0 0 d_clk_grp_1_ctrl_1
flabel metal3 118618 79234 118618 79234 1 FreeSans 3200 0 0 0 d_clk_grp_1_ctrl_0
flabel metal3 119176 85292 119176 85292 1 FreeSans 3200 0 0 0 debug
flabel metal3 118902 92728 118902 92728 1 FreeSans 3200 0 0 0 a_mod_grp_ctrl_0
flabel metal3 119190 100140 119190 100140 1 FreeSans 3200 0 0 0 a_mod_grp_ctrl_1
flabel metal3 68190 113976 68190 113996 1 FreeSans 3200 0 0 0 i_bias_2
flabel metal3 40188 113976 40188 113976 1 FreeSans 3200 0 0 0 a_probe_1
<< end >>
