* SPICE3 file created from transmission_gate_flat.ext - technology: sky130A

.subckt transmission_gate_flat in out en en_b
X0 out en in VSS sky130_fd_pr__nfet_01v8 ad=1.537e+12p pd=1.118e+07u as=1.537e+12p ps=1.118e+07u w=5.3e+06u l=150000u
X1 out en_b in VDD sky130_fd_pr__pfet_01v8 ad=3.973e+12p pd=2.798e+07u as=3.973e+12p ps=2.798e+07u w=1.37e+07u l=150000u
C0 VDD in 1.80fF
C1 en_b in 0.11fF
C2 in en 0.54fF
C3 out VDD 2.10fF
C4 en_b out 0.06fF
C5 out en 0.12fF
C6 en_b VDD 0.34fF
C7 VDD en 0.01fF
C8 en_b en 0.04fF
C9 out in 5.94fF
C10 en VSS 0.59fF
C11 in VSS 1.74fF
C12 en_b VSS 0.09fF
C13 out VSS 1.58fF
C14 VDD VSS 4.69fF **FLOATING
.ends
