* SPICE3 file created from transmission_gate_flat.ext - technology: sky130A

.subckt transmission_gate_flat in out en en_b VDD VSS
X0 out en in VSS sky130_fd_pr__nfet_01v8 ad=1.537e+12p pd=1.118e+07u as=1.537e+12p ps=1.118e+07u w=5.3e+06u l=150000u
X1 out en_b in VDD sky130_fd_pr__pfet_01v8 ad=3.973e+12p pd=2.798e+07u as=3.973e+12p ps=2.798e+07u w=1.37e+07u l=150000u
C0 VDD in 1.80fF
C1 en_b in 0.11fF
C2 in en 0.54fF
C3 out VDD 2.10fF
C4 en_b out 0.06fF
C5 out en 0.12fF
C6 en_b VDD 0.34fF
C7 VDD en 0.01fF
C8 en_b en 0.04fF
C9 out in 5.94fF
C10 en VSS 0.59fF
C11 in VSS 1.74fF
C12 en_b VSS 0.09fF
C13 out VSS 1.58fF
C14 VDD VSS 4.69fF
.ends
**.subckt transmission_gate_tb
x2 clk GND GND VDD VDD net1 sky130_fd_sc_hd__inv_4
V2 VDD GND 1.8
V3 clk GND 1.8
V1 in GND DC 0.9
x1 in n1 clk net1 VDD VSS transmission_gate_flat
x3 __UNCONNECTED_PIN__0 out clk net1 VDD VSS transmission_gate_flat
C1 out GND 1p m=1
XM1 n1 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
**** begin user architecture code


.options savecurrents
.control
op
print v(n1)
write transmission_gate_tb_sim_post.raw
.endc



** opencircuitdesign pdks install
.lib /farmshare/home/classes/ee/372/PDKs/open_pdks_1.0.310/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc /farmshare/home/classes/ee/372/PDKs/open_pdks_1.0.310/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=4
* sym_path:
*+ /home/users/yaqingx/EE372/incremental_delta_sigma_adc/design/analog_modulator/schematic/transmission_gate.sym
* sch_path:
*+ /home/users/yaqingx/EE372/incremental_delta_sigma_adc/design/analog_modulator/schematic/transmission_gate.sch
*.subckt transmission_gate  in out en en_b  VDD  VSS     N=1 W_N=5.3 L_N=0.15 W_P=13.7 L_P=0.15
*.iopin in
*.iopin out
*.ipin en
*.ipin en_b
*XM1 out en in VSS sky130_fd_pr__nfet_01v8 L='L_N' W='W_N' nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
*+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
*+ sa=0 sb=0 sd=0 mult='N' m='N' 
*XM2 out en_b in VDD sky130_fd_pr__pfet_01v8 L='L_P' W='W_P' nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
*+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
*+ sa=0 sb=0 sd=0 mult='N' m='N' 
*.ends

.GLOBAL GND
.GLOBAL VDD
** flattened .save nodes
.end
