
x2 clk GND GND VDD VDD net1 sky130_fd_sc_hd__inv_4
V2 VDD GND 1.8
V3 clk GND DC 0 PULSE(0 1.8 1n 10p 10p 1 1)
V1 in GND DC 1.8
x1 in out clk net1 VDD VSS transmission_gate_flat
C1 out GND 1p m=1

.options savecurrents
.ic v(out)=0
.control
tran 0.05n 3n
plot v(out)
write transmission_gate_tb.raw
.endc

.lib /farmshare/home/classes/ee/372/PDKs/open_pdks_1.0.310/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc /farmshare/home/classes/ee/372/PDKs/open_pdks_1.0.310/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


.GLOBAL GND
.GLOBAL VDD
.end
