* NGSPICE file created from comparator_flat.ext - technology: sky130A

.subckt comparator_flat clk ip in outp outn VDD VSS
X0 VSS outp a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=3.6639e+12p pd=3.788e+07u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1 VDD sky130_fd_sc_hd__nand2_4_1/A outn VDD sky130_fd_pr__pfet_01v8_hvt ad=5.351e+12p pd=5.194e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X2 VDD a_177_3251# sky130_fd_sc_hd__nand2_4_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 outn sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=6.375e+11p pd=6.55e+06u as=0p ps=0u w=500000u l=150000u
X5 VDD clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.4e+11p ps=6.56e+06u w=500000u l=150000u
X6 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=3.24e+06u as=8.05e+11p ps=8.22e+06u w=500000u l=150000u
X7 a_282_408# in a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=1.5015e+12p pd=1.504e+07u as=8.05e+11p ps=8.22e+06u w=500000u l=150000u
X8 VSS outp a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VDD sky130_fd_sc_hd__buf_2_0/A a_721_3251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11 a_1067_3524# sky130_fd_sc_hd__nand2_4_1/A outn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X12 outp sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X13 VSS a_177_3251# sky130_fd_sc_hd__nand2_4_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X15 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=3.24e+06u as=0p ps=0u w=500000u l=150000u
X16 VDD outp outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 outn outp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 outp sky130_fd_sc_hd__nand2_4_0/A a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X19 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X20 outn outp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VDD sky130_fd_sc_hd__buf_2_1/A a_177_3251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X23 a_475_1219# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X24 VDD outn outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VDD sky130_fd_sc_hd__nand2_4_1/A outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VSS a_721_3251# sky130_fd_sc_hd__nand2_4_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X27 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X29 a_282_408# ip a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X30 a_282_408# ip a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X31 a_n16_2554# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X32 a_475_1219# in a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X33 a_282_408# in a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X34 VSS VSS a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X35 a_203_3524# outn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X37 a_n16_2554# ip a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X38 outn sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VDD sky130_fd_sc_hd__nand2_4_0/A outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VSS sky130_fd_sc_hd__buf_2_1/A a_177_3251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X42 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X43 outp sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 sky130_fd_sc_hd__buf_2_1/A clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X45 sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X46 VDD a_721_3251# sky130_fd_sc_hd__nand2_4_1/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X47 VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X48 a_203_3524# sky130_fd_sc_hd__nand2_4_0/A outp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 VDD clk a_n16_2554# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
X50 a_475_1219# clk VDD VDD sky130_fd_pr__pfet_01v8 ad=1.425e+11p pd=1.57e+06u as=0p ps=0u w=500000u l=150000u
X51 a_n16_2554# ip a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X52 outp sky130_fd_sc_hd__nand2_4_0/A a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X53 a_1067_3524# outp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X54 outp outn VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 VDD outn outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 outn sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X58 VSS VSS a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X59 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X60 a_n16_2554# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X61 outp outn VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 VSS outn a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X63 a_203_3524# outn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X64 VDD sky130_fd_sc_hd__nand2_4_0/A outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_1067_3524# sky130_fd_sc_hd__nand2_4_1/A outn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X66 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X67 VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X68 outn sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X69 a_282_408# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X70 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X71 VDD outp outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 VSS outn a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X73 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 VDD VDD sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X75 a_475_1219# in a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X76 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X77 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X78 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X79 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X80 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X81 a_203_3524# sky130_fd_sc_hd__nand2_4_0/A outp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X82 a_475_1219# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X83 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X84 a_1067_3524# outp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X85 VSS sky130_fd_sc_hd__buf_2_0/A a_721_3251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X86 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X87 VSS VSS a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
.ends

