magic
tech sky130A
magscale 1 2
timestamp 1654725802
<< nwell >>
rect 162 468 2977 1118
<< pwell >>
rect 162 6 2977 468
rect 1430 4 1686 6
<< nmos >>
rect 362 216 392 320
rect 458 216 488 320
rect 554 216 584 320
rect 650 216 680 320
rect 746 216 776 320
rect 842 216 872 320
rect 938 216 968 320
rect 1034 216 1064 320
rect 1130 216 1160 320
rect 1226 216 1256 320
rect 1538 222 1568 322
rect 1883 216 1913 320
rect 1979 216 2009 320
rect 2075 216 2105 320
rect 2171 216 2201 320
rect 2267 216 2297 320
rect 2363 216 2393 320
rect 2459 216 2489 320
rect 2555 216 2585 320
rect 2651 216 2681 320
rect 2747 216 2777 320
<< pmos >>
rect 362 626 392 898
rect 458 626 488 898
rect 554 626 584 898
rect 650 626 680 898
rect 746 626 776 898
rect 842 626 872 898
rect 938 626 968 898
rect 1034 626 1064 898
rect 1130 626 1160 898
rect 1226 626 1256 898
rect 1883 626 1913 898
rect 1979 626 2009 898
rect 2075 626 2105 898
rect 2171 626 2201 898
rect 2267 626 2297 898
rect 2363 626 2393 898
rect 2459 626 2489 898
rect 2555 626 2585 898
rect 2651 626 2681 898
rect 2747 626 2777 898
<< ndiff >>
rect 300 308 362 320
rect 300 228 312 308
rect 346 228 362 308
rect 300 216 362 228
rect 392 308 458 320
rect 392 228 408 308
rect 442 228 458 308
rect 392 216 458 228
rect 488 308 554 320
rect 488 228 504 308
rect 538 228 554 308
rect 488 216 554 228
rect 584 308 650 320
rect 584 228 600 308
rect 634 228 650 308
rect 584 216 650 228
rect 680 308 746 320
rect 680 228 696 308
rect 730 228 746 308
rect 680 216 746 228
rect 776 308 842 320
rect 776 228 792 308
rect 826 228 842 308
rect 776 216 842 228
rect 872 308 938 320
rect 872 228 888 308
rect 922 228 938 308
rect 872 216 938 228
rect 968 308 1034 320
rect 968 228 984 308
rect 1018 228 1034 308
rect 968 216 1034 228
rect 1064 308 1130 320
rect 1064 228 1080 308
rect 1114 228 1130 308
rect 1064 216 1130 228
rect 1160 308 1226 320
rect 1160 228 1176 308
rect 1210 228 1226 308
rect 1160 216 1226 228
rect 1256 308 1318 320
rect 1256 228 1272 308
rect 1306 228 1318 308
rect 1256 216 1318 228
rect 1480 310 1538 322
rect 1480 234 1492 310
rect 1526 234 1538 310
rect 1480 222 1538 234
rect 1568 310 1626 322
rect 1568 234 1580 310
rect 1614 234 1626 310
rect 1568 222 1626 234
rect 1821 308 1883 320
rect 1821 228 1833 308
rect 1867 228 1883 308
rect 1821 216 1883 228
rect 1913 308 1979 320
rect 1913 228 1929 308
rect 1963 228 1979 308
rect 1913 216 1979 228
rect 2009 308 2075 320
rect 2009 228 2025 308
rect 2059 228 2075 308
rect 2009 216 2075 228
rect 2105 308 2171 320
rect 2105 228 2121 308
rect 2155 228 2171 308
rect 2105 216 2171 228
rect 2201 308 2267 320
rect 2201 228 2217 308
rect 2251 228 2267 308
rect 2201 216 2267 228
rect 2297 308 2363 320
rect 2297 228 2313 308
rect 2347 228 2363 308
rect 2297 216 2363 228
rect 2393 308 2459 320
rect 2393 228 2409 308
rect 2443 228 2459 308
rect 2393 216 2459 228
rect 2489 308 2555 320
rect 2489 228 2505 308
rect 2539 228 2555 308
rect 2489 216 2555 228
rect 2585 308 2651 320
rect 2585 228 2601 308
rect 2635 228 2651 308
rect 2585 216 2651 228
rect 2681 308 2747 320
rect 2681 228 2697 308
rect 2731 228 2747 308
rect 2681 216 2747 228
rect 2777 308 2839 320
rect 2777 228 2793 308
rect 2827 228 2839 308
rect 2777 216 2839 228
<< pdiff >>
rect 300 886 362 898
rect 300 638 312 886
rect 346 638 362 886
rect 300 626 362 638
rect 392 886 458 898
rect 392 638 408 886
rect 442 638 458 886
rect 392 626 458 638
rect 488 886 554 898
rect 488 638 504 886
rect 538 638 554 886
rect 488 626 554 638
rect 584 886 650 898
rect 584 638 600 886
rect 634 638 650 886
rect 584 626 650 638
rect 680 886 746 898
rect 680 638 696 886
rect 730 638 746 886
rect 680 626 746 638
rect 776 886 842 898
rect 776 638 792 886
rect 826 638 842 886
rect 776 626 842 638
rect 872 886 938 898
rect 872 638 888 886
rect 922 638 938 886
rect 872 626 938 638
rect 968 886 1034 898
rect 968 638 984 886
rect 1018 638 1034 886
rect 968 626 1034 638
rect 1064 886 1130 898
rect 1064 638 1080 886
rect 1114 638 1130 886
rect 1064 626 1130 638
rect 1160 886 1226 898
rect 1160 638 1176 886
rect 1210 638 1226 886
rect 1160 626 1226 638
rect 1256 886 1318 898
rect 1256 638 1272 886
rect 1306 638 1318 886
rect 1256 626 1318 638
rect 1821 886 1883 898
rect 1821 638 1833 886
rect 1867 638 1883 886
rect 1821 626 1883 638
rect 1913 886 1979 898
rect 1913 638 1929 886
rect 1963 638 1979 886
rect 1913 626 1979 638
rect 2009 886 2075 898
rect 2009 638 2025 886
rect 2059 638 2075 886
rect 2009 626 2075 638
rect 2105 886 2171 898
rect 2105 638 2121 886
rect 2155 638 2171 886
rect 2105 626 2171 638
rect 2201 886 2267 898
rect 2201 638 2217 886
rect 2251 638 2267 886
rect 2201 626 2267 638
rect 2297 886 2363 898
rect 2297 638 2313 886
rect 2347 638 2363 886
rect 2297 626 2363 638
rect 2393 886 2459 898
rect 2393 638 2409 886
rect 2443 638 2459 886
rect 2393 626 2459 638
rect 2489 886 2555 898
rect 2489 638 2505 886
rect 2539 638 2555 886
rect 2489 626 2555 638
rect 2585 886 2651 898
rect 2585 638 2601 886
rect 2635 638 2651 886
rect 2585 626 2651 638
rect 2681 886 2747 898
rect 2681 638 2697 886
rect 2731 638 2747 886
rect 2681 626 2747 638
rect 2777 886 2839 898
rect 2777 638 2793 886
rect 2827 638 2839 886
rect 2777 626 2839 638
<< ndiffc >>
rect 312 228 346 308
rect 408 228 442 308
rect 504 228 538 308
rect 600 228 634 308
rect 696 228 730 308
rect 792 228 826 308
rect 888 228 922 308
rect 984 228 1018 308
rect 1080 228 1114 308
rect 1176 228 1210 308
rect 1272 228 1306 308
rect 1492 234 1526 310
rect 1580 234 1614 310
rect 1833 228 1867 308
rect 1929 228 1963 308
rect 2025 228 2059 308
rect 2121 228 2155 308
rect 2217 228 2251 308
rect 2313 228 2347 308
rect 2409 228 2443 308
rect 2505 228 2539 308
rect 2601 228 2635 308
rect 2697 228 2731 308
rect 2793 228 2827 308
<< pdiffc >>
rect 312 638 346 886
rect 408 638 442 886
rect 504 638 538 886
rect 600 638 634 886
rect 696 638 730 886
rect 792 638 826 886
rect 888 638 922 886
rect 984 638 1018 886
rect 1080 638 1114 886
rect 1176 638 1210 886
rect 1272 638 1306 886
rect 1833 638 1867 886
rect 1929 638 1963 886
rect 2025 638 2059 886
rect 2121 638 2155 886
rect 2217 638 2251 886
rect 2313 638 2347 886
rect 2409 638 2443 886
rect 2505 638 2539 886
rect 2601 638 2635 886
rect 2697 638 2731 886
rect 2793 638 2827 886
<< psubdiff >>
rect 198 398 294 432
rect 1324 398 1420 432
rect 198 336 232 398
rect 1386 336 1420 398
rect 1719 398 1815 432
rect 2845 398 2941 432
rect 198 76 232 138
rect 1719 336 1753 398
rect 1386 76 1420 138
rect 198 42 294 76
rect 1324 42 1420 76
rect 2907 336 2941 398
rect 1719 76 1753 138
rect 2907 76 2941 138
rect 1719 42 1815 76
rect 2845 42 2941 76
<< nsubdiff >>
rect 198 1048 294 1082
rect 1324 1048 1420 1082
rect 198 986 232 1048
rect 1386 986 1420 1048
rect 198 538 232 600
rect 1386 538 1420 600
rect 198 504 294 538
rect 1324 504 1420 538
rect 1719 1048 1815 1082
rect 2845 1048 2941 1082
rect 1719 986 1753 1048
rect 2907 986 2941 1048
rect 1719 538 1753 600
rect 2907 538 2941 600
rect 1719 504 1815 538
rect 2845 504 2941 538
<< psubdiffcont >>
rect 294 398 1324 432
rect 198 138 232 336
rect 1815 398 2845 432
rect 1386 138 1420 336
rect 294 42 1324 76
rect 1719 138 1753 336
rect 2907 138 2941 336
rect 1815 42 2845 76
<< nsubdiffcont >>
rect 294 1048 1324 1082
rect 198 600 232 986
rect 1386 600 1420 986
rect 294 504 1324 538
rect 1815 1048 2845 1082
rect 1719 600 1753 986
rect 2907 600 2941 986
rect 1815 504 2845 538
<< poly >>
rect 296 980 1322 996
rect 296 946 312 980
rect 346 946 504 980
rect 538 946 696 980
rect 730 946 888 980
rect 922 946 1080 980
rect 1114 946 1272 980
rect 1306 946 1322 980
rect 296 930 1322 946
rect 362 898 392 930
rect 458 898 488 930
rect 554 898 584 930
rect 650 898 680 930
rect 746 898 776 930
rect 842 898 872 930
rect 938 898 968 930
rect 1034 898 1064 930
rect 1130 898 1160 930
rect 1226 898 1256 930
rect 362 600 392 626
rect 458 600 488 626
rect 554 600 584 626
rect 650 600 680 626
rect 746 600 776 626
rect 842 600 872 626
rect 938 600 968 626
rect 1034 600 1064 626
rect 1130 600 1160 626
rect 1226 600 1256 626
rect 1817 980 2843 996
rect 1817 946 1833 980
rect 1867 946 2025 980
rect 2059 946 2217 980
rect 2251 946 2409 980
rect 2443 946 2601 980
rect 2635 946 2793 980
rect 2827 946 2843 980
rect 1817 930 2843 946
rect 1883 898 1913 930
rect 1979 898 2009 930
rect 2075 898 2105 930
rect 2171 898 2201 930
rect 2267 898 2297 930
rect 2363 898 2393 930
rect 2459 898 2489 930
rect 2555 898 2585 930
rect 2651 898 2681 930
rect 2747 898 2777 930
rect 1883 600 1913 626
rect 1979 600 2009 626
rect 2075 600 2105 626
rect 2171 600 2201 626
rect 2267 600 2297 626
rect 2363 600 2393 626
rect 2459 600 2489 626
rect 2555 600 2585 626
rect 2651 600 2681 626
rect 2747 600 2777 626
rect 362 320 392 346
rect 458 320 488 346
rect 554 320 584 346
rect 650 320 680 346
rect 746 320 776 346
rect 842 320 872 346
rect 938 320 968 346
rect 1034 320 1064 346
rect 1130 320 1160 346
rect 1226 320 1256 346
rect 1520 394 1586 410
rect 1520 360 1536 394
rect 1570 360 1586 394
rect 1520 344 1586 360
rect 362 185 392 216
rect 458 185 488 216
rect 554 185 584 216
rect 650 185 680 216
rect 746 185 776 216
rect 842 185 872 216
rect 938 185 968 216
rect 1034 185 1064 216
rect 1130 185 1160 216
rect 1226 185 1256 216
rect 296 169 1322 185
rect 296 135 312 169
rect 346 135 504 169
rect 538 135 696 169
rect 730 135 888 169
rect 922 135 1080 169
rect 1114 135 1272 169
rect 1306 135 1322 169
rect 296 119 1322 135
rect 1538 322 1568 344
rect 1538 196 1568 222
rect 1883 320 1913 346
rect 1979 320 2009 346
rect 2075 320 2105 346
rect 2171 320 2201 346
rect 2267 320 2297 346
rect 2363 320 2393 346
rect 2459 320 2489 346
rect 2555 320 2585 346
rect 2651 320 2681 346
rect 2747 320 2777 346
rect 1883 185 1913 216
rect 1979 185 2009 216
rect 2075 185 2105 216
rect 2171 185 2201 216
rect 2267 185 2297 216
rect 2363 185 2393 216
rect 2459 185 2489 216
rect 2555 185 2585 216
rect 2651 185 2681 216
rect 2747 185 2777 216
rect 1817 169 2843 185
rect 1817 135 1833 169
rect 1867 135 2025 169
rect 2059 135 2217 169
rect 2251 135 2409 169
rect 2443 135 2601 169
rect 2635 135 2793 169
rect 2827 135 2843 169
rect 1817 119 2843 135
<< polycont >>
rect 312 946 346 980
rect 504 946 538 980
rect 696 946 730 980
rect 888 946 922 980
rect 1080 946 1114 980
rect 1272 946 1306 980
rect 1833 946 1867 980
rect 2025 946 2059 980
rect 2217 946 2251 980
rect 2409 946 2443 980
rect 2601 946 2635 980
rect 2793 946 2827 980
rect 1536 360 1570 394
rect 312 135 346 169
rect 504 135 538 169
rect 696 135 730 169
rect 888 135 922 169
rect 1080 135 1114 169
rect 1272 135 1306 169
rect 1833 135 1867 169
rect 2025 135 2059 169
rect 2217 135 2251 169
rect 2409 135 2443 169
rect 2601 135 2635 169
rect 2793 135 2827 169
<< locali >>
rect 198 1048 294 1082
rect 1324 1048 1815 1082
rect 2845 1048 2941 1082
rect 198 986 232 1048
rect 1386 1014 1759 1048
rect 296 980 1322 988
rect 296 946 312 980
rect 346 946 504 980
rect 538 946 696 980
rect 730 946 888 980
rect 922 946 1080 980
rect 1114 946 1272 980
rect 1306 946 1322 980
rect 296 938 1322 946
rect 1386 986 1420 1014
rect 312 886 346 902
rect 312 622 346 638
rect 408 886 442 902
rect 408 622 442 638
rect 504 886 538 902
rect 504 622 538 638
rect 600 886 634 902
rect 600 622 634 638
rect 696 886 730 902
rect 696 622 730 638
rect 792 886 826 902
rect 792 622 826 638
rect 888 886 922 902
rect 888 622 922 638
rect 984 886 1018 902
rect 984 622 1018 638
rect 1080 886 1114 902
rect 1080 622 1114 638
rect 1176 886 1210 902
rect 1176 622 1210 638
rect 1272 886 1306 902
rect 1272 622 1306 638
rect 198 538 232 600
rect 1386 538 1420 600
rect 198 504 294 538
rect 1324 504 1420 538
rect 1719 986 1753 1014
rect 1817 980 2843 988
rect 1817 946 1833 980
rect 1867 946 2025 980
rect 2059 946 2217 980
rect 2251 946 2409 980
rect 2443 946 2601 980
rect 2635 946 2793 980
rect 2827 946 2843 980
rect 1817 938 2843 946
rect 2907 986 2941 1048
rect 1833 886 1867 902
rect 1833 622 1867 638
rect 1929 886 1963 902
rect 1929 622 1963 638
rect 2025 886 2059 902
rect 2025 622 2059 638
rect 2121 886 2155 902
rect 2121 622 2155 638
rect 2217 886 2251 902
rect 2217 622 2251 638
rect 2313 886 2347 902
rect 2313 622 2347 638
rect 2409 886 2443 902
rect 2409 622 2443 638
rect 2505 886 2539 902
rect 2505 622 2539 638
rect 2601 886 2635 902
rect 2601 622 2635 638
rect 2697 886 2731 902
rect 2697 622 2731 638
rect 2793 886 2827 902
rect 2793 622 2827 638
rect 1719 538 1753 600
rect 2907 538 2941 600
rect 1719 504 1815 538
rect 2845 504 2941 538
rect 198 398 294 432
rect 1324 398 1420 432
rect 198 336 232 398
rect 1386 336 1420 398
rect 1719 398 1815 432
rect 2845 398 2941 432
rect 1520 360 1536 394
rect 1570 360 1586 394
rect 312 308 346 324
rect 312 212 346 228
rect 408 308 442 324
rect 408 212 442 228
rect 504 308 538 324
rect 504 212 538 228
rect 600 308 634 324
rect 600 212 634 228
rect 696 308 730 324
rect 696 212 730 228
rect 792 308 826 324
rect 792 212 826 228
rect 888 308 922 324
rect 888 212 922 228
rect 984 308 1018 324
rect 984 212 1018 228
rect 1080 308 1114 324
rect 1080 212 1114 228
rect 1176 308 1210 324
rect 1176 212 1210 228
rect 1272 308 1306 324
rect 1272 212 1306 228
rect 1719 336 1753 398
rect 198 76 232 138
rect 296 169 1322 177
rect 296 135 312 169
rect 346 135 504 169
rect 538 135 696 169
rect 730 135 888 169
rect 922 135 1080 169
rect 1114 135 1272 169
rect 1306 135 1322 169
rect 296 127 1322 135
rect 1492 310 1526 326
rect 1492 218 1526 234
rect 1580 310 1614 326
rect 1580 218 1614 234
rect 1386 108 1420 138
rect 2907 336 2941 398
rect 1833 308 1867 324
rect 1833 212 1867 228
rect 1929 308 1963 324
rect 1929 212 1963 228
rect 2025 308 2059 324
rect 2025 212 2059 228
rect 2121 308 2155 324
rect 2121 212 2155 228
rect 2217 308 2251 324
rect 2217 212 2251 228
rect 2313 308 2347 324
rect 2313 212 2347 228
rect 2409 308 2443 324
rect 2409 212 2443 228
rect 2505 308 2539 324
rect 2505 212 2539 228
rect 2601 308 2635 324
rect 2601 212 2635 228
rect 2697 308 2731 324
rect 2697 212 2731 228
rect 2793 308 2827 324
rect 2793 212 2827 228
rect 1719 108 1753 138
rect 1817 169 2843 177
rect 1817 135 1833 169
rect 1867 135 2025 169
rect 2059 135 2217 169
rect 2251 135 2409 169
rect 2443 135 2601 169
rect 2635 135 2793 169
rect 2827 135 2843 169
rect 1817 127 2843 135
rect 1386 76 1753 108
rect 2907 76 2941 138
rect 198 42 294 76
rect 1324 42 1815 76
rect 2845 42 2941 76
rect 1368 40 1766 42
<< viali >>
rect 312 946 346 980
rect 1272 946 1306 980
rect 312 638 346 886
rect 408 638 442 886
rect 504 638 538 886
rect 600 638 634 886
rect 696 638 730 886
rect 792 638 826 886
rect 888 638 922 886
rect 984 638 1018 886
rect 1080 638 1114 886
rect 1176 638 1210 886
rect 1272 638 1306 886
rect 1833 946 1867 980
rect 2793 946 2827 980
rect 1833 638 1867 886
rect 1929 638 1963 886
rect 2025 638 2059 886
rect 2121 638 2155 886
rect 2217 638 2251 886
rect 2313 638 2347 886
rect 2409 638 2443 886
rect 2505 638 2539 886
rect 2601 638 2635 886
rect 2697 638 2731 886
rect 2793 638 2827 886
rect 1536 360 1570 394
rect 312 228 346 308
rect 408 228 442 308
rect 504 228 538 308
rect 600 228 634 308
rect 696 228 730 308
rect 792 228 826 308
rect 888 228 922 308
rect 984 228 1018 308
rect 1080 228 1114 308
rect 1176 228 1210 308
rect 1272 228 1306 308
rect 1386 223 1420 323
rect 312 135 346 169
rect 1272 135 1306 169
rect 1492 234 1526 310
rect 1580 234 1614 310
rect 1833 228 1867 308
rect 1929 228 1963 308
rect 2025 228 2059 308
rect 2121 228 2155 308
rect 2217 228 2251 308
rect 2313 228 2347 308
rect 2409 228 2443 308
rect 2505 228 2539 308
rect 2601 228 2635 308
rect 2697 228 2731 308
rect 2793 228 2827 308
rect 1833 135 1867 169
rect 2793 135 2827 169
<< metal1 >>
rect 162 1048 1210 1082
rect 162 493 196 1048
rect 293 937 303 989
rect 355 937 365 989
rect 408 898 442 1048
rect 600 898 634 1048
rect 792 898 826 1048
rect 984 898 1018 1048
rect 1176 898 1210 1048
rect 1683 1048 2731 1082
rect 1252 938 1262 990
rect 1314 938 1324 990
rect 306 886 352 898
rect 306 638 312 886
rect 346 638 352 886
rect 306 626 352 638
rect 402 886 448 898
rect 402 638 408 886
rect 442 638 448 886
rect 402 626 448 638
rect 498 886 544 898
rect 498 638 504 886
rect 538 638 544 886
rect 498 626 544 638
rect 594 886 640 898
rect 594 638 600 886
rect 634 638 640 886
rect 594 626 640 638
rect 690 886 736 898
rect 690 638 696 886
rect 730 638 736 886
rect 690 626 736 638
rect 786 886 832 898
rect 786 638 792 886
rect 826 638 832 886
rect 786 626 832 638
rect 882 886 928 898
rect 882 638 888 886
rect 922 638 928 886
rect 882 626 928 638
rect 978 886 1024 898
rect 978 638 984 886
rect 1018 638 1024 886
rect 978 626 1024 638
rect 1074 886 1120 898
rect 1074 638 1080 886
rect 1114 638 1120 886
rect 1074 626 1120 638
rect 1170 886 1216 898
rect 1170 638 1176 886
rect 1210 638 1216 886
rect 1170 626 1216 638
rect 1266 886 1312 898
rect 1266 638 1272 886
rect 1306 638 1312 886
rect 1266 626 1312 638
rect 92 441 196 493
rect 162 74 196 441
rect 312 485 346 626
rect 504 485 538 626
rect 696 485 730 626
rect 888 485 922 626
rect 1080 485 1114 626
rect 1272 485 1306 626
rect 1683 485 1717 1048
rect 1813 938 1823 990
rect 1875 938 1885 990
rect 1929 898 1963 1048
rect 2121 898 2155 1048
rect 2313 898 2347 1048
rect 2505 898 2539 1048
rect 2697 898 2731 1048
rect 2773 938 2783 990
rect 2835 938 2845 990
rect 1827 886 1873 898
rect 1827 638 1833 886
rect 1867 638 1873 886
rect 1827 626 1873 638
rect 1923 886 1969 898
rect 1923 638 1929 886
rect 1963 638 1969 886
rect 1923 626 1969 638
rect 2019 886 2065 898
rect 2019 638 2025 886
rect 2059 638 2065 886
rect 2019 626 2065 638
rect 2115 886 2161 898
rect 2115 638 2121 886
rect 2155 638 2161 886
rect 2115 626 2161 638
rect 2211 886 2257 898
rect 2211 638 2217 886
rect 2251 638 2257 886
rect 2211 626 2257 638
rect 2307 886 2353 898
rect 2307 638 2313 886
rect 2347 638 2353 886
rect 2307 626 2353 638
rect 2403 886 2449 898
rect 2403 638 2409 886
rect 2443 638 2449 886
rect 2403 626 2449 638
rect 2499 886 2545 898
rect 2499 638 2505 886
rect 2539 638 2545 886
rect 2499 626 2545 638
rect 2595 886 2641 898
rect 2595 638 2601 886
rect 2635 638 2641 886
rect 2595 626 2641 638
rect 2691 886 2737 898
rect 2691 638 2697 886
rect 2731 638 2737 886
rect 2691 626 2737 638
rect 2787 886 2833 898
rect 2787 638 2793 886
rect 2827 638 2833 886
rect 2787 626 2833 638
rect 312 451 1717 485
rect 312 320 346 451
rect 504 320 538 451
rect 696 320 730 451
rect 888 320 922 451
rect 1080 320 1114 451
rect 1272 320 1306 451
rect 1517 361 1527 413
rect 1579 361 1589 413
rect 1524 360 1536 361
rect 1570 360 1582 361
rect 1524 354 1582 360
rect 1380 323 1426 335
rect 1683 323 1717 451
rect 306 308 352 320
rect 306 228 312 308
rect 346 228 352 308
rect 306 216 352 228
rect 402 308 448 320
rect 402 228 408 308
rect 442 228 448 308
rect 402 216 448 228
rect 498 308 544 320
rect 498 228 504 308
rect 538 228 544 308
rect 498 216 544 228
rect 594 308 640 320
rect 594 228 600 308
rect 634 228 640 308
rect 594 216 640 228
rect 690 308 736 320
rect 690 228 696 308
rect 730 228 736 308
rect 690 216 736 228
rect 786 308 832 320
rect 786 228 792 308
rect 826 228 832 308
rect 786 216 832 228
rect 882 308 928 320
rect 882 228 888 308
rect 922 228 928 308
rect 882 216 928 228
rect 978 308 1024 320
rect 978 228 984 308
rect 1018 228 1024 308
rect 978 216 1024 228
rect 1074 308 1120 320
rect 1074 228 1080 308
rect 1114 228 1120 308
rect 1074 216 1120 228
rect 1170 308 1216 320
rect 1170 228 1176 308
rect 1210 228 1216 308
rect 1170 216 1216 228
rect 1266 308 1312 320
rect 1266 228 1272 308
rect 1306 228 1312 308
rect 1266 216 1312 228
rect 1380 223 1386 323
rect 1420 322 1526 323
rect 1580 322 1717 323
rect 1420 310 1532 322
rect 1420 234 1492 310
rect 1526 234 1532 310
rect 1420 223 1532 234
rect 292 124 302 176
rect 354 124 364 176
rect 408 74 442 216
rect 600 74 634 216
rect 792 74 826 216
rect 984 74 1018 216
rect 1176 74 1210 216
rect 1380 211 1426 223
rect 1486 222 1532 223
rect 1574 310 1717 322
rect 1833 485 1867 626
rect 2025 485 2059 626
rect 2217 485 2251 626
rect 2409 485 2443 626
rect 2601 485 2635 626
rect 2793 485 2827 626
rect 1833 451 2942 485
rect 1833 320 1867 451
rect 2025 320 2059 451
rect 2217 320 2251 451
rect 2409 320 2443 451
rect 2601 320 2635 451
rect 2793 320 2827 451
rect 1574 234 1580 310
rect 1614 234 1717 310
rect 1574 223 1717 234
rect 1574 222 1620 223
rect 1254 126 1264 178
rect 1316 126 1326 178
rect 162 40 1210 74
rect 1683 74 1717 223
rect 1827 308 1873 320
rect 1827 228 1833 308
rect 1867 228 1873 308
rect 1827 216 1873 228
rect 1923 308 1969 320
rect 1923 228 1929 308
rect 1963 228 1969 308
rect 1923 216 1969 228
rect 2019 308 2065 320
rect 2019 228 2025 308
rect 2059 228 2065 308
rect 2019 216 2065 228
rect 2115 308 2161 320
rect 2115 228 2121 308
rect 2155 228 2161 308
rect 2115 216 2161 228
rect 2211 308 2257 320
rect 2211 228 2217 308
rect 2251 228 2257 308
rect 2211 216 2257 228
rect 2307 308 2353 320
rect 2307 228 2313 308
rect 2347 228 2353 308
rect 2307 216 2353 228
rect 2403 308 2449 320
rect 2403 228 2409 308
rect 2443 228 2449 308
rect 2403 216 2449 228
rect 2499 308 2545 320
rect 2499 228 2505 308
rect 2539 228 2545 308
rect 2499 216 2545 228
rect 2595 308 2641 320
rect 2595 228 2601 308
rect 2635 228 2641 308
rect 2595 216 2641 228
rect 2691 308 2737 320
rect 2691 228 2697 308
rect 2731 228 2737 308
rect 2691 216 2737 228
rect 2787 308 2833 320
rect 2787 228 2793 308
rect 2827 228 2833 308
rect 2787 216 2833 228
rect 1815 126 1825 178
rect 1877 126 1887 178
rect 1929 74 1963 216
rect 2121 74 2155 216
rect 2313 74 2347 216
rect 2505 74 2539 216
rect 2697 74 2731 216
rect 2775 126 2785 178
rect 2837 126 2847 178
rect 1683 40 2731 74
<< via1 >>
rect 303 980 355 989
rect 303 946 312 980
rect 312 946 346 980
rect 346 946 355 980
rect 303 937 355 946
rect 1262 980 1314 990
rect 1262 946 1272 980
rect 1272 946 1306 980
rect 1306 946 1314 980
rect 1262 938 1314 946
rect 1823 980 1875 990
rect 1823 946 1833 980
rect 1833 946 1867 980
rect 1867 946 1875 980
rect 1823 938 1875 946
rect 2783 980 2835 990
rect 2783 946 2793 980
rect 2793 946 2827 980
rect 2827 946 2835 980
rect 2783 938 2835 946
rect 1527 394 1579 413
rect 1527 361 1536 394
rect 1536 361 1570 394
rect 1570 361 1579 394
rect 302 169 354 176
rect 302 135 312 169
rect 312 135 346 169
rect 346 135 354 169
rect 302 124 354 135
rect 1264 169 1316 178
rect 1264 135 1272 169
rect 1272 135 1306 169
rect 1306 135 1316 169
rect 1264 126 1316 135
rect 1825 169 1877 178
rect 1825 135 1833 169
rect 1833 135 1867 169
rect 1867 135 1877 169
rect 1825 126 1877 135
rect 2785 169 2837 178
rect 2785 135 2793 169
rect 2793 135 2827 169
rect 2827 135 2837 169
rect 2785 126 2837 135
<< metal2 >>
rect 303 990 355 999
rect 1262 990 1314 1000
rect 1823 990 1875 1000
rect 2783 990 2835 1000
rect 101 989 1262 990
rect 101 938 303 989
rect 355 938 1262 989
rect 1314 938 1823 990
rect 1875 938 2783 990
rect 2835 938 2849 990
rect 303 927 355 937
rect 1262 928 1314 938
rect 1527 413 1579 938
rect 1823 928 1875 938
rect 2783 928 2835 938
rect 1527 351 1579 361
rect 302 183 354 186
rect 394 183 460 185
rect 1264 183 1316 188
rect 1825 183 1877 188
rect 2785 183 2837 188
rect 92 178 2837 183
rect 92 176 1264 178
rect 92 131 302 176
rect 354 131 1264 176
rect 302 114 354 124
rect 394 119 460 131
rect 1316 131 1825 178
rect 1264 116 1316 126
rect 1877 131 2785 178
rect 1825 116 1877 126
rect 2785 116 2837 126
<< labels >>
flabel locali 1553 1056 1553 1056 1 FreeSans 400 0 0 0 VDD
port 5 n power bidirectional
flabel locali 1553 66 1553 66 1 FreeSans 400 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 114 469 114 469 1 FreeSans 400 0 0 0 in
port 1 n
flabel metal2 120 965 120 965 1 FreeSans 400 0 0 0 en_b
port 4 n
flabel metal2 114 158 114 158 1 FreeSans 400 0 0 0 en
port 3 n
flabel metal1 2927 465 2927 465 1 FreeSans 400 0 0 0 out
port 2 n
<< end >>
