magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< nwell >>
rect -7664 -7309 3823 -1120
<< pwell >>
rect -7631 -7647 13745 -7495
rect -7631 -17433 -7479 -7647
rect 13593 -17433 13745 -7647
rect -7631 -17585 -7297 -17433
rect 13358 -17585 13745 -17433
<< psubdiff >>
rect -7605 -7554 13719 -7521
rect -7605 -7588 -7264 -7554
rect -7230 -7588 -7196 -7554
rect -7162 -7588 -7128 -7554
rect -7094 -7588 -7060 -7554
rect -7026 -7588 -6992 -7554
rect -6958 -7588 -6924 -7554
rect -6890 -7588 -6856 -7554
rect -6822 -7588 -6788 -7554
rect -6754 -7588 -6720 -7554
rect -6686 -7588 -6652 -7554
rect -6618 -7588 -6584 -7554
rect -6550 -7588 -6516 -7554
rect -6482 -7588 -6448 -7554
rect -6414 -7588 -6380 -7554
rect -6346 -7588 -6312 -7554
rect -6278 -7588 -6244 -7554
rect -6210 -7588 -6176 -7554
rect -6142 -7588 -6108 -7554
rect -6074 -7588 -6040 -7554
rect -6006 -7588 -5972 -7554
rect -5938 -7588 -5904 -7554
rect -5870 -7588 -5836 -7554
rect -5802 -7588 -5768 -7554
rect -5734 -7588 -5700 -7554
rect -5666 -7588 -5632 -7554
rect -5598 -7588 -5564 -7554
rect -5530 -7588 -5496 -7554
rect -5462 -7588 -5428 -7554
rect -5394 -7588 -5360 -7554
rect -5326 -7588 -5292 -7554
rect -5258 -7588 -5224 -7554
rect -5190 -7588 -5156 -7554
rect -5122 -7588 -5088 -7554
rect -5054 -7588 -5020 -7554
rect -4986 -7588 -4952 -7554
rect -4918 -7588 -4884 -7554
rect -4850 -7588 -4816 -7554
rect -4782 -7588 -4748 -7554
rect -4714 -7588 -4680 -7554
rect -4646 -7588 -4612 -7554
rect -4578 -7588 -4544 -7554
rect -4510 -7588 -4476 -7554
rect -4442 -7588 -4408 -7554
rect -4374 -7588 -4340 -7554
rect -4306 -7588 -4272 -7554
rect -4238 -7588 -4204 -7554
rect -4170 -7588 -4136 -7554
rect -4102 -7588 -4068 -7554
rect -4034 -7588 -4000 -7554
rect -3966 -7588 -3932 -7554
rect -3898 -7588 -3864 -7554
rect -3830 -7588 -3796 -7554
rect -3762 -7588 -3728 -7554
rect -3694 -7588 -3660 -7554
rect -3626 -7588 -3592 -7554
rect -3558 -7588 -3524 -7554
rect -3490 -7588 -3456 -7554
rect -3422 -7588 -3388 -7554
rect -3354 -7588 -3320 -7554
rect -3286 -7588 -3252 -7554
rect -3218 -7588 -3184 -7554
rect -3150 -7588 -3116 -7554
rect -3082 -7588 -3048 -7554
rect -3014 -7588 -2980 -7554
rect -2946 -7588 -2912 -7554
rect -2878 -7588 -2844 -7554
rect -2810 -7588 -2776 -7554
rect -2742 -7588 -2708 -7554
rect -2674 -7588 -2640 -7554
rect -2606 -7588 -2572 -7554
rect -2538 -7588 -2504 -7554
rect -2470 -7588 -2436 -7554
rect -2402 -7588 -2368 -7554
rect -2334 -7588 -2300 -7554
rect -2266 -7588 -2232 -7554
rect -2198 -7588 -2164 -7554
rect -2130 -7588 -2096 -7554
rect -2062 -7588 -2028 -7554
rect -1994 -7588 -1960 -7554
rect -1926 -7588 -1892 -7554
rect -1858 -7588 -1824 -7554
rect -1790 -7588 -1756 -7554
rect -1722 -7588 -1688 -7554
rect -1654 -7588 -1620 -7554
rect -1586 -7588 -1552 -7554
rect -1518 -7588 -1484 -7554
rect -1450 -7588 -1416 -7554
rect -1382 -7588 -1348 -7554
rect -1314 -7588 -1280 -7554
rect -1246 -7588 -1212 -7554
rect -1178 -7588 -1144 -7554
rect -1110 -7588 -1076 -7554
rect -1042 -7588 -1008 -7554
rect -974 -7588 -940 -7554
rect -906 -7588 -872 -7554
rect -838 -7588 -804 -7554
rect -770 -7588 -736 -7554
rect -702 -7588 -668 -7554
rect -634 -7588 -600 -7554
rect -566 -7588 -532 -7554
rect -498 -7588 -464 -7554
rect -430 -7588 -396 -7554
rect -362 -7588 -328 -7554
rect -294 -7588 -260 -7554
rect -226 -7588 -192 -7554
rect -158 -7588 -124 -7554
rect -90 -7588 -56 -7554
rect -22 -7588 12 -7554
rect 46 -7588 80 -7554
rect 114 -7588 148 -7554
rect 182 -7588 216 -7554
rect 250 -7588 284 -7554
rect 318 -7588 352 -7554
rect 386 -7588 420 -7554
rect 454 -7588 488 -7554
rect 522 -7588 556 -7554
rect 590 -7588 624 -7554
rect 658 -7588 692 -7554
rect 726 -7588 760 -7554
rect 794 -7588 828 -7554
rect 862 -7588 896 -7554
rect 930 -7588 964 -7554
rect 998 -7588 1032 -7554
rect 1066 -7588 1100 -7554
rect 1134 -7588 1168 -7554
rect 1202 -7588 1236 -7554
rect 1270 -7588 1304 -7554
rect 1338 -7588 1372 -7554
rect 1406 -7588 1440 -7554
rect 1474 -7588 1508 -7554
rect 1542 -7588 1576 -7554
rect 1610 -7588 1644 -7554
rect 1678 -7588 1712 -7554
rect 1746 -7588 1780 -7554
rect 1814 -7588 1848 -7554
rect 1882 -7588 1916 -7554
rect 1950 -7588 1984 -7554
rect 2018 -7588 2052 -7554
rect 2086 -7588 2120 -7554
rect 2154 -7588 2188 -7554
rect 2222 -7588 2256 -7554
rect 2290 -7588 2324 -7554
rect 2358 -7588 2392 -7554
rect 2426 -7588 2460 -7554
rect 2494 -7588 2528 -7554
rect 2562 -7588 2596 -7554
rect 2630 -7588 2664 -7554
rect 2698 -7588 2732 -7554
rect 2766 -7588 2800 -7554
rect 2834 -7588 2868 -7554
rect 2902 -7588 2936 -7554
rect 2970 -7588 3004 -7554
rect 3038 -7588 3072 -7554
rect 3106 -7588 3140 -7554
rect 3174 -7588 3208 -7554
rect 3242 -7588 3276 -7554
rect 3310 -7588 3344 -7554
rect 3378 -7588 3412 -7554
rect 3446 -7588 3480 -7554
rect 3514 -7588 3548 -7554
rect 3582 -7588 3616 -7554
rect 3650 -7588 3684 -7554
rect 3718 -7588 3752 -7554
rect 3786 -7588 3820 -7554
rect 3854 -7588 3888 -7554
rect 3922 -7588 3956 -7554
rect 3990 -7588 4024 -7554
rect 4058 -7588 4092 -7554
rect 4126 -7588 4160 -7554
rect 4194 -7588 4228 -7554
rect 4262 -7588 4296 -7554
rect 4330 -7588 4364 -7554
rect 4398 -7588 4432 -7554
rect 4466 -7588 4500 -7554
rect 4534 -7588 4568 -7554
rect 4602 -7588 4636 -7554
rect 4670 -7588 4704 -7554
rect 4738 -7588 4772 -7554
rect 4806 -7588 4840 -7554
rect 4874 -7588 4908 -7554
rect 4942 -7588 4976 -7554
rect 5010 -7588 5044 -7554
rect 5078 -7588 5112 -7554
rect 5146 -7588 5180 -7554
rect 5214 -7588 5248 -7554
rect 5282 -7588 5316 -7554
rect 5350 -7588 5384 -7554
rect 5418 -7588 5452 -7554
rect 5486 -7588 5520 -7554
rect 5554 -7588 5588 -7554
rect 5622 -7588 5656 -7554
rect 5690 -7588 5724 -7554
rect 5758 -7588 5792 -7554
rect 5826 -7588 5860 -7554
rect 5894 -7588 5928 -7554
rect 5962 -7588 5996 -7554
rect 6030 -7588 6064 -7554
rect 6098 -7588 6132 -7554
rect 6166 -7588 6200 -7554
rect 6234 -7588 6268 -7554
rect 6302 -7588 6336 -7554
rect 6370 -7588 6404 -7554
rect 6438 -7588 6472 -7554
rect 6506 -7588 6540 -7554
rect 6574 -7588 6608 -7554
rect 6642 -7588 6676 -7554
rect 6710 -7588 6744 -7554
rect 6778 -7588 6812 -7554
rect 6846 -7588 6880 -7554
rect 6914 -7588 6948 -7554
rect 6982 -7588 7016 -7554
rect 7050 -7588 7084 -7554
rect 7118 -7588 7152 -7554
rect 7186 -7588 7220 -7554
rect 7254 -7588 7288 -7554
rect 7322 -7588 7356 -7554
rect 7390 -7588 7424 -7554
rect 7458 -7588 7492 -7554
rect 7526 -7588 7560 -7554
rect 7594 -7588 7628 -7554
rect 7662 -7588 7696 -7554
rect 7730 -7588 7764 -7554
rect 7798 -7588 7832 -7554
rect 7866 -7588 7900 -7554
rect 7934 -7588 7968 -7554
rect 8002 -7588 8036 -7554
rect 8070 -7588 8104 -7554
rect 8138 -7588 8172 -7554
rect 8206 -7588 8240 -7554
rect 8274 -7588 8308 -7554
rect 8342 -7588 8376 -7554
rect 8410 -7588 8444 -7554
rect 8478 -7588 8512 -7554
rect 8546 -7588 8580 -7554
rect 8614 -7588 8648 -7554
rect 8682 -7588 8716 -7554
rect 8750 -7588 8784 -7554
rect 8818 -7588 8852 -7554
rect 8886 -7588 8920 -7554
rect 8954 -7588 8988 -7554
rect 9022 -7588 9056 -7554
rect 9090 -7588 9124 -7554
rect 9158 -7588 9192 -7554
rect 9226 -7588 9260 -7554
rect 9294 -7588 9328 -7554
rect 9362 -7588 9396 -7554
rect 9430 -7588 9464 -7554
rect 9498 -7588 9532 -7554
rect 9566 -7588 9600 -7554
rect 9634 -7588 9668 -7554
rect 9702 -7588 9736 -7554
rect 9770 -7588 9804 -7554
rect 9838 -7588 9872 -7554
rect 9906 -7588 9940 -7554
rect 9974 -7588 10008 -7554
rect 10042 -7588 10076 -7554
rect 10110 -7588 10144 -7554
rect 10178 -7588 10212 -7554
rect 10246 -7588 10280 -7554
rect 10314 -7588 10348 -7554
rect 10382 -7588 10416 -7554
rect 10450 -7588 10484 -7554
rect 10518 -7588 10552 -7554
rect 10586 -7588 10620 -7554
rect 10654 -7588 10688 -7554
rect 10722 -7588 10756 -7554
rect 10790 -7588 10824 -7554
rect 10858 -7588 10892 -7554
rect 10926 -7588 10960 -7554
rect 10994 -7588 11028 -7554
rect 11062 -7588 11096 -7554
rect 11130 -7588 11164 -7554
rect 11198 -7588 11232 -7554
rect 11266 -7588 11300 -7554
rect 11334 -7588 11368 -7554
rect 11402 -7588 11436 -7554
rect 11470 -7588 11504 -7554
rect 11538 -7588 11572 -7554
rect 11606 -7588 11640 -7554
rect 11674 -7588 11708 -7554
rect 11742 -7588 11776 -7554
rect 11810 -7588 11844 -7554
rect 11878 -7588 11912 -7554
rect 11946 -7588 11980 -7554
rect 12014 -7588 12048 -7554
rect 12082 -7588 12116 -7554
rect 12150 -7588 12184 -7554
rect 12218 -7588 12252 -7554
rect 12286 -7588 12320 -7554
rect 12354 -7588 12388 -7554
rect 12422 -7588 12456 -7554
rect 12490 -7588 12524 -7554
rect 12558 -7588 12592 -7554
rect 12626 -7588 12660 -7554
rect 12694 -7588 12728 -7554
rect 12762 -7588 12796 -7554
rect 12830 -7588 12864 -7554
rect 12898 -7588 12932 -7554
rect 12966 -7588 13000 -7554
rect 13034 -7588 13068 -7554
rect 13102 -7588 13136 -7554
rect 13170 -7588 13204 -7554
rect 13238 -7588 13272 -7554
rect 13306 -7588 13340 -7554
rect 13374 -7588 13408 -7554
rect 13442 -7588 13719 -7554
rect -7605 -7621 13719 -7588
rect -7605 -7850 -7505 -7621
rect -7605 -7884 -7572 -7850
rect -7538 -7884 -7505 -7850
rect -7605 -7918 -7505 -7884
rect -7605 -7952 -7572 -7918
rect -7538 -7952 -7505 -7918
rect -7605 -7986 -7505 -7952
rect -7605 -8020 -7572 -7986
rect -7538 -8020 -7505 -7986
rect -7605 -8054 -7505 -8020
rect -7605 -8088 -7572 -8054
rect -7538 -8088 -7505 -8054
rect -7605 -8122 -7505 -8088
rect -7605 -8156 -7572 -8122
rect -7538 -8156 -7505 -8122
rect -7605 -8190 -7505 -8156
rect -7605 -8224 -7572 -8190
rect -7538 -8224 -7505 -8190
rect -7605 -8258 -7505 -8224
rect -7605 -8292 -7572 -8258
rect -7538 -8292 -7505 -8258
rect -7605 -8326 -7505 -8292
rect -7605 -8360 -7572 -8326
rect -7538 -8360 -7505 -8326
rect -7605 -8394 -7505 -8360
rect -7605 -8428 -7572 -8394
rect -7538 -8428 -7505 -8394
rect -7605 -8462 -7505 -8428
rect -7605 -8496 -7572 -8462
rect -7538 -8496 -7505 -8462
rect -7605 -8530 -7505 -8496
rect -7605 -8564 -7572 -8530
rect -7538 -8564 -7505 -8530
rect -7605 -8598 -7505 -8564
rect -7605 -8632 -7572 -8598
rect -7538 -8632 -7505 -8598
rect -7605 -8666 -7505 -8632
rect -7605 -8700 -7572 -8666
rect -7538 -8700 -7505 -8666
rect -7605 -8734 -7505 -8700
rect -7605 -8768 -7572 -8734
rect -7538 -8768 -7505 -8734
rect -7605 -8802 -7505 -8768
rect -7605 -8836 -7572 -8802
rect -7538 -8836 -7505 -8802
rect -7605 -8870 -7505 -8836
rect -7605 -8904 -7572 -8870
rect -7538 -8904 -7505 -8870
rect -7605 -8938 -7505 -8904
rect -7605 -8972 -7572 -8938
rect -7538 -8972 -7505 -8938
rect -7605 -9006 -7505 -8972
rect -7605 -9040 -7572 -9006
rect -7538 -9040 -7505 -9006
rect -7605 -9074 -7505 -9040
rect -7605 -9108 -7572 -9074
rect -7538 -9108 -7505 -9074
rect -7605 -9142 -7505 -9108
rect -7605 -9176 -7572 -9142
rect -7538 -9176 -7505 -9142
rect -7605 -9210 -7505 -9176
rect -7605 -9244 -7572 -9210
rect -7538 -9244 -7505 -9210
rect -7605 -9278 -7505 -9244
rect -7605 -9312 -7572 -9278
rect -7538 -9312 -7505 -9278
rect -7605 -9346 -7505 -9312
rect -7605 -9380 -7572 -9346
rect -7538 -9380 -7505 -9346
rect -7605 -9414 -7505 -9380
rect -7605 -9448 -7572 -9414
rect -7538 -9448 -7505 -9414
rect -7605 -9482 -7505 -9448
rect -7605 -9516 -7572 -9482
rect -7538 -9516 -7505 -9482
rect -7605 -9550 -7505 -9516
rect -7605 -9584 -7572 -9550
rect -7538 -9584 -7505 -9550
rect -7605 -9618 -7505 -9584
rect -7605 -9652 -7572 -9618
rect -7538 -9652 -7505 -9618
rect -7605 -9686 -7505 -9652
rect -7605 -9720 -7572 -9686
rect -7538 -9720 -7505 -9686
rect -7605 -9754 -7505 -9720
rect -7605 -9788 -7572 -9754
rect -7538 -9788 -7505 -9754
rect -7605 -9822 -7505 -9788
rect -7605 -9856 -7572 -9822
rect -7538 -9856 -7505 -9822
rect -7605 -9890 -7505 -9856
rect -7605 -9924 -7572 -9890
rect -7538 -9924 -7505 -9890
rect -7605 -9958 -7505 -9924
rect -7605 -9992 -7572 -9958
rect -7538 -9992 -7505 -9958
rect -7605 -10026 -7505 -9992
rect -7605 -10060 -7572 -10026
rect -7538 -10060 -7505 -10026
rect -7605 -10094 -7505 -10060
rect -7605 -10128 -7572 -10094
rect -7538 -10128 -7505 -10094
rect -7605 -10162 -7505 -10128
rect -7605 -10196 -7572 -10162
rect -7538 -10196 -7505 -10162
rect -7605 -10230 -7505 -10196
rect -7605 -10264 -7572 -10230
rect -7538 -10264 -7505 -10230
rect -7605 -10298 -7505 -10264
rect -7605 -10332 -7572 -10298
rect -7538 -10332 -7505 -10298
rect -7605 -10366 -7505 -10332
rect -7605 -10400 -7572 -10366
rect -7538 -10400 -7505 -10366
rect -7605 -10434 -7505 -10400
rect -7605 -10468 -7572 -10434
rect -7538 -10468 -7505 -10434
rect -7605 -10502 -7505 -10468
rect -7605 -10536 -7572 -10502
rect -7538 -10536 -7505 -10502
rect -7605 -10570 -7505 -10536
rect -7605 -10604 -7572 -10570
rect -7538 -10604 -7505 -10570
rect -7605 -10638 -7505 -10604
rect -7605 -10672 -7572 -10638
rect -7538 -10672 -7505 -10638
rect -7605 -10706 -7505 -10672
rect -7605 -10740 -7572 -10706
rect -7538 -10740 -7505 -10706
rect -7605 -10774 -7505 -10740
rect -7605 -10808 -7572 -10774
rect -7538 -10808 -7505 -10774
rect -7605 -10842 -7505 -10808
rect -7605 -10876 -7572 -10842
rect -7538 -10876 -7505 -10842
rect -7605 -10910 -7505 -10876
rect -7605 -10944 -7572 -10910
rect -7538 -10944 -7505 -10910
rect -7605 -10978 -7505 -10944
rect -7605 -11012 -7572 -10978
rect -7538 -11012 -7505 -10978
rect -7605 -11046 -7505 -11012
rect -7605 -11080 -7572 -11046
rect -7538 -11080 -7505 -11046
rect -7605 -11114 -7505 -11080
rect -7605 -11148 -7572 -11114
rect -7538 -11148 -7505 -11114
rect -7605 -11182 -7505 -11148
rect -7605 -11216 -7572 -11182
rect -7538 -11216 -7505 -11182
rect -7605 -11250 -7505 -11216
rect -7605 -11284 -7572 -11250
rect -7538 -11284 -7505 -11250
rect -7605 -11318 -7505 -11284
rect -7605 -11352 -7572 -11318
rect -7538 -11352 -7505 -11318
rect -7605 -11386 -7505 -11352
rect -7605 -11420 -7572 -11386
rect -7538 -11420 -7505 -11386
rect -7605 -11454 -7505 -11420
rect -7605 -11488 -7572 -11454
rect -7538 -11488 -7505 -11454
rect -7605 -11522 -7505 -11488
rect -7605 -11556 -7572 -11522
rect -7538 -11556 -7505 -11522
rect -7605 -11590 -7505 -11556
rect -7605 -11624 -7572 -11590
rect -7538 -11624 -7505 -11590
rect -7605 -11658 -7505 -11624
rect -7605 -11692 -7572 -11658
rect -7538 -11692 -7505 -11658
rect -7605 -11726 -7505 -11692
rect -7605 -11760 -7572 -11726
rect -7538 -11760 -7505 -11726
rect -7605 -11794 -7505 -11760
rect -7605 -11828 -7572 -11794
rect -7538 -11828 -7505 -11794
rect -7605 -11862 -7505 -11828
rect -7605 -11896 -7572 -11862
rect -7538 -11896 -7505 -11862
rect -7605 -11930 -7505 -11896
rect -7605 -11964 -7572 -11930
rect -7538 -11964 -7505 -11930
rect -7605 -11998 -7505 -11964
rect -7605 -12032 -7572 -11998
rect -7538 -12032 -7505 -11998
rect -7605 -12066 -7505 -12032
rect -7605 -12100 -7572 -12066
rect -7538 -12100 -7505 -12066
rect -7605 -12134 -7505 -12100
rect -7605 -12168 -7572 -12134
rect -7538 -12168 -7505 -12134
rect -7605 -12202 -7505 -12168
rect -7605 -12236 -7572 -12202
rect -7538 -12236 -7505 -12202
rect -7605 -12270 -7505 -12236
rect -7605 -12304 -7572 -12270
rect -7538 -12304 -7505 -12270
rect -7605 -12338 -7505 -12304
rect -7605 -12372 -7572 -12338
rect -7538 -12372 -7505 -12338
rect -7605 -12406 -7505 -12372
rect -7605 -12440 -7572 -12406
rect -7538 -12440 -7505 -12406
rect -7605 -12474 -7505 -12440
rect -7605 -12508 -7572 -12474
rect -7538 -12508 -7505 -12474
rect -7605 -12542 -7505 -12508
rect -7605 -12576 -7572 -12542
rect -7538 -12576 -7505 -12542
rect -7605 -12610 -7505 -12576
rect -7605 -12644 -7572 -12610
rect -7538 -12644 -7505 -12610
rect -7605 -12678 -7505 -12644
rect -7605 -12712 -7572 -12678
rect -7538 -12712 -7505 -12678
rect -7605 -12746 -7505 -12712
rect -7605 -12780 -7572 -12746
rect -7538 -12780 -7505 -12746
rect -7605 -12814 -7505 -12780
rect -7605 -12848 -7572 -12814
rect -7538 -12848 -7505 -12814
rect -7605 -12882 -7505 -12848
rect -7605 -12916 -7572 -12882
rect -7538 -12916 -7505 -12882
rect -7605 -12950 -7505 -12916
rect -7605 -12984 -7572 -12950
rect -7538 -12984 -7505 -12950
rect -7605 -13018 -7505 -12984
rect -7605 -13052 -7572 -13018
rect -7538 -13052 -7505 -13018
rect -7605 -13086 -7505 -13052
rect -7605 -13120 -7572 -13086
rect -7538 -13120 -7505 -13086
rect -7605 -13154 -7505 -13120
rect -7605 -13188 -7572 -13154
rect -7538 -13188 -7505 -13154
rect -7605 -13222 -7505 -13188
rect -7605 -13256 -7572 -13222
rect -7538 -13256 -7505 -13222
rect -7605 -13290 -7505 -13256
rect -7605 -13324 -7572 -13290
rect -7538 -13324 -7505 -13290
rect -7605 -13358 -7505 -13324
rect -7605 -13392 -7572 -13358
rect -7538 -13392 -7505 -13358
rect -7605 -13426 -7505 -13392
rect -7605 -13460 -7572 -13426
rect -7538 -13460 -7505 -13426
rect -7605 -13494 -7505 -13460
rect -7605 -13528 -7572 -13494
rect -7538 -13528 -7505 -13494
rect -7605 -13562 -7505 -13528
rect -7605 -13596 -7572 -13562
rect -7538 -13596 -7505 -13562
rect -7605 -13630 -7505 -13596
rect -7605 -13664 -7572 -13630
rect -7538 -13664 -7505 -13630
rect -7605 -13698 -7505 -13664
rect -7605 -13732 -7572 -13698
rect -7538 -13732 -7505 -13698
rect -7605 -13766 -7505 -13732
rect -7605 -13800 -7572 -13766
rect -7538 -13800 -7505 -13766
rect -7605 -13834 -7505 -13800
rect -7605 -13868 -7572 -13834
rect -7538 -13868 -7505 -13834
rect -7605 -13902 -7505 -13868
rect -7605 -13936 -7572 -13902
rect -7538 -13936 -7505 -13902
rect -7605 -13970 -7505 -13936
rect -7605 -14004 -7572 -13970
rect -7538 -14004 -7505 -13970
rect -7605 -14038 -7505 -14004
rect -7605 -14072 -7572 -14038
rect -7538 -14072 -7505 -14038
rect -7605 -14106 -7505 -14072
rect -7605 -14140 -7572 -14106
rect -7538 -14140 -7505 -14106
rect -7605 -14174 -7505 -14140
rect -7605 -14208 -7572 -14174
rect -7538 -14208 -7505 -14174
rect -7605 -14242 -7505 -14208
rect -7605 -14276 -7572 -14242
rect -7538 -14276 -7505 -14242
rect -7605 -14310 -7505 -14276
rect -7605 -14344 -7572 -14310
rect -7538 -14344 -7505 -14310
rect -7605 -14378 -7505 -14344
rect -7605 -14412 -7572 -14378
rect -7538 -14412 -7505 -14378
rect -7605 -14446 -7505 -14412
rect -7605 -14480 -7572 -14446
rect -7538 -14480 -7505 -14446
rect -7605 -14514 -7505 -14480
rect -7605 -14548 -7572 -14514
rect -7538 -14548 -7505 -14514
rect -7605 -14582 -7505 -14548
rect -7605 -14616 -7572 -14582
rect -7538 -14616 -7505 -14582
rect -7605 -14650 -7505 -14616
rect -7605 -14684 -7572 -14650
rect -7538 -14684 -7505 -14650
rect -7605 -14718 -7505 -14684
rect -7605 -14752 -7572 -14718
rect -7538 -14752 -7505 -14718
rect -7605 -14786 -7505 -14752
rect -7605 -14820 -7572 -14786
rect -7538 -14820 -7505 -14786
rect -7605 -14854 -7505 -14820
rect -7605 -14888 -7572 -14854
rect -7538 -14888 -7505 -14854
rect -7605 -14922 -7505 -14888
rect -7605 -14956 -7572 -14922
rect -7538 -14956 -7505 -14922
rect -7605 -14990 -7505 -14956
rect -7605 -15024 -7572 -14990
rect -7538 -15024 -7505 -14990
rect -7605 -15058 -7505 -15024
rect -7605 -15092 -7572 -15058
rect -7538 -15092 -7505 -15058
rect -7605 -15126 -7505 -15092
rect -7605 -15160 -7572 -15126
rect -7538 -15160 -7505 -15126
rect -7605 -15194 -7505 -15160
rect -7605 -15228 -7572 -15194
rect -7538 -15228 -7505 -15194
rect -7605 -15262 -7505 -15228
rect -7605 -15296 -7572 -15262
rect -7538 -15296 -7505 -15262
rect -7605 -15330 -7505 -15296
rect -7605 -15364 -7572 -15330
rect -7538 -15364 -7505 -15330
rect -7605 -15398 -7505 -15364
rect -7605 -15432 -7572 -15398
rect -7538 -15432 -7505 -15398
rect -7605 -15466 -7505 -15432
rect -7605 -15500 -7572 -15466
rect -7538 -15500 -7505 -15466
rect -7605 -15534 -7505 -15500
rect -7605 -15568 -7572 -15534
rect -7538 -15568 -7505 -15534
rect -7605 -15602 -7505 -15568
rect -7605 -15636 -7572 -15602
rect -7538 -15636 -7505 -15602
rect -7605 -15670 -7505 -15636
rect -7605 -15704 -7572 -15670
rect -7538 -15704 -7505 -15670
rect -7605 -15738 -7505 -15704
rect -7605 -15772 -7572 -15738
rect -7538 -15772 -7505 -15738
rect -7605 -15806 -7505 -15772
rect -7605 -15840 -7572 -15806
rect -7538 -15840 -7505 -15806
rect -7605 -15874 -7505 -15840
rect -7605 -15908 -7572 -15874
rect -7538 -15908 -7505 -15874
rect -7605 -15942 -7505 -15908
rect -7605 -15976 -7572 -15942
rect -7538 -15976 -7505 -15942
rect -7605 -16010 -7505 -15976
rect -7605 -16044 -7572 -16010
rect -7538 -16044 -7505 -16010
rect -7605 -16078 -7505 -16044
rect -7605 -16112 -7572 -16078
rect -7538 -16112 -7505 -16078
rect -7605 -16146 -7505 -16112
rect -7605 -16180 -7572 -16146
rect -7538 -16180 -7505 -16146
rect -7605 -16214 -7505 -16180
rect -7605 -16248 -7572 -16214
rect -7538 -16248 -7505 -16214
rect -7605 -16282 -7505 -16248
rect -7605 -16316 -7572 -16282
rect -7538 -16316 -7505 -16282
rect -7605 -16350 -7505 -16316
rect -7605 -16384 -7572 -16350
rect -7538 -16384 -7505 -16350
rect -7605 -16418 -7505 -16384
rect -7605 -16452 -7572 -16418
rect -7538 -16452 -7505 -16418
rect -7605 -16486 -7505 -16452
rect -7605 -16520 -7572 -16486
rect -7538 -16520 -7505 -16486
rect -7605 -16554 -7505 -16520
rect -7605 -16588 -7572 -16554
rect -7538 -16588 -7505 -16554
rect -7605 -16622 -7505 -16588
rect -7605 -16656 -7572 -16622
rect -7538 -16656 -7505 -16622
rect -7605 -16690 -7505 -16656
rect -7605 -16724 -7572 -16690
rect -7538 -16724 -7505 -16690
rect -7605 -16758 -7505 -16724
rect -7605 -16792 -7572 -16758
rect -7538 -16792 -7505 -16758
rect -7605 -16826 -7505 -16792
rect -7605 -16860 -7572 -16826
rect -7538 -16860 -7505 -16826
rect -7605 -16894 -7505 -16860
rect -7605 -16928 -7572 -16894
rect -7538 -16928 -7505 -16894
rect -7605 -16962 -7505 -16928
rect -7605 -16996 -7572 -16962
rect -7538 -16996 -7505 -16962
rect -7605 -17030 -7505 -16996
rect -7605 -17064 -7572 -17030
rect -7538 -17064 -7505 -17030
rect -7605 -17098 -7505 -17064
rect -7605 -17132 -7572 -17098
rect -7538 -17132 -7505 -17098
rect -7605 -17166 -7505 -17132
rect -7605 -17200 -7572 -17166
rect -7538 -17200 -7505 -17166
rect -7605 -17234 -7505 -17200
rect -7605 -17268 -7572 -17234
rect -7538 -17268 -7505 -17234
rect -7605 -17459 -7505 -17268
rect 13619 -7731 13719 -7621
rect 13619 -7765 13652 -7731
rect 13686 -7765 13719 -7731
rect 13619 -7799 13719 -7765
rect 13619 -7833 13652 -7799
rect 13686 -7833 13719 -7799
rect 13619 -7867 13719 -7833
rect 13619 -7901 13652 -7867
rect 13686 -7901 13719 -7867
rect 13619 -7935 13719 -7901
rect 13619 -7969 13652 -7935
rect 13686 -7969 13719 -7935
rect 13619 -8003 13719 -7969
rect 13619 -8037 13652 -8003
rect 13686 -8037 13719 -8003
rect 13619 -8071 13719 -8037
rect 13619 -8105 13652 -8071
rect 13686 -8105 13719 -8071
rect 13619 -8139 13719 -8105
rect 13619 -8173 13652 -8139
rect 13686 -8173 13719 -8139
rect 13619 -8207 13719 -8173
rect 13619 -8241 13652 -8207
rect 13686 -8241 13719 -8207
rect 13619 -8275 13719 -8241
rect 13619 -8309 13652 -8275
rect 13686 -8309 13719 -8275
rect 13619 -8343 13719 -8309
rect 13619 -8377 13652 -8343
rect 13686 -8377 13719 -8343
rect 13619 -8411 13719 -8377
rect 13619 -8445 13652 -8411
rect 13686 -8445 13719 -8411
rect 13619 -8479 13719 -8445
rect 13619 -8513 13652 -8479
rect 13686 -8513 13719 -8479
rect 13619 -8547 13719 -8513
rect 13619 -8581 13652 -8547
rect 13686 -8581 13719 -8547
rect 13619 -8615 13719 -8581
rect 13619 -8649 13652 -8615
rect 13686 -8649 13719 -8615
rect 13619 -8683 13719 -8649
rect 13619 -8717 13652 -8683
rect 13686 -8717 13719 -8683
rect 13619 -8751 13719 -8717
rect 13619 -8785 13652 -8751
rect 13686 -8785 13719 -8751
rect 13619 -8819 13719 -8785
rect 13619 -8853 13652 -8819
rect 13686 -8853 13719 -8819
rect 13619 -8887 13719 -8853
rect 13619 -8921 13652 -8887
rect 13686 -8921 13719 -8887
rect 13619 -8955 13719 -8921
rect 13619 -8989 13652 -8955
rect 13686 -8989 13719 -8955
rect 13619 -9023 13719 -8989
rect 13619 -9057 13652 -9023
rect 13686 -9057 13719 -9023
rect 13619 -9091 13719 -9057
rect 13619 -9125 13652 -9091
rect 13686 -9125 13719 -9091
rect 13619 -9159 13719 -9125
rect 13619 -9193 13652 -9159
rect 13686 -9193 13719 -9159
rect 13619 -9227 13719 -9193
rect 13619 -9261 13652 -9227
rect 13686 -9261 13719 -9227
rect 13619 -9295 13719 -9261
rect 13619 -9329 13652 -9295
rect 13686 -9329 13719 -9295
rect 13619 -9363 13719 -9329
rect 13619 -9397 13652 -9363
rect 13686 -9397 13719 -9363
rect 13619 -9431 13719 -9397
rect 13619 -9465 13652 -9431
rect 13686 -9465 13719 -9431
rect 13619 -9499 13719 -9465
rect 13619 -9533 13652 -9499
rect 13686 -9533 13719 -9499
rect 13619 -9567 13719 -9533
rect 13619 -9601 13652 -9567
rect 13686 -9601 13719 -9567
rect 13619 -9635 13719 -9601
rect 13619 -9669 13652 -9635
rect 13686 -9669 13719 -9635
rect 13619 -9703 13719 -9669
rect 13619 -9737 13652 -9703
rect 13686 -9737 13719 -9703
rect 13619 -9771 13719 -9737
rect 13619 -9805 13652 -9771
rect 13686 -9805 13719 -9771
rect 13619 -9839 13719 -9805
rect 13619 -9873 13652 -9839
rect 13686 -9873 13719 -9839
rect 13619 -9907 13719 -9873
rect 13619 -9941 13652 -9907
rect 13686 -9941 13719 -9907
rect 13619 -9975 13719 -9941
rect 13619 -10009 13652 -9975
rect 13686 -10009 13719 -9975
rect 13619 -10043 13719 -10009
rect 13619 -10077 13652 -10043
rect 13686 -10077 13719 -10043
rect 13619 -10111 13719 -10077
rect 13619 -10145 13652 -10111
rect 13686 -10145 13719 -10111
rect 13619 -10179 13719 -10145
rect 13619 -10213 13652 -10179
rect 13686 -10213 13719 -10179
rect 13619 -10247 13719 -10213
rect 13619 -10281 13652 -10247
rect 13686 -10281 13719 -10247
rect 13619 -10315 13719 -10281
rect 13619 -10349 13652 -10315
rect 13686 -10349 13719 -10315
rect 13619 -10383 13719 -10349
rect 13619 -10417 13652 -10383
rect 13686 -10417 13719 -10383
rect 13619 -10451 13719 -10417
rect 13619 -10485 13652 -10451
rect 13686 -10485 13719 -10451
rect 13619 -10519 13719 -10485
rect 13619 -10553 13652 -10519
rect 13686 -10553 13719 -10519
rect 13619 -10587 13719 -10553
rect 13619 -10621 13652 -10587
rect 13686 -10621 13719 -10587
rect 13619 -10655 13719 -10621
rect 13619 -10689 13652 -10655
rect 13686 -10689 13719 -10655
rect 13619 -10723 13719 -10689
rect 13619 -10757 13652 -10723
rect 13686 -10757 13719 -10723
rect 13619 -10791 13719 -10757
rect 13619 -10825 13652 -10791
rect 13686 -10825 13719 -10791
rect 13619 -10859 13719 -10825
rect 13619 -10893 13652 -10859
rect 13686 -10893 13719 -10859
rect 13619 -10927 13719 -10893
rect 13619 -10961 13652 -10927
rect 13686 -10961 13719 -10927
rect 13619 -10995 13719 -10961
rect 13619 -11029 13652 -10995
rect 13686 -11029 13719 -10995
rect 13619 -11063 13719 -11029
rect 13619 -11097 13652 -11063
rect 13686 -11097 13719 -11063
rect 13619 -11131 13719 -11097
rect 13619 -11165 13652 -11131
rect 13686 -11165 13719 -11131
rect 13619 -11199 13719 -11165
rect 13619 -11233 13652 -11199
rect 13686 -11233 13719 -11199
rect 13619 -11267 13719 -11233
rect 13619 -11301 13652 -11267
rect 13686 -11301 13719 -11267
rect 13619 -11335 13719 -11301
rect 13619 -11369 13652 -11335
rect 13686 -11369 13719 -11335
rect 13619 -11403 13719 -11369
rect 13619 -11437 13652 -11403
rect 13686 -11437 13719 -11403
rect 13619 -11471 13719 -11437
rect 13619 -11505 13652 -11471
rect 13686 -11505 13719 -11471
rect 13619 -11539 13719 -11505
rect 13619 -11573 13652 -11539
rect 13686 -11573 13719 -11539
rect 13619 -11607 13719 -11573
rect 13619 -11641 13652 -11607
rect 13686 -11641 13719 -11607
rect 13619 -11675 13719 -11641
rect 13619 -11709 13652 -11675
rect 13686 -11709 13719 -11675
rect 13619 -11743 13719 -11709
rect 13619 -11777 13652 -11743
rect 13686 -11777 13719 -11743
rect 13619 -11811 13719 -11777
rect 13619 -11845 13652 -11811
rect 13686 -11845 13719 -11811
rect 13619 -11879 13719 -11845
rect 13619 -11913 13652 -11879
rect 13686 -11913 13719 -11879
rect 13619 -11947 13719 -11913
rect 13619 -11981 13652 -11947
rect 13686 -11981 13719 -11947
rect 13619 -12015 13719 -11981
rect 13619 -12049 13652 -12015
rect 13686 -12049 13719 -12015
rect 13619 -12083 13719 -12049
rect 13619 -12117 13652 -12083
rect 13686 -12117 13719 -12083
rect 13619 -12151 13719 -12117
rect 13619 -12185 13652 -12151
rect 13686 -12185 13719 -12151
rect 13619 -12219 13719 -12185
rect 13619 -12253 13652 -12219
rect 13686 -12253 13719 -12219
rect 13619 -12287 13719 -12253
rect 13619 -12321 13652 -12287
rect 13686 -12321 13719 -12287
rect 13619 -12355 13719 -12321
rect 13619 -12389 13652 -12355
rect 13686 -12389 13719 -12355
rect 13619 -12423 13719 -12389
rect 13619 -12457 13652 -12423
rect 13686 -12457 13719 -12423
rect 13619 -12491 13719 -12457
rect 13619 -12525 13652 -12491
rect 13686 -12525 13719 -12491
rect 13619 -12559 13719 -12525
rect 13619 -12593 13652 -12559
rect 13686 -12593 13719 -12559
rect 13619 -12627 13719 -12593
rect 13619 -12661 13652 -12627
rect 13686 -12661 13719 -12627
rect 13619 -12695 13719 -12661
rect 13619 -12729 13652 -12695
rect 13686 -12729 13719 -12695
rect 13619 -12763 13719 -12729
rect 13619 -12797 13652 -12763
rect 13686 -12797 13719 -12763
rect 13619 -12831 13719 -12797
rect 13619 -12865 13652 -12831
rect 13686 -12865 13719 -12831
rect 13619 -12899 13719 -12865
rect 13619 -12933 13652 -12899
rect 13686 -12933 13719 -12899
rect 13619 -12967 13719 -12933
rect 13619 -13001 13652 -12967
rect 13686 -13001 13719 -12967
rect 13619 -13035 13719 -13001
rect 13619 -13069 13652 -13035
rect 13686 -13069 13719 -13035
rect 13619 -13103 13719 -13069
rect 13619 -13137 13652 -13103
rect 13686 -13137 13719 -13103
rect 13619 -13171 13719 -13137
rect 13619 -13205 13652 -13171
rect 13686 -13205 13719 -13171
rect 13619 -13239 13719 -13205
rect 13619 -13273 13652 -13239
rect 13686 -13273 13719 -13239
rect 13619 -13307 13719 -13273
rect 13619 -13341 13652 -13307
rect 13686 -13341 13719 -13307
rect 13619 -13375 13719 -13341
rect 13619 -13409 13652 -13375
rect 13686 -13409 13719 -13375
rect 13619 -13443 13719 -13409
rect 13619 -13477 13652 -13443
rect 13686 -13477 13719 -13443
rect 13619 -13511 13719 -13477
rect 13619 -13545 13652 -13511
rect 13686 -13545 13719 -13511
rect 13619 -13579 13719 -13545
rect 13619 -13613 13652 -13579
rect 13686 -13613 13719 -13579
rect 13619 -13647 13719 -13613
rect 13619 -13681 13652 -13647
rect 13686 -13681 13719 -13647
rect 13619 -13715 13719 -13681
rect 13619 -13749 13652 -13715
rect 13686 -13749 13719 -13715
rect 13619 -13783 13719 -13749
rect 13619 -13817 13652 -13783
rect 13686 -13817 13719 -13783
rect 13619 -13851 13719 -13817
rect 13619 -13885 13652 -13851
rect 13686 -13885 13719 -13851
rect 13619 -13919 13719 -13885
rect 13619 -13953 13652 -13919
rect 13686 -13953 13719 -13919
rect 13619 -13987 13719 -13953
rect 13619 -14021 13652 -13987
rect 13686 -14021 13719 -13987
rect 13619 -14055 13719 -14021
rect 13619 -14089 13652 -14055
rect 13686 -14089 13719 -14055
rect 13619 -14123 13719 -14089
rect 13619 -14157 13652 -14123
rect 13686 -14157 13719 -14123
rect 13619 -14191 13719 -14157
rect 13619 -14225 13652 -14191
rect 13686 -14225 13719 -14191
rect 13619 -14259 13719 -14225
rect 13619 -14293 13652 -14259
rect 13686 -14293 13719 -14259
rect 13619 -14327 13719 -14293
rect 13619 -14361 13652 -14327
rect 13686 -14361 13719 -14327
rect 13619 -14395 13719 -14361
rect 13619 -14429 13652 -14395
rect 13686 -14429 13719 -14395
rect 13619 -14463 13719 -14429
rect 13619 -14497 13652 -14463
rect 13686 -14497 13719 -14463
rect 13619 -14531 13719 -14497
rect 13619 -14565 13652 -14531
rect 13686 -14565 13719 -14531
rect 13619 -14599 13719 -14565
rect 13619 -14633 13652 -14599
rect 13686 -14633 13719 -14599
rect 13619 -14667 13719 -14633
rect 13619 -14701 13652 -14667
rect 13686 -14701 13719 -14667
rect 13619 -14735 13719 -14701
rect 13619 -14769 13652 -14735
rect 13686 -14769 13719 -14735
rect 13619 -14803 13719 -14769
rect 13619 -14837 13652 -14803
rect 13686 -14837 13719 -14803
rect 13619 -14871 13719 -14837
rect 13619 -14905 13652 -14871
rect 13686 -14905 13719 -14871
rect 13619 -14939 13719 -14905
rect 13619 -14973 13652 -14939
rect 13686 -14973 13719 -14939
rect 13619 -15007 13719 -14973
rect 13619 -15041 13652 -15007
rect 13686 -15041 13719 -15007
rect 13619 -15075 13719 -15041
rect 13619 -15109 13652 -15075
rect 13686 -15109 13719 -15075
rect 13619 -15143 13719 -15109
rect 13619 -15177 13652 -15143
rect 13686 -15177 13719 -15143
rect 13619 -15211 13719 -15177
rect 13619 -15245 13652 -15211
rect 13686 -15245 13719 -15211
rect 13619 -15279 13719 -15245
rect 13619 -15313 13652 -15279
rect 13686 -15313 13719 -15279
rect 13619 -15347 13719 -15313
rect 13619 -15381 13652 -15347
rect 13686 -15381 13719 -15347
rect 13619 -15415 13719 -15381
rect 13619 -15449 13652 -15415
rect 13686 -15449 13719 -15415
rect 13619 -15483 13719 -15449
rect 13619 -15517 13652 -15483
rect 13686 -15517 13719 -15483
rect 13619 -15551 13719 -15517
rect 13619 -15585 13652 -15551
rect 13686 -15585 13719 -15551
rect 13619 -15619 13719 -15585
rect 13619 -15653 13652 -15619
rect 13686 -15653 13719 -15619
rect 13619 -15687 13719 -15653
rect 13619 -15721 13652 -15687
rect 13686 -15721 13719 -15687
rect 13619 -15755 13719 -15721
rect 13619 -15789 13652 -15755
rect 13686 -15789 13719 -15755
rect 13619 -15823 13719 -15789
rect 13619 -15857 13652 -15823
rect 13686 -15857 13719 -15823
rect 13619 -15891 13719 -15857
rect 13619 -15925 13652 -15891
rect 13686 -15925 13719 -15891
rect 13619 -15959 13719 -15925
rect 13619 -15993 13652 -15959
rect 13686 -15993 13719 -15959
rect 13619 -16027 13719 -15993
rect 13619 -16061 13652 -16027
rect 13686 -16061 13719 -16027
rect 13619 -16095 13719 -16061
rect 13619 -16129 13652 -16095
rect 13686 -16129 13719 -16095
rect 13619 -16163 13719 -16129
rect 13619 -16197 13652 -16163
rect 13686 -16197 13719 -16163
rect 13619 -16231 13719 -16197
rect 13619 -16265 13652 -16231
rect 13686 -16265 13719 -16231
rect 13619 -16299 13719 -16265
rect 13619 -16333 13652 -16299
rect 13686 -16333 13719 -16299
rect 13619 -16367 13719 -16333
rect 13619 -16401 13652 -16367
rect 13686 -16401 13719 -16367
rect 13619 -16435 13719 -16401
rect 13619 -16469 13652 -16435
rect 13686 -16469 13719 -16435
rect 13619 -16503 13719 -16469
rect 13619 -16537 13652 -16503
rect 13686 -16537 13719 -16503
rect 13619 -16571 13719 -16537
rect 13619 -16605 13652 -16571
rect 13686 -16605 13719 -16571
rect 13619 -16639 13719 -16605
rect 13619 -16673 13652 -16639
rect 13686 -16673 13719 -16639
rect 13619 -16707 13719 -16673
rect 13619 -16741 13652 -16707
rect 13686 -16741 13719 -16707
rect 13619 -16775 13719 -16741
rect 13619 -16809 13652 -16775
rect 13686 -16809 13719 -16775
rect 13619 -16843 13719 -16809
rect 13619 -16877 13652 -16843
rect 13686 -16877 13719 -16843
rect 13619 -16911 13719 -16877
rect 13619 -16945 13652 -16911
rect 13686 -16945 13719 -16911
rect 13619 -16979 13719 -16945
rect 13619 -17013 13652 -16979
rect 13686 -17013 13719 -16979
rect 13619 -17047 13719 -17013
rect 13619 -17081 13652 -17047
rect 13686 -17081 13719 -17047
rect 13619 -17115 13719 -17081
rect 13619 -17149 13652 -17115
rect 13686 -17149 13719 -17115
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< nsubdiff >>
rect -7606 -1290 3703 -1260
rect -7606 -1324 -7346 -1290
rect -7312 -1324 -7278 -1290
rect -7244 -1324 -7210 -1290
rect -7176 -1324 -7142 -1290
rect -7108 -1324 -7074 -1290
rect -7040 -1324 -7006 -1290
rect -6972 -1324 -6938 -1290
rect -6904 -1324 -6870 -1290
rect -6836 -1324 -6802 -1290
rect -6768 -1324 -6734 -1290
rect -6700 -1324 -6666 -1290
rect -6632 -1324 -6598 -1290
rect -6564 -1324 -6530 -1290
rect -6496 -1324 -6462 -1290
rect -6428 -1324 -6394 -1290
rect -6360 -1324 -6326 -1290
rect -6292 -1324 -6258 -1290
rect -6224 -1324 -6190 -1290
rect -6156 -1324 -6122 -1290
rect -6088 -1324 -6054 -1290
rect -6020 -1324 -5986 -1290
rect -5952 -1324 -5918 -1290
rect -5884 -1324 -5850 -1290
rect -5816 -1324 -5782 -1290
rect -5748 -1324 -5714 -1290
rect -5680 -1324 -5646 -1290
rect -5612 -1324 -5578 -1290
rect -5544 -1324 -5510 -1290
rect -5476 -1324 -5442 -1290
rect -5408 -1324 -5374 -1290
rect -5340 -1324 -5306 -1290
rect -5272 -1324 -5238 -1290
rect -5204 -1324 -5170 -1290
rect -5136 -1324 -5102 -1290
rect -5068 -1324 -5034 -1290
rect -5000 -1324 -4966 -1290
rect -4932 -1324 -4898 -1290
rect -4864 -1324 -4830 -1290
rect -4796 -1324 -4762 -1290
rect -4728 -1324 -4694 -1290
rect -4660 -1324 -4626 -1290
rect -4592 -1324 -4558 -1290
rect -4524 -1324 -4490 -1290
rect -4456 -1324 -4422 -1290
rect -4388 -1324 -4354 -1290
rect -4320 -1324 -4286 -1290
rect -4252 -1324 -4218 -1290
rect -4184 -1324 -4150 -1290
rect -4116 -1324 -4082 -1290
rect -4048 -1324 -4014 -1290
rect -3980 -1324 -3946 -1290
rect -3912 -1324 -3878 -1290
rect -3844 -1324 -3810 -1290
rect -3776 -1324 -3742 -1290
rect -3708 -1324 -3674 -1290
rect -3640 -1324 -3606 -1290
rect -3572 -1324 -3538 -1290
rect -3504 -1324 -3470 -1290
rect -3436 -1324 -3402 -1290
rect -3368 -1324 -3334 -1290
rect -3300 -1324 -3266 -1290
rect -3232 -1324 -3198 -1290
rect -3164 -1324 -3130 -1290
rect -3096 -1324 -3062 -1290
rect -3028 -1324 -2994 -1290
rect -2960 -1324 -2926 -1290
rect -2892 -1324 -2858 -1290
rect -2824 -1324 -2790 -1290
rect -2756 -1324 -2722 -1290
rect -2688 -1324 -2654 -1290
rect -2620 -1324 -2586 -1290
rect -2552 -1324 -2518 -1290
rect -2484 -1324 -2450 -1290
rect -2416 -1324 -2382 -1290
rect -2348 -1324 -2314 -1290
rect -2280 -1324 -2246 -1290
rect -2212 -1324 -2178 -1290
rect -2144 -1324 -2110 -1290
rect -2076 -1324 -2042 -1290
rect -2008 -1324 -1974 -1290
rect -1940 -1324 -1906 -1290
rect -1872 -1324 -1838 -1290
rect -1804 -1324 -1770 -1290
rect -1736 -1324 -1702 -1290
rect -1668 -1324 -1634 -1290
rect -1600 -1324 -1566 -1290
rect -1532 -1324 -1498 -1290
rect -1464 -1324 -1430 -1290
rect -1396 -1324 -1362 -1290
rect -1328 -1324 -1294 -1290
rect -1260 -1324 -1226 -1290
rect -1192 -1324 -1158 -1290
rect -1124 -1324 -1090 -1290
rect -1056 -1324 -1022 -1290
rect -988 -1324 -954 -1290
rect -920 -1324 -886 -1290
rect -852 -1324 -818 -1290
rect -784 -1324 -750 -1290
rect -716 -1324 -682 -1290
rect -648 -1324 -614 -1290
rect -580 -1324 -546 -1290
rect -512 -1324 -478 -1290
rect -444 -1324 -410 -1290
rect -376 -1324 -342 -1290
rect -308 -1324 -274 -1290
rect -240 -1324 -206 -1290
rect -172 -1324 -138 -1290
rect -104 -1324 -70 -1290
rect -36 -1324 -2 -1290
rect 32 -1324 66 -1290
rect 100 -1324 134 -1290
rect 168 -1324 202 -1290
rect 236 -1324 270 -1290
rect 304 -1324 338 -1290
rect 372 -1324 406 -1290
rect 440 -1324 474 -1290
rect 508 -1324 542 -1290
rect 576 -1324 610 -1290
rect 644 -1324 678 -1290
rect 712 -1324 746 -1290
rect 780 -1324 814 -1290
rect 848 -1324 882 -1290
rect 916 -1324 950 -1290
rect 984 -1324 1018 -1290
rect 1052 -1324 1086 -1290
rect 1120 -1324 1154 -1290
rect 1188 -1324 1222 -1290
rect 1256 -1324 1290 -1290
rect 1324 -1324 1358 -1290
rect 1392 -1324 1426 -1290
rect 1460 -1324 1494 -1290
rect 1528 -1324 1562 -1290
rect 1596 -1324 1630 -1290
rect 1664 -1324 1698 -1290
rect 1732 -1324 1766 -1290
rect 1800 -1324 1834 -1290
rect 1868 -1324 1902 -1290
rect 1936 -1324 1970 -1290
rect 2004 -1324 2038 -1290
rect 2072 -1324 2106 -1290
rect 2140 -1324 2174 -1290
rect 2208 -1324 2242 -1290
rect 2276 -1324 2310 -1290
rect 2344 -1324 2378 -1290
rect 2412 -1324 2446 -1290
rect 2480 -1324 2514 -1290
rect 2548 -1324 2582 -1290
rect 2616 -1324 2650 -1290
rect 2684 -1324 2718 -1290
rect 2752 -1324 2786 -1290
rect 2820 -1324 2854 -1290
rect 2888 -1324 2922 -1290
rect 2956 -1324 2990 -1290
rect 3024 -1324 3058 -1290
rect 3092 -1324 3126 -1290
rect 3160 -1324 3194 -1290
rect 3228 -1324 3262 -1290
rect 3296 -1324 3703 -1290
rect -7606 -1353 3703 -1324
rect -7605 -1539 -7512 -1353
rect -7605 -1573 -7576 -1539
rect -7542 -1573 -7512 -1539
rect -7605 -1607 -7512 -1573
rect -7605 -1641 -7576 -1607
rect -7542 -1641 -7512 -1607
rect -7605 -1675 -7512 -1641
rect -7605 -1709 -7576 -1675
rect -7542 -1709 -7512 -1675
rect -7605 -1743 -7512 -1709
rect -7605 -1777 -7576 -1743
rect -7542 -1777 -7512 -1743
rect -7605 -1811 -7512 -1777
rect -7605 -1845 -7576 -1811
rect -7542 -1845 -7512 -1811
rect -7605 -1879 -7512 -1845
rect -7605 -1913 -7576 -1879
rect -7542 -1913 -7512 -1879
rect -7605 -1947 -7512 -1913
rect -7605 -1981 -7576 -1947
rect -7542 -1981 -7512 -1947
rect -7605 -2015 -7512 -1981
rect -7605 -2049 -7576 -2015
rect -7542 -2049 -7512 -2015
rect -7605 -2083 -7512 -2049
rect -7605 -2117 -7576 -2083
rect -7542 -2117 -7512 -2083
rect -7605 -2151 -7512 -2117
rect -7605 -2185 -7576 -2151
rect -7542 -2185 -7512 -2151
rect -7605 -2219 -7512 -2185
rect -7605 -2253 -7576 -2219
rect -7542 -2253 -7512 -2219
rect -7605 -2287 -7512 -2253
rect -7605 -2321 -7576 -2287
rect -7542 -2321 -7512 -2287
rect -7605 -2355 -7512 -2321
rect -7605 -2389 -7576 -2355
rect -7542 -2389 -7512 -2355
rect -7605 -2423 -7512 -2389
rect -7605 -2457 -7576 -2423
rect -7542 -2457 -7512 -2423
rect -7605 -2491 -7512 -2457
rect -7605 -2525 -7576 -2491
rect -7542 -2525 -7512 -2491
rect -7605 -2559 -7512 -2525
rect -7605 -2593 -7576 -2559
rect -7542 -2593 -7512 -2559
rect -7605 -2627 -7512 -2593
rect -7605 -2661 -7576 -2627
rect -7542 -2661 -7512 -2627
rect -7605 -2695 -7512 -2661
rect -7605 -2729 -7576 -2695
rect -7542 -2729 -7512 -2695
rect -7605 -2763 -7512 -2729
rect -7605 -2797 -7576 -2763
rect -7542 -2797 -7512 -2763
rect -7605 -2831 -7512 -2797
rect -7605 -2865 -7576 -2831
rect -7542 -2865 -7512 -2831
rect -7605 -2899 -7512 -2865
rect -7605 -2933 -7576 -2899
rect -7542 -2933 -7512 -2899
rect -7605 -2967 -7512 -2933
rect -7605 -3001 -7576 -2967
rect -7542 -3001 -7512 -2967
rect -7605 -3035 -7512 -3001
rect -7605 -3069 -7576 -3035
rect -7542 -3069 -7512 -3035
rect -7605 -3103 -7512 -3069
rect -7605 -3137 -7576 -3103
rect -7542 -3137 -7512 -3103
rect -7605 -3171 -7512 -3137
rect -7605 -3205 -7576 -3171
rect -7542 -3205 -7512 -3171
rect -7605 -3239 -7512 -3205
rect -7605 -3273 -7576 -3239
rect -7542 -3273 -7512 -3239
rect -7605 -3307 -7512 -3273
rect -7605 -3341 -7576 -3307
rect -7542 -3341 -7512 -3307
rect -7605 -3375 -7512 -3341
rect -7605 -3409 -7576 -3375
rect -7542 -3409 -7512 -3375
rect -7605 -3443 -7512 -3409
rect -7605 -3477 -7576 -3443
rect -7542 -3477 -7512 -3443
rect -7605 -3511 -7512 -3477
rect -7605 -3545 -7576 -3511
rect -7542 -3545 -7512 -3511
rect -7605 -3579 -7512 -3545
rect -7605 -3613 -7576 -3579
rect -7542 -3613 -7512 -3579
rect -7605 -3647 -7512 -3613
rect -7605 -3681 -7576 -3647
rect -7542 -3681 -7512 -3647
rect -7605 -3715 -7512 -3681
rect -7605 -3749 -7576 -3715
rect -7542 -3749 -7512 -3715
rect -7605 -3783 -7512 -3749
rect -7605 -3817 -7576 -3783
rect -7542 -3817 -7512 -3783
rect -7605 -3851 -7512 -3817
rect -7605 -3885 -7576 -3851
rect -7542 -3885 -7512 -3851
rect -7605 -3919 -7512 -3885
rect -7605 -3953 -7576 -3919
rect -7542 -3953 -7512 -3919
rect -7605 -3987 -7512 -3953
rect -7605 -4021 -7576 -3987
rect -7542 -4021 -7512 -3987
rect -7605 -4055 -7512 -4021
rect -7605 -4089 -7576 -4055
rect -7542 -4089 -7512 -4055
rect -7605 -4123 -7512 -4089
rect -7605 -4157 -7576 -4123
rect -7542 -4157 -7512 -4123
rect -7605 -4191 -7512 -4157
rect -7605 -4225 -7576 -4191
rect -7542 -4225 -7512 -4191
rect -7605 -4259 -7512 -4225
rect -7605 -4293 -7576 -4259
rect -7542 -4293 -7512 -4259
rect -7605 -4327 -7512 -4293
rect -7605 -4361 -7576 -4327
rect -7542 -4361 -7512 -4327
rect -7605 -4395 -7512 -4361
rect -7605 -4429 -7576 -4395
rect -7542 -4429 -7512 -4395
rect -7605 -4463 -7512 -4429
rect -7605 -4497 -7576 -4463
rect -7542 -4497 -7512 -4463
rect -7605 -4531 -7512 -4497
rect -7605 -4565 -7576 -4531
rect -7542 -4565 -7512 -4531
rect -7605 -4599 -7512 -4565
rect -7605 -4633 -7576 -4599
rect -7542 -4633 -7512 -4599
rect -7605 -4667 -7512 -4633
rect -7605 -4701 -7576 -4667
rect -7542 -4701 -7512 -4667
rect -7605 -4735 -7512 -4701
rect -7605 -4769 -7576 -4735
rect -7542 -4769 -7512 -4735
rect -7605 -4803 -7512 -4769
rect -7605 -4837 -7576 -4803
rect -7542 -4837 -7512 -4803
rect -7605 -4871 -7512 -4837
rect -7605 -4905 -7576 -4871
rect -7542 -4905 -7512 -4871
rect -7605 -4939 -7512 -4905
rect -7605 -4973 -7576 -4939
rect -7542 -4973 -7512 -4939
rect -7605 -5007 -7512 -4973
rect -7605 -5041 -7576 -5007
rect -7542 -5041 -7512 -5007
rect -7605 -5075 -7512 -5041
rect -7605 -5109 -7576 -5075
rect -7542 -5109 -7512 -5075
rect -7605 -5143 -7512 -5109
rect -7605 -5177 -7576 -5143
rect -7542 -5177 -7512 -5143
rect -7605 -5211 -7512 -5177
rect -7605 -5245 -7576 -5211
rect -7542 -5245 -7512 -5211
rect -7605 -5279 -7512 -5245
rect -7605 -5313 -7576 -5279
rect -7542 -5313 -7512 -5279
rect -7605 -5347 -7512 -5313
rect -7605 -5381 -7576 -5347
rect -7542 -5381 -7512 -5347
rect -7605 -5415 -7512 -5381
rect -7605 -5449 -7576 -5415
rect -7542 -5449 -7512 -5415
rect -7605 -5483 -7512 -5449
rect -7605 -5517 -7576 -5483
rect -7542 -5517 -7512 -5483
rect -7605 -5551 -7512 -5517
rect -7605 -5585 -7576 -5551
rect -7542 -5585 -7512 -5551
rect -7605 -5619 -7512 -5585
rect -7605 -5653 -7576 -5619
rect -7542 -5653 -7512 -5619
rect -7605 -5687 -7512 -5653
rect -7605 -5721 -7576 -5687
rect -7542 -5721 -7512 -5687
rect -7605 -5755 -7512 -5721
rect -7605 -5789 -7576 -5755
rect -7542 -5789 -7512 -5755
rect -7605 -5823 -7512 -5789
rect -7605 -5857 -7576 -5823
rect -7542 -5857 -7512 -5823
rect -7605 -5891 -7512 -5857
rect -7605 -5925 -7576 -5891
rect -7542 -5925 -7512 -5891
rect -7605 -5959 -7512 -5925
rect -7605 -5993 -7576 -5959
rect -7542 -5993 -7512 -5959
rect -7605 -6027 -7512 -5993
rect -7605 -6061 -7576 -6027
rect -7542 -6061 -7512 -6027
rect -7605 -6095 -7512 -6061
rect -7605 -6129 -7576 -6095
rect -7542 -6129 -7512 -6095
rect -7605 -6163 -7512 -6129
rect -7605 -6197 -7576 -6163
rect -7542 -6197 -7512 -6163
rect -7605 -6231 -7512 -6197
rect -7605 -6265 -7576 -6231
rect -7542 -6265 -7512 -6231
rect -7605 -6299 -7512 -6265
rect -7605 -6333 -7576 -6299
rect -7542 -6333 -7512 -6299
rect -7605 -6367 -7512 -6333
rect -7605 -6401 -7576 -6367
rect -7542 -6401 -7512 -6367
rect -7605 -6435 -7512 -6401
rect -7605 -6469 -7576 -6435
rect -7542 -6469 -7512 -6435
rect -7605 -6503 -7512 -6469
rect -7605 -6537 -7576 -6503
rect -7542 -6537 -7512 -6503
rect -7605 -6571 -7512 -6537
rect -7605 -6605 -7576 -6571
rect -7542 -6605 -7512 -6571
rect -7605 -6639 -7512 -6605
rect -7605 -6673 -7576 -6639
rect -7542 -6673 -7512 -6639
rect -7605 -6707 -7512 -6673
rect -7605 -6741 -7576 -6707
rect -7542 -6741 -7512 -6707
rect -7605 -6775 -7512 -6741
rect -7605 -6809 -7576 -6775
rect -7542 -6809 -7512 -6775
rect -7605 -6843 -7512 -6809
rect -7605 -6877 -7576 -6843
rect -7542 -6877 -7512 -6843
rect -7605 -6911 -7512 -6877
rect -7605 -6945 -7576 -6911
rect -7542 -6945 -7512 -6911
rect -7605 -7140 -7512 -6945
rect 3610 -1552 3703 -1353
rect 3610 -1586 3639 -1552
rect 3673 -1586 3703 -1552
rect 3610 -1620 3703 -1586
rect 3610 -1654 3639 -1620
rect 3673 -1654 3703 -1620
rect 3610 -1688 3703 -1654
rect 3610 -1722 3639 -1688
rect 3673 -1722 3703 -1688
rect 3610 -1756 3703 -1722
rect 3610 -1790 3639 -1756
rect 3673 -1790 3703 -1756
rect 3610 -1824 3703 -1790
rect 3610 -1858 3639 -1824
rect 3673 -1858 3703 -1824
rect 3610 -1892 3703 -1858
rect 3610 -1926 3639 -1892
rect 3673 -1926 3703 -1892
rect 3610 -1960 3703 -1926
rect 3610 -1994 3639 -1960
rect 3673 -1994 3703 -1960
rect 3610 -2028 3703 -1994
rect 3610 -2062 3639 -2028
rect 3673 -2062 3703 -2028
rect 3610 -2096 3703 -2062
rect 3610 -2130 3639 -2096
rect 3673 -2130 3703 -2096
rect 3610 -2164 3703 -2130
rect 3610 -2198 3639 -2164
rect 3673 -2198 3703 -2164
rect 3610 -2232 3703 -2198
rect 3610 -2266 3639 -2232
rect 3673 -2266 3703 -2232
rect 3610 -2300 3703 -2266
rect 3610 -2334 3639 -2300
rect 3673 -2334 3703 -2300
rect 3610 -2368 3703 -2334
rect 3610 -2402 3639 -2368
rect 3673 -2402 3703 -2368
rect 3610 -2436 3703 -2402
rect 3610 -2470 3639 -2436
rect 3673 -2470 3703 -2436
rect 3610 -2504 3703 -2470
rect 3610 -2538 3639 -2504
rect 3673 -2538 3703 -2504
rect 3610 -2572 3703 -2538
rect 3610 -2606 3639 -2572
rect 3673 -2606 3703 -2572
rect 3610 -2640 3703 -2606
rect 3610 -2674 3639 -2640
rect 3673 -2674 3703 -2640
rect 3610 -2708 3703 -2674
rect 3610 -2742 3639 -2708
rect 3673 -2742 3703 -2708
rect 3610 -2776 3703 -2742
rect 3610 -2810 3639 -2776
rect 3673 -2810 3703 -2776
rect 3610 -2844 3703 -2810
rect 3610 -2878 3639 -2844
rect 3673 -2878 3703 -2844
rect 3610 -2912 3703 -2878
rect 3610 -2946 3639 -2912
rect 3673 -2946 3703 -2912
rect 3610 -2980 3703 -2946
rect 3610 -3014 3639 -2980
rect 3673 -3014 3703 -2980
rect 3610 -3048 3703 -3014
rect 3610 -3082 3639 -3048
rect 3673 -3082 3703 -3048
rect 3610 -3116 3703 -3082
rect 3610 -3150 3639 -3116
rect 3673 -3150 3703 -3116
rect 3610 -3184 3703 -3150
rect 3610 -3218 3639 -3184
rect 3673 -3218 3703 -3184
rect 3610 -3252 3703 -3218
rect 3610 -3286 3639 -3252
rect 3673 -3286 3703 -3252
rect 3610 -3320 3703 -3286
rect 3610 -3354 3639 -3320
rect 3673 -3354 3703 -3320
rect 3610 -3388 3703 -3354
rect 3610 -3422 3639 -3388
rect 3673 -3422 3703 -3388
rect 3610 -3456 3703 -3422
rect 3610 -3490 3639 -3456
rect 3673 -3490 3703 -3456
rect 3610 -3524 3703 -3490
rect 3610 -3558 3639 -3524
rect 3673 -3558 3703 -3524
rect 3610 -3592 3703 -3558
rect 3610 -3626 3639 -3592
rect 3673 -3626 3703 -3592
rect 3610 -3660 3703 -3626
rect 3610 -3694 3639 -3660
rect 3673 -3694 3703 -3660
rect 3610 -3728 3703 -3694
rect 3610 -3762 3639 -3728
rect 3673 -3762 3703 -3728
rect 3610 -3796 3703 -3762
rect 3610 -3830 3639 -3796
rect 3673 -3830 3703 -3796
rect 3610 -3864 3703 -3830
rect 3610 -3898 3639 -3864
rect 3673 -3898 3703 -3864
rect 3610 -3932 3703 -3898
rect 3610 -3966 3639 -3932
rect 3673 -3966 3703 -3932
rect 3610 -4000 3703 -3966
rect 3610 -4034 3639 -4000
rect 3673 -4034 3703 -4000
rect 3610 -4068 3703 -4034
rect 3610 -4102 3639 -4068
rect 3673 -4102 3703 -4068
rect 3610 -4136 3703 -4102
rect 3610 -4170 3639 -4136
rect 3673 -4170 3703 -4136
rect 3610 -4204 3703 -4170
rect 3610 -4238 3639 -4204
rect 3673 -4238 3703 -4204
rect 3610 -4272 3703 -4238
rect 3610 -4306 3639 -4272
rect 3673 -4306 3703 -4272
rect 3610 -4340 3703 -4306
rect 3610 -4374 3639 -4340
rect 3673 -4374 3703 -4340
rect 3610 -4408 3703 -4374
rect 3610 -4442 3639 -4408
rect 3673 -4442 3703 -4408
rect 3610 -4476 3703 -4442
rect 3610 -4510 3639 -4476
rect 3673 -4510 3703 -4476
rect 3610 -4544 3703 -4510
rect 3610 -4578 3639 -4544
rect 3673 -4578 3703 -4544
rect 3610 -4612 3703 -4578
rect 3610 -4646 3639 -4612
rect 3673 -4646 3703 -4612
rect 3610 -4680 3703 -4646
rect 3610 -4714 3639 -4680
rect 3673 -4714 3703 -4680
rect 3610 -4748 3703 -4714
rect 3610 -4782 3639 -4748
rect 3673 -4782 3703 -4748
rect 3610 -4816 3703 -4782
rect 3610 -4850 3639 -4816
rect 3673 -4850 3703 -4816
rect 3610 -4884 3703 -4850
rect 3610 -4918 3639 -4884
rect 3673 -4918 3703 -4884
rect 3610 -4952 3703 -4918
rect 3610 -4986 3639 -4952
rect 3673 -4986 3703 -4952
rect 3610 -5020 3703 -4986
rect 3610 -5054 3639 -5020
rect 3673 -5054 3703 -5020
rect 3610 -5088 3703 -5054
rect 3610 -5122 3639 -5088
rect 3673 -5122 3703 -5088
rect 3610 -5156 3703 -5122
rect 3610 -5190 3639 -5156
rect 3673 -5190 3703 -5156
rect 3610 -5224 3703 -5190
rect 3610 -5258 3639 -5224
rect 3673 -5258 3703 -5224
rect 3610 -5292 3703 -5258
rect 3610 -5326 3639 -5292
rect 3673 -5326 3703 -5292
rect 3610 -5360 3703 -5326
rect 3610 -5394 3639 -5360
rect 3673 -5394 3703 -5360
rect 3610 -5428 3703 -5394
rect 3610 -5462 3639 -5428
rect 3673 -5462 3703 -5428
rect 3610 -5496 3703 -5462
rect 3610 -5530 3639 -5496
rect 3673 -5530 3703 -5496
rect 3610 -5564 3703 -5530
rect 3610 -5598 3639 -5564
rect 3673 -5598 3703 -5564
rect 3610 -5632 3703 -5598
rect 3610 -5666 3639 -5632
rect 3673 -5666 3703 -5632
rect 3610 -5700 3703 -5666
rect 3610 -5734 3639 -5700
rect 3673 -5734 3703 -5700
rect 3610 -5768 3703 -5734
rect 3610 -5802 3639 -5768
rect 3673 -5802 3703 -5768
rect 3610 -5836 3703 -5802
rect 3610 -5870 3639 -5836
rect 3673 -5870 3703 -5836
rect 3610 -5904 3703 -5870
rect 3610 -5938 3639 -5904
rect 3673 -5938 3703 -5904
rect 3610 -5972 3703 -5938
rect 3610 -6006 3639 -5972
rect 3673 -6006 3703 -5972
rect 3610 -6040 3703 -6006
rect 3610 -6074 3639 -6040
rect 3673 -6074 3703 -6040
rect 3610 -6108 3703 -6074
rect 3610 -6142 3639 -6108
rect 3673 -6142 3703 -6108
rect 3610 -6176 3703 -6142
rect 3610 -6210 3639 -6176
rect 3673 -6210 3703 -6176
rect 3610 -6244 3703 -6210
rect 3610 -6278 3639 -6244
rect 3673 -6278 3703 -6244
rect 3610 -6312 3703 -6278
rect 3610 -6346 3639 -6312
rect 3673 -6346 3703 -6312
rect 3610 -6380 3703 -6346
rect 3610 -6414 3639 -6380
rect 3673 -6414 3703 -6380
rect 3610 -6448 3703 -6414
rect 3610 -6482 3639 -6448
rect 3673 -6482 3703 -6448
rect 3610 -6516 3703 -6482
rect 3610 -6550 3639 -6516
rect 3673 -6550 3703 -6516
rect 3610 -6584 3703 -6550
rect 3610 -6618 3639 -6584
rect 3673 -6618 3703 -6584
rect 3610 -6652 3703 -6618
rect 3610 -6686 3639 -6652
rect 3673 -6686 3703 -6652
rect 3610 -6720 3703 -6686
rect 3610 -6754 3639 -6720
rect 3673 -6754 3703 -6720
rect 3610 -6788 3703 -6754
rect 3610 -6822 3639 -6788
rect 3673 -6822 3703 -6788
rect 3610 -6856 3703 -6822
rect 3610 -6890 3639 -6856
rect 3673 -6890 3703 -6856
rect 3610 -6924 3703 -6890
rect 3610 -6958 3639 -6924
rect 3673 -6958 3703 -6924
rect 3610 -7140 3703 -6958
rect -7605 -7170 3703 -7140
rect -7605 -7204 -7249 -7170
rect -7215 -7204 -7181 -7170
rect -7147 -7204 -7113 -7170
rect -7079 -7204 -7045 -7170
rect -7011 -7204 -6977 -7170
rect -6943 -7204 -6909 -7170
rect -6875 -7204 -6841 -7170
rect -6807 -7204 -6773 -7170
rect -6739 -7204 -6705 -7170
rect -6671 -7204 -6637 -7170
rect -6603 -7204 -6569 -7170
rect -6535 -7204 -6501 -7170
rect -6467 -7204 -6433 -7170
rect -6399 -7204 -6365 -7170
rect -6331 -7204 -6297 -7170
rect -6263 -7204 -6229 -7170
rect -6195 -7204 -6161 -7170
rect -6127 -7204 -6093 -7170
rect -6059 -7204 -6025 -7170
rect -5991 -7204 -5957 -7170
rect -5923 -7204 -5889 -7170
rect -5855 -7204 -5821 -7170
rect -5787 -7204 -5753 -7170
rect -5719 -7204 -5685 -7170
rect -5651 -7204 -5617 -7170
rect -5583 -7204 -5549 -7170
rect -5515 -7204 -5481 -7170
rect -5447 -7204 -5413 -7170
rect -5379 -7204 -5345 -7170
rect -5311 -7204 -5277 -7170
rect -5243 -7204 -5209 -7170
rect -5175 -7204 -5141 -7170
rect -5107 -7204 -5073 -7170
rect -5039 -7204 -5005 -7170
rect -4971 -7204 -4937 -7170
rect -4903 -7204 -4869 -7170
rect -4835 -7204 -4801 -7170
rect -4767 -7204 -4733 -7170
rect -4699 -7204 -4665 -7170
rect -4631 -7204 -4597 -7170
rect -4563 -7204 -4529 -7170
rect -4495 -7204 -4461 -7170
rect -4427 -7204 -4393 -7170
rect -4359 -7204 -4325 -7170
rect -4291 -7204 -4257 -7170
rect -4223 -7204 -4189 -7170
rect -4155 -7204 -4121 -7170
rect -4087 -7204 -4053 -7170
rect -4019 -7204 -3985 -7170
rect -3951 -7204 -3917 -7170
rect -3883 -7204 -3849 -7170
rect -3815 -7204 -3781 -7170
rect -3747 -7204 -3713 -7170
rect -3679 -7204 -3645 -7170
rect -3611 -7204 -3577 -7170
rect -3543 -7204 -3509 -7170
rect -3475 -7204 -3441 -7170
rect -3407 -7204 -3373 -7170
rect -3339 -7204 -3305 -7170
rect -3271 -7204 -3237 -7170
rect -3203 -7204 -3169 -7170
rect -3135 -7204 -3101 -7170
rect -3067 -7204 -3033 -7170
rect -2999 -7204 -2965 -7170
rect -2931 -7204 -2897 -7170
rect -2863 -7204 -2829 -7170
rect -2795 -7204 -2761 -7170
rect -2727 -7204 -2693 -7170
rect -2659 -7204 -2625 -7170
rect -2591 -7204 -2557 -7170
rect -2523 -7204 -2489 -7170
rect -2455 -7204 -2421 -7170
rect -2387 -7204 -2353 -7170
rect -2319 -7204 -2285 -7170
rect -2251 -7204 -2217 -7170
rect -2183 -7204 -2149 -7170
rect -2115 -7204 -2081 -7170
rect -2047 -7204 -2013 -7170
rect -1979 -7204 -1945 -7170
rect -1911 -7204 -1877 -7170
rect -1843 -7204 -1809 -7170
rect -1775 -7204 -1741 -7170
rect -1707 -7204 -1673 -7170
rect -1639 -7204 -1605 -7170
rect -1571 -7204 -1537 -7170
rect -1503 -7204 -1469 -7170
rect -1435 -7204 -1401 -7170
rect -1367 -7204 -1333 -7170
rect -1299 -7204 -1265 -7170
rect -1231 -7204 -1197 -7170
rect -1163 -7204 -1129 -7170
rect -1095 -7204 -1061 -7170
rect -1027 -7204 -993 -7170
rect -959 -7204 -925 -7170
rect -891 -7204 -857 -7170
rect -823 -7204 -789 -7170
rect -755 -7204 -721 -7170
rect -687 -7204 -653 -7170
rect -619 -7204 -585 -7170
rect -551 -7204 -517 -7170
rect -483 -7204 -449 -7170
rect -415 -7204 -381 -7170
rect -347 -7204 -313 -7170
rect -279 -7204 -245 -7170
rect -211 -7204 -177 -7170
rect -143 -7204 -109 -7170
rect -75 -7204 -41 -7170
rect -7 -7204 27 -7170
rect 61 -7204 95 -7170
rect 129 -7204 163 -7170
rect 197 -7204 231 -7170
rect 265 -7204 299 -7170
rect 333 -7204 367 -7170
rect 401 -7204 435 -7170
rect 469 -7204 503 -7170
rect 537 -7204 571 -7170
rect 605 -7204 639 -7170
rect 673 -7204 707 -7170
rect 741 -7204 775 -7170
rect 809 -7204 843 -7170
rect 877 -7204 911 -7170
rect 945 -7204 979 -7170
rect 1013 -7204 1047 -7170
rect 1081 -7204 1115 -7170
rect 1149 -7204 1183 -7170
rect 1217 -7204 1251 -7170
rect 1285 -7204 1319 -7170
rect 1353 -7204 1387 -7170
rect 1421 -7204 1455 -7170
rect 1489 -7204 1523 -7170
rect 1557 -7204 1591 -7170
rect 1625 -7204 1659 -7170
rect 1693 -7204 1727 -7170
rect 1761 -7204 1795 -7170
rect 1829 -7204 1863 -7170
rect 1897 -7204 1931 -7170
rect 1965 -7204 1999 -7170
rect 2033 -7204 2067 -7170
rect 2101 -7204 2135 -7170
rect 2169 -7204 2203 -7170
rect 2237 -7204 2271 -7170
rect 2305 -7204 2339 -7170
rect 2373 -7204 2407 -7170
rect 2441 -7204 2475 -7170
rect 2509 -7204 2543 -7170
rect 2577 -7204 2611 -7170
rect 2645 -7204 2679 -7170
rect 2713 -7204 2747 -7170
rect 2781 -7204 2815 -7170
rect 2849 -7204 2883 -7170
rect 2917 -7204 2951 -7170
rect 2985 -7204 3019 -7170
rect 3053 -7204 3087 -7170
rect 3121 -7204 3155 -7170
rect 3189 -7204 3223 -7170
rect 3257 -7204 3291 -7170
rect 3325 -7204 3359 -7170
rect 3393 -7204 3703 -7170
rect -7605 -7233 3703 -7204
<< psubdiffcont >>
rect -7264 -7588 -7230 -7554
rect -7196 -7588 -7162 -7554
rect -7128 -7588 -7094 -7554
rect -7060 -7588 -7026 -7554
rect -6992 -7588 -6958 -7554
rect -6924 -7588 -6890 -7554
rect -6856 -7588 -6822 -7554
rect -6788 -7588 -6754 -7554
rect -6720 -7588 -6686 -7554
rect -6652 -7588 -6618 -7554
rect -6584 -7588 -6550 -7554
rect -6516 -7588 -6482 -7554
rect -6448 -7588 -6414 -7554
rect -6380 -7588 -6346 -7554
rect -6312 -7588 -6278 -7554
rect -6244 -7588 -6210 -7554
rect -6176 -7588 -6142 -7554
rect -6108 -7588 -6074 -7554
rect -6040 -7588 -6006 -7554
rect -5972 -7588 -5938 -7554
rect -5904 -7588 -5870 -7554
rect -5836 -7588 -5802 -7554
rect -5768 -7588 -5734 -7554
rect -5700 -7588 -5666 -7554
rect -5632 -7588 -5598 -7554
rect -5564 -7588 -5530 -7554
rect -5496 -7588 -5462 -7554
rect -5428 -7588 -5394 -7554
rect -5360 -7588 -5326 -7554
rect -5292 -7588 -5258 -7554
rect -5224 -7588 -5190 -7554
rect -5156 -7588 -5122 -7554
rect -5088 -7588 -5054 -7554
rect -5020 -7588 -4986 -7554
rect -4952 -7588 -4918 -7554
rect -4884 -7588 -4850 -7554
rect -4816 -7588 -4782 -7554
rect -4748 -7588 -4714 -7554
rect -4680 -7588 -4646 -7554
rect -4612 -7588 -4578 -7554
rect -4544 -7588 -4510 -7554
rect -4476 -7588 -4442 -7554
rect -4408 -7588 -4374 -7554
rect -4340 -7588 -4306 -7554
rect -4272 -7588 -4238 -7554
rect -4204 -7588 -4170 -7554
rect -4136 -7588 -4102 -7554
rect -4068 -7588 -4034 -7554
rect -4000 -7588 -3966 -7554
rect -3932 -7588 -3898 -7554
rect -3864 -7588 -3830 -7554
rect -3796 -7588 -3762 -7554
rect -3728 -7588 -3694 -7554
rect -3660 -7588 -3626 -7554
rect -3592 -7588 -3558 -7554
rect -3524 -7588 -3490 -7554
rect -3456 -7588 -3422 -7554
rect -3388 -7588 -3354 -7554
rect -3320 -7588 -3286 -7554
rect -3252 -7588 -3218 -7554
rect -3184 -7588 -3150 -7554
rect -3116 -7588 -3082 -7554
rect -3048 -7588 -3014 -7554
rect -2980 -7588 -2946 -7554
rect -2912 -7588 -2878 -7554
rect -2844 -7588 -2810 -7554
rect -2776 -7588 -2742 -7554
rect -2708 -7588 -2674 -7554
rect -2640 -7588 -2606 -7554
rect -2572 -7588 -2538 -7554
rect -2504 -7588 -2470 -7554
rect -2436 -7588 -2402 -7554
rect -2368 -7588 -2334 -7554
rect -2300 -7588 -2266 -7554
rect -2232 -7588 -2198 -7554
rect -2164 -7588 -2130 -7554
rect -2096 -7588 -2062 -7554
rect -2028 -7588 -1994 -7554
rect -1960 -7588 -1926 -7554
rect -1892 -7588 -1858 -7554
rect -1824 -7588 -1790 -7554
rect -1756 -7588 -1722 -7554
rect -1688 -7588 -1654 -7554
rect -1620 -7588 -1586 -7554
rect -1552 -7588 -1518 -7554
rect -1484 -7588 -1450 -7554
rect -1416 -7588 -1382 -7554
rect -1348 -7588 -1314 -7554
rect -1280 -7588 -1246 -7554
rect -1212 -7588 -1178 -7554
rect -1144 -7588 -1110 -7554
rect -1076 -7588 -1042 -7554
rect -1008 -7588 -974 -7554
rect -940 -7588 -906 -7554
rect -872 -7588 -838 -7554
rect -804 -7588 -770 -7554
rect -736 -7588 -702 -7554
rect -668 -7588 -634 -7554
rect -600 -7588 -566 -7554
rect -532 -7588 -498 -7554
rect -464 -7588 -430 -7554
rect -396 -7588 -362 -7554
rect -328 -7588 -294 -7554
rect -260 -7588 -226 -7554
rect -192 -7588 -158 -7554
rect -124 -7588 -90 -7554
rect -56 -7588 -22 -7554
rect 12 -7588 46 -7554
rect 80 -7588 114 -7554
rect 148 -7588 182 -7554
rect 216 -7588 250 -7554
rect 284 -7588 318 -7554
rect 352 -7588 386 -7554
rect 420 -7588 454 -7554
rect 488 -7588 522 -7554
rect 556 -7588 590 -7554
rect 624 -7588 658 -7554
rect 692 -7588 726 -7554
rect 760 -7588 794 -7554
rect 828 -7588 862 -7554
rect 896 -7588 930 -7554
rect 964 -7588 998 -7554
rect 1032 -7588 1066 -7554
rect 1100 -7588 1134 -7554
rect 1168 -7588 1202 -7554
rect 1236 -7588 1270 -7554
rect 1304 -7588 1338 -7554
rect 1372 -7588 1406 -7554
rect 1440 -7588 1474 -7554
rect 1508 -7588 1542 -7554
rect 1576 -7588 1610 -7554
rect 1644 -7588 1678 -7554
rect 1712 -7588 1746 -7554
rect 1780 -7588 1814 -7554
rect 1848 -7588 1882 -7554
rect 1916 -7588 1950 -7554
rect 1984 -7588 2018 -7554
rect 2052 -7588 2086 -7554
rect 2120 -7588 2154 -7554
rect 2188 -7588 2222 -7554
rect 2256 -7588 2290 -7554
rect 2324 -7588 2358 -7554
rect 2392 -7588 2426 -7554
rect 2460 -7588 2494 -7554
rect 2528 -7588 2562 -7554
rect 2596 -7588 2630 -7554
rect 2664 -7588 2698 -7554
rect 2732 -7588 2766 -7554
rect 2800 -7588 2834 -7554
rect 2868 -7588 2902 -7554
rect 2936 -7588 2970 -7554
rect 3004 -7588 3038 -7554
rect 3072 -7588 3106 -7554
rect 3140 -7588 3174 -7554
rect 3208 -7588 3242 -7554
rect 3276 -7588 3310 -7554
rect 3344 -7588 3378 -7554
rect 3412 -7588 3446 -7554
rect 3480 -7588 3514 -7554
rect 3548 -7588 3582 -7554
rect 3616 -7588 3650 -7554
rect 3684 -7588 3718 -7554
rect 3752 -7588 3786 -7554
rect 3820 -7588 3854 -7554
rect 3888 -7588 3922 -7554
rect 3956 -7588 3990 -7554
rect 4024 -7588 4058 -7554
rect 4092 -7588 4126 -7554
rect 4160 -7588 4194 -7554
rect 4228 -7588 4262 -7554
rect 4296 -7588 4330 -7554
rect 4364 -7588 4398 -7554
rect 4432 -7588 4466 -7554
rect 4500 -7588 4534 -7554
rect 4568 -7588 4602 -7554
rect 4636 -7588 4670 -7554
rect 4704 -7588 4738 -7554
rect 4772 -7588 4806 -7554
rect 4840 -7588 4874 -7554
rect 4908 -7588 4942 -7554
rect 4976 -7588 5010 -7554
rect 5044 -7588 5078 -7554
rect 5112 -7588 5146 -7554
rect 5180 -7588 5214 -7554
rect 5248 -7588 5282 -7554
rect 5316 -7588 5350 -7554
rect 5384 -7588 5418 -7554
rect 5452 -7588 5486 -7554
rect 5520 -7588 5554 -7554
rect 5588 -7588 5622 -7554
rect 5656 -7588 5690 -7554
rect 5724 -7588 5758 -7554
rect 5792 -7588 5826 -7554
rect 5860 -7588 5894 -7554
rect 5928 -7588 5962 -7554
rect 5996 -7588 6030 -7554
rect 6064 -7588 6098 -7554
rect 6132 -7588 6166 -7554
rect 6200 -7588 6234 -7554
rect 6268 -7588 6302 -7554
rect 6336 -7588 6370 -7554
rect 6404 -7588 6438 -7554
rect 6472 -7588 6506 -7554
rect 6540 -7588 6574 -7554
rect 6608 -7588 6642 -7554
rect 6676 -7588 6710 -7554
rect 6744 -7588 6778 -7554
rect 6812 -7588 6846 -7554
rect 6880 -7588 6914 -7554
rect 6948 -7588 6982 -7554
rect 7016 -7588 7050 -7554
rect 7084 -7588 7118 -7554
rect 7152 -7588 7186 -7554
rect 7220 -7588 7254 -7554
rect 7288 -7588 7322 -7554
rect 7356 -7588 7390 -7554
rect 7424 -7588 7458 -7554
rect 7492 -7588 7526 -7554
rect 7560 -7588 7594 -7554
rect 7628 -7588 7662 -7554
rect 7696 -7588 7730 -7554
rect 7764 -7588 7798 -7554
rect 7832 -7588 7866 -7554
rect 7900 -7588 7934 -7554
rect 7968 -7588 8002 -7554
rect 8036 -7588 8070 -7554
rect 8104 -7588 8138 -7554
rect 8172 -7588 8206 -7554
rect 8240 -7588 8274 -7554
rect 8308 -7588 8342 -7554
rect 8376 -7588 8410 -7554
rect 8444 -7588 8478 -7554
rect 8512 -7588 8546 -7554
rect 8580 -7588 8614 -7554
rect 8648 -7588 8682 -7554
rect 8716 -7588 8750 -7554
rect 8784 -7588 8818 -7554
rect 8852 -7588 8886 -7554
rect 8920 -7588 8954 -7554
rect 8988 -7588 9022 -7554
rect 9056 -7588 9090 -7554
rect 9124 -7588 9158 -7554
rect 9192 -7588 9226 -7554
rect 9260 -7588 9294 -7554
rect 9328 -7588 9362 -7554
rect 9396 -7588 9430 -7554
rect 9464 -7588 9498 -7554
rect 9532 -7588 9566 -7554
rect 9600 -7588 9634 -7554
rect 9668 -7588 9702 -7554
rect 9736 -7588 9770 -7554
rect 9804 -7588 9838 -7554
rect 9872 -7588 9906 -7554
rect 9940 -7588 9974 -7554
rect 10008 -7588 10042 -7554
rect 10076 -7588 10110 -7554
rect 10144 -7588 10178 -7554
rect 10212 -7588 10246 -7554
rect 10280 -7588 10314 -7554
rect 10348 -7588 10382 -7554
rect 10416 -7588 10450 -7554
rect 10484 -7588 10518 -7554
rect 10552 -7588 10586 -7554
rect 10620 -7588 10654 -7554
rect 10688 -7588 10722 -7554
rect 10756 -7588 10790 -7554
rect 10824 -7588 10858 -7554
rect 10892 -7588 10926 -7554
rect 10960 -7588 10994 -7554
rect 11028 -7588 11062 -7554
rect 11096 -7588 11130 -7554
rect 11164 -7588 11198 -7554
rect 11232 -7588 11266 -7554
rect 11300 -7588 11334 -7554
rect 11368 -7588 11402 -7554
rect 11436 -7588 11470 -7554
rect 11504 -7588 11538 -7554
rect 11572 -7588 11606 -7554
rect 11640 -7588 11674 -7554
rect 11708 -7588 11742 -7554
rect 11776 -7588 11810 -7554
rect 11844 -7588 11878 -7554
rect 11912 -7588 11946 -7554
rect 11980 -7588 12014 -7554
rect 12048 -7588 12082 -7554
rect 12116 -7588 12150 -7554
rect 12184 -7588 12218 -7554
rect 12252 -7588 12286 -7554
rect 12320 -7588 12354 -7554
rect 12388 -7588 12422 -7554
rect 12456 -7588 12490 -7554
rect 12524 -7588 12558 -7554
rect 12592 -7588 12626 -7554
rect 12660 -7588 12694 -7554
rect 12728 -7588 12762 -7554
rect 12796 -7588 12830 -7554
rect 12864 -7588 12898 -7554
rect 12932 -7588 12966 -7554
rect 13000 -7588 13034 -7554
rect 13068 -7588 13102 -7554
rect 13136 -7588 13170 -7554
rect 13204 -7588 13238 -7554
rect 13272 -7588 13306 -7554
rect 13340 -7588 13374 -7554
rect 13408 -7588 13442 -7554
rect -7572 -7884 -7538 -7850
rect -7572 -7952 -7538 -7918
rect -7572 -8020 -7538 -7986
rect -7572 -8088 -7538 -8054
rect -7572 -8156 -7538 -8122
rect -7572 -8224 -7538 -8190
rect -7572 -8292 -7538 -8258
rect -7572 -8360 -7538 -8326
rect -7572 -8428 -7538 -8394
rect -7572 -8496 -7538 -8462
rect -7572 -8564 -7538 -8530
rect -7572 -8632 -7538 -8598
rect -7572 -8700 -7538 -8666
rect -7572 -8768 -7538 -8734
rect -7572 -8836 -7538 -8802
rect -7572 -8904 -7538 -8870
rect -7572 -8972 -7538 -8938
rect -7572 -9040 -7538 -9006
rect -7572 -9108 -7538 -9074
rect -7572 -9176 -7538 -9142
rect -7572 -9244 -7538 -9210
rect -7572 -9312 -7538 -9278
rect -7572 -9380 -7538 -9346
rect -7572 -9448 -7538 -9414
rect -7572 -9516 -7538 -9482
rect -7572 -9584 -7538 -9550
rect -7572 -9652 -7538 -9618
rect -7572 -9720 -7538 -9686
rect -7572 -9788 -7538 -9754
rect -7572 -9856 -7538 -9822
rect -7572 -9924 -7538 -9890
rect -7572 -9992 -7538 -9958
rect -7572 -10060 -7538 -10026
rect -7572 -10128 -7538 -10094
rect -7572 -10196 -7538 -10162
rect -7572 -10264 -7538 -10230
rect -7572 -10332 -7538 -10298
rect -7572 -10400 -7538 -10366
rect -7572 -10468 -7538 -10434
rect -7572 -10536 -7538 -10502
rect -7572 -10604 -7538 -10570
rect -7572 -10672 -7538 -10638
rect -7572 -10740 -7538 -10706
rect -7572 -10808 -7538 -10774
rect -7572 -10876 -7538 -10842
rect -7572 -10944 -7538 -10910
rect -7572 -11012 -7538 -10978
rect -7572 -11080 -7538 -11046
rect -7572 -11148 -7538 -11114
rect -7572 -11216 -7538 -11182
rect -7572 -11284 -7538 -11250
rect -7572 -11352 -7538 -11318
rect -7572 -11420 -7538 -11386
rect -7572 -11488 -7538 -11454
rect -7572 -11556 -7538 -11522
rect -7572 -11624 -7538 -11590
rect -7572 -11692 -7538 -11658
rect -7572 -11760 -7538 -11726
rect -7572 -11828 -7538 -11794
rect -7572 -11896 -7538 -11862
rect -7572 -11964 -7538 -11930
rect -7572 -12032 -7538 -11998
rect -7572 -12100 -7538 -12066
rect -7572 -12168 -7538 -12134
rect -7572 -12236 -7538 -12202
rect -7572 -12304 -7538 -12270
rect -7572 -12372 -7538 -12338
rect -7572 -12440 -7538 -12406
rect -7572 -12508 -7538 -12474
rect -7572 -12576 -7538 -12542
rect -7572 -12644 -7538 -12610
rect -7572 -12712 -7538 -12678
rect -7572 -12780 -7538 -12746
rect -7572 -12848 -7538 -12814
rect -7572 -12916 -7538 -12882
rect -7572 -12984 -7538 -12950
rect -7572 -13052 -7538 -13018
rect -7572 -13120 -7538 -13086
rect -7572 -13188 -7538 -13154
rect -7572 -13256 -7538 -13222
rect -7572 -13324 -7538 -13290
rect -7572 -13392 -7538 -13358
rect -7572 -13460 -7538 -13426
rect -7572 -13528 -7538 -13494
rect -7572 -13596 -7538 -13562
rect -7572 -13664 -7538 -13630
rect -7572 -13732 -7538 -13698
rect -7572 -13800 -7538 -13766
rect -7572 -13868 -7538 -13834
rect -7572 -13936 -7538 -13902
rect -7572 -14004 -7538 -13970
rect -7572 -14072 -7538 -14038
rect -7572 -14140 -7538 -14106
rect -7572 -14208 -7538 -14174
rect -7572 -14276 -7538 -14242
rect -7572 -14344 -7538 -14310
rect -7572 -14412 -7538 -14378
rect -7572 -14480 -7538 -14446
rect -7572 -14548 -7538 -14514
rect -7572 -14616 -7538 -14582
rect -7572 -14684 -7538 -14650
rect -7572 -14752 -7538 -14718
rect -7572 -14820 -7538 -14786
rect -7572 -14888 -7538 -14854
rect -7572 -14956 -7538 -14922
rect -7572 -15024 -7538 -14990
rect -7572 -15092 -7538 -15058
rect -7572 -15160 -7538 -15126
rect -7572 -15228 -7538 -15194
rect -7572 -15296 -7538 -15262
rect -7572 -15364 -7538 -15330
rect -7572 -15432 -7538 -15398
rect -7572 -15500 -7538 -15466
rect -7572 -15568 -7538 -15534
rect -7572 -15636 -7538 -15602
rect -7572 -15704 -7538 -15670
rect -7572 -15772 -7538 -15738
rect -7572 -15840 -7538 -15806
rect -7572 -15908 -7538 -15874
rect -7572 -15976 -7538 -15942
rect -7572 -16044 -7538 -16010
rect -7572 -16112 -7538 -16078
rect -7572 -16180 -7538 -16146
rect -7572 -16248 -7538 -16214
rect -7572 -16316 -7538 -16282
rect -7572 -16384 -7538 -16350
rect -7572 -16452 -7538 -16418
rect -7572 -16520 -7538 -16486
rect -7572 -16588 -7538 -16554
rect -7572 -16656 -7538 -16622
rect -7572 -16724 -7538 -16690
rect -7572 -16792 -7538 -16758
rect -7572 -16860 -7538 -16826
rect -7572 -16928 -7538 -16894
rect -7572 -16996 -7538 -16962
rect -7572 -17064 -7538 -17030
rect -7572 -17132 -7538 -17098
rect -7572 -17200 -7538 -17166
rect -7572 -17268 -7538 -17234
rect 13652 -7765 13686 -7731
rect 13652 -7833 13686 -7799
rect 13652 -7901 13686 -7867
rect 13652 -7969 13686 -7935
rect 13652 -8037 13686 -8003
rect 13652 -8105 13686 -8071
rect 13652 -8173 13686 -8139
rect 13652 -8241 13686 -8207
rect 13652 -8309 13686 -8275
rect 13652 -8377 13686 -8343
rect 13652 -8445 13686 -8411
rect 13652 -8513 13686 -8479
rect 13652 -8581 13686 -8547
rect 13652 -8649 13686 -8615
rect 13652 -8717 13686 -8683
rect 13652 -8785 13686 -8751
rect 13652 -8853 13686 -8819
rect 13652 -8921 13686 -8887
rect 13652 -8989 13686 -8955
rect 13652 -9057 13686 -9023
rect 13652 -9125 13686 -9091
rect 13652 -9193 13686 -9159
rect 13652 -9261 13686 -9227
rect 13652 -9329 13686 -9295
rect 13652 -9397 13686 -9363
rect 13652 -9465 13686 -9431
rect 13652 -9533 13686 -9499
rect 13652 -9601 13686 -9567
rect 13652 -9669 13686 -9635
rect 13652 -9737 13686 -9703
rect 13652 -9805 13686 -9771
rect 13652 -9873 13686 -9839
rect 13652 -9941 13686 -9907
rect 13652 -10009 13686 -9975
rect 13652 -10077 13686 -10043
rect 13652 -10145 13686 -10111
rect 13652 -10213 13686 -10179
rect 13652 -10281 13686 -10247
rect 13652 -10349 13686 -10315
rect 13652 -10417 13686 -10383
rect 13652 -10485 13686 -10451
rect 13652 -10553 13686 -10519
rect 13652 -10621 13686 -10587
rect 13652 -10689 13686 -10655
rect 13652 -10757 13686 -10723
rect 13652 -10825 13686 -10791
rect 13652 -10893 13686 -10859
rect 13652 -10961 13686 -10927
rect 13652 -11029 13686 -10995
rect 13652 -11097 13686 -11063
rect 13652 -11165 13686 -11131
rect 13652 -11233 13686 -11199
rect 13652 -11301 13686 -11267
rect 13652 -11369 13686 -11335
rect 13652 -11437 13686 -11403
rect 13652 -11505 13686 -11471
rect 13652 -11573 13686 -11539
rect 13652 -11641 13686 -11607
rect 13652 -11709 13686 -11675
rect 13652 -11777 13686 -11743
rect 13652 -11845 13686 -11811
rect 13652 -11913 13686 -11879
rect 13652 -11981 13686 -11947
rect 13652 -12049 13686 -12015
rect 13652 -12117 13686 -12083
rect 13652 -12185 13686 -12151
rect 13652 -12253 13686 -12219
rect 13652 -12321 13686 -12287
rect 13652 -12389 13686 -12355
rect 13652 -12457 13686 -12423
rect 13652 -12525 13686 -12491
rect 13652 -12593 13686 -12559
rect 13652 -12661 13686 -12627
rect 13652 -12729 13686 -12695
rect 13652 -12797 13686 -12763
rect 13652 -12865 13686 -12831
rect 13652 -12933 13686 -12899
rect 13652 -13001 13686 -12967
rect 13652 -13069 13686 -13035
rect 13652 -13137 13686 -13103
rect 13652 -13205 13686 -13171
rect 13652 -13273 13686 -13239
rect 13652 -13341 13686 -13307
rect 13652 -13409 13686 -13375
rect 13652 -13477 13686 -13443
rect 13652 -13545 13686 -13511
rect 13652 -13613 13686 -13579
rect 13652 -13681 13686 -13647
rect 13652 -13749 13686 -13715
rect 13652 -13817 13686 -13783
rect 13652 -13885 13686 -13851
rect 13652 -13953 13686 -13919
rect 13652 -14021 13686 -13987
rect 13652 -14089 13686 -14055
rect 13652 -14157 13686 -14123
rect 13652 -14225 13686 -14191
rect 13652 -14293 13686 -14259
rect 13652 -14361 13686 -14327
rect 13652 -14429 13686 -14395
rect 13652 -14497 13686 -14463
rect 13652 -14565 13686 -14531
rect 13652 -14633 13686 -14599
rect 13652 -14701 13686 -14667
rect 13652 -14769 13686 -14735
rect 13652 -14837 13686 -14803
rect 13652 -14905 13686 -14871
rect 13652 -14973 13686 -14939
rect 13652 -15041 13686 -15007
rect 13652 -15109 13686 -15075
rect 13652 -15177 13686 -15143
rect 13652 -15245 13686 -15211
rect 13652 -15313 13686 -15279
rect 13652 -15381 13686 -15347
rect 13652 -15449 13686 -15415
rect 13652 -15517 13686 -15483
rect 13652 -15585 13686 -15551
rect 13652 -15653 13686 -15619
rect 13652 -15721 13686 -15687
rect 13652 -15789 13686 -15755
rect 13652 -15857 13686 -15823
rect 13652 -15925 13686 -15891
rect 13652 -15993 13686 -15959
rect 13652 -16061 13686 -16027
rect 13652 -16129 13686 -16095
rect 13652 -16197 13686 -16163
rect 13652 -16265 13686 -16231
rect 13652 -16333 13686 -16299
rect 13652 -16401 13686 -16367
rect 13652 -16469 13686 -16435
rect 13652 -16537 13686 -16503
rect 13652 -16605 13686 -16571
rect 13652 -16673 13686 -16639
rect 13652 -16741 13686 -16707
rect 13652 -16809 13686 -16775
rect 13652 -16877 13686 -16843
rect 13652 -16945 13686 -16911
rect 13652 -17013 13686 -16979
rect 13652 -17081 13686 -17047
rect 13652 -17149 13686 -17115
<< nsubdiffcont >>
rect -7346 -1324 -7312 -1290
rect -7278 -1324 -7244 -1290
rect -7210 -1324 -7176 -1290
rect -7142 -1324 -7108 -1290
rect -7074 -1324 -7040 -1290
rect -7006 -1324 -6972 -1290
rect -6938 -1324 -6904 -1290
rect -6870 -1324 -6836 -1290
rect -6802 -1324 -6768 -1290
rect -6734 -1324 -6700 -1290
rect -6666 -1324 -6632 -1290
rect -6598 -1324 -6564 -1290
rect -6530 -1324 -6496 -1290
rect -6462 -1324 -6428 -1290
rect -6394 -1324 -6360 -1290
rect -6326 -1324 -6292 -1290
rect -6258 -1324 -6224 -1290
rect -6190 -1324 -6156 -1290
rect -6122 -1324 -6088 -1290
rect -6054 -1324 -6020 -1290
rect -5986 -1324 -5952 -1290
rect -5918 -1324 -5884 -1290
rect -5850 -1324 -5816 -1290
rect -5782 -1324 -5748 -1290
rect -5714 -1324 -5680 -1290
rect -5646 -1324 -5612 -1290
rect -5578 -1324 -5544 -1290
rect -5510 -1324 -5476 -1290
rect -5442 -1324 -5408 -1290
rect -5374 -1324 -5340 -1290
rect -5306 -1324 -5272 -1290
rect -5238 -1324 -5204 -1290
rect -5170 -1324 -5136 -1290
rect -5102 -1324 -5068 -1290
rect -5034 -1324 -5000 -1290
rect -4966 -1324 -4932 -1290
rect -4898 -1324 -4864 -1290
rect -4830 -1324 -4796 -1290
rect -4762 -1324 -4728 -1290
rect -4694 -1324 -4660 -1290
rect -4626 -1324 -4592 -1290
rect -4558 -1324 -4524 -1290
rect -4490 -1324 -4456 -1290
rect -4422 -1324 -4388 -1290
rect -4354 -1324 -4320 -1290
rect -4286 -1324 -4252 -1290
rect -4218 -1324 -4184 -1290
rect -4150 -1324 -4116 -1290
rect -4082 -1324 -4048 -1290
rect -4014 -1324 -3980 -1290
rect -3946 -1324 -3912 -1290
rect -3878 -1324 -3844 -1290
rect -3810 -1324 -3776 -1290
rect -3742 -1324 -3708 -1290
rect -3674 -1324 -3640 -1290
rect -3606 -1324 -3572 -1290
rect -3538 -1324 -3504 -1290
rect -3470 -1324 -3436 -1290
rect -3402 -1324 -3368 -1290
rect -3334 -1324 -3300 -1290
rect -3266 -1324 -3232 -1290
rect -3198 -1324 -3164 -1290
rect -3130 -1324 -3096 -1290
rect -3062 -1324 -3028 -1290
rect -2994 -1324 -2960 -1290
rect -2926 -1324 -2892 -1290
rect -2858 -1324 -2824 -1290
rect -2790 -1324 -2756 -1290
rect -2722 -1324 -2688 -1290
rect -2654 -1324 -2620 -1290
rect -2586 -1324 -2552 -1290
rect -2518 -1324 -2484 -1290
rect -2450 -1324 -2416 -1290
rect -2382 -1324 -2348 -1290
rect -2314 -1324 -2280 -1290
rect -2246 -1324 -2212 -1290
rect -2178 -1324 -2144 -1290
rect -2110 -1324 -2076 -1290
rect -2042 -1324 -2008 -1290
rect -1974 -1324 -1940 -1290
rect -1906 -1324 -1872 -1290
rect -1838 -1324 -1804 -1290
rect -1770 -1324 -1736 -1290
rect -1702 -1324 -1668 -1290
rect -1634 -1324 -1600 -1290
rect -1566 -1324 -1532 -1290
rect -1498 -1324 -1464 -1290
rect -1430 -1324 -1396 -1290
rect -1362 -1324 -1328 -1290
rect -1294 -1324 -1260 -1290
rect -1226 -1324 -1192 -1290
rect -1158 -1324 -1124 -1290
rect -1090 -1324 -1056 -1290
rect -1022 -1324 -988 -1290
rect -954 -1324 -920 -1290
rect -886 -1324 -852 -1290
rect -818 -1324 -784 -1290
rect -750 -1324 -716 -1290
rect -682 -1324 -648 -1290
rect -614 -1324 -580 -1290
rect -546 -1324 -512 -1290
rect -478 -1324 -444 -1290
rect -410 -1324 -376 -1290
rect -342 -1324 -308 -1290
rect -274 -1324 -240 -1290
rect -206 -1324 -172 -1290
rect -138 -1324 -104 -1290
rect -70 -1324 -36 -1290
rect -2 -1324 32 -1290
rect 66 -1324 100 -1290
rect 134 -1324 168 -1290
rect 202 -1324 236 -1290
rect 270 -1324 304 -1290
rect 338 -1324 372 -1290
rect 406 -1324 440 -1290
rect 474 -1324 508 -1290
rect 542 -1324 576 -1290
rect 610 -1324 644 -1290
rect 678 -1324 712 -1290
rect 746 -1324 780 -1290
rect 814 -1324 848 -1290
rect 882 -1324 916 -1290
rect 950 -1324 984 -1290
rect 1018 -1324 1052 -1290
rect 1086 -1324 1120 -1290
rect 1154 -1324 1188 -1290
rect 1222 -1324 1256 -1290
rect 1290 -1324 1324 -1290
rect 1358 -1324 1392 -1290
rect 1426 -1324 1460 -1290
rect 1494 -1324 1528 -1290
rect 1562 -1324 1596 -1290
rect 1630 -1324 1664 -1290
rect 1698 -1324 1732 -1290
rect 1766 -1324 1800 -1290
rect 1834 -1324 1868 -1290
rect 1902 -1324 1936 -1290
rect 1970 -1324 2004 -1290
rect 2038 -1324 2072 -1290
rect 2106 -1324 2140 -1290
rect 2174 -1324 2208 -1290
rect 2242 -1324 2276 -1290
rect 2310 -1324 2344 -1290
rect 2378 -1324 2412 -1290
rect 2446 -1324 2480 -1290
rect 2514 -1324 2548 -1290
rect 2582 -1324 2616 -1290
rect 2650 -1324 2684 -1290
rect 2718 -1324 2752 -1290
rect 2786 -1324 2820 -1290
rect 2854 -1324 2888 -1290
rect 2922 -1324 2956 -1290
rect 2990 -1324 3024 -1290
rect 3058 -1324 3092 -1290
rect 3126 -1324 3160 -1290
rect 3194 -1324 3228 -1290
rect 3262 -1324 3296 -1290
rect -7576 -1573 -7542 -1539
rect -7576 -1641 -7542 -1607
rect -7576 -1709 -7542 -1675
rect -7576 -1777 -7542 -1743
rect -7576 -1845 -7542 -1811
rect -7576 -1913 -7542 -1879
rect -7576 -1981 -7542 -1947
rect -7576 -2049 -7542 -2015
rect -7576 -2117 -7542 -2083
rect -7576 -2185 -7542 -2151
rect -7576 -2253 -7542 -2219
rect -7576 -2321 -7542 -2287
rect -7576 -2389 -7542 -2355
rect -7576 -2457 -7542 -2423
rect -7576 -2525 -7542 -2491
rect -7576 -2593 -7542 -2559
rect -7576 -2661 -7542 -2627
rect -7576 -2729 -7542 -2695
rect -7576 -2797 -7542 -2763
rect -7576 -2865 -7542 -2831
rect -7576 -2933 -7542 -2899
rect -7576 -3001 -7542 -2967
rect -7576 -3069 -7542 -3035
rect -7576 -3137 -7542 -3103
rect -7576 -3205 -7542 -3171
rect -7576 -3273 -7542 -3239
rect -7576 -3341 -7542 -3307
rect -7576 -3409 -7542 -3375
rect -7576 -3477 -7542 -3443
rect -7576 -3545 -7542 -3511
rect -7576 -3613 -7542 -3579
rect -7576 -3681 -7542 -3647
rect -7576 -3749 -7542 -3715
rect -7576 -3817 -7542 -3783
rect -7576 -3885 -7542 -3851
rect -7576 -3953 -7542 -3919
rect -7576 -4021 -7542 -3987
rect -7576 -4089 -7542 -4055
rect -7576 -4157 -7542 -4123
rect -7576 -4225 -7542 -4191
rect -7576 -4293 -7542 -4259
rect -7576 -4361 -7542 -4327
rect -7576 -4429 -7542 -4395
rect -7576 -4497 -7542 -4463
rect -7576 -4565 -7542 -4531
rect -7576 -4633 -7542 -4599
rect -7576 -4701 -7542 -4667
rect -7576 -4769 -7542 -4735
rect -7576 -4837 -7542 -4803
rect -7576 -4905 -7542 -4871
rect -7576 -4973 -7542 -4939
rect -7576 -5041 -7542 -5007
rect -7576 -5109 -7542 -5075
rect -7576 -5177 -7542 -5143
rect -7576 -5245 -7542 -5211
rect -7576 -5313 -7542 -5279
rect -7576 -5381 -7542 -5347
rect -7576 -5449 -7542 -5415
rect -7576 -5517 -7542 -5483
rect -7576 -5585 -7542 -5551
rect -7576 -5653 -7542 -5619
rect -7576 -5721 -7542 -5687
rect -7576 -5789 -7542 -5755
rect -7576 -5857 -7542 -5823
rect -7576 -5925 -7542 -5891
rect -7576 -5993 -7542 -5959
rect -7576 -6061 -7542 -6027
rect -7576 -6129 -7542 -6095
rect -7576 -6197 -7542 -6163
rect -7576 -6265 -7542 -6231
rect -7576 -6333 -7542 -6299
rect -7576 -6401 -7542 -6367
rect -7576 -6469 -7542 -6435
rect -7576 -6537 -7542 -6503
rect -7576 -6605 -7542 -6571
rect -7576 -6673 -7542 -6639
rect -7576 -6741 -7542 -6707
rect -7576 -6809 -7542 -6775
rect -7576 -6877 -7542 -6843
rect -7576 -6945 -7542 -6911
rect 3639 -1586 3673 -1552
rect 3639 -1654 3673 -1620
rect 3639 -1722 3673 -1688
rect 3639 -1790 3673 -1756
rect 3639 -1858 3673 -1824
rect 3639 -1926 3673 -1892
rect 3639 -1994 3673 -1960
rect 3639 -2062 3673 -2028
rect 3639 -2130 3673 -2096
rect 3639 -2198 3673 -2164
rect 3639 -2266 3673 -2232
rect 3639 -2334 3673 -2300
rect 3639 -2402 3673 -2368
rect 3639 -2470 3673 -2436
rect 3639 -2538 3673 -2504
rect 3639 -2606 3673 -2572
rect 3639 -2674 3673 -2640
rect 3639 -2742 3673 -2708
rect 3639 -2810 3673 -2776
rect 3639 -2878 3673 -2844
rect 3639 -2946 3673 -2912
rect 3639 -3014 3673 -2980
rect 3639 -3082 3673 -3048
rect 3639 -3150 3673 -3116
rect 3639 -3218 3673 -3184
rect 3639 -3286 3673 -3252
rect 3639 -3354 3673 -3320
rect 3639 -3422 3673 -3388
rect 3639 -3490 3673 -3456
rect 3639 -3558 3673 -3524
rect 3639 -3626 3673 -3592
rect 3639 -3694 3673 -3660
rect 3639 -3762 3673 -3728
rect 3639 -3830 3673 -3796
rect 3639 -3898 3673 -3864
rect 3639 -3966 3673 -3932
rect 3639 -4034 3673 -4000
rect 3639 -4102 3673 -4068
rect 3639 -4170 3673 -4136
rect 3639 -4238 3673 -4204
rect 3639 -4306 3673 -4272
rect 3639 -4374 3673 -4340
rect 3639 -4442 3673 -4408
rect 3639 -4510 3673 -4476
rect 3639 -4578 3673 -4544
rect 3639 -4646 3673 -4612
rect 3639 -4714 3673 -4680
rect 3639 -4782 3673 -4748
rect 3639 -4850 3673 -4816
rect 3639 -4918 3673 -4884
rect 3639 -4986 3673 -4952
rect 3639 -5054 3673 -5020
rect 3639 -5122 3673 -5088
rect 3639 -5190 3673 -5156
rect 3639 -5258 3673 -5224
rect 3639 -5326 3673 -5292
rect 3639 -5394 3673 -5360
rect 3639 -5462 3673 -5428
rect 3639 -5530 3673 -5496
rect 3639 -5598 3673 -5564
rect 3639 -5666 3673 -5632
rect 3639 -5734 3673 -5700
rect 3639 -5802 3673 -5768
rect 3639 -5870 3673 -5836
rect 3639 -5938 3673 -5904
rect 3639 -6006 3673 -5972
rect 3639 -6074 3673 -6040
rect 3639 -6142 3673 -6108
rect 3639 -6210 3673 -6176
rect 3639 -6278 3673 -6244
rect 3639 -6346 3673 -6312
rect 3639 -6414 3673 -6380
rect 3639 -6482 3673 -6448
rect 3639 -6550 3673 -6516
rect 3639 -6618 3673 -6584
rect 3639 -6686 3673 -6652
rect 3639 -6754 3673 -6720
rect 3639 -6822 3673 -6788
rect 3639 -6890 3673 -6856
rect 3639 -6958 3673 -6924
rect -7249 -7204 -7215 -7170
rect -7181 -7204 -7147 -7170
rect -7113 -7204 -7079 -7170
rect -7045 -7204 -7011 -7170
rect -6977 -7204 -6943 -7170
rect -6909 -7204 -6875 -7170
rect -6841 -7204 -6807 -7170
rect -6773 -7204 -6739 -7170
rect -6705 -7204 -6671 -7170
rect -6637 -7204 -6603 -7170
rect -6569 -7204 -6535 -7170
rect -6501 -7204 -6467 -7170
rect -6433 -7204 -6399 -7170
rect -6365 -7204 -6331 -7170
rect -6297 -7204 -6263 -7170
rect -6229 -7204 -6195 -7170
rect -6161 -7204 -6127 -7170
rect -6093 -7204 -6059 -7170
rect -6025 -7204 -5991 -7170
rect -5957 -7204 -5923 -7170
rect -5889 -7204 -5855 -7170
rect -5821 -7204 -5787 -7170
rect -5753 -7204 -5719 -7170
rect -5685 -7204 -5651 -7170
rect -5617 -7204 -5583 -7170
rect -5549 -7204 -5515 -7170
rect -5481 -7204 -5447 -7170
rect -5413 -7204 -5379 -7170
rect -5345 -7204 -5311 -7170
rect -5277 -7204 -5243 -7170
rect -5209 -7204 -5175 -7170
rect -5141 -7204 -5107 -7170
rect -5073 -7204 -5039 -7170
rect -5005 -7204 -4971 -7170
rect -4937 -7204 -4903 -7170
rect -4869 -7204 -4835 -7170
rect -4801 -7204 -4767 -7170
rect -4733 -7204 -4699 -7170
rect -4665 -7204 -4631 -7170
rect -4597 -7204 -4563 -7170
rect -4529 -7204 -4495 -7170
rect -4461 -7204 -4427 -7170
rect -4393 -7204 -4359 -7170
rect -4325 -7204 -4291 -7170
rect -4257 -7204 -4223 -7170
rect -4189 -7204 -4155 -7170
rect -4121 -7204 -4087 -7170
rect -4053 -7204 -4019 -7170
rect -3985 -7204 -3951 -7170
rect -3917 -7204 -3883 -7170
rect -3849 -7204 -3815 -7170
rect -3781 -7204 -3747 -7170
rect -3713 -7204 -3679 -7170
rect -3645 -7204 -3611 -7170
rect -3577 -7204 -3543 -7170
rect -3509 -7204 -3475 -7170
rect -3441 -7204 -3407 -7170
rect -3373 -7204 -3339 -7170
rect -3305 -7204 -3271 -7170
rect -3237 -7204 -3203 -7170
rect -3169 -7204 -3135 -7170
rect -3101 -7204 -3067 -7170
rect -3033 -7204 -2999 -7170
rect -2965 -7204 -2931 -7170
rect -2897 -7204 -2863 -7170
rect -2829 -7204 -2795 -7170
rect -2761 -7204 -2727 -7170
rect -2693 -7204 -2659 -7170
rect -2625 -7204 -2591 -7170
rect -2557 -7204 -2523 -7170
rect -2489 -7204 -2455 -7170
rect -2421 -7204 -2387 -7170
rect -2353 -7204 -2319 -7170
rect -2285 -7204 -2251 -7170
rect -2217 -7204 -2183 -7170
rect -2149 -7204 -2115 -7170
rect -2081 -7204 -2047 -7170
rect -2013 -7204 -1979 -7170
rect -1945 -7204 -1911 -7170
rect -1877 -7204 -1843 -7170
rect -1809 -7204 -1775 -7170
rect -1741 -7204 -1707 -7170
rect -1673 -7204 -1639 -7170
rect -1605 -7204 -1571 -7170
rect -1537 -7204 -1503 -7170
rect -1469 -7204 -1435 -7170
rect -1401 -7204 -1367 -7170
rect -1333 -7204 -1299 -7170
rect -1265 -7204 -1231 -7170
rect -1197 -7204 -1163 -7170
rect -1129 -7204 -1095 -7170
rect -1061 -7204 -1027 -7170
rect -993 -7204 -959 -7170
rect -925 -7204 -891 -7170
rect -857 -7204 -823 -7170
rect -789 -7204 -755 -7170
rect -721 -7204 -687 -7170
rect -653 -7204 -619 -7170
rect -585 -7204 -551 -7170
rect -517 -7204 -483 -7170
rect -449 -7204 -415 -7170
rect -381 -7204 -347 -7170
rect -313 -7204 -279 -7170
rect -245 -7204 -211 -7170
rect -177 -7204 -143 -7170
rect -109 -7204 -75 -7170
rect -41 -7204 -7 -7170
rect 27 -7204 61 -7170
rect 95 -7204 129 -7170
rect 163 -7204 197 -7170
rect 231 -7204 265 -7170
rect 299 -7204 333 -7170
rect 367 -7204 401 -7170
rect 435 -7204 469 -7170
rect 503 -7204 537 -7170
rect 571 -7204 605 -7170
rect 639 -7204 673 -7170
rect 707 -7204 741 -7170
rect 775 -7204 809 -7170
rect 843 -7204 877 -7170
rect 911 -7204 945 -7170
rect 979 -7204 1013 -7170
rect 1047 -7204 1081 -7170
rect 1115 -7204 1149 -7170
rect 1183 -7204 1217 -7170
rect 1251 -7204 1285 -7170
rect 1319 -7204 1353 -7170
rect 1387 -7204 1421 -7170
rect 1455 -7204 1489 -7170
rect 1523 -7204 1557 -7170
rect 1591 -7204 1625 -7170
rect 1659 -7204 1693 -7170
rect 1727 -7204 1761 -7170
rect 1795 -7204 1829 -7170
rect 1863 -7204 1897 -7170
rect 1931 -7204 1965 -7170
rect 1999 -7204 2033 -7170
rect 2067 -7204 2101 -7170
rect 2135 -7204 2169 -7170
rect 2203 -7204 2237 -7170
rect 2271 -7204 2305 -7170
rect 2339 -7204 2373 -7170
rect 2407 -7204 2441 -7170
rect 2475 -7204 2509 -7170
rect 2543 -7204 2577 -7170
rect 2611 -7204 2645 -7170
rect 2679 -7204 2713 -7170
rect 2747 -7204 2781 -7170
rect 2815 -7204 2849 -7170
rect 2883 -7204 2917 -7170
rect 2951 -7204 2985 -7170
rect 3019 -7204 3053 -7170
rect 3087 -7204 3121 -7170
rect 3155 -7204 3189 -7170
rect 3223 -7204 3257 -7170
rect 3291 -7204 3325 -7170
rect 3359 -7204 3393 -7170
<< locali >>
rect -7606 -1290 3703 -1260
rect -7606 -1324 -7370 -1290
rect -7312 -1324 -7298 -1290
rect -7244 -1324 -7226 -1290
rect -7176 -1324 -7154 -1290
rect -7108 -1324 -7082 -1290
rect -7040 -1324 -7010 -1290
rect -6972 -1324 -6938 -1290
rect -6904 -1324 -6870 -1290
rect -6832 -1324 -6802 -1290
rect -6760 -1324 -6734 -1290
rect -6688 -1324 -6666 -1290
rect -6616 -1324 -6598 -1290
rect -6544 -1324 -6530 -1290
rect -6472 -1324 -6462 -1290
rect -6400 -1324 -6394 -1290
rect -6328 -1324 -6326 -1290
rect -6292 -1324 -6290 -1290
rect -6224 -1324 -6218 -1290
rect -6156 -1324 -6146 -1290
rect -6088 -1324 -6074 -1290
rect -6020 -1324 -6002 -1290
rect -5952 -1324 -5930 -1290
rect -5884 -1324 -5858 -1290
rect -5816 -1324 -5786 -1290
rect -5748 -1324 -5714 -1290
rect -5680 -1324 -5646 -1290
rect -5608 -1324 -5578 -1290
rect -5536 -1324 -5510 -1290
rect -5464 -1324 -5442 -1290
rect -5392 -1324 -5374 -1290
rect -5320 -1324 -5306 -1290
rect -5248 -1324 -5238 -1290
rect -5176 -1324 -5170 -1290
rect -5104 -1324 -5102 -1290
rect -5068 -1324 -5066 -1290
rect -5000 -1324 -4994 -1290
rect -4932 -1324 -4922 -1290
rect -4864 -1324 -4850 -1290
rect -4796 -1324 -4778 -1290
rect -4728 -1324 -4706 -1290
rect -4660 -1324 -4634 -1290
rect -4592 -1324 -4562 -1290
rect -4524 -1324 -4490 -1290
rect -4456 -1324 -4422 -1290
rect -4384 -1324 -4354 -1290
rect -4312 -1324 -4286 -1290
rect -4240 -1324 -4218 -1290
rect -4168 -1324 -4150 -1290
rect -4096 -1324 -4082 -1290
rect -4024 -1324 -4014 -1290
rect -3952 -1324 -3946 -1290
rect -3880 -1324 -3878 -1290
rect -3844 -1324 -3842 -1290
rect -3776 -1324 -3770 -1290
rect -3708 -1324 -3698 -1290
rect -3640 -1324 -3626 -1290
rect -3572 -1324 -3554 -1290
rect -3504 -1324 -3482 -1290
rect -3436 -1324 -3410 -1290
rect -3368 -1324 -3338 -1290
rect -3300 -1324 -3266 -1290
rect -3232 -1324 -3198 -1290
rect -3160 -1324 -3130 -1290
rect -3088 -1324 -3062 -1290
rect -3016 -1324 -2994 -1290
rect -2944 -1324 -2926 -1290
rect -2872 -1324 -2858 -1290
rect -2800 -1324 -2790 -1290
rect -2728 -1324 -2722 -1290
rect -2656 -1324 -2654 -1290
rect -2620 -1324 -2618 -1290
rect -2552 -1324 -2546 -1290
rect -2484 -1324 -2474 -1290
rect -2416 -1324 -2402 -1290
rect -2348 -1324 -2330 -1290
rect -2280 -1324 -2258 -1290
rect -2212 -1324 -2186 -1290
rect -2144 -1324 -2114 -1290
rect -2076 -1324 -2042 -1290
rect -2008 -1324 -1974 -1290
rect -1936 -1324 -1906 -1290
rect -1864 -1324 -1838 -1290
rect -1792 -1324 -1770 -1290
rect -1720 -1324 -1702 -1290
rect -1648 -1324 -1634 -1290
rect -1576 -1324 -1566 -1290
rect -1504 -1324 -1498 -1290
rect -1432 -1324 -1430 -1290
rect -1396 -1324 -1394 -1290
rect -1328 -1324 -1322 -1290
rect -1260 -1324 -1250 -1290
rect -1192 -1324 -1178 -1290
rect -1124 -1324 -1106 -1290
rect -1056 -1324 -1034 -1290
rect -988 -1324 -962 -1290
rect -920 -1324 -890 -1290
rect -852 -1324 -818 -1290
rect -784 -1324 -750 -1290
rect -712 -1324 -682 -1290
rect -640 -1324 -614 -1290
rect -568 -1324 -546 -1290
rect -496 -1324 -478 -1290
rect -424 -1324 -410 -1290
rect -352 -1324 -342 -1290
rect -280 -1324 -274 -1290
rect -208 -1324 -206 -1290
rect -172 -1324 -170 -1290
rect -104 -1324 -98 -1290
rect -36 -1324 -26 -1290
rect 32 -1324 46 -1290
rect 100 -1324 118 -1290
rect 168 -1324 190 -1290
rect 236 -1324 262 -1290
rect 304 -1324 334 -1290
rect 372 -1324 406 -1290
rect 440 -1324 474 -1290
rect 512 -1324 542 -1290
rect 584 -1324 610 -1290
rect 656 -1324 678 -1290
rect 728 -1324 746 -1290
rect 800 -1324 814 -1290
rect 872 -1324 882 -1290
rect 944 -1324 950 -1290
rect 1016 -1324 1018 -1290
rect 1052 -1324 1054 -1290
rect 1120 -1324 1126 -1290
rect 1188 -1324 1198 -1290
rect 1256 -1324 1270 -1290
rect 1324 -1324 1342 -1290
rect 1392 -1324 1414 -1290
rect 1460 -1324 1486 -1290
rect 1528 -1324 1558 -1290
rect 1596 -1324 1630 -1290
rect 1664 -1324 1698 -1290
rect 1736 -1324 1766 -1290
rect 1808 -1324 1834 -1290
rect 1880 -1324 1902 -1290
rect 1952 -1324 1970 -1290
rect 2024 -1324 2038 -1290
rect 2096 -1324 2106 -1290
rect 2168 -1324 2174 -1290
rect 2240 -1324 2242 -1290
rect 2276 -1324 2278 -1290
rect 2344 -1324 2350 -1290
rect 2412 -1324 2422 -1290
rect 2480 -1324 2494 -1290
rect 2548 -1324 2566 -1290
rect 2616 -1324 2638 -1290
rect 2684 -1324 2710 -1290
rect 2752 -1324 2782 -1290
rect 2820 -1324 2854 -1290
rect 2888 -1324 2922 -1290
rect 2960 -1324 2990 -1290
rect 3032 -1324 3058 -1290
rect 3104 -1324 3126 -1290
rect 3176 -1324 3194 -1290
rect 3248 -1324 3262 -1290
rect 3320 -1324 3703 -1290
rect -7606 -1353 3703 -1324
rect -7605 -1539 -7512 -1353
rect -7605 -1573 -7576 -1539
rect -7542 -1573 -7512 -1539
rect -7605 -1607 -7512 -1573
rect -7605 -1641 -7576 -1607
rect -7542 -1641 -7512 -1607
rect -7605 -1675 -7512 -1641
rect -7605 -1709 -7576 -1675
rect -7542 -1709 -7512 -1675
rect -7605 -1743 -7512 -1709
rect -7605 -1777 -7576 -1743
rect -7542 -1777 -7512 -1743
rect -7605 -1811 -7512 -1777
rect -7605 -1845 -7576 -1811
rect -7542 -1845 -7512 -1811
rect -7605 -1879 -7512 -1845
rect -7605 -1913 -7576 -1879
rect -7542 -1913 -7512 -1879
rect -7605 -1947 -7512 -1913
rect -7605 -1981 -7576 -1947
rect -7542 -1981 -7512 -1947
rect -7605 -2015 -7512 -1981
rect -7605 -2049 -7576 -2015
rect -7542 -2049 -7512 -2015
rect -7605 -2083 -7512 -2049
rect -7605 -2117 -7576 -2083
rect -7542 -2117 -7512 -2083
rect -7605 -2151 -7512 -2117
rect -7605 -2185 -7576 -2151
rect -7542 -2185 -7512 -2151
rect -7605 -2219 -7512 -2185
rect -7605 -2253 -7576 -2219
rect -7542 -2253 -7512 -2219
rect -7605 -2287 -7512 -2253
rect -7605 -2321 -7576 -2287
rect -7542 -2321 -7512 -2287
rect -7605 -2355 -7512 -2321
rect -7605 -2389 -7576 -2355
rect -7542 -2389 -7512 -2355
rect -7605 -2423 -7512 -2389
rect -7605 -2457 -7576 -2423
rect -7542 -2457 -7512 -2423
rect -7605 -2491 -7512 -2457
rect -7605 -2525 -7576 -2491
rect -7542 -2525 -7512 -2491
rect -7605 -2559 -7512 -2525
rect -7605 -2593 -7576 -2559
rect -7542 -2593 -7512 -2559
rect -7605 -2627 -7512 -2593
rect -7605 -2661 -7576 -2627
rect -7542 -2661 -7512 -2627
rect -7605 -2695 -7512 -2661
rect -7605 -2729 -7576 -2695
rect -7542 -2729 -7512 -2695
rect -7605 -2763 -7512 -2729
rect -7605 -2797 -7576 -2763
rect -7542 -2797 -7512 -2763
rect -7605 -2831 -7512 -2797
rect -7605 -2865 -7576 -2831
rect -7542 -2865 -7512 -2831
rect -7605 -2899 -7512 -2865
rect -7605 -2933 -7576 -2899
rect -7542 -2933 -7512 -2899
rect -7605 -2967 -7512 -2933
rect -7605 -3001 -7576 -2967
rect -7542 -3001 -7512 -2967
rect -7605 -3035 -7512 -3001
rect -7605 -3069 -7576 -3035
rect -7542 -3069 -7512 -3035
rect -7605 -3103 -7512 -3069
rect -7605 -3137 -7576 -3103
rect -7542 -3137 -7512 -3103
rect -7605 -3171 -7512 -3137
rect -7605 -3205 -7576 -3171
rect -7542 -3205 -7512 -3171
rect -7605 -3239 -7512 -3205
rect -7605 -3273 -7576 -3239
rect -7542 -3273 -7512 -3239
rect -7605 -3307 -7512 -3273
rect -7605 -3341 -7576 -3307
rect -7542 -3341 -7512 -3307
rect -7605 -3375 -7512 -3341
rect -7605 -3409 -7576 -3375
rect -7542 -3409 -7512 -3375
rect -7605 -3443 -7512 -3409
rect -7605 -3477 -7576 -3443
rect -7542 -3477 -7512 -3443
rect -7605 -3511 -7512 -3477
rect -7605 -3545 -7576 -3511
rect -7542 -3545 -7512 -3511
rect -7605 -3579 -7512 -3545
rect -7605 -3613 -7576 -3579
rect -7542 -3613 -7512 -3579
rect -7605 -3647 -7512 -3613
rect -7605 -3681 -7576 -3647
rect -7542 -3681 -7512 -3647
rect -7605 -3715 -7512 -3681
rect -7605 -3749 -7576 -3715
rect -7542 -3749 -7512 -3715
rect -7605 -3783 -7512 -3749
rect -7605 -3817 -7576 -3783
rect -7542 -3817 -7512 -3783
rect -7605 -3851 -7512 -3817
rect -7605 -3885 -7576 -3851
rect -7542 -3885 -7512 -3851
rect -7605 -3919 -7512 -3885
rect -7605 -3953 -7576 -3919
rect -7542 -3953 -7512 -3919
rect -7605 -3987 -7512 -3953
rect -7605 -4021 -7576 -3987
rect -7542 -4021 -7512 -3987
rect -7605 -4055 -7512 -4021
rect -7605 -4089 -7576 -4055
rect -7542 -4089 -7512 -4055
rect -7605 -4123 -7512 -4089
rect -7605 -4157 -7576 -4123
rect -7542 -4157 -7512 -4123
rect -7605 -4191 -7512 -4157
rect -7605 -4225 -7576 -4191
rect -7542 -4225 -7512 -4191
rect -7605 -4259 -7512 -4225
rect -7605 -4293 -7576 -4259
rect -7542 -4293 -7512 -4259
rect -7605 -4327 -7512 -4293
rect -7605 -4361 -7576 -4327
rect -7542 -4361 -7512 -4327
rect -7605 -4395 -7512 -4361
rect -7605 -4429 -7576 -4395
rect -7542 -4429 -7512 -4395
rect -7605 -4463 -7512 -4429
rect -7605 -4497 -7576 -4463
rect -7542 -4497 -7512 -4463
rect -7605 -4531 -7512 -4497
rect -7605 -4565 -7576 -4531
rect -7542 -4565 -7512 -4531
rect -7605 -4599 -7512 -4565
rect -7605 -4633 -7576 -4599
rect -7542 -4633 -7512 -4599
rect -7605 -4667 -7512 -4633
rect -7605 -4701 -7576 -4667
rect -7542 -4701 -7512 -4667
rect -7605 -4735 -7512 -4701
rect -7605 -4769 -7576 -4735
rect -7542 -4769 -7512 -4735
rect -7605 -4803 -7512 -4769
rect -7605 -4837 -7576 -4803
rect -7542 -4837 -7512 -4803
rect -7605 -4871 -7512 -4837
rect -7605 -4905 -7576 -4871
rect -7542 -4905 -7512 -4871
rect -7605 -4939 -7512 -4905
rect -7605 -4973 -7576 -4939
rect -7542 -4973 -7512 -4939
rect -7605 -5007 -7512 -4973
rect -7605 -5041 -7576 -5007
rect -7542 -5041 -7512 -5007
rect -7605 -5075 -7512 -5041
rect -7605 -5109 -7576 -5075
rect -7542 -5109 -7512 -5075
rect -7605 -5143 -7512 -5109
rect -7605 -5177 -7576 -5143
rect -7542 -5177 -7512 -5143
rect -7605 -5211 -7512 -5177
rect -7605 -5245 -7576 -5211
rect -7542 -5245 -7512 -5211
rect -7605 -5279 -7512 -5245
rect -7605 -5313 -7576 -5279
rect -7542 -5313 -7512 -5279
rect -7605 -5347 -7512 -5313
rect -7605 -5381 -7576 -5347
rect -7542 -5381 -7512 -5347
rect -7605 -5415 -7512 -5381
rect -7605 -5449 -7576 -5415
rect -7542 -5449 -7512 -5415
rect -7605 -5483 -7512 -5449
rect -7605 -5517 -7576 -5483
rect -7542 -5517 -7512 -5483
rect -7605 -5551 -7512 -5517
rect -7605 -5585 -7576 -5551
rect -7542 -5585 -7512 -5551
rect -7605 -5619 -7512 -5585
rect -7605 -5653 -7576 -5619
rect -7542 -5653 -7512 -5619
rect -7605 -5687 -7512 -5653
rect -7605 -5721 -7576 -5687
rect -7542 -5721 -7512 -5687
rect -7605 -5755 -7512 -5721
rect -7605 -5789 -7576 -5755
rect -7542 -5789 -7512 -5755
rect -7605 -5823 -7512 -5789
rect -7605 -5857 -7576 -5823
rect -7542 -5857 -7512 -5823
rect -7605 -5891 -7512 -5857
rect -7605 -5925 -7576 -5891
rect -7542 -5925 -7512 -5891
rect -7605 -5959 -7512 -5925
rect -7605 -5993 -7576 -5959
rect -7542 -5993 -7512 -5959
rect -7605 -6027 -7512 -5993
rect -7605 -6061 -7576 -6027
rect -7542 -6061 -7512 -6027
rect -7605 -6095 -7512 -6061
rect -7605 -6129 -7576 -6095
rect -7542 -6129 -7512 -6095
rect -7605 -6163 -7512 -6129
rect -7605 -6197 -7576 -6163
rect -7542 -6197 -7512 -6163
rect -7605 -6231 -7512 -6197
rect -7605 -6265 -7576 -6231
rect -7542 -6265 -7512 -6231
rect -7605 -6299 -7512 -6265
rect -7605 -6333 -7576 -6299
rect -7542 -6333 -7512 -6299
rect -7605 -6367 -7512 -6333
rect -7605 -6401 -7576 -6367
rect -7542 -6401 -7512 -6367
rect -7605 -6435 -7512 -6401
rect -7605 -6469 -7576 -6435
rect -7542 -6469 -7512 -6435
rect -7605 -6503 -7512 -6469
rect -7605 -6537 -7576 -6503
rect -7542 -6537 -7512 -6503
rect -7605 -6571 -7512 -6537
rect -7605 -6605 -7576 -6571
rect -7542 -6605 -7512 -6571
rect -7605 -6639 -7512 -6605
rect -7605 -6673 -7576 -6639
rect -7542 -6673 -7512 -6639
rect -7605 -6707 -7512 -6673
rect -7605 -6741 -7576 -6707
rect -7542 -6741 -7512 -6707
rect -7605 -6775 -7512 -6741
rect -7605 -6809 -7576 -6775
rect -7542 -6809 -7512 -6775
rect -7605 -6843 -7512 -6809
rect -7605 -6877 -7576 -6843
rect -7542 -6877 -7512 -6843
rect -7605 -6911 -7512 -6877
rect -7605 -6945 -7576 -6911
rect -7542 -6945 -7512 -6911
rect -7605 -7140 -7512 -6945
rect 3610 -1552 3703 -1353
rect 3610 -1586 3639 -1552
rect 3673 -1586 3703 -1552
rect 3610 -1620 3703 -1586
rect 3610 -1654 3639 -1620
rect 3673 -1654 3703 -1620
rect 3610 -1688 3703 -1654
rect 3610 -1722 3639 -1688
rect 3673 -1722 3703 -1688
rect 3610 -1756 3703 -1722
rect 3610 -1790 3639 -1756
rect 3673 -1790 3703 -1756
rect 3610 -1824 3703 -1790
rect 3610 -1858 3639 -1824
rect 3673 -1858 3703 -1824
rect 3610 -1892 3703 -1858
rect 3610 -1926 3639 -1892
rect 3673 -1926 3703 -1892
rect 3610 -1960 3703 -1926
rect 3610 -1994 3639 -1960
rect 3673 -1994 3703 -1960
rect 3610 -2028 3703 -1994
rect 3610 -2062 3639 -2028
rect 3673 -2062 3703 -2028
rect 3610 -2096 3703 -2062
rect 3610 -2130 3639 -2096
rect 3673 -2130 3703 -2096
rect 3610 -2164 3703 -2130
rect 3610 -2198 3639 -2164
rect 3673 -2198 3703 -2164
rect 3610 -2232 3703 -2198
rect 3610 -2266 3639 -2232
rect 3673 -2266 3703 -2232
rect 3610 -2300 3703 -2266
rect 3610 -2334 3639 -2300
rect 3673 -2334 3703 -2300
rect 3610 -2368 3703 -2334
rect 3610 -2402 3639 -2368
rect 3673 -2402 3703 -2368
rect 3610 -2436 3703 -2402
rect 3610 -2470 3639 -2436
rect 3673 -2470 3703 -2436
rect 3610 -2504 3703 -2470
rect 3610 -2538 3639 -2504
rect 3673 -2538 3703 -2504
rect 3610 -2572 3703 -2538
rect 3610 -2606 3639 -2572
rect 3673 -2606 3703 -2572
rect 3610 -2640 3703 -2606
rect 3610 -2674 3639 -2640
rect 3673 -2674 3703 -2640
rect 3610 -2708 3703 -2674
rect 3610 -2742 3639 -2708
rect 3673 -2742 3703 -2708
rect 3610 -2776 3703 -2742
rect 3610 -2810 3639 -2776
rect 3673 -2810 3703 -2776
rect 3610 -2844 3703 -2810
rect 3610 -2878 3639 -2844
rect 3673 -2878 3703 -2844
rect 3610 -2912 3703 -2878
rect 3610 -2946 3639 -2912
rect 3673 -2946 3703 -2912
rect 3610 -2980 3703 -2946
rect 3610 -3014 3639 -2980
rect 3673 -3014 3703 -2980
rect 3610 -3048 3703 -3014
rect 3610 -3082 3639 -3048
rect 3673 -3082 3703 -3048
rect 3610 -3116 3703 -3082
rect 3610 -3150 3639 -3116
rect 3673 -3150 3703 -3116
rect 3610 -3184 3703 -3150
rect 3610 -3218 3639 -3184
rect 3673 -3218 3703 -3184
rect 3610 -3252 3703 -3218
rect 3610 -3286 3639 -3252
rect 3673 -3286 3703 -3252
rect 3610 -3320 3703 -3286
rect 3610 -3354 3639 -3320
rect 3673 -3354 3703 -3320
rect 3610 -3388 3703 -3354
rect 3610 -3422 3639 -3388
rect 3673 -3422 3703 -3388
rect 3610 -3456 3703 -3422
rect 3610 -3490 3639 -3456
rect 3673 -3490 3703 -3456
rect 3610 -3524 3703 -3490
rect 3610 -3558 3639 -3524
rect 3673 -3558 3703 -3524
rect 3610 -3592 3703 -3558
rect 3610 -3626 3639 -3592
rect 3673 -3626 3703 -3592
rect 3610 -3660 3703 -3626
rect 3610 -3694 3639 -3660
rect 3673 -3694 3703 -3660
rect 3610 -3728 3703 -3694
rect 3610 -3762 3639 -3728
rect 3673 -3762 3703 -3728
rect 3610 -3796 3703 -3762
rect 3610 -3830 3639 -3796
rect 3673 -3830 3703 -3796
rect 3610 -3864 3703 -3830
rect 3610 -3898 3639 -3864
rect 3673 -3898 3703 -3864
rect 3610 -3932 3703 -3898
rect 3610 -3966 3639 -3932
rect 3673 -3966 3703 -3932
rect 3610 -4000 3703 -3966
rect 3610 -4034 3639 -4000
rect 3673 -4034 3703 -4000
rect 3610 -4068 3703 -4034
rect 3610 -4102 3639 -4068
rect 3673 -4102 3703 -4068
rect 3610 -4136 3703 -4102
rect 3610 -4170 3639 -4136
rect 3673 -4170 3703 -4136
rect 3610 -4204 3703 -4170
rect 3610 -4238 3639 -4204
rect 3673 -4238 3703 -4204
rect 3610 -4272 3703 -4238
rect 3610 -4306 3639 -4272
rect 3673 -4306 3703 -4272
rect 3610 -4340 3703 -4306
rect 3610 -4374 3639 -4340
rect 3673 -4374 3703 -4340
rect 3610 -4408 3703 -4374
rect 3610 -4442 3639 -4408
rect 3673 -4442 3703 -4408
rect 3610 -4476 3703 -4442
rect 3610 -4510 3639 -4476
rect 3673 -4510 3703 -4476
rect 3610 -4544 3703 -4510
rect 3610 -4578 3639 -4544
rect 3673 -4578 3703 -4544
rect 3610 -4612 3703 -4578
rect 3610 -4646 3639 -4612
rect 3673 -4646 3703 -4612
rect 3610 -4680 3703 -4646
rect 3610 -4714 3639 -4680
rect 3673 -4714 3703 -4680
rect 3610 -4748 3703 -4714
rect 3610 -4782 3639 -4748
rect 3673 -4782 3703 -4748
rect 3610 -4816 3703 -4782
rect 3610 -4850 3639 -4816
rect 3673 -4850 3703 -4816
rect 3610 -4884 3703 -4850
rect 3610 -4918 3639 -4884
rect 3673 -4918 3703 -4884
rect 3610 -4952 3703 -4918
rect 3610 -4986 3639 -4952
rect 3673 -4986 3703 -4952
rect 3610 -5020 3703 -4986
rect 3610 -5054 3639 -5020
rect 3673 -5054 3703 -5020
rect 3610 -5088 3703 -5054
rect 3610 -5122 3639 -5088
rect 3673 -5122 3703 -5088
rect 3610 -5156 3703 -5122
rect 3610 -5190 3639 -5156
rect 3673 -5190 3703 -5156
rect 3610 -5224 3703 -5190
rect 3610 -5258 3639 -5224
rect 3673 -5258 3703 -5224
rect 3610 -5292 3703 -5258
rect 3610 -5326 3639 -5292
rect 3673 -5326 3703 -5292
rect 3610 -5360 3703 -5326
rect 3610 -5394 3639 -5360
rect 3673 -5394 3703 -5360
rect 3610 -5428 3703 -5394
rect 3610 -5462 3639 -5428
rect 3673 -5462 3703 -5428
rect 3610 -5496 3703 -5462
rect 3610 -5530 3639 -5496
rect 3673 -5530 3703 -5496
rect 3610 -5564 3703 -5530
rect 3610 -5598 3639 -5564
rect 3673 -5598 3703 -5564
rect 3610 -5632 3703 -5598
rect 3610 -5666 3639 -5632
rect 3673 -5666 3703 -5632
rect 3610 -5700 3703 -5666
rect 3610 -5734 3639 -5700
rect 3673 -5734 3703 -5700
rect 3610 -5768 3703 -5734
rect 3610 -5802 3639 -5768
rect 3673 -5802 3703 -5768
rect 3610 -5836 3703 -5802
rect 3610 -5870 3639 -5836
rect 3673 -5870 3703 -5836
rect 3610 -5904 3703 -5870
rect 3610 -5938 3639 -5904
rect 3673 -5938 3703 -5904
rect 3610 -5972 3703 -5938
rect 3610 -6006 3639 -5972
rect 3673 -6006 3703 -5972
rect 3610 -6040 3703 -6006
rect 3610 -6074 3639 -6040
rect 3673 -6074 3703 -6040
rect 3610 -6108 3703 -6074
rect 3610 -6142 3639 -6108
rect 3673 -6142 3703 -6108
rect 3610 -6176 3703 -6142
rect 3610 -6210 3639 -6176
rect 3673 -6210 3703 -6176
rect 3610 -6244 3703 -6210
rect 3610 -6278 3639 -6244
rect 3673 -6278 3703 -6244
rect 3610 -6312 3703 -6278
rect 3610 -6346 3639 -6312
rect 3673 -6346 3703 -6312
rect 3610 -6380 3703 -6346
rect 3610 -6414 3639 -6380
rect 3673 -6414 3703 -6380
rect 3610 -6448 3703 -6414
rect 3610 -6482 3639 -6448
rect 3673 -6482 3703 -6448
rect 3610 -6516 3703 -6482
rect 3610 -6550 3639 -6516
rect 3673 -6550 3703 -6516
rect 3610 -6584 3703 -6550
rect 3610 -6618 3639 -6584
rect 3673 -6618 3703 -6584
rect 3610 -6652 3703 -6618
rect 3610 -6686 3639 -6652
rect 3673 -6686 3703 -6652
rect 3610 -6720 3703 -6686
rect 3610 -6754 3639 -6720
rect 3673 -6754 3703 -6720
rect 3610 -6788 3703 -6754
rect 3610 -6822 3639 -6788
rect 3673 -6822 3703 -6788
rect 3610 -6856 3703 -6822
rect 3610 -6890 3639 -6856
rect 3673 -6890 3703 -6856
rect 3610 -6924 3703 -6890
rect 3610 -6958 3639 -6924
rect 3673 -6958 3703 -6924
rect 3610 -7140 3703 -6958
rect -7605 -7170 3703 -7140
rect -7605 -7204 -7249 -7170
rect -7215 -7204 -7181 -7170
rect -7147 -7204 -7113 -7170
rect -7079 -7204 -7045 -7170
rect -7011 -7204 -6977 -7170
rect -6943 -7204 -6909 -7170
rect -6875 -7204 -6841 -7170
rect -6807 -7204 -6773 -7170
rect -6739 -7204 -6705 -7170
rect -6671 -7204 -6637 -7170
rect -6603 -7204 -6569 -7170
rect -6535 -7204 -6501 -7170
rect -6467 -7204 -6433 -7170
rect -6399 -7204 -6365 -7170
rect -6331 -7204 -6297 -7170
rect -6263 -7204 -6229 -7170
rect -6195 -7204 -6161 -7170
rect -6127 -7204 -6093 -7170
rect -6059 -7204 -6025 -7170
rect -5991 -7204 -5957 -7170
rect -5923 -7204 -5889 -7170
rect -5855 -7204 -5821 -7170
rect -5787 -7204 -5753 -7170
rect -5719 -7204 -5685 -7170
rect -5651 -7204 -5617 -7170
rect -5583 -7204 -5549 -7170
rect -5515 -7204 -5481 -7170
rect -5447 -7204 -5413 -7170
rect -5379 -7204 -5345 -7170
rect -5311 -7204 -5277 -7170
rect -5243 -7204 -5209 -7170
rect -5175 -7204 -5141 -7170
rect -5107 -7204 -5073 -7170
rect -5039 -7204 -5005 -7170
rect -4971 -7204 -4937 -7170
rect -4903 -7204 -4869 -7170
rect -4835 -7204 -4801 -7170
rect -4767 -7204 -4733 -7170
rect -4699 -7204 -4665 -7170
rect -4631 -7204 -4597 -7170
rect -4563 -7204 -4529 -7170
rect -4495 -7204 -4461 -7170
rect -4427 -7204 -4393 -7170
rect -4359 -7204 -4325 -7170
rect -4291 -7204 -4257 -7170
rect -4223 -7204 -4189 -7170
rect -4155 -7204 -4121 -7170
rect -4087 -7204 -4053 -7170
rect -4019 -7204 -3985 -7170
rect -3951 -7204 -3917 -7170
rect -3883 -7204 -3849 -7170
rect -3815 -7204 -3781 -7170
rect -3747 -7204 -3713 -7170
rect -3679 -7204 -3645 -7170
rect -3611 -7204 -3577 -7170
rect -3543 -7204 -3509 -7170
rect -3475 -7204 -3441 -7170
rect -3407 -7204 -3373 -7170
rect -3339 -7204 -3305 -7170
rect -3271 -7204 -3237 -7170
rect -3203 -7204 -3169 -7170
rect -3135 -7204 -3101 -7170
rect -3067 -7204 -3033 -7170
rect -2999 -7204 -2965 -7170
rect -2931 -7204 -2897 -7170
rect -2863 -7204 -2829 -7170
rect -2795 -7204 -2761 -7170
rect -2727 -7204 -2693 -7170
rect -2659 -7204 -2625 -7170
rect -2591 -7204 -2557 -7170
rect -2523 -7204 -2489 -7170
rect -2455 -7204 -2421 -7170
rect -2387 -7204 -2353 -7170
rect -2319 -7204 -2285 -7170
rect -2251 -7204 -2217 -7170
rect -2183 -7204 -2149 -7170
rect -2115 -7204 -2081 -7170
rect -2047 -7204 -2013 -7170
rect -1979 -7204 -1945 -7170
rect -1911 -7204 -1877 -7170
rect -1843 -7204 -1809 -7170
rect -1775 -7204 -1741 -7170
rect -1707 -7204 -1673 -7170
rect -1639 -7204 -1605 -7170
rect -1571 -7204 -1537 -7170
rect -1503 -7204 -1469 -7170
rect -1435 -7204 -1401 -7170
rect -1367 -7204 -1333 -7170
rect -1299 -7204 -1265 -7170
rect -1231 -7204 -1197 -7170
rect -1163 -7204 -1129 -7170
rect -1095 -7204 -1061 -7170
rect -1027 -7204 -993 -7170
rect -959 -7204 -925 -7170
rect -891 -7204 -857 -7170
rect -823 -7204 -789 -7170
rect -755 -7204 -721 -7170
rect -687 -7204 -653 -7170
rect -619 -7204 -585 -7170
rect -551 -7204 -517 -7170
rect -483 -7204 -449 -7170
rect -415 -7204 -381 -7170
rect -347 -7204 -313 -7170
rect -279 -7204 -245 -7170
rect -211 -7204 -177 -7170
rect -143 -7204 -109 -7170
rect -75 -7204 -41 -7170
rect -7 -7204 27 -7170
rect 61 -7204 95 -7170
rect 129 -7204 163 -7170
rect 197 -7204 231 -7170
rect 265 -7204 299 -7170
rect 333 -7204 367 -7170
rect 401 -7204 435 -7170
rect 469 -7204 503 -7170
rect 537 -7204 571 -7170
rect 605 -7204 639 -7170
rect 673 -7204 707 -7170
rect 741 -7204 775 -7170
rect 809 -7204 843 -7170
rect 877 -7204 911 -7170
rect 945 -7204 979 -7170
rect 1013 -7204 1047 -7170
rect 1081 -7204 1115 -7170
rect 1149 -7204 1183 -7170
rect 1217 -7204 1251 -7170
rect 1285 -7204 1319 -7170
rect 1353 -7204 1387 -7170
rect 1421 -7204 1455 -7170
rect 1489 -7204 1523 -7170
rect 1557 -7204 1591 -7170
rect 1625 -7204 1659 -7170
rect 1693 -7204 1727 -7170
rect 1761 -7204 1795 -7170
rect 1829 -7204 1863 -7170
rect 1897 -7204 1931 -7170
rect 1965 -7204 1999 -7170
rect 2033 -7204 2067 -7170
rect 2101 -7204 2135 -7170
rect 2169 -7204 2203 -7170
rect 2237 -7204 2271 -7170
rect 2305 -7204 2339 -7170
rect 2373 -7204 2407 -7170
rect 2441 -7204 2475 -7170
rect 2509 -7204 2543 -7170
rect 2577 -7204 2611 -7170
rect 2645 -7204 2679 -7170
rect 2713 -7204 2747 -7170
rect 2781 -7204 2815 -7170
rect 2849 -7204 2883 -7170
rect 2917 -7204 2951 -7170
rect 2985 -7204 3019 -7170
rect 3053 -7204 3087 -7170
rect 3121 -7204 3155 -7170
rect 3189 -7204 3223 -7170
rect 3257 -7204 3291 -7170
rect 3325 -7204 3359 -7170
rect 3393 -7204 3703 -7170
rect -7605 -7233 3703 -7204
rect -7605 -7554 13719 -7521
rect -7605 -7588 -7264 -7554
rect -7230 -7588 -7196 -7554
rect -7162 -7588 -7128 -7554
rect -7094 -7588 -7060 -7554
rect -7026 -7588 -6992 -7554
rect -6958 -7588 -6924 -7554
rect -6890 -7588 -6856 -7554
rect -6822 -7588 -6788 -7554
rect -6754 -7588 -6720 -7554
rect -6686 -7588 -6652 -7554
rect -6618 -7588 -6584 -7554
rect -6550 -7588 -6516 -7554
rect -6482 -7588 -6448 -7554
rect -6414 -7588 -6380 -7554
rect -6346 -7588 -6312 -7554
rect -6278 -7588 -6244 -7554
rect -6210 -7588 -6176 -7554
rect -6142 -7588 -6108 -7554
rect -6074 -7588 -6040 -7554
rect -6006 -7588 -5972 -7554
rect -5938 -7588 -5904 -7554
rect -5870 -7588 -5836 -7554
rect -5802 -7588 -5768 -7554
rect -5734 -7588 -5700 -7554
rect -5666 -7588 -5632 -7554
rect -5598 -7588 -5564 -7554
rect -5530 -7588 -5496 -7554
rect -5462 -7588 -5428 -7554
rect -5394 -7588 -5360 -7554
rect -5326 -7588 -5292 -7554
rect -5258 -7588 -5224 -7554
rect -5190 -7588 -5156 -7554
rect -5122 -7588 -5088 -7554
rect -5054 -7588 -5020 -7554
rect -4986 -7588 -4952 -7554
rect -4918 -7588 -4884 -7554
rect -4850 -7588 -4816 -7554
rect -4782 -7588 -4748 -7554
rect -4714 -7588 -4680 -7554
rect -4646 -7588 -4612 -7554
rect -4578 -7588 -4544 -7554
rect -4510 -7588 -4476 -7554
rect -4442 -7588 -4408 -7554
rect -4374 -7588 -4340 -7554
rect -4306 -7588 -4272 -7554
rect -4238 -7588 -4204 -7554
rect -4170 -7588 -4136 -7554
rect -4102 -7588 -4068 -7554
rect -4034 -7588 -4000 -7554
rect -3966 -7588 -3932 -7554
rect -3898 -7588 -3864 -7554
rect -3830 -7588 -3796 -7554
rect -3762 -7588 -3728 -7554
rect -3694 -7588 -3660 -7554
rect -3626 -7588 -3592 -7554
rect -3558 -7588 -3524 -7554
rect -3490 -7588 -3456 -7554
rect -3422 -7588 -3388 -7554
rect -3354 -7588 -3320 -7554
rect -3286 -7588 -3252 -7554
rect -3218 -7588 -3184 -7554
rect -3150 -7588 -3116 -7554
rect -3082 -7588 -3048 -7554
rect -3014 -7588 -2980 -7554
rect -2946 -7588 -2912 -7554
rect -2878 -7588 -2844 -7554
rect -2810 -7588 -2776 -7554
rect -2742 -7588 -2708 -7554
rect -2674 -7588 -2640 -7554
rect -2606 -7588 -2572 -7554
rect -2538 -7588 -2504 -7554
rect -2470 -7588 -2436 -7554
rect -2402 -7588 -2368 -7554
rect -2334 -7588 -2300 -7554
rect -2266 -7588 -2232 -7554
rect -2198 -7588 -2164 -7554
rect -2130 -7588 -2096 -7554
rect -2062 -7588 -2028 -7554
rect -1994 -7588 -1960 -7554
rect -1926 -7588 -1892 -7554
rect -1858 -7588 -1824 -7554
rect -1790 -7588 -1756 -7554
rect -1722 -7588 -1688 -7554
rect -1654 -7588 -1620 -7554
rect -1586 -7588 -1552 -7554
rect -1518 -7588 -1484 -7554
rect -1450 -7588 -1416 -7554
rect -1382 -7588 -1348 -7554
rect -1314 -7588 -1280 -7554
rect -1246 -7588 -1212 -7554
rect -1178 -7588 -1144 -7554
rect -1110 -7588 -1076 -7554
rect -1042 -7588 -1008 -7554
rect -974 -7588 -940 -7554
rect -906 -7588 -872 -7554
rect -838 -7588 -804 -7554
rect -770 -7588 -736 -7554
rect -702 -7588 -668 -7554
rect -634 -7588 -600 -7554
rect -566 -7588 -532 -7554
rect -498 -7588 -464 -7554
rect -430 -7588 -396 -7554
rect -362 -7588 -328 -7554
rect -294 -7588 -260 -7554
rect -226 -7588 -192 -7554
rect -158 -7588 -124 -7554
rect -90 -7588 -56 -7554
rect -22 -7588 12 -7554
rect 46 -7588 80 -7554
rect 114 -7588 148 -7554
rect 182 -7588 216 -7554
rect 250 -7588 284 -7554
rect 318 -7588 352 -7554
rect 386 -7588 420 -7554
rect 454 -7588 488 -7554
rect 522 -7588 556 -7554
rect 590 -7588 624 -7554
rect 658 -7588 692 -7554
rect 726 -7588 760 -7554
rect 794 -7588 828 -7554
rect 862 -7588 896 -7554
rect 930 -7588 964 -7554
rect 998 -7588 1032 -7554
rect 1066 -7588 1100 -7554
rect 1134 -7588 1168 -7554
rect 1202 -7588 1236 -7554
rect 1270 -7588 1304 -7554
rect 1338 -7588 1372 -7554
rect 1406 -7588 1440 -7554
rect 1474 -7588 1508 -7554
rect 1542 -7588 1576 -7554
rect 1610 -7588 1644 -7554
rect 1678 -7588 1712 -7554
rect 1746 -7588 1780 -7554
rect 1814 -7588 1848 -7554
rect 1882 -7588 1916 -7554
rect 1950 -7588 1984 -7554
rect 2018 -7588 2052 -7554
rect 2086 -7588 2120 -7554
rect 2154 -7588 2188 -7554
rect 2222 -7588 2256 -7554
rect 2290 -7588 2324 -7554
rect 2358 -7588 2392 -7554
rect 2426 -7588 2460 -7554
rect 2494 -7588 2528 -7554
rect 2562 -7588 2596 -7554
rect 2630 -7588 2664 -7554
rect 2698 -7588 2732 -7554
rect 2766 -7588 2800 -7554
rect 2834 -7588 2868 -7554
rect 2902 -7588 2936 -7554
rect 2970 -7588 3004 -7554
rect 3038 -7588 3072 -7554
rect 3106 -7588 3140 -7554
rect 3174 -7588 3208 -7554
rect 3242 -7588 3276 -7554
rect 3310 -7588 3344 -7554
rect 3378 -7588 3412 -7554
rect 3446 -7588 3480 -7554
rect 3514 -7588 3548 -7554
rect 3582 -7588 3616 -7554
rect 3650 -7588 3684 -7554
rect 3718 -7588 3752 -7554
rect 3786 -7588 3820 -7554
rect 3854 -7588 3888 -7554
rect 3922 -7588 3956 -7554
rect 3990 -7588 4024 -7554
rect 4058 -7588 4092 -7554
rect 4126 -7588 4160 -7554
rect 4194 -7588 4228 -7554
rect 4262 -7588 4296 -7554
rect 4330 -7588 4364 -7554
rect 4398 -7588 4432 -7554
rect 4466 -7588 4500 -7554
rect 4534 -7588 4568 -7554
rect 4602 -7588 4636 -7554
rect 4670 -7588 4704 -7554
rect 4738 -7588 4772 -7554
rect 4806 -7588 4840 -7554
rect 4874 -7588 4908 -7554
rect 4942 -7588 4976 -7554
rect 5010 -7588 5044 -7554
rect 5078 -7588 5112 -7554
rect 5146 -7588 5180 -7554
rect 5214 -7588 5248 -7554
rect 5282 -7588 5316 -7554
rect 5350 -7588 5384 -7554
rect 5418 -7588 5452 -7554
rect 5486 -7588 5520 -7554
rect 5554 -7588 5588 -7554
rect 5622 -7588 5656 -7554
rect 5690 -7588 5724 -7554
rect 5758 -7588 5792 -7554
rect 5826 -7588 5860 -7554
rect 5894 -7588 5928 -7554
rect 5962 -7588 5996 -7554
rect 6030 -7588 6064 -7554
rect 6098 -7588 6132 -7554
rect 6166 -7588 6200 -7554
rect 6234 -7588 6268 -7554
rect 6302 -7588 6336 -7554
rect 6370 -7588 6404 -7554
rect 6438 -7588 6472 -7554
rect 6506 -7588 6540 -7554
rect 6574 -7588 6608 -7554
rect 6642 -7588 6676 -7554
rect 6710 -7588 6744 -7554
rect 6778 -7588 6812 -7554
rect 6846 -7588 6880 -7554
rect 6914 -7588 6948 -7554
rect 6982 -7588 7016 -7554
rect 7050 -7588 7084 -7554
rect 7118 -7588 7152 -7554
rect 7186 -7588 7220 -7554
rect 7254 -7588 7288 -7554
rect 7322 -7588 7356 -7554
rect 7390 -7588 7424 -7554
rect 7458 -7588 7492 -7554
rect 7526 -7588 7560 -7554
rect 7594 -7588 7628 -7554
rect 7662 -7588 7696 -7554
rect 7730 -7588 7764 -7554
rect 7798 -7588 7832 -7554
rect 7866 -7588 7900 -7554
rect 7934 -7588 7968 -7554
rect 8002 -7588 8036 -7554
rect 8070 -7588 8104 -7554
rect 8138 -7588 8172 -7554
rect 8206 -7588 8240 -7554
rect 8274 -7588 8308 -7554
rect 8342 -7588 8376 -7554
rect 8410 -7588 8444 -7554
rect 8478 -7588 8512 -7554
rect 8546 -7588 8580 -7554
rect 8614 -7588 8648 -7554
rect 8682 -7588 8716 -7554
rect 8750 -7588 8784 -7554
rect 8818 -7588 8852 -7554
rect 8886 -7588 8920 -7554
rect 8954 -7588 8988 -7554
rect 9022 -7588 9056 -7554
rect 9090 -7588 9124 -7554
rect 9158 -7588 9192 -7554
rect 9226 -7588 9260 -7554
rect 9294 -7588 9328 -7554
rect 9362 -7588 9396 -7554
rect 9430 -7588 9464 -7554
rect 9498 -7588 9532 -7554
rect 9566 -7588 9600 -7554
rect 9634 -7588 9668 -7554
rect 9702 -7588 9736 -7554
rect 9770 -7588 9804 -7554
rect 9838 -7588 9872 -7554
rect 9906 -7588 9940 -7554
rect 9974 -7588 10008 -7554
rect 10042 -7588 10076 -7554
rect 10110 -7588 10144 -7554
rect 10178 -7588 10212 -7554
rect 10246 -7588 10280 -7554
rect 10314 -7588 10348 -7554
rect 10382 -7588 10416 -7554
rect 10450 -7588 10484 -7554
rect 10518 -7588 10552 -7554
rect 10586 -7588 10620 -7554
rect 10654 -7588 10688 -7554
rect 10722 -7588 10756 -7554
rect 10790 -7588 10824 -7554
rect 10858 -7588 10892 -7554
rect 10926 -7588 10960 -7554
rect 10994 -7588 11028 -7554
rect 11062 -7588 11096 -7554
rect 11130 -7588 11164 -7554
rect 11198 -7588 11232 -7554
rect 11266 -7588 11300 -7554
rect 11334 -7588 11368 -7554
rect 11402 -7588 11436 -7554
rect 11470 -7588 11504 -7554
rect 11538 -7588 11572 -7554
rect 11606 -7588 11640 -7554
rect 11674 -7588 11708 -7554
rect 11742 -7588 11776 -7554
rect 11810 -7588 11844 -7554
rect 11878 -7588 11912 -7554
rect 11946 -7588 11980 -7554
rect 12014 -7588 12048 -7554
rect 12082 -7588 12116 -7554
rect 12150 -7588 12184 -7554
rect 12218 -7588 12252 -7554
rect 12286 -7588 12320 -7554
rect 12354 -7588 12388 -7554
rect 12422 -7588 12456 -7554
rect 12490 -7588 12524 -7554
rect 12558 -7588 12592 -7554
rect 12626 -7588 12660 -7554
rect 12694 -7588 12728 -7554
rect 12762 -7588 12796 -7554
rect 12830 -7588 12864 -7554
rect 12898 -7588 12932 -7554
rect 12966 -7588 13000 -7554
rect 13034 -7588 13068 -7554
rect 13102 -7588 13136 -7554
rect 13170 -7588 13204 -7554
rect 13238 -7588 13272 -7554
rect 13306 -7588 13340 -7554
rect 13374 -7588 13408 -7554
rect 13442 -7588 13719 -7554
rect -7605 -7621 13719 -7588
rect -7605 -7850 -7505 -7621
rect -7605 -7884 -7572 -7850
rect -7538 -7884 -7505 -7850
rect -7605 -7918 -7505 -7884
rect -7605 -7952 -7572 -7918
rect -7538 -7952 -7505 -7918
rect -7605 -7986 -7505 -7952
rect -7605 -8020 -7572 -7986
rect -7538 -8020 -7505 -7986
rect -7605 -8054 -7505 -8020
rect -7605 -8088 -7572 -8054
rect -7538 -8088 -7505 -8054
rect -7605 -8122 -7505 -8088
rect -7605 -8156 -7572 -8122
rect -7538 -8156 -7505 -8122
rect -7605 -8190 -7505 -8156
rect -7605 -8224 -7572 -8190
rect -7538 -8224 -7505 -8190
rect -7605 -8258 -7505 -8224
rect -7605 -8292 -7572 -8258
rect -7538 -8292 -7505 -8258
rect -7605 -8326 -7505 -8292
rect -7605 -8360 -7572 -8326
rect -7538 -8360 -7505 -8326
rect -7605 -8394 -7505 -8360
rect -7605 -8428 -7572 -8394
rect -7538 -8428 -7505 -8394
rect -7605 -8462 -7505 -8428
rect -7605 -8496 -7572 -8462
rect -7538 -8496 -7505 -8462
rect -7605 -8530 -7505 -8496
rect -7605 -8564 -7572 -8530
rect -7538 -8564 -7505 -8530
rect -7605 -8598 -7505 -8564
rect -7605 -8632 -7572 -8598
rect -7538 -8632 -7505 -8598
rect -7605 -8666 -7505 -8632
rect -7605 -8700 -7572 -8666
rect -7538 -8700 -7505 -8666
rect -7605 -8734 -7505 -8700
rect -7605 -8768 -7572 -8734
rect -7538 -8768 -7505 -8734
rect -7605 -8802 -7505 -8768
rect -7605 -8836 -7572 -8802
rect -7538 -8836 -7505 -8802
rect -7605 -8870 -7505 -8836
rect -7605 -8904 -7572 -8870
rect -7538 -8904 -7505 -8870
rect -7605 -8938 -7505 -8904
rect -7605 -8972 -7572 -8938
rect -7538 -8972 -7505 -8938
rect -7605 -9006 -7505 -8972
rect -7605 -9040 -7572 -9006
rect -7538 -9040 -7505 -9006
rect -7605 -9074 -7505 -9040
rect -7605 -9108 -7572 -9074
rect -7538 -9108 -7505 -9074
rect -7605 -9142 -7505 -9108
rect -7605 -9176 -7572 -9142
rect -7538 -9176 -7505 -9142
rect -7605 -9210 -7505 -9176
rect -7605 -9244 -7572 -9210
rect -7538 -9244 -7505 -9210
rect -7605 -9278 -7505 -9244
rect -7605 -9312 -7572 -9278
rect -7538 -9312 -7505 -9278
rect -7605 -9346 -7505 -9312
rect -7605 -9380 -7572 -9346
rect -7538 -9380 -7505 -9346
rect -7605 -9414 -7505 -9380
rect -7605 -9448 -7572 -9414
rect -7538 -9448 -7505 -9414
rect -7605 -9482 -7505 -9448
rect -7605 -9516 -7572 -9482
rect -7538 -9516 -7505 -9482
rect -7605 -9550 -7505 -9516
rect -7605 -9584 -7572 -9550
rect -7538 -9584 -7505 -9550
rect -7605 -9618 -7505 -9584
rect -7605 -9652 -7572 -9618
rect -7538 -9652 -7505 -9618
rect -7605 -9686 -7505 -9652
rect -7605 -9720 -7572 -9686
rect -7538 -9720 -7505 -9686
rect -7605 -9754 -7505 -9720
rect -7605 -9788 -7572 -9754
rect -7538 -9788 -7505 -9754
rect -7605 -9822 -7505 -9788
rect -7605 -9856 -7572 -9822
rect -7538 -9856 -7505 -9822
rect -7605 -9890 -7505 -9856
rect -7605 -9924 -7572 -9890
rect -7538 -9924 -7505 -9890
rect -7605 -9958 -7505 -9924
rect -7605 -9992 -7572 -9958
rect -7538 -9992 -7505 -9958
rect -7605 -10026 -7505 -9992
rect -7605 -10060 -7572 -10026
rect -7538 -10060 -7505 -10026
rect -7605 -10094 -7505 -10060
rect -7605 -10128 -7572 -10094
rect -7538 -10128 -7505 -10094
rect -7605 -10162 -7505 -10128
rect -7605 -10196 -7572 -10162
rect -7538 -10196 -7505 -10162
rect -7605 -10230 -7505 -10196
rect -7605 -10264 -7572 -10230
rect -7538 -10264 -7505 -10230
rect -7605 -10298 -7505 -10264
rect -7605 -10332 -7572 -10298
rect -7538 -10332 -7505 -10298
rect -7605 -10366 -7505 -10332
rect -7605 -10400 -7572 -10366
rect -7538 -10400 -7505 -10366
rect -7605 -10434 -7505 -10400
rect -7605 -10468 -7572 -10434
rect -7538 -10468 -7505 -10434
rect -7605 -10502 -7505 -10468
rect -7605 -10536 -7572 -10502
rect -7538 -10536 -7505 -10502
rect -7605 -10570 -7505 -10536
rect -7605 -10604 -7572 -10570
rect -7538 -10604 -7505 -10570
rect -7605 -10638 -7505 -10604
rect -7605 -10672 -7572 -10638
rect -7538 -10672 -7505 -10638
rect -7605 -10706 -7505 -10672
rect -7605 -10740 -7572 -10706
rect -7538 -10740 -7505 -10706
rect -7605 -10774 -7505 -10740
rect -7605 -10808 -7572 -10774
rect -7538 -10808 -7505 -10774
rect -7605 -10842 -7505 -10808
rect -7605 -10876 -7572 -10842
rect -7538 -10876 -7505 -10842
rect -7605 -10910 -7505 -10876
rect -7605 -10944 -7572 -10910
rect -7538 -10944 -7505 -10910
rect -7605 -10978 -7505 -10944
rect -7605 -11012 -7572 -10978
rect -7538 -11012 -7505 -10978
rect -7605 -11046 -7505 -11012
rect -7605 -11080 -7572 -11046
rect -7538 -11080 -7505 -11046
rect -7605 -11114 -7505 -11080
rect -7605 -11148 -7572 -11114
rect -7538 -11148 -7505 -11114
rect -7605 -11182 -7505 -11148
rect -7605 -11216 -7572 -11182
rect -7538 -11216 -7505 -11182
rect -7605 -11250 -7505 -11216
rect -7605 -11284 -7572 -11250
rect -7538 -11284 -7505 -11250
rect -7605 -11318 -7505 -11284
rect -7605 -11352 -7572 -11318
rect -7538 -11352 -7505 -11318
rect -7605 -11386 -7505 -11352
rect -7605 -11420 -7572 -11386
rect -7538 -11420 -7505 -11386
rect -7605 -11454 -7505 -11420
rect -7605 -11488 -7572 -11454
rect -7538 -11488 -7505 -11454
rect -7605 -11522 -7505 -11488
rect -7605 -11556 -7572 -11522
rect -7538 -11556 -7505 -11522
rect -7605 -11590 -7505 -11556
rect -7605 -11624 -7572 -11590
rect -7538 -11624 -7505 -11590
rect -7605 -11658 -7505 -11624
rect -7605 -11692 -7572 -11658
rect -7538 -11692 -7505 -11658
rect -7605 -11726 -7505 -11692
rect -7605 -11760 -7572 -11726
rect -7538 -11760 -7505 -11726
rect -7605 -11794 -7505 -11760
rect -7605 -11828 -7572 -11794
rect -7538 -11828 -7505 -11794
rect -7605 -11862 -7505 -11828
rect -7605 -11896 -7572 -11862
rect -7538 -11896 -7505 -11862
rect -7605 -11930 -7505 -11896
rect -7605 -11964 -7572 -11930
rect -7538 -11964 -7505 -11930
rect -7605 -11998 -7505 -11964
rect -7605 -12032 -7572 -11998
rect -7538 -12032 -7505 -11998
rect -7605 -12066 -7505 -12032
rect -7605 -12100 -7572 -12066
rect -7538 -12100 -7505 -12066
rect -7605 -12134 -7505 -12100
rect -7605 -12168 -7572 -12134
rect -7538 -12168 -7505 -12134
rect -7605 -12202 -7505 -12168
rect -7605 -12236 -7572 -12202
rect -7538 -12236 -7505 -12202
rect -7605 -12270 -7505 -12236
rect -7605 -12304 -7572 -12270
rect -7538 -12304 -7505 -12270
rect -7605 -12338 -7505 -12304
rect -7605 -12372 -7572 -12338
rect -7538 -12372 -7505 -12338
rect -7605 -12406 -7505 -12372
rect -7605 -12440 -7572 -12406
rect -7538 -12440 -7505 -12406
rect -7605 -12474 -7505 -12440
rect -7605 -12508 -7572 -12474
rect -7538 -12508 -7505 -12474
rect -7605 -12542 -7505 -12508
rect -7605 -12576 -7572 -12542
rect -7538 -12576 -7505 -12542
rect -7605 -12610 -7505 -12576
rect -7605 -12644 -7572 -12610
rect -7538 -12644 -7505 -12610
rect -7605 -12678 -7505 -12644
rect -7605 -12712 -7572 -12678
rect -7538 -12712 -7505 -12678
rect -7605 -12746 -7505 -12712
rect -7605 -12780 -7572 -12746
rect -7538 -12780 -7505 -12746
rect -7605 -12814 -7505 -12780
rect -7605 -12848 -7572 -12814
rect -7538 -12848 -7505 -12814
rect -7605 -12882 -7505 -12848
rect -7605 -12916 -7572 -12882
rect -7538 -12916 -7505 -12882
rect -7605 -12950 -7505 -12916
rect -7605 -12984 -7572 -12950
rect -7538 -12984 -7505 -12950
rect -7605 -13018 -7505 -12984
rect -7605 -13052 -7572 -13018
rect -7538 -13052 -7505 -13018
rect -7605 -13086 -7505 -13052
rect -7605 -13120 -7572 -13086
rect -7538 -13120 -7505 -13086
rect -7605 -13154 -7505 -13120
rect -7605 -13188 -7572 -13154
rect -7538 -13188 -7505 -13154
rect -7605 -13222 -7505 -13188
rect -7605 -13256 -7572 -13222
rect -7538 -13256 -7505 -13222
rect -7605 -13290 -7505 -13256
rect -7605 -13324 -7572 -13290
rect -7538 -13324 -7505 -13290
rect -7605 -13358 -7505 -13324
rect -7605 -13392 -7572 -13358
rect -7538 -13392 -7505 -13358
rect -7605 -13426 -7505 -13392
rect -7605 -13460 -7572 -13426
rect -7538 -13460 -7505 -13426
rect -7605 -13494 -7505 -13460
rect -7605 -13528 -7572 -13494
rect -7538 -13528 -7505 -13494
rect -7605 -13562 -7505 -13528
rect -7605 -13596 -7572 -13562
rect -7538 -13596 -7505 -13562
rect -7605 -13630 -7505 -13596
rect -7605 -13664 -7572 -13630
rect -7538 -13664 -7505 -13630
rect -7605 -13698 -7505 -13664
rect -7605 -13732 -7572 -13698
rect -7538 -13732 -7505 -13698
rect -7605 -13766 -7505 -13732
rect -7605 -13800 -7572 -13766
rect -7538 -13800 -7505 -13766
rect -7605 -13834 -7505 -13800
rect -7605 -13868 -7572 -13834
rect -7538 -13868 -7505 -13834
rect -7605 -13902 -7505 -13868
rect -7605 -13936 -7572 -13902
rect -7538 -13936 -7505 -13902
rect -7605 -13970 -7505 -13936
rect -7605 -14004 -7572 -13970
rect -7538 -14004 -7505 -13970
rect -7605 -14038 -7505 -14004
rect -7605 -14072 -7572 -14038
rect -7538 -14072 -7505 -14038
rect -7605 -14106 -7505 -14072
rect -7605 -14140 -7572 -14106
rect -7538 -14140 -7505 -14106
rect -7605 -14174 -7505 -14140
rect -7605 -14208 -7572 -14174
rect -7538 -14208 -7505 -14174
rect -7605 -14242 -7505 -14208
rect -7605 -14276 -7572 -14242
rect -7538 -14276 -7505 -14242
rect -7605 -14310 -7505 -14276
rect -7605 -14344 -7572 -14310
rect -7538 -14344 -7505 -14310
rect -7605 -14378 -7505 -14344
rect -7605 -14412 -7572 -14378
rect -7538 -14412 -7505 -14378
rect -7605 -14446 -7505 -14412
rect -7605 -14480 -7572 -14446
rect -7538 -14480 -7505 -14446
rect -7605 -14514 -7505 -14480
rect -7605 -14548 -7572 -14514
rect -7538 -14548 -7505 -14514
rect -7605 -14582 -7505 -14548
rect -7605 -14616 -7572 -14582
rect -7538 -14616 -7505 -14582
rect -7605 -14650 -7505 -14616
rect -7605 -14684 -7572 -14650
rect -7538 -14684 -7505 -14650
rect -7605 -14718 -7505 -14684
rect -7605 -14752 -7572 -14718
rect -7538 -14752 -7505 -14718
rect -7605 -14786 -7505 -14752
rect -7605 -14820 -7572 -14786
rect -7538 -14820 -7505 -14786
rect -7605 -14854 -7505 -14820
rect -7605 -14888 -7572 -14854
rect -7538 -14888 -7505 -14854
rect -7605 -14922 -7505 -14888
rect -7605 -14956 -7572 -14922
rect -7538 -14956 -7505 -14922
rect -7605 -14990 -7505 -14956
rect -7605 -15024 -7572 -14990
rect -7538 -15024 -7505 -14990
rect -7605 -15058 -7505 -15024
rect -7605 -15092 -7572 -15058
rect -7538 -15092 -7505 -15058
rect -7605 -15126 -7505 -15092
rect -7605 -15160 -7572 -15126
rect -7538 -15160 -7505 -15126
rect -7605 -15194 -7505 -15160
rect -7605 -15228 -7572 -15194
rect -7538 -15228 -7505 -15194
rect -7605 -15262 -7505 -15228
rect -7605 -15296 -7572 -15262
rect -7538 -15296 -7505 -15262
rect -7605 -15330 -7505 -15296
rect -7605 -15364 -7572 -15330
rect -7538 -15364 -7505 -15330
rect -7605 -15398 -7505 -15364
rect -7605 -15432 -7572 -15398
rect -7538 -15432 -7505 -15398
rect -7605 -15466 -7505 -15432
rect -7605 -15500 -7572 -15466
rect -7538 -15500 -7505 -15466
rect -7605 -15534 -7505 -15500
rect -7605 -15568 -7572 -15534
rect -7538 -15568 -7505 -15534
rect -7605 -15602 -7505 -15568
rect -7605 -15636 -7572 -15602
rect -7538 -15636 -7505 -15602
rect -7605 -15670 -7505 -15636
rect -7605 -15704 -7572 -15670
rect -7538 -15704 -7505 -15670
rect -7605 -15738 -7505 -15704
rect -7605 -15772 -7572 -15738
rect -7538 -15772 -7505 -15738
rect -7605 -15806 -7505 -15772
rect -7605 -15840 -7572 -15806
rect -7538 -15840 -7505 -15806
rect -7605 -15874 -7505 -15840
rect -7605 -15908 -7572 -15874
rect -7538 -15908 -7505 -15874
rect -7605 -15942 -7505 -15908
rect -7605 -15976 -7572 -15942
rect -7538 -15976 -7505 -15942
rect -7605 -16010 -7505 -15976
rect -7605 -16044 -7572 -16010
rect -7538 -16044 -7505 -16010
rect -7605 -16078 -7505 -16044
rect -7605 -16112 -7572 -16078
rect -7538 -16112 -7505 -16078
rect -7605 -16146 -7505 -16112
rect -7605 -16180 -7572 -16146
rect -7538 -16180 -7505 -16146
rect -7605 -16214 -7505 -16180
rect -7605 -16248 -7572 -16214
rect -7538 -16248 -7505 -16214
rect -7605 -16282 -7505 -16248
rect -7605 -16316 -7572 -16282
rect -7538 -16316 -7505 -16282
rect -7605 -16350 -7505 -16316
rect -7605 -16384 -7572 -16350
rect -7538 -16384 -7505 -16350
rect -7605 -16418 -7505 -16384
rect -7605 -16452 -7572 -16418
rect -7538 -16452 -7505 -16418
rect -7605 -16486 -7505 -16452
rect -7605 -16520 -7572 -16486
rect -7538 -16520 -7505 -16486
rect -7605 -16554 -7505 -16520
rect -7605 -16588 -7572 -16554
rect -7538 -16588 -7505 -16554
rect -7605 -16622 -7505 -16588
rect -7605 -16656 -7572 -16622
rect -7538 -16656 -7505 -16622
rect -7605 -16690 -7505 -16656
rect -7605 -16724 -7572 -16690
rect -7538 -16724 -7505 -16690
rect -7605 -16758 -7505 -16724
rect -7605 -16792 -7572 -16758
rect -7538 -16792 -7505 -16758
rect -7605 -16826 -7505 -16792
rect -7605 -16860 -7572 -16826
rect -7538 -16860 -7505 -16826
rect -7605 -16894 -7505 -16860
rect -7605 -16928 -7572 -16894
rect -7538 -16928 -7505 -16894
rect -7605 -16962 -7505 -16928
rect -7605 -16996 -7572 -16962
rect -7538 -16996 -7505 -16962
rect -7605 -17030 -7505 -16996
rect -7605 -17064 -7572 -17030
rect -7538 -17064 -7505 -17030
rect -7605 -17098 -7505 -17064
rect -7605 -17132 -7572 -17098
rect -7538 -17132 -7505 -17098
rect -7605 -17166 -7505 -17132
rect -7605 -17200 -7572 -17166
rect -7538 -17200 -7505 -17166
rect -7605 -17234 -7505 -17200
rect -7605 -17268 -7572 -17234
rect -7538 -17268 -7505 -17234
rect -7605 -17459 -7505 -17268
rect 13619 -7731 13719 -7621
rect 13619 -7765 13652 -7731
rect 13686 -7765 13719 -7731
rect 13619 -7799 13719 -7765
rect 13619 -7833 13652 -7799
rect 13686 -7833 13719 -7799
rect 13619 -7867 13719 -7833
rect 13619 -7901 13652 -7867
rect 13686 -7901 13719 -7867
rect 13619 -7935 13719 -7901
rect 13619 -7969 13652 -7935
rect 13686 -7969 13719 -7935
rect 13619 -8003 13719 -7969
rect 13619 -8037 13652 -8003
rect 13686 -8037 13719 -8003
rect 13619 -8071 13719 -8037
rect 13619 -8105 13652 -8071
rect 13686 -8105 13719 -8071
rect 13619 -8139 13719 -8105
rect 13619 -8173 13652 -8139
rect 13686 -8173 13719 -8139
rect 13619 -8207 13719 -8173
rect 13619 -8241 13652 -8207
rect 13686 -8241 13719 -8207
rect 13619 -8275 13719 -8241
rect 13619 -8309 13652 -8275
rect 13686 -8309 13719 -8275
rect 13619 -8343 13719 -8309
rect 13619 -8377 13652 -8343
rect 13686 -8377 13719 -8343
rect 13619 -8411 13719 -8377
rect 13619 -8445 13652 -8411
rect 13686 -8445 13719 -8411
rect 13619 -8479 13719 -8445
rect 13619 -8513 13652 -8479
rect 13686 -8513 13719 -8479
rect 13619 -8547 13719 -8513
rect 13619 -8581 13652 -8547
rect 13686 -8581 13719 -8547
rect 13619 -8615 13719 -8581
rect 13619 -8649 13652 -8615
rect 13686 -8649 13719 -8615
rect 13619 -8683 13719 -8649
rect 13619 -8717 13652 -8683
rect 13686 -8717 13719 -8683
rect 13619 -8751 13719 -8717
rect 13619 -8785 13652 -8751
rect 13686 -8785 13719 -8751
rect 13619 -8819 13719 -8785
rect 13619 -8853 13652 -8819
rect 13686 -8853 13719 -8819
rect 13619 -8887 13719 -8853
rect 13619 -8921 13652 -8887
rect 13686 -8921 13719 -8887
rect 13619 -8955 13719 -8921
rect 13619 -8989 13652 -8955
rect 13686 -8989 13719 -8955
rect 13619 -9023 13719 -8989
rect 13619 -9057 13652 -9023
rect 13686 -9057 13719 -9023
rect 13619 -9091 13719 -9057
rect 13619 -9125 13652 -9091
rect 13686 -9125 13719 -9091
rect 13619 -9159 13719 -9125
rect 13619 -9193 13652 -9159
rect 13686 -9193 13719 -9159
rect 13619 -9227 13719 -9193
rect 13619 -9261 13652 -9227
rect 13686 -9261 13719 -9227
rect 13619 -9295 13719 -9261
rect 13619 -9329 13652 -9295
rect 13686 -9329 13719 -9295
rect 13619 -9363 13719 -9329
rect 13619 -9397 13652 -9363
rect 13686 -9397 13719 -9363
rect 13619 -9431 13719 -9397
rect 13619 -9465 13652 -9431
rect 13686 -9465 13719 -9431
rect 13619 -9499 13719 -9465
rect 13619 -9533 13652 -9499
rect 13686 -9533 13719 -9499
rect 13619 -9567 13719 -9533
rect 13619 -9601 13652 -9567
rect 13686 -9601 13719 -9567
rect 13619 -9635 13719 -9601
rect 13619 -9669 13652 -9635
rect 13686 -9669 13719 -9635
rect 13619 -9703 13719 -9669
rect 13619 -9737 13652 -9703
rect 13686 -9737 13719 -9703
rect 13619 -9771 13719 -9737
rect 13619 -9805 13652 -9771
rect 13686 -9805 13719 -9771
rect 13619 -9839 13719 -9805
rect 13619 -9873 13652 -9839
rect 13686 -9873 13719 -9839
rect 13619 -9907 13719 -9873
rect 13619 -9941 13652 -9907
rect 13686 -9941 13719 -9907
rect 13619 -9975 13719 -9941
rect 13619 -10009 13652 -9975
rect 13686 -10009 13719 -9975
rect 13619 -10043 13719 -10009
rect 13619 -10077 13652 -10043
rect 13686 -10077 13719 -10043
rect 13619 -10111 13719 -10077
rect 13619 -10145 13652 -10111
rect 13686 -10145 13719 -10111
rect 13619 -10179 13719 -10145
rect 13619 -10213 13652 -10179
rect 13686 -10213 13719 -10179
rect 13619 -10247 13719 -10213
rect 13619 -10281 13652 -10247
rect 13686 -10281 13719 -10247
rect 13619 -10315 13719 -10281
rect 13619 -10349 13652 -10315
rect 13686 -10349 13719 -10315
rect 13619 -10383 13719 -10349
rect 13619 -10417 13652 -10383
rect 13686 -10417 13719 -10383
rect 13619 -10451 13719 -10417
rect 13619 -10485 13652 -10451
rect 13686 -10485 13719 -10451
rect 13619 -10519 13719 -10485
rect 13619 -10553 13652 -10519
rect 13686 -10553 13719 -10519
rect 13619 -10587 13719 -10553
rect 13619 -10621 13652 -10587
rect 13686 -10621 13719 -10587
rect 13619 -10655 13719 -10621
rect 13619 -10689 13652 -10655
rect 13686 -10689 13719 -10655
rect 13619 -10723 13719 -10689
rect 13619 -10757 13652 -10723
rect 13686 -10757 13719 -10723
rect 13619 -10791 13719 -10757
rect 13619 -10825 13652 -10791
rect 13686 -10825 13719 -10791
rect 13619 -10859 13719 -10825
rect 13619 -10893 13652 -10859
rect 13686 -10893 13719 -10859
rect 13619 -10927 13719 -10893
rect 13619 -10961 13652 -10927
rect 13686 -10961 13719 -10927
rect 13619 -10995 13719 -10961
rect 13619 -11029 13652 -10995
rect 13686 -11029 13719 -10995
rect 13619 -11063 13719 -11029
rect 13619 -11097 13652 -11063
rect 13686 -11097 13719 -11063
rect 13619 -11131 13719 -11097
rect 13619 -11165 13652 -11131
rect 13686 -11165 13719 -11131
rect 13619 -11199 13719 -11165
rect 13619 -11233 13652 -11199
rect 13686 -11233 13719 -11199
rect 13619 -11267 13719 -11233
rect 13619 -11301 13652 -11267
rect 13686 -11301 13719 -11267
rect 13619 -11335 13719 -11301
rect 13619 -11369 13652 -11335
rect 13686 -11369 13719 -11335
rect 13619 -11403 13719 -11369
rect 13619 -11437 13652 -11403
rect 13686 -11437 13719 -11403
rect 13619 -11471 13719 -11437
rect 13619 -11505 13652 -11471
rect 13686 -11505 13719 -11471
rect 13619 -11539 13719 -11505
rect 13619 -11573 13652 -11539
rect 13686 -11573 13719 -11539
rect 13619 -11607 13719 -11573
rect 13619 -11641 13652 -11607
rect 13686 -11641 13719 -11607
rect 13619 -11675 13719 -11641
rect 13619 -11709 13652 -11675
rect 13686 -11709 13719 -11675
rect 13619 -11743 13719 -11709
rect 13619 -11777 13652 -11743
rect 13686 -11777 13719 -11743
rect 13619 -11811 13719 -11777
rect 13619 -11845 13652 -11811
rect 13686 -11845 13719 -11811
rect 13619 -11879 13719 -11845
rect 13619 -11913 13652 -11879
rect 13686 -11913 13719 -11879
rect 13619 -11947 13719 -11913
rect 13619 -11981 13652 -11947
rect 13686 -11981 13719 -11947
rect 13619 -12015 13719 -11981
rect 13619 -12049 13652 -12015
rect 13686 -12049 13719 -12015
rect 13619 -12083 13719 -12049
rect 13619 -12117 13652 -12083
rect 13686 -12117 13719 -12083
rect 13619 -12151 13719 -12117
rect 13619 -12185 13652 -12151
rect 13686 -12185 13719 -12151
rect 13619 -12219 13719 -12185
rect 13619 -12253 13652 -12219
rect 13686 -12253 13719 -12219
rect 13619 -12287 13719 -12253
rect 13619 -12321 13652 -12287
rect 13686 -12321 13719 -12287
rect 13619 -12355 13719 -12321
rect 13619 -12389 13652 -12355
rect 13686 -12389 13719 -12355
rect 13619 -12423 13719 -12389
rect 13619 -12457 13652 -12423
rect 13686 -12457 13719 -12423
rect 13619 -12491 13719 -12457
rect 13619 -12525 13652 -12491
rect 13686 -12525 13719 -12491
rect 13619 -12559 13719 -12525
rect 13619 -12593 13652 -12559
rect 13686 -12593 13719 -12559
rect 13619 -12627 13719 -12593
rect 13619 -12661 13652 -12627
rect 13686 -12661 13719 -12627
rect 13619 -12695 13719 -12661
rect 13619 -12729 13652 -12695
rect 13686 -12729 13719 -12695
rect 13619 -12763 13719 -12729
rect 13619 -12797 13652 -12763
rect 13686 -12797 13719 -12763
rect 13619 -12831 13719 -12797
rect 13619 -12865 13652 -12831
rect 13686 -12865 13719 -12831
rect 13619 -12899 13719 -12865
rect 13619 -12933 13652 -12899
rect 13686 -12933 13719 -12899
rect 13619 -12967 13719 -12933
rect 13619 -13001 13652 -12967
rect 13686 -13001 13719 -12967
rect 13619 -13035 13719 -13001
rect 13619 -13069 13652 -13035
rect 13686 -13069 13719 -13035
rect 13619 -13103 13719 -13069
rect 13619 -13137 13652 -13103
rect 13686 -13137 13719 -13103
rect 13619 -13171 13719 -13137
rect 13619 -13205 13652 -13171
rect 13686 -13205 13719 -13171
rect 13619 -13239 13719 -13205
rect 13619 -13273 13652 -13239
rect 13686 -13273 13719 -13239
rect 13619 -13307 13719 -13273
rect 13619 -13341 13652 -13307
rect 13686 -13341 13719 -13307
rect 13619 -13375 13719 -13341
rect 13619 -13409 13652 -13375
rect 13686 -13409 13719 -13375
rect 13619 -13443 13719 -13409
rect 13619 -13477 13652 -13443
rect 13686 -13477 13719 -13443
rect 13619 -13511 13719 -13477
rect 13619 -13545 13652 -13511
rect 13686 -13545 13719 -13511
rect 13619 -13579 13719 -13545
rect 13619 -13613 13652 -13579
rect 13686 -13613 13719 -13579
rect 13619 -13647 13719 -13613
rect 13619 -13681 13652 -13647
rect 13686 -13681 13719 -13647
rect 13619 -13715 13719 -13681
rect 13619 -13749 13652 -13715
rect 13686 -13749 13719 -13715
rect 13619 -13783 13719 -13749
rect 13619 -13817 13652 -13783
rect 13686 -13817 13719 -13783
rect 13619 -13851 13719 -13817
rect 13619 -13885 13652 -13851
rect 13686 -13885 13719 -13851
rect 13619 -13919 13719 -13885
rect 13619 -13953 13652 -13919
rect 13686 -13953 13719 -13919
rect 13619 -13987 13719 -13953
rect 13619 -14021 13652 -13987
rect 13686 -14021 13719 -13987
rect 13619 -14055 13719 -14021
rect 13619 -14089 13652 -14055
rect 13686 -14089 13719 -14055
rect 13619 -14123 13719 -14089
rect 13619 -14157 13652 -14123
rect 13686 -14157 13719 -14123
rect 13619 -14191 13719 -14157
rect 13619 -14225 13652 -14191
rect 13686 -14225 13719 -14191
rect 13619 -14259 13719 -14225
rect 13619 -14293 13652 -14259
rect 13686 -14293 13719 -14259
rect 13619 -14327 13719 -14293
rect 13619 -14361 13652 -14327
rect 13686 -14361 13719 -14327
rect 13619 -14395 13719 -14361
rect 13619 -14429 13652 -14395
rect 13686 -14429 13719 -14395
rect 13619 -14463 13719 -14429
rect 13619 -14497 13652 -14463
rect 13686 -14497 13719 -14463
rect 13619 -14531 13719 -14497
rect 13619 -14565 13652 -14531
rect 13686 -14565 13719 -14531
rect 13619 -14599 13719 -14565
rect 13619 -14633 13652 -14599
rect 13686 -14633 13719 -14599
rect 13619 -14667 13719 -14633
rect 13619 -14701 13652 -14667
rect 13686 -14701 13719 -14667
rect 13619 -14735 13719 -14701
rect 13619 -14769 13652 -14735
rect 13686 -14769 13719 -14735
rect 13619 -14803 13719 -14769
rect 13619 -14837 13652 -14803
rect 13686 -14837 13719 -14803
rect 13619 -14871 13719 -14837
rect 13619 -14905 13652 -14871
rect 13686 -14905 13719 -14871
rect 13619 -14939 13719 -14905
rect 13619 -14973 13652 -14939
rect 13686 -14973 13719 -14939
rect 13619 -15007 13719 -14973
rect 13619 -15041 13652 -15007
rect 13686 -15041 13719 -15007
rect 13619 -15075 13719 -15041
rect 13619 -15109 13652 -15075
rect 13686 -15109 13719 -15075
rect 13619 -15143 13719 -15109
rect 13619 -15177 13652 -15143
rect 13686 -15177 13719 -15143
rect 13619 -15211 13719 -15177
rect 13619 -15245 13652 -15211
rect 13686 -15245 13719 -15211
rect 13619 -15279 13719 -15245
rect 13619 -15313 13652 -15279
rect 13686 -15313 13719 -15279
rect 13619 -15347 13719 -15313
rect 13619 -15381 13652 -15347
rect 13686 -15381 13719 -15347
rect 13619 -15415 13719 -15381
rect 13619 -15449 13652 -15415
rect 13686 -15449 13719 -15415
rect 13619 -15483 13719 -15449
rect 13619 -15517 13652 -15483
rect 13686 -15517 13719 -15483
rect 13619 -15551 13719 -15517
rect 13619 -15585 13652 -15551
rect 13686 -15585 13719 -15551
rect 13619 -15619 13719 -15585
rect 13619 -15653 13652 -15619
rect 13686 -15653 13719 -15619
rect 13619 -15687 13719 -15653
rect 13619 -15721 13652 -15687
rect 13686 -15721 13719 -15687
rect 13619 -15755 13719 -15721
rect 13619 -15789 13652 -15755
rect 13686 -15789 13719 -15755
rect 13619 -15823 13719 -15789
rect 13619 -15857 13652 -15823
rect 13686 -15857 13719 -15823
rect 13619 -15891 13719 -15857
rect 13619 -15925 13652 -15891
rect 13686 -15925 13719 -15891
rect 13619 -15959 13719 -15925
rect 13619 -15993 13652 -15959
rect 13686 -15993 13719 -15959
rect 13619 -16027 13719 -15993
rect 13619 -16061 13652 -16027
rect 13686 -16061 13719 -16027
rect 13619 -16095 13719 -16061
rect 13619 -16129 13652 -16095
rect 13686 -16129 13719 -16095
rect 13619 -16163 13719 -16129
rect 13619 -16197 13652 -16163
rect 13686 -16197 13719 -16163
rect 13619 -16231 13719 -16197
rect 13619 -16265 13652 -16231
rect 13686 -16265 13719 -16231
rect 13619 -16299 13719 -16265
rect 13619 -16333 13652 -16299
rect 13686 -16333 13719 -16299
rect 13619 -16367 13719 -16333
rect 13619 -16401 13652 -16367
rect 13686 -16401 13719 -16367
rect 13619 -16435 13719 -16401
rect 13619 -16469 13652 -16435
rect 13686 -16469 13719 -16435
rect 13619 -16503 13719 -16469
rect 13619 -16537 13652 -16503
rect 13686 -16537 13719 -16503
rect 13619 -16571 13719 -16537
rect 13619 -16605 13652 -16571
rect 13686 -16605 13719 -16571
rect 13619 -16639 13719 -16605
rect 13619 -16673 13652 -16639
rect 13686 -16673 13719 -16639
rect 13619 -16707 13719 -16673
rect 13619 -16741 13652 -16707
rect 13686 -16741 13719 -16707
rect 13619 -16775 13719 -16741
rect 13619 -16809 13652 -16775
rect 13686 -16809 13719 -16775
rect 13619 -16843 13719 -16809
rect 13619 -16877 13652 -16843
rect 13686 -16877 13719 -16843
rect 13619 -16911 13719 -16877
rect 13619 -16945 13652 -16911
rect 13686 -16945 13719 -16911
rect 13619 -16979 13719 -16945
rect 13619 -17013 13652 -16979
rect 13686 -17013 13719 -16979
rect 13619 -17047 13719 -17013
rect 13619 -17081 13652 -17047
rect 13686 -17081 13719 -17047
rect 13619 -17115 13719 -17081
rect 13619 -17149 13652 -17115
rect 13686 -17149 13719 -17115
rect 13619 -17459 13719 -17149
rect -7605 -17492 13719 -17459
rect -7605 -17526 -7319 -17492
rect -7285 -17526 -7247 -17492
rect -7213 -17526 -7175 -17492
rect -7141 -17526 -7103 -17492
rect -7069 -17526 -7031 -17492
rect -6997 -17526 -6959 -17492
rect -6925 -17526 -6887 -17492
rect -6853 -17526 -6815 -17492
rect -6781 -17526 -6743 -17492
rect -6709 -17526 -6671 -17492
rect -6637 -17526 -6599 -17492
rect -6565 -17526 -6527 -17492
rect -6493 -17526 -6455 -17492
rect -6421 -17526 -6383 -17492
rect -6349 -17526 -6311 -17492
rect -6277 -17526 -6239 -17492
rect -6205 -17526 -6167 -17492
rect -6133 -17526 -6095 -17492
rect -6061 -17526 -6023 -17492
rect -5989 -17526 -5951 -17492
rect -5917 -17526 -5879 -17492
rect -5845 -17526 -5807 -17492
rect -5773 -17526 -5735 -17492
rect -5701 -17526 -5663 -17492
rect -5629 -17526 -5591 -17492
rect -5557 -17526 -5519 -17492
rect -5485 -17526 -5447 -17492
rect -5413 -17526 -5375 -17492
rect -5341 -17526 -5303 -17492
rect -5269 -17526 -5231 -17492
rect -5197 -17526 -5159 -17492
rect -5125 -17526 -5087 -17492
rect -5053 -17526 -5015 -17492
rect -4981 -17526 -4943 -17492
rect -4909 -17526 -4871 -17492
rect -4837 -17526 -4799 -17492
rect -4765 -17526 -4727 -17492
rect -4693 -17526 -4655 -17492
rect -4621 -17526 -4583 -17492
rect -4549 -17526 -4511 -17492
rect -4477 -17526 -4439 -17492
rect -4405 -17526 -4367 -17492
rect -4333 -17526 -4295 -17492
rect -4261 -17526 -4223 -17492
rect -4189 -17526 -4151 -17492
rect -4117 -17526 -4079 -17492
rect -4045 -17526 -4007 -17492
rect -3973 -17526 -3935 -17492
rect -3901 -17526 -3863 -17492
rect -3829 -17526 -3791 -17492
rect -3757 -17526 -3719 -17492
rect -3685 -17526 -3647 -17492
rect -3613 -17526 -3575 -17492
rect -3541 -17526 -3503 -17492
rect -3469 -17526 -3431 -17492
rect -3397 -17526 -3359 -17492
rect -3325 -17526 -3287 -17492
rect -3253 -17526 -3215 -17492
rect -3181 -17526 -3143 -17492
rect -3109 -17526 -3071 -17492
rect -3037 -17526 -2999 -17492
rect -2965 -17526 -2927 -17492
rect -2893 -17526 -2855 -17492
rect -2821 -17526 -2783 -17492
rect -2749 -17526 -2711 -17492
rect -2677 -17526 -2639 -17492
rect -2605 -17526 -2567 -17492
rect -2533 -17526 -2495 -17492
rect -2461 -17526 -2423 -17492
rect -2389 -17526 -2351 -17492
rect -2317 -17526 -2279 -17492
rect -2245 -17526 -2207 -17492
rect -2173 -17526 -2135 -17492
rect -2101 -17526 -2063 -17492
rect -2029 -17526 -1991 -17492
rect -1957 -17526 -1919 -17492
rect -1885 -17526 -1847 -17492
rect -1813 -17526 -1775 -17492
rect -1741 -17526 -1703 -17492
rect -1669 -17526 -1631 -17492
rect -1597 -17526 -1559 -17492
rect -1525 -17526 -1487 -17492
rect -1453 -17526 -1415 -17492
rect -1381 -17526 -1343 -17492
rect -1309 -17526 -1271 -17492
rect -1237 -17526 -1199 -17492
rect -1165 -17526 -1127 -17492
rect -1093 -17526 -1055 -17492
rect -1021 -17526 -983 -17492
rect -949 -17526 -911 -17492
rect -877 -17526 -839 -17492
rect -805 -17526 -767 -17492
rect -733 -17526 -695 -17492
rect -661 -17526 -623 -17492
rect -589 -17526 -551 -17492
rect -517 -17526 -479 -17492
rect -445 -17526 -407 -17492
rect -373 -17526 -335 -17492
rect -301 -17526 -263 -17492
rect -229 -17526 -191 -17492
rect -157 -17526 -119 -17492
rect -85 -17526 -47 -17492
rect -13 -17526 25 -17492
rect 59 -17526 97 -17492
rect 131 -17526 169 -17492
rect 203 -17526 241 -17492
rect 275 -17526 313 -17492
rect 347 -17526 385 -17492
rect 419 -17526 457 -17492
rect 491 -17526 529 -17492
rect 563 -17526 601 -17492
rect 635 -17526 673 -17492
rect 707 -17526 745 -17492
rect 779 -17526 817 -17492
rect 851 -17526 889 -17492
rect 923 -17526 961 -17492
rect 995 -17526 1033 -17492
rect 1067 -17526 1105 -17492
rect 1139 -17526 1177 -17492
rect 1211 -17526 1249 -17492
rect 1283 -17526 1321 -17492
rect 1355 -17526 1393 -17492
rect 1427 -17526 1465 -17492
rect 1499 -17526 1537 -17492
rect 1571 -17526 1609 -17492
rect 1643 -17526 1681 -17492
rect 1715 -17526 1753 -17492
rect 1787 -17526 1825 -17492
rect 1859 -17526 1897 -17492
rect 1931 -17526 1969 -17492
rect 2003 -17526 2041 -17492
rect 2075 -17526 2113 -17492
rect 2147 -17526 2185 -17492
rect 2219 -17526 2257 -17492
rect 2291 -17526 2329 -17492
rect 2363 -17526 2401 -17492
rect 2435 -17526 2473 -17492
rect 2507 -17526 2545 -17492
rect 2579 -17526 2617 -17492
rect 2651 -17526 2689 -17492
rect 2723 -17526 2761 -17492
rect 2795 -17526 2833 -17492
rect 2867 -17526 2905 -17492
rect 2939 -17526 2977 -17492
rect 3011 -17526 3049 -17492
rect 3083 -17526 3121 -17492
rect 3155 -17526 3193 -17492
rect 3227 -17526 3265 -17492
rect 3299 -17526 3337 -17492
rect 3371 -17526 3409 -17492
rect 3443 -17526 3481 -17492
rect 3515 -17526 3553 -17492
rect 3587 -17526 3625 -17492
rect 3659 -17526 3697 -17492
rect 3731 -17526 3769 -17492
rect 3803 -17526 3841 -17492
rect 3875 -17526 3913 -17492
rect 3947 -17526 3985 -17492
rect 4019 -17526 4057 -17492
rect 4091 -17526 4129 -17492
rect 4163 -17526 4201 -17492
rect 4235 -17526 4273 -17492
rect 4307 -17526 4345 -17492
rect 4379 -17526 4417 -17492
rect 4451 -17526 4489 -17492
rect 4523 -17526 4561 -17492
rect 4595 -17526 4633 -17492
rect 4667 -17526 4705 -17492
rect 4739 -17526 4777 -17492
rect 4811 -17526 4849 -17492
rect 4883 -17526 4921 -17492
rect 4955 -17526 4993 -17492
rect 5027 -17526 5065 -17492
rect 5099 -17526 5137 -17492
rect 5171 -17526 5209 -17492
rect 5243 -17526 5281 -17492
rect 5315 -17526 5353 -17492
rect 5387 -17526 5425 -17492
rect 5459 -17526 5497 -17492
rect 5531 -17526 5569 -17492
rect 5603 -17526 5641 -17492
rect 5675 -17526 5713 -17492
rect 5747 -17526 5785 -17492
rect 5819 -17526 5857 -17492
rect 5891 -17526 5929 -17492
rect 5963 -17526 6001 -17492
rect 6035 -17526 6073 -17492
rect 6107 -17526 6145 -17492
rect 6179 -17526 6217 -17492
rect 6251 -17526 6289 -17492
rect 6323 -17526 6361 -17492
rect 6395 -17526 6433 -17492
rect 6467 -17526 6505 -17492
rect 6539 -17526 6577 -17492
rect 6611 -17526 6649 -17492
rect 6683 -17526 6721 -17492
rect 6755 -17526 6793 -17492
rect 6827 -17526 6865 -17492
rect 6899 -17526 6937 -17492
rect 6971 -17526 7009 -17492
rect 7043 -17526 7081 -17492
rect 7115 -17526 7153 -17492
rect 7187 -17526 7225 -17492
rect 7259 -17526 7297 -17492
rect 7331 -17526 7369 -17492
rect 7403 -17526 7441 -17492
rect 7475 -17526 7513 -17492
rect 7547 -17526 7585 -17492
rect 7619 -17526 7657 -17492
rect 7691 -17526 7729 -17492
rect 7763 -17526 7801 -17492
rect 7835 -17526 7873 -17492
rect 7907 -17526 7945 -17492
rect 7979 -17526 8017 -17492
rect 8051 -17526 8089 -17492
rect 8123 -17526 8161 -17492
rect 8195 -17526 8233 -17492
rect 8267 -17526 8305 -17492
rect 8339 -17526 8377 -17492
rect 8411 -17526 8449 -17492
rect 8483 -17526 8521 -17492
rect 8555 -17526 8593 -17492
rect 8627 -17526 8665 -17492
rect 8699 -17526 8737 -17492
rect 8771 -17526 8809 -17492
rect 8843 -17526 8881 -17492
rect 8915 -17526 8953 -17492
rect 8987 -17526 9025 -17492
rect 9059 -17526 9097 -17492
rect 9131 -17526 9169 -17492
rect 9203 -17526 9241 -17492
rect 9275 -17526 9313 -17492
rect 9347 -17526 9385 -17492
rect 9419 -17526 9457 -17492
rect 9491 -17526 9529 -17492
rect 9563 -17526 9601 -17492
rect 9635 -17526 9673 -17492
rect 9707 -17526 9745 -17492
rect 9779 -17526 9817 -17492
rect 9851 -17526 9889 -17492
rect 9923 -17526 9961 -17492
rect 9995 -17526 10033 -17492
rect 10067 -17526 10105 -17492
rect 10139 -17526 10177 -17492
rect 10211 -17526 10249 -17492
rect 10283 -17526 10321 -17492
rect 10355 -17526 10393 -17492
rect 10427 -17526 10465 -17492
rect 10499 -17526 10537 -17492
rect 10571 -17526 10609 -17492
rect 10643 -17526 10681 -17492
rect 10715 -17526 10753 -17492
rect 10787 -17526 10825 -17492
rect 10859 -17526 10897 -17492
rect 10931 -17526 10969 -17492
rect 11003 -17526 11041 -17492
rect 11075 -17526 11113 -17492
rect 11147 -17526 11185 -17492
rect 11219 -17526 11257 -17492
rect 11291 -17526 11329 -17492
rect 11363 -17526 11401 -17492
rect 11435 -17526 11473 -17492
rect 11507 -17526 11545 -17492
rect 11579 -17526 11617 -17492
rect 11651 -17526 11689 -17492
rect 11723 -17526 11761 -17492
rect 11795 -17526 11833 -17492
rect 11867 -17526 11905 -17492
rect 11939 -17526 11977 -17492
rect 12011 -17526 12049 -17492
rect 12083 -17526 12121 -17492
rect 12155 -17526 12193 -17492
rect 12227 -17526 12265 -17492
rect 12299 -17526 12337 -17492
rect 12371 -17526 12409 -17492
rect 12443 -17526 12481 -17492
rect 12515 -17526 12553 -17492
rect 12587 -17526 12625 -17492
rect 12659 -17526 12697 -17492
rect 12731 -17526 12769 -17492
rect 12803 -17526 12841 -17492
rect 12875 -17526 12913 -17492
rect 12947 -17526 12985 -17492
rect 13019 -17526 13057 -17492
rect 13091 -17526 13129 -17492
rect 13163 -17526 13201 -17492
rect 13235 -17526 13273 -17492
rect 13307 -17526 13345 -17492
rect 13379 -17526 13719 -17492
rect -7605 -17559 13719 -17526
<< viali >>
rect -7370 -1324 -7346 -1290
rect -7346 -1324 -7336 -1290
rect -7298 -1324 -7278 -1290
rect -7278 -1324 -7264 -1290
rect -7226 -1324 -7210 -1290
rect -7210 -1324 -7192 -1290
rect -7154 -1324 -7142 -1290
rect -7142 -1324 -7120 -1290
rect -7082 -1324 -7074 -1290
rect -7074 -1324 -7048 -1290
rect -7010 -1324 -7006 -1290
rect -7006 -1324 -6976 -1290
rect -6938 -1324 -6904 -1290
rect -6866 -1324 -6836 -1290
rect -6836 -1324 -6832 -1290
rect -6794 -1324 -6768 -1290
rect -6768 -1324 -6760 -1290
rect -6722 -1324 -6700 -1290
rect -6700 -1324 -6688 -1290
rect -6650 -1324 -6632 -1290
rect -6632 -1324 -6616 -1290
rect -6578 -1324 -6564 -1290
rect -6564 -1324 -6544 -1290
rect -6506 -1324 -6496 -1290
rect -6496 -1324 -6472 -1290
rect -6434 -1324 -6428 -1290
rect -6428 -1324 -6400 -1290
rect -6362 -1324 -6360 -1290
rect -6360 -1324 -6328 -1290
rect -6290 -1324 -6258 -1290
rect -6258 -1324 -6256 -1290
rect -6218 -1324 -6190 -1290
rect -6190 -1324 -6184 -1290
rect -6146 -1324 -6122 -1290
rect -6122 -1324 -6112 -1290
rect -6074 -1324 -6054 -1290
rect -6054 -1324 -6040 -1290
rect -6002 -1324 -5986 -1290
rect -5986 -1324 -5968 -1290
rect -5930 -1324 -5918 -1290
rect -5918 -1324 -5896 -1290
rect -5858 -1324 -5850 -1290
rect -5850 -1324 -5824 -1290
rect -5786 -1324 -5782 -1290
rect -5782 -1324 -5752 -1290
rect -5714 -1324 -5680 -1290
rect -5642 -1324 -5612 -1290
rect -5612 -1324 -5608 -1290
rect -5570 -1324 -5544 -1290
rect -5544 -1324 -5536 -1290
rect -5498 -1324 -5476 -1290
rect -5476 -1324 -5464 -1290
rect -5426 -1324 -5408 -1290
rect -5408 -1324 -5392 -1290
rect -5354 -1324 -5340 -1290
rect -5340 -1324 -5320 -1290
rect -5282 -1324 -5272 -1290
rect -5272 -1324 -5248 -1290
rect -5210 -1324 -5204 -1290
rect -5204 -1324 -5176 -1290
rect -5138 -1324 -5136 -1290
rect -5136 -1324 -5104 -1290
rect -5066 -1324 -5034 -1290
rect -5034 -1324 -5032 -1290
rect -4994 -1324 -4966 -1290
rect -4966 -1324 -4960 -1290
rect -4922 -1324 -4898 -1290
rect -4898 -1324 -4888 -1290
rect -4850 -1324 -4830 -1290
rect -4830 -1324 -4816 -1290
rect -4778 -1324 -4762 -1290
rect -4762 -1324 -4744 -1290
rect -4706 -1324 -4694 -1290
rect -4694 -1324 -4672 -1290
rect -4634 -1324 -4626 -1290
rect -4626 -1324 -4600 -1290
rect -4562 -1324 -4558 -1290
rect -4558 -1324 -4528 -1290
rect -4490 -1324 -4456 -1290
rect -4418 -1324 -4388 -1290
rect -4388 -1324 -4384 -1290
rect -4346 -1324 -4320 -1290
rect -4320 -1324 -4312 -1290
rect -4274 -1324 -4252 -1290
rect -4252 -1324 -4240 -1290
rect -4202 -1324 -4184 -1290
rect -4184 -1324 -4168 -1290
rect -4130 -1324 -4116 -1290
rect -4116 -1324 -4096 -1290
rect -4058 -1324 -4048 -1290
rect -4048 -1324 -4024 -1290
rect -3986 -1324 -3980 -1290
rect -3980 -1324 -3952 -1290
rect -3914 -1324 -3912 -1290
rect -3912 -1324 -3880 -1290
rect -3842 -1324 -3810 -1290
rect -3810 -1324 -3808 -1290
rect -3770 -1324 -3742 -1290
rect -3742 -1324 -3736 -1290
rect -3698 -1324 -3674 -1290
rect -3674 -1324 -3664 -1290
rect -3626 -1324 -3606 -1290
rect -3606 -1324 -3592 -1290
rect -3554 -1324 -3538 -1290
rect -3538 -1324 -3520 -1290
rect -3482 -1324 -3470 -1290
rect -3470 -1324 -3448 -1290
rect -3410 -1324 -3402 -1290
rect -3402 -1324 -3376 -1290
rect -3338 -1324 -3334 -1290
rect -3334 -1324 -3304 -1290
rect -3266 -1324 -3232 -1290
rect -3194 -1324 -3164 -1290
rect -3164 -1324 -3160 -1290
rect -3122 -1324 -3096 -1290
rect -3096 -1324 -3088 -1290
rect -3050 -1324 -3028 -1290
rect -3028 -1324 -3016 -1290
rect -2978 -1324 -2960 -1290
rect -2960 -1324 -2944 -1290
rect -2906 -1324 -2892 -1290
rect -2892 -1324 -2872 -1290
rect -2834 -1324 -2824 -1290
rect -2824 -1324 -2800 -1290
rect -2762 -1324 -2756 -1290
rect -2756 -1324 -2728 -1290
rect -2690 -1324 -2688 -1290
rect -2688 -1324 -2656 -1290
rect -2618 -1324 -2586 -1290
rect -2586 -1324 -2584 -1290
rect -2546 -1324 -2518 -1290
rect -2518 -1324 -2512 -1290
rect -2474 -1324 -2450 -1290
rect -2450 -1324 -2440 -1290
rect -2402 -1324 -2382 -1290
rect -2382 -1324 -2368 -1290
rect -2330 -1324 -2314 -1290
rect -2314 -1324 -2296 -1290
rect -2258 -1324 -2246 -1290
rect -2246 -1324 -2224 -1290
rect -2186 -1324 -2178 -1290
rect -2178 -1324 -2152 -1290
rect -2114 -1324 -2110 -1290
rect -2110 -1324 -2080 -1290
rect -2042 -1324 -2008 -1290
rect -1970 -1324 -1940 -1290
rect -1940 -1324 -1936 -1290
rect -1898 -1324 -1872 -1290
rect -1872 -1324 -1864 -1290
rect -1826 -1324 -1804 -1290
rect -1804 -1324 -1792 -1290
rect -1754 -1324 -1736 -1290
rect -1736 -1324 -1720 -1290
rect -1682 -1324 -1668 -1290
rect -1668 -1324 -1648 -1290
rect -1610 -1324 -1600 -1290
rect -1600 -1324 -1576 -1290
rect -1538 -1324 -1532 -1290
rect -1532 -1324 -1504 -1290
rect -1466 -1324 -1464 -1290
rect -1464 -1324 -1432 -1290
rect -1394 -1324 -1362 -1290
rect -1362 -1324 -1360 -1290
rect -1322 -1324 -1294 -1290
rect -1294 -1324 -1288 -1290
rect -1250 -1324 -1226 -1290
rect -1226 -1324 -1216 -1290
rect -1178 -1324 -1158 -1290
rect -1158 -1324 -1144 -1290
rect -1106 -1324 -1090 -1290
rect -1090 -1324 -1072 -1290
rect -1034 -1324 -1022 -1290
rect -1022 -1324 -1000 -1290
rect -962 -1324 -954 -1290
rect -954 -1324 -928 -1290
rect -890 -1324 -886 -1290
rect -886 -1324 -856 -1290
rect -818 -1324 -784 -1290
rect -746 -1324 -716 -1290
rect -716 -1324 -712 -1290
rect -674 -1324 -648 -1290
rect -648 -1324 -640 -1290
rect -602 -1324 -580 -1290
rect -580 -1324 -568 -1290
rect -530 -1324 -512 -1290
rect -512 -1324 -496 -1290
rect -458 -1324 -444 -1290
rect -444 -1324 -424 -1290
rect -386 -1324 -376 -1290
rect -376 -1324 -352 -1290
rect -314 -1324 -308 -1290
rect -308 -1324 -280 -1290
rect -242 -1324 -240 -1290
rect -240 -1324 -208 -1290
rect -170 -1324 -138 -1290
rect -138 -1324 -136 -1290
rect -98 -1324 -70 -1290
rect -70 -1324 -64 -1290
rect -26 -1324 -2 -1290
rect -2 -1324 8 -1290
rect 46 -1324 66 -1290
rect 66 -1324 80 -1290
rect 118 -1324 134 -1290
rect 134 -1324 152 -1290
rect 190 -1324 202 -1290
rect 202 -1324 224 -1290
rect 262 -1324 270 -1290
rect 270 -1324 296 -1290
rect 334 -1324 338 -1290
rect 338 -1324 368 -1290
rect 406 -1324 440 -1290
rect 478 -1324 508 -1290
rect 508 -1324 512 -1290
rect 550 -1324 576 -1290
rect 576 -1324 584 -1290
rect 622 -1324 644 -1290
rect 644 -1324 656 -1290
rect 694 -1324 712 -1290
rect 712 -1324 728 -1290
rect 766 -1324 780 -1290
rect 780 -1324 800 -1290
rect 838 -1324 848 -1290
rect 848 -1324 872 -1290
rect 910 -1324 916 -1290
rect 916 -1324 944 -1290
rect 982 -1324 984 -1290
rect 984 -1324 1016 -1290
rect 1054 -1324 1086 -1290
rect 1086 -1324 1088 -1290
rect 1126 -1324 1154 -1290
rect 1154 -1324 1160 -1290
rect 1198 -1324 1222 -1290
rect 1222 -1324 1232 -1290
rect 1270 -1324 1290 -1290
rect 1290 -1324 1304 -1290
rect 1342 -1324 1358 -1290
rect 1358 -1324 1376 -1290
rect 1414 -1324 1426 -1290
rect 1426 -1324 1448 -1290
rect 1486 -1324 1494 -1290
rect 1494 -1324 1520 -1290
rect 1558 -1324 1562 -1290
rect 1562 -1324 1592 -1290
rect 1630 -1324 1664 -1290
rect 1702 -1324 1732 -1290
rect 1732 -1324 1736 -1290
rect 1774 -1324 1800 -1290
rect 1800 -1324 1808 -1290
rect 1846 -1324 1868 -1290
rect 1868 -1324 1880 -1290
rect 1918 -1324 1936 -1290
rect 1936 -1324 1952 -1290
rect 1990 -1324 2004 -1290
rect 2004 -1324 2024 -1290
rect 2062 -1324 2072 -1290
rect 2072 -1324 2096 -1290
rect 2134 -1324 2140 -1290
rect 2140 -1324 2168 -1290
rect 2206 -1324 2208 -1290
rect 2208 -1324 2240 -1290
rect 2278 -1324 2310 -1290
rect 2310 -1324 2312 -1290
rect 2350 -1324 2378 -1290
rect 2378 -1324 2384 -1290
rect 2422 -1324 2446 -1290
rect 2446 -1324 2456 -1290
rect 2494 -1324 2514 -1290
rect 2514 -1324 2528 -1290
rect 2566 -1324 2582 -1290
rect 2582 -1324 2600 -1290
rect 2638 -1324 2650 -1290
rect 2650 -1324 2672 -1290
rect 2710 -1324 2718 -1290
rect 2718 -1324 2744 -1290
rect 2782 -1324 2786 -1290
rect 2786 -1324 2816 -1290
rect 2854 -1324 2888 -1290
rect 2926 -1324 2956 -1290
rect 2956 -1324 2960 -1290
rect 2998 -1324 3024 -1290
rect 3024 -1324 3032 -1290
rect 3070 -1324 3092 -1290
rect 3092 -1324 3104 -1290
rect 3142 -1324 3160 -1290
rect 3160 -1324 3176 -1290
rect 3214 -1324 3228 -1290
rect 3228 -1324 3248 -1290
rect 3286 -1324 3296 -1290
rect 3296 -1324 3320 -1290
rect -7319 -17526 -7285 -17492
rect -7247 -17526 -7213 -17492
rect -7175 -17526 -7141 -17492
rect -7103 -17526 -7069 -17492
rect -7031 -17526 -6997 -17492
rect -6959 -17526 -6925 -17492
rect -6887 -17526 -6853 -17492
rect -6815 -17526 -6781 -17492
rect -6743 -17526 -6709 -17492
rect -6671 -17526 -6637 -17492
rect -6599 -17526 -6565 -17492
rect -6527 -17526 -6493 -17492
rect -6455 -17526 -6421 -17492
rect -6383 -17526 -6349 -17492
rect -6311 -17526 -6277 -17492
rect -6239 -17526 -6205 -17492
rect -6167 -17526 -6133 -17492
rect -6095 -17526 -6061 -17492
rect -6023 -17526 -5989 -17492
rect -5951 -17526 -5917 -17492
rect -5879 -17526 -5845 -17492
rect -5807 -17526 -5773 -17492
rect -5735 -17526 -5701 -17492
rect -5663 -17526 -5629 -17492
rect -5591 -17526 -5557 -17492
rect -5519 -17526 -5485 -17492
rect -5447 -17526 -5413 -17492
rect -5375 -17526 -5341 -17492
rect -5303 -17526 -5269 -17492
rect -5231 -17526 -5197 -17492
rect -5159 -17526 -5125 -17492
rect -5087 -17526 -5053 -17492
rect -5015 -17526 -4981 -17492
rect -4943 -17526 -4909 -17492
rect -4871 -17526 -4837 -17492
rect -4799 -17526 -4765 -17492
rect -4727 -17526 -4693 -17492
rect -4655 -17526 -4621 -17492
rect -4583 -17526 -4549 -17492
rect -4511 -17526 -4477 -17492
rect -4439 -17526 -4405 -17492
rect -4367 -17526 -4333 -17492
rect -4295 -17526 -4261 -17492
rect -4223 -17526 -4189 -17492
rect -4151 -17526 -4117 -17492
rect -4079 -17526 -4045 -17492
rect -4007 -17526 -3973 -17492
rect -3935 -17526 -3901 -17492
rect -3863 -17526 -3829 -17492
rect -3791 -17526 -3757 -17492
rect -3719 -17526 -3685 -17492
rect -3647 -17526 -3613 -17492
rect -3575 -17526 -3541 -17492
rect -3503 -17526 -3469 -17492
rect -3431 -17526 -3397 -17492
rect -3359 -17526 -3325 -17492
rect -3287 -17526 -3253 -17492
rect -3215 -17526 -3181 -17492
rect -3143 -17526 -3109 -17492
rect -3071 -17526 -3037 -17492
rect -2999 -17526 -2965 -17492
rect -2927 -17526 -2893 -17492
rect -2855 -17526 -2821 -17492
rect -2783 -17526 -2749 -17492
rect -2711 -17526 -2677 -17492
rect -2639 -17526 -2605 -17492
rect -2567 -17526 -2533 -17492
rect -2495 -17526 -2461 -17492
rect -2423 -17526 -2389 -17492
rect -2351 -17526 -2317 -17492
rect -2279 -17526 -2245 -17492
rect -2207 -17526 -2173 -17492
rect -2135 -17526 -2101 -17492
rect -2063 -17526 -2029 -17492
rect -1991 -17526 -1957 -17492
rect -1919 -17526 -1885 -17492
rect -1847 -17526 -1813 -17492
rect -1775 -17526 -1741 -17492
rect -1703 -17526 -1669 -17492
rect -1631 -17526 -1597 -17492
rect -1559 -17526 -1525 -17492
rect -1487 -17526 -1453 -17492
rect -1415 -17526 -1381 -17492
rect -1343 -17526 -1309 -17492
rect -1271 -17526 -1237 -17492
rect -1199 -17526 -1165 -17492
rect -1127 -17526 -1093 -17492
rect -1055 -17526 -1021 -17492
rect -983 -17526 -949 -17492
rect -911 -17526 -877 -17492
rect -839 -17526 -805 -17492
rect -767 -17526 -733 -17492
rect -695 -17526 -661 -17492
rect -623 -17526 -589 -17492
rect -551 -17526 -517 -17492
rect -479 -17526 -445 -17492
rect -407 -17526 -373 -17492
rect -335 -17526 -301 -17492
rect -263 -17526 -229 -17492
rect -191 -17526 -157 -17492
rect -119 -17526 -85 -17492
rect -47 -17526 -13 -17492
rect 25 -17526 59 -17492
rect 97 -17526 131 -17492
rect 169 -17526 203 -17492
rect 241 -17526 275 -17492
rect 313 -17526 347 -17492
rect 385 -17526 419 -17492
rect 457 -17526 491 -17492
rect 529 -17526 563 -17492
rect 601 -17526 635 -17492
rect 673 -17526 707 -17492
rect 745 -17526 779 -17492
rect 817 -17526 851 -17492
rect 889 -17526 923 -17492
rect 961 -17526 995 -17492
rect 1033 -17526 1067 -17492
rect 1105 -17526 1139 -17492
rect 1177 -17526 1211 -17492
rect 1249 -17526 1283 -17492
rect 1321 -17526 1355 -17492
rect 1393 -17526 1427 -17492
rect 1465 -17526 1499 -17492
rect 1537 -17526 1571 -17492
rect 1609 -17526 1643 -17492
rect 1681 -17526 1715 -17492
rect 1753 -17526 1787 -17492
rect 1825 -17526 1859 -17492
rect 1897 -17526 1931 -17492
rect 1969 -17526 2003 -17492
rect 2041 -17526 2075 -17492
rect 2113 -17526 2147 -17492
rect 2185 -17526 2219 -17492
rect 2257 -17526 2291 -17492
rect 2329 -17526 2363 -17492
rect 2401 -17526 2435 -17492
rect 2473 -17526 2507 -17492
rect 2545 -17526 2579 -17492
rect 2617 -17526 2651 -17492
rect 2689 -17526 2723 -17492
rect 2761 -17526 2795 -17492
rect 2833 -17526 2867 -17492
rect 2905 -17526 2939 -17492
rect 2977 -17526 3011 -17492
rect 3049 -17526 3083 -17492
rect 3121 -17526 3155 -17492
rect 3193 -17526 3227 -17492
rect 3265 -17526 3299 -17492
rect 3337 -17526 3371 -17492
rect 3409 -17526 3443 -17492
rect 3481 -17526 3515 -17492
rect 3553 -17526 3587 -17492
rect 3625 -17526 3659 -17492
rect 3697 -17526 3731 -17492
rect 3769 -17526 3803 -17492
rect 3841 -17526 3875 -17492
rect 3913 -17526 3947 -17492
rect 3985 -17526 4019 -17492
rect 4057 -17526 4091 -17492
rect 4129 -17526 4163 -17492
rect 4201 -17526 4235 -17492
rect 4273 -17526 4307 -17492
rect 4345 -17526 4379 -17492
rect 4417 -17526 4451 -17492
rect 4489 -17526 4523 -17492
rect 4561 -17526 4595 -17492
rect 4633 -17526 4667 -17492
rect 4705 -17526 4739 -17492
rect 4777 -17526 4811 -17492
rect 4849 -17526 4883 -17492
rect 4921 -17526 4955 -17492
rect 4993 -17526 5027 -17492
rect 5065 -17526 5099 -17492
rect 5137 -17526 5171 -17492
rect 5209 -17526 5243 -17492
rect 5281 -17526 5315 -17492
rect 5353 -17526 5387 -17492
rect 5425 -17526 5459 -17492
rect 5497 -17526 5531 -17492
rect 5569 -17526 5603 -17492
rect 5641 -17526 5675 -17492
rect 5713 -17526 5747 -17492
rect 5785 -17526 5819 -17492
rect 5857 -17526 5891 -17492
rect 5929 -17526 5963 -17492
rect 6001 -17526 6035 -17492
rect 6073 -17526 6107 -17492
rect 6145 -17526 6179 -17492
rect 6217 -17526 6251 -17492
rect 6289 -17526 6323 -17492
rect 6361 -17526 6395 -17492
rect 6433 -17526 6467 -17492
rect 6505 -17526 6539 -17492
rect 6577 -17526 6611 -17492
rect 6649 -17526 6683 -17492
rect 6721 -17526 6755 -17492
rect 6793 -17526 6827 -17492
rect 6865 -17526 6899 -17492
rect 6937 -17526 6971 -17492
rect 7009 -17526 7043 -17492
rect 7081 -17526 7115 -17492
rect 7153 -17526 7187 -17492
rect 7225 -17526 7259 -17492
rect 7297 -17526 7331 -17492
rect 7369 -17526 7403 -17492
rect 7441 -17526 7475 -17492
rect 7513 -17526 7547 -17492
rect 7585 -17526 7619 -17492
rect 7657 -17526 7691 -17492
rect 7729 -17526 7763 -17492
rect 7801 -17526 7835 -17492
rect 7873 -17526 7907 -17492
rect 7945 -17526 7979 -17492
rect 8017 -17526 8051 -17492
rect 8089 -17526 8123 -17492
rect 8161 -17526 8195 -17492
rect 8233 -17526 8267 -17492
rect 8305 -17526 8339 -17492
rect 8377 -17526 8411 -17492
rect 8449 -17526 8483 -17492
rect 8521 -17526 8555 -17492
rect 8593 -17526 8627 -17492
rect 8665 -17526 8699 -17492
rect 8737 -17526 8771 -17492
rect 8809 -17526 8843 -17492
rect 8881 -17526 8915 -17492
rect 8953 -17526 8987 -17492
rect 9025 -17526 9059 -17492
rect 9097 -17526 9131 -17492
rect 9169 -17526 9203 -17492
rect 9241 -17526 9275 -17492
rect 9313 -17526 9347 -17492
rect 9385 -17526 9419 -17492
rect 9457 -17526 9491 -17492
rect 9529 -17526 9563 -17492
rect 9601 -17526 9635 -17492
rect 9673 -17526 9707 -17492
rect 9745 -17526 9779 -17492
rect 9817 -17526 9851 -17492
rect 9889 -17526 9923 -17492
rect 9961 -17526 9995 -17492
rect 10033 -17526 10067 -17492
rect 10105 -17526 10139 -17492
rect 10177 -17526 10211 -17492
rect 10249 -17526 10283 -17492
rect 10321 -17526 10355 -17492
rect 10393 -17526 10427 -17492
rect 10465 -17526 10499 -17492
rect 10537 -17526 10571 -17492
rect 10609 -17526 10643 -17492
rect 10681 -17526 10715 -17492
rect 10753 -17526 10787 -17492
rect 10825 -17526 10859 -17492
rect 10897 -17526 10931 -17492
rect 10969 -17526 11003 -17492
rect 11041 -17526 11075 -17492
rect 11113 -17526 11147 -17492
rect 11185 -17526 11219 -17492
rect 11257 -17526 11291 -17492
rect 11329 -17526 11363 -17492
rect 11401 -17526 11435 -17492
rect 11473 -17526 11507 -17492
rect 11545 -17526 11579 -17492
rect 11617 -17526 11651 -17492
rect 11689 -17526 11723 -17492
rect 11761 -17526 11795 -17492
rect 11833 -17526 11867 -17492
rect 11905 -17526 11939 -17492
rect 11977 -17526 12011 -17492
rect 12049 -17526 12083 -17492
rect 12121 -17526 12155 -17492
rect 12193 -17526 12227 -17492
rect 12265 -17526 12299 -17492
rect 12337 -17526 12371 -17492
rect 12409 -17526 12443 -17492
rect 12481 -17526 12515 -17492
rect 12553 -17526 12587 -17492
rect 12625 -17526 12659 -17492
rect 12697 -17526 12731 -17492
rect 12769 -17526 12803 -17492
rect 12841 -17526 12875 -17492
rect 12913 -17526 12947 -17492
rect 12985 -17526 13019 -17492
rect 13057 -17526 13091 -17492
rect 13129 -17526 13163 -17492
rect 13201 -17526 13235 -17492
rect 13273 -17526 13307 -17492
rect 13345 -17526 13379 -17492
<< metal1 >>
rect 7034 2713 7080 2891
rect 16034 2713 16080 2891
rect 7034 1691 7080 1863
rect 16034 1691 16080 1863
rect 7034 913 7080 1091
rect 16034 913 16080 1091
rect 7034 -109 7080 63
rect 16034 -109 16080 63
rect 7034 -887 7080 -709
rect 16034 -887 16080 -709
rect -7605 -1290 3704 -1200
rect -7605 -1324 -7370 -1290
rect -7336 -1324 -7298 -1290
rect -7264 -1324 -7226 -1290
rect -7192 -1324 -7154 -1290
rect -7120 -1324 -7082 -1290
rect -7048 -1324 -7010 -1290
rect -6976 -1324 -6938 -1290
rect -6904 -1324 -6866 -1290
rect -6832 -1324 -6794 -1290
rect -6760 -1324 -6722 -1290
rect -6688 -1324 -6650 -1290
rect -6616 -1324 -6578 -1290
rect -6544 -1324 -6506 -1290
rect -6472 -1324 -6434 -1290
rect -6400 -1324 -6362 -1290
rect -6328 -1324 -6290 -1290
rect -6256 -1324 -6218 -1290
rect -6184 -1324 -6146 -1290
rect -6112 -1324 -6074 -1290
rect -6040 -1324 -6002 -1290
rect -5968 -1324 -5930 -1290
rect -5896 -1324 -5858 -1290
rect -5824 -1324 -5786 -1290
rect -5752 -1324 -5714 -1290
rect -5680 -1324 -5642 -1290
rect -5608 -1324 -5570 -1290
rect -5536 -1324 -5498 -1290
rect -5464 -1324 -5426 -1290
rect -5392 -1324 -5354 -1290
rect -5320 -1324 -5282 -1290
rect -5248 -1324 -5210 -1290
rect -5176 -1324 -5138 -1290
rect -5104 -1324 -5066 -1290
rect -5032 -1324 -4994 -1290
rect -4960 -1324 -4922 -1290
rect -4888 -1324 -4850 -1290
rect -4816 -1324 -4778 -1290
rect -4744 -1324 -4706 -1290
rect -4672 -1324 -4634 -1290
rect -4600 -1324 -4562 -1290
rect -4528 -1324 -4490 -1290
rect -4456 -1324 -4418 -1290
rect -4384 -1324 -4346 -1290
rect -4312 -1324 -4274 -1290
rect -4240 -1324 -4202 -1290
rect -4168 -1324 -4130 -1290
rect -4096 -1324 -4058 -1290
rect -4024 -1324 -3986 -1290
rect -3952 -1324 -3914 -1290
rect -3880 -1324 -3842 -1290
rect -3808 -1324 -3770 -1290
rect -3736 -1324 -3698 -1290
rect -3664 -1324 -3626 -1290
rect -3592 -1324 -3554 -1290
rect -3520 -1324 -3482 -1290
rect -3448 -1324 -3410 -1290
rect -3376 -1324 -3338 -1290
rect -3304 -1324 -3266 -1290
rect -3232 -1324 -3194 -1290
rect -3160 -1324 -3122 -1290
rect -3088 -1324 -3050 -1290
rect -3016 -1324 -2978 -1290
rect -2944 -1324 -2906 -1290
rect -2872 -1324 -2834 -1290
rect -2800 -1324 -2762 -1290
rect -2728 -1324 -2690 -1290
rect -2656 -1324 -2618 -1290
rect -2584 -1324 -2546 -1290
rect -2512 -1324 -2474 -1290
rect -2440 -1324 -2402 -1290
rect -2368 -1324 -2330 -1290
rect -2296 -1324 -2258 -1290
rect -2224 -1324 -2186 -1290
rect -2152 -1324 -2114 -1290
rect -2080 -1324 -2042 -1290
rect -2008 -1324 -1970 -1290
rect -1936 -1324 -1898 -1290
rect -1864 -1324 -1826 -1290
rect -1792 -1324 -1754 -1290
rect -1720 -1324 -1682 -1290
rect -1648 -1324 -1610 -1290
rect -1576 -1324 -1538 -1290
rect -1504 -1324 -1466 -1290
rect -1432 -1324 -1394 -1290
rect -1360 -1324 -1322 -1290
rect -1288 -1324 -1250 -1290
rect -1216 -1324 -1178 -1290
rect -1144 -1324 -1106 -1290
rect -1072 -1324 -1034 -1290
rect -1000 -1324 -962 -1290
rect -928 -1324 -890 -1290
rect -856 -1324 -818 -1290
rect -784 -1324 -746 -1290
rect -712 -1324 -674 -1290
rect -640 -1324 -602 -1290
rect -568 -1324 -530 -1290
rect -496 -1324 -458 -1290
rect -424 -1324 -386 -1290
rect -352 -1324 -314 -1290
rect -280 -1324 -242 -1290
rect -208 -1324 -170 -1290
rect -136 -1324 -98 -1290
rect -64 -1324 -26 -1290
rect 8 -1324 46 -1290
rect 80 -1324 118 -1290
rect 152 -1324 190 -1290
rect 224 -1324 262 -1290
rect 296 -1324 334 -1290
rect 368 -1324 406 -1290
rect 440 -1324 478 -1290
rect 512 -1324 550 -1290
rect 584 -1324 622 -1290
rect 656 -1324 694 -1290
rect 728 -1324 766 -1290
rect 800 -1324 838 -1290
rect 872 -1324 910 -1290
rect 944 -1324 982 -1290
rect 1016 -1324 1054 -1290
rect 1088 -1324 1126 -1290
rect 1160 -1324 1198 -1290
rect 1232 -1324 1270 -1290
rect 1304 -1324 1342 -1290
rect 1376 -1324 1414 -1290
rect 1448 -1324 1486 -1290
rect 1520 -1324 1558 -1290
rect 1592 -1324 1630 -1290
rect 1664 -1324 1702 -1290
rect 1736 -1324 1774 -1290
rect 1808 -1324 1846 -1290
rect 1880 -1324 1918 -1290
rect 1952 -1324 1990 -1290
rect 2024 -1324 2062 -1290
rect 2096 -1324 2134 -1290
rect 2168 -1324 2206 -1290
rect 2240 -1324 2278 -1290
rect 2312 -1324 2350 -1290
rect 2384 -1324 2422 -1290
rect 2456 -1324 2494 -1290
rect 2528 -1324 2566 -1290
rect 2600 -1324 2638 -1290
rect 2672 -1324 2710 -1290
rect 2744 -1324 2782 -1290
rect 2816 -1324 2854 -1290
rect 2888 -1324 2926 -1290
rect 2960 -1324 2998 -1290
rect 3032 -1324 3070 -1290
rect 3104 -1324 3142 -1290
rect 3176 -1324 3214 -1290
rect 3248 -1324 3286 -1290
rect 3320 -1324 3704 -1290
rect -7605 -1467 3704 -1324
rect -5132 -1741 -4948 -1467
rect -5945 -1841 -3776 -1741
rect -5945 -2039 -5911 -1841
rect -5877 -1911 -5804 -1910
rect -5877 -1963 -5867 -1911
rect -5815 -1963 -5804 -1911
rect -5699 -1911 -5626 -1910
rect -5699 -1963 -5689 -1911
rect -5637 -1963 -5626 -1911
rect -5520 -1911 -5447 -1910
rect -5520 -1963 -5510 -1911
rect -5458 -1963 -5447 -1911
rect -5343 -1911 -5270 -1910
rect -5343 -1963 -5333 -1911
rect -5281 -1963 -5270 -1911
rect -5165 -1911 -5092 -1910
rect -5165 -1963 -5155 -1911
rect -5103 -1963 -5092 -1911
rect -4986 -1911 -4913 -1910
rect -4986 -1963 -4976 -1911
rect -4924 -1963 -4913 -1911
rect -4809 -1911 -4736 -1910
rect -4809 -1963 -4799 -1911
rect -4747 -1963 -4736 -1911
rect -4631 -1911 -4558 -1910
rect -4631 -1963 -4621 -1911
rect -4569 -1963 -4558 -1911
rect -4453 -1911 -4380 -1910
rect -4453 -1963 -4443 -1911
rect -4391 -1963 -4380 -1911
rect -4275 -1911 -4202 -1910
rect -4275 -1963 -4265 -1911
rect -4213 -1963 -4202 -1911
rect -4096 -1911 -4023 -1910
rect -4096 -1963 -4086 -1911
rect -4034 -1963 -4023 -1911
rect -3919 -1911 -3846 -1910
rect -3919 -1963 -3909 -1911
rect -3857 -1963 -3846 -1911
rect -6302 -2073 -5911 -2039
rect -6302 -2135 -6268 -2073
rect -6126 -2150 -6092 -2073
rect -5945 -2132 -5911 -2073
rect -5857 -2079 -5823 -1963
rect -5679 -2079 -5645 -1963
rect -5501 -2079 -5467 -1963
rect -5322 -2079 -5288 -1963
rect -5145 -2079 -5111 -1963
rect -4967 -2079 -4933 -1963
rect -4789 -2079 -4755 -1963
rect -4611 -2079 -4577 -1963
rect -4433 -2079 -4399 -1963
rect -4255 -2079 -4221 -1963
rect -4077 -2079 -4043 -1963
rect -3898 -2079 -3864 -1963
rect -3810 -2133 -3776 -1841
rect -1119 -1911 -1046 -1910
rect -1119 -1963 -1109 -1911
rect -1057 -1963 -1046 -1911
rect -6508 -2530 -6435 -2529
rect -6508 -2582 -6498 -2530
rect -6446 -2582 -6435 -2530
rect -6635 -3402 -6562 -3401
rect -6635 -3454 -6625 -3402
rect -6573 -3454 -6562 -3402
rect -6625 -5322 -6572 -3454
rect -6498 -3640 -6445 -2582
rect -6054 -2781 -5981 -2780
rect -6054 -2833 -6044 -2781
rect -5992 -2833 -5981 -2781
rect -6302 -2945 -6090 -2911
rect -6302 -3020 -6268 -2945
rect -6124 -3022 -6090 -2945
rect -6035 -2949 -6001 -2833
rect -6124 -3401 -6090 -3259
rect -6144 -3402 -6071 -3401
rect -6144 -3454 -6134 -3402
rect -6082 -3454 -6071 -3402
rect -6508 -3641 -6435 -3640
rect -6508 -3693 -6498 -3641
rect -6446 -3693 -6435 -3641
rect -6498 -4271 -6445 -3693
rect -6302 -3812 -6090 -3778
rect -6302 -3889 -6268 -3812
rect -6124 -3888 -6090 -3812
rect -6035 -3819 -6001 -3311
rect -6508 -4272 -6435 -4271
rect -6508 -4324 -6498 -4272
rect -6446 -4324 -6435 -4272
rect -6498 -5141 -6445 -4324
rect -6124 -4390 -6090 -4128
rect -6144 -4391 -6071 -4390
rect -6144 -4443 -6134 -4391
rect -6082 -4443 -6071 -4391
rect -6302 -4683 -6090 -4649
rect -6302 -4763 -6268 -4683
rect -6124 -4761 -6090 -4683
rect -6035 -4689 -6001 -4181
rect -6508 -5142 -6435 -5141
rect -6508 -5194 -6498 -5142
rect -6446 -5194 -6435 -5142
rect -6635 -5323 -6562 -5322
rect -6635 -5375 -6625 -5323
rect -6573 -5375 -6562 -5323
rect -6498 -6248 -6445 -5194
rect -6124 -5232 -6090 -4998
rect -6144 -5233 -6071 -5232
rect -6144 -5285 -6134 -5233
rect -6082 -5285 -6071 -5233
rect -6301 -5519 -6091 -5518
rect -5946 -5519 -5912 -2388
rect -5856 -2780 -5822 -2447
rect -5768 -2530 -5734 -2389
rect -5787 -2531 -5714 -2530
rect -5787 -2583 -5777 -2531
rect -5725 -2583 -5714 -2531
rect -5876 -2781 -5803 -2780
rect -5876 -2833 -5866 -2781
rect -5814 -2833 -5803 -2781
rect -5856 -2943 -5822 -2833
rect -5679 -2949 -5645 -2447
rect -5857 -3819 -5823 -3311
rect -5768 -3516 -5734 -3258
rect -5787 -3517 -5714 -3516
rect -5787 -3569 -5777 -3517
rect -5725 -3569 -5714 -3517
rect -5679 -3819 -5645 -3311
rect -5857 -4689 -5823 -4181
rect -5768 -4271 -5734 -4128
rect -5788 -4272 -5715 -4271
rect -5788 -4324 -5778 -4272
rect -5726 -4324 -5715 -4272
rect -5679 -4689 -5645 -4181
rect -6301 -5552 -5912 -5519
rect -6301 -5636 -6267 -5552
rect -6125 -5553 -5912 -5552
rect -6125 -5639 -6091 -5553
rect -5946 -5612 -5912 -5553
rect -5857 -5559 -5823 -5051
rect -5768 -5415 -5734 -4999
rect -5787 -5416 -5714 -5415
rect -5787 -5468 -5777 -5416
rect -5725 -5468 -5714 -5416
rect -5679 -5559 -5645 -5051
rect -5590 -5612 -5556 -2388
rect -5501 -2949 -5467 -2441
rect -5412 -2668 -5378 -2388
rect -5431 -2669 -5358 -2668
rect -5431 -2721 -5421 -2669
rect -5369 -2721 -5358 -2669
rect -5323 -2949 -5289 -2441
rect -5501 -3819 -5467 -3311
rect -5412 -3640 -5378 -3258
rect -5432 -3641 -5359 -3640
rect -5432 -3693 -5422 -3641
rect -5370 -3693 -5359 -3641
rect -5323 -3819 -5289 -3311
rect -5501 -4689 -5467 -4181
rect -5412 -4506 -5378 -4128
rect -5432 -4507 -5359 -4506
rect -5432 -4559 -5422 -4507
rect -5370 -4559 -5359 -4507
rect -5323 -4689 -5289 -4181
rect -5501 -5559 -5467 -5051
rect -5412 -5141 -5378 -4998
rect -5432 -5142 -5359 -5141
rect -5432 -5194 -5422 -5142
rect -5370 -5194 -5359 -5142
rect -5323 -5559 -5289 -5051
rect -5234 -5612 -5200 -2388
rect -5145 -2949 -5111 -2441
rect -5056 -2530 -5022 -2388
rect -5076 -2531 -5003 -2530
rect -5076 -2583 -5066 -2531
rect -5014 -2583 -5003 -2531
rect -4967 -2949 -4933 -2441
rect -5145 -3819 -5111 -3311
rect -5056 -3401 -5022 -3259
rect -5076 -3402 -5003 -3401
rect -5076 -3454 -5066 -3402
rect -5014 -3454 -5003 -3402
rect -4967 -3819 -4933 -3311
rect -5145 -4689 -5111 -4181
rect -5056 -4390 -5022 -4127
rect -5076 -4391 -5003 -4390
rect -5076 -4443 -5066 -4391
rect -5014 -4443 -5003 -4391
rect -4967 -4689 -4933 -4181
rect -5145 -5559 -5111 -5051
rect -5056 -5233 -5022 -4998
rect -5076 -5234 -5003 -5233
rect -5076 -5286 -5066 -5234
rect -5014 -5286 -5003 -5234
rect -4967 -5559 -4933 -5051
rect -4878 -5612 -4844 -2388
rect -4789 -2949 -4755 -2441
rect -4700 -2668 -4666 -2388
rect -4720 -2669 -4647 -2668
rect -4720 -2721 -4710 -2669
rect -4658 -2721 -4647 -2669
rect -4611 -2949 -4577 -2441
rect -4789 -3819 -4755 -3311
rect -4700 -3401 -4666 -3258
rect -4720 -3402 -4647 -3401
rect -4720 -3454 -4710 -3402
rect -4658 -3454 -4647 -3402
rect -4611 -3819 -4577 -3311
rect -4789 -4689 -4755 -4181
rect -4700 -4390 -4666 -4128
rect -4719 -4391 -4646 -4390
rect -4719 -4443 -4709 -4391
rect -4657 -4443 -4646 -4391
rect -4611 -4689 -4577 -4181
rect -4789 -5559 -4755 -5051
rect -4700 -5322 -4666 -4998
rect -4720 -5323 -4647 -5322
rect -4720 -5375 -4710 -5323
rect -4658 -5375 -4647 -5323
rect -4611 -5559 -4577 -5051
rect -4522 -5612 -4488 -2388
rect -4433 -2949 -4399 -2441
rect -4344 -2530 -4310 -2388
rect -4364 -2531 -4291 -2530
rect -4364 -2583 -4354 -2531
rect -4302 -2583 -4291 -2531
rect -4255 -2949 -4221 -2441
rect -4433 -3819 -4399 -3311
rect -4344 -3640 -4310 -3258
rect -4363 -3641 -4290 -3640
rect -4363 -3693 -4353 -3641
rect -4301 -3693 -4290 -3641
rect -4254 -3819 -4220 -3311
rect -4433 -4689 -4399 -4181
rect -4344 -4506 -4310 -4128
rect -4363 -4507 -4290 -4506
rect -4363 -4559 -4353 -4507
rect -4301 -4559 -4290 -4507
rect -4255 -4689 -4221 -4181
rect -4433 -5559 -4399 -5051
rect -4344 -5141 -4310 -4998
rect -4363 -5142 -4290 -5141
rect -4363 -5194 -4353 -5142
rect -4301 -5194 -4290 -5142
rect -4255 -5559 -4221 -5051
rect -4166 -5612 -4132 -2388
rect -4077 -2949 -4043 -2441
rect -3988 -2668 -3954 -2388
rect -4008 -2669 -3935 -2668
rect -4008 -2721 -3998 -2669
rect -3946 -2721 -3935 -2669
rect -3899 -2780 -3865 -2441
rect -3810 -2446 -3776 -2388
rect -3633 -2446 -3599 -2364
rect -3454 -2446 -3420 -2370
rect -1099 -2425 -1065 -1963
rect -3810 -2480 -3420 -2446
rect -1119 -2426 -1046 -2425
rect -1119 -2478 -1109 -2426
rect -1057 -2478 -1046 -2426
rect -762 -2426 -689 -2425
rect -762 -2478 -752 -2426
rect -700 -2478 -689 -2426
rect -3918 -2781 -3845 -2780
rect -3918 -2833 -3908 -2781
rect -3856 -2833 -3845 -2781
rect -3899 -2949 -3865 -2833
rect -4077 -3819 -4043 -3311
rect -3988 -3516 -3954 -3258
rect -4008 -3517 -3935 -3516
rect -4008 -3569 -3998 -3517
rect -3946 -3569 -3935 -3517
rect -3899 -3819 -3865 -3311
rect -4077 -4689 -4043 -4181
rect -3988 -4271 -3954 -4128
rect -4008 -4272 -3935 -4271
rect -4008 -4324 -3998 -4272
rect -3946 -4324 -3935 -4272
rect -3899 -4689 -3865 -4181
rect -4077 -5559 -4043 -5051
rect -3988 -5415 -3954 -4998
rect -4007 -5416 -3934 -5415
rect -4007 -5468 -3997 -5416
rect -3945 -5468 -3934 -5416
rect -3899 -5559 -3865 -5051
rect -3810 -5612 -3776 -2480
rect -2634 -2559 -2561 -2558
rect -2634 -2611 -2624 -2559
rect -2572 -2611 -2561 -2559
rect -1295 -2559 -1222 -2558
rect -1295 -2611 -1285 -2559
rect -1233 -2611 -1222 -2559
rect -3308 -2669 -3235 -2668
rect -3308 -2721 -3298 -2669
rect -3246 -2721 -3235 -2669
rect -3741 -2781 -3668 -2780
rect -3741 -2833 -3731 -2781
rect -3679 -2833 -3668 -2781
rect -3721 -2949 -3687 -2833
rect -3721 -3819 -3687 -3311
rect -3632 -3316 -3598 -3258
rect -3454 -3316 -3420 -3234
rect -3632 -3350 -3420 -3316
rect -3632 -3401 -3598 -3350
rect -3652 -3402 -3579 -3401
rect -3652 -3454 -3642 -3402
rect -3590 -3454 -3579 -3402
rect -3298 -3516 -3245 -2721
rect -3141 -3402 -3068 -3401
rect -3141 -3454 -3131 -3402
rect -3079 -3454 -3068 -3402
rect -3308 -3517 -3235 -3516
rect -3308 -3569 -3298 -3517
rect -3246 -3569 -3235 -3517
rect -3721 -4689 -3687 -4181
rect -3632 -4186 -3598 -4128
rect -3453 -4186 -3419 -4076
rect -3632 -4220 -3419 -4186
rect -3632 -4390 -3598 -4220
rect -3652 -4391 -3579 -4390
rect -3652 -4443 -3642 -4391
rect -3590 -4443 -3579 -4391
rect -3298 -4506 -3245 -3569
rect -3308 -4507 -3235 -4506
rect -3308 -4559 -3298 -4507
rect -3246 -4559 -3235 -4507
rect -3632 -5056 -3598 -4999
rect -3453 -5056 -3419 -4946
rect -3632 -5090 -3419 -5056
rect -3632 -5319 -3598 -5090
rect -3652 -5320 -3579 -5319
rect -3652 -5372 -3642 -5320
rect -3590 -5372 -3579 -5320
rect -3298 -5416 -3245 -4559
rect -3130 -5233 -3077 -3454
rect -3140 -5234 -3067 -5233
rect -3140 -5286 -3130 -5234
rect -3078 -5286 -3067 -5234
rect -2624 -5324 -2571 -2611
rect -1276 -2885 -1242 -2611
rect -1207 -2666 -1134 -2665
rect -1207 -2718 -1197 -2666
rect -1145 -2718 -1134 -2666
rect -1187 -2825 -1153 -2718
rect -1099 -2884 -1065 -2478
rect -940 -2559 -867 -2558
rect -940 -2611 -930 -2559
rect -878 -2611 -867 -2559
rect -1029 -2666 -956 -2665
rect -1029 -2718 -1019 -2666
rect -967 -2718 -956 -2666
rect -1009 -2831 -975 -2718
rect -920 -2886 -886 -2611
rect -851 -2666 -778 -2665
rect -851 -2718 -841 -2666
rect -789 -2718 -778 -2666
rect -831 -2831 -797 -2718
rect -742 -2884 -708 -2478
rect -208 -2605 182 -2571
rect -208 -2883 -174 -2605
rect -139 -2666 -66 -2665
rect -139 -2718 -129 -2666
rect -77 -2718 -66 -2666
rect 40 -2666 113 -2665
rect 40 -2718 50 -2666
rect 102 -2718 113 -2666
rect -119 -2831 -85 -2718
rect 59 -2831 93 -2718
rect 148 -2886 182 -2605
rect 217 -2666 290 -2665
rect 217 -2718 227 -2666
rect 279 -2718 290 -2666
rect 237 -2831 271 -2718
rect 594 -2825 628 -1467
rect 7034 -1909 7080 -1737
rect 16034 -1909 16080 -1737
rect 6670 -2205 6754 -2199
rect 5327 -2206 5400 -2205
rect 5327 -2258 5337 -2206
rect 5389 -2258 5400 -2206
rect 6670 -2257 6686 -2205
rect 6738 -2257 6754 -2205
rect 1909 -2427 1982 -2426
rect 1909 -2479 1919 -2427
rect 1971 -2479 1982 -2427
rect 2265 -2427 2338 -2426
rect 2265 -2479 2275 -2427
rect 2327 -2479 2338 -2427
rect 3183 -2428 3256 -2427
rect 1038 -2611 1428 -2577
rect 930 -2666 1003 -2665
rect 930 -2718 940 -2666
rect 992 -2718 1003 -2666
rect 949 -2831 983 -2718
rect 1038 -2886 1072 -2611
rect 1107 -2666 1180 -2665
rect 1107 -2718 1117 -2666
rect 1169 -2718 1180 -2666
rect 1285 -2666 1358 -2665
rect 1285 -2718 1295 -2666
rect 1347 -2718 1358 -2666
rect 1127 -2831 1161 -2718
rect 1305 -2831 1339 -2718
rect -1454 -3282 -1420 -3140
rect -1365 -3282 -1331 -3199
rect -1276 -3282 -1242 -3141
rect -1454 -3316 -1242 -3282
rect -1454 -3317 -1420 -3316
rect -1655 -3454 -1574 -3449
rect -1655 -3506 -1641 -3454
rect -1589 -3506 -1574 -3454
rect -1655 -3510 -1574 -3506
rect -2014 -4413 -1941 -4412
rect -2014 -4465 -2004 -4413
rect -1952 -4465 -1941 -4413
rect -2003 -4517 -1950 -4465
rect -2634 -5325 -2561 -5324
rect -2634 -5377 -2624 -5325
rect -2572 -5377 -2561 -5325
rect -3308 -5417 -3235 -5416
rect -3308 -5469 -3298 -5417
rect -3246 -5469 -3235 -5417
rect -5946 -6016 -5912 -5869
rect -5966 -6017 -5893 -6016
rect -5966 -6069 -5956 -6017
rect -5904 -6069 -5893 -6017
rect -5768 -6131 -5734 -5868
rect -5590 -6016 -5556 -5868
rect -5611 -6017 -5538 -6016
rect -5611 -6069 -5601 -6017
rect -5549 -6069 -5538 -6017
rect -5788 -6132 -5715 -6131
rect -5788 -6184 -5778 -6132
rect -5726 -6184 -5715 -6132
rect -5412 -6248 -5378 -5868
rect -5234 -6016 -5200 -5868
rect -5254 -6017 -5181 -6016
rect -5254 -6069 -5244 -6017
rect -5192 -6069 -5181 -6017
rect -5056 -6131 -5022 -5869
rect -5075 -6132 -5002 -6131
rect -5075 -6184 -5065 -6132
rect -5013 -6184 -5002 -6132
rect -6508 -6249 -6435 -6248
rect -6508 -6301 -6498 -6249
rect -6446 -6301 -6435 -6249
rect -5431 -6249 -5358 -6248
rect -5431 -6301 -5421 -6249
rect -5369 -6301 -5358 -6249
rect -4967 -6376 -4933 -5927
rect -4878 -6016 -4844 -5868
rect -4898 -6017 -4825 -6016
rect -4898 -6069 -4888 -6017
rect -4836 -6069 -4825 -6017
rect -4700 -6248 -4666 -5868
rect -4720 -6249 -4647 -6248
rect -4720 -6301 -4710 -6249
rect -4658 -6301 -4647 -6249
rect -4613 -6376 -4579 -5921
rect -4522 -6016 -4488 -5868
rect -4542 -6017 -4469 -6016
rect -4542 -6069 -4532 -6017
rect -4480 -6069 -4469 -6017
rect -4344 -6131 -4310 -5868
rect -4166 -6016 -4132 -5868
rect -4185 -6017 -4112 -6016
rect -4185 -6069 -4175 -6017
rect -4123 -6069 -4112 -6017
rect -4364 -6132 -4291 -6131
rect -4364 -6184 -4354 -6132
rect -4302 -6184 -4291 -6132
rect -3988 -6247 -3954 -5868
rect -3810 -5928 -3776 -5868
rect -3632 -5928 -3598 -5836
rect -3455 -5928 -3421 -5814
rect -3810 -5962 -3421 -5928
rect -3810 -6016 -3776 -5962
rect -3830 -6017 -3757 -6016
rect -3830 -6069 -3820 -6017
rect -3768 -6069 -3757 -6017
rect -3298 -6131 -3245 -5469
rect -2624 -6007 -2571 -5377
rect -2634 -6008 -2561 -6007
rect -2634 -6060 -2624 -6008
rect -2572 -6060 -2561 -6008
rect -3308 -6132 -3235 -6131
rect -3308 -6184 -3298 -6132
rect -3246 -6184 -3235 -6132
rect -4008 -6248 -3935 -6247
rect -4008 -6300 -3998 -6248
rect -3946 -6300 -3935 -6248
rect -3988 -6301 -3954 -6300
rect -4967 -6379 -4579 -6376
rect -4967 -6410 -4786 -6379
rect -4796 -6431 -4786 -6410
rect -4734 -6410 -4579 -6379
rect -4734 -6431 -4723 -6410
rect -2002 -6714 -1950 -4517
rect -1886 -5233 -1813 -5232
rect -1886 -5285 -1876 -5233
rect -1824 -5285 -1813 -5233
rect -1646 -5278 -1585 -3510
rect -1296 -3572 -1223 -3571
rect -1296 -3624 -1286 -3572
rect -1234 -3624 -1223 -3572
rect -1276 -3784 -1242 -3624
rect -1186 -3724 -1152 -3200
rect -1118 -3457 -1045 -3456
rect -1118 -3509 -1108 -3457
rect -1056 -3509 -1045 -3457
rect -1098 -3784 -1064 -3509
rect -1009 -3724 -975 -3200
rect -939 -3572 -866 -3571
rect -939 -3624 -929 -3572
rect -877 -3624 -866 -3572
rect -919 -3784 -885 -3624
rect -831 -3724 -797 -3200
rect -653 -3282 -619 -3199
rect -563 -3282 -529 -3140
rect -474 -3282 -440 -3199
rect -385 -3282 -351 -3140
rect -295 -3282 -261 -3199
rect -653 -3302 -261 -3282
rect -653 -3316 -484 -3302
rect -494 -3354 -484 -3316
rect -432 -3316 -261 -3302
rect -432 -3354 -421 -3316
rect -760 -3457 -687 -3456
rect -760 -3509 -750 -3457
rect -698 -3509 -687 -3457
rect -406 -3457 -333 -3456
rect -406 -3509 -396 -3457
rect -344 -3509 -333 -3457
rect -742 -3784 -708 -3509
rect -583 -3572 -510 -3571
rect -583 -3624 -573 -3572
rect -521 -3624 -510 -3572
rect -564 -3784 -530 -3624
rect -386 -3784 -352 -3509
rect -208 -3571 -174 -3140
rect -227 -3572 -154 -3571
rect -227 -3624 -217 -3572
rect -165 -3624 -154 -3572
rect -208 -3784 -174 -3624
rect -119 -3724 -85 -3200
rect -30 -3456 4 -3138
rect 327 -3456 361 -3139
rect 414 -3283 448 -3199
rect 504 -3283 538 -3141
rect 592 -3283 626 -3199
rect 682 -3283 716 -3141
rect 771 -3283 805 -3199
rect 414 -3302 805 -3283
rect 414 -3317 583 -3302
rect 573 -3354 583 -3317
rect 635 -3317 805 -3302
rect 635 -3354 646 -3317
rect -49 -3457 24 -3456
rect -49 -3509 -39 -3457
rect 13 -3509 24 -3457
rect 307 -3457 380 -3456
rect 307 -3509 317 -3457
rect 369 -3509 380 -3457
rect -30 -3784 4 -3509
rect 589 -3598 623 -3354
rect 860 -3456 894 -3139
rect 1216 -3456 1250 -3136
rect 840 -3457 913 -3456
rect 840 -3509 850 -3457
rect 902 -3509 913 -3457
rect 1196 -3457 1269 -3456
rect 1196 -3509 1206 -3457
rect 1258 -3509 1269 -3457
rect 59 -3632 1160 -3598
rect 59 -3725 93 -3632
rect 149 -3633 271 -3632
rect 149 -3784 183 -3633
rect 237 -3725 271 -3633
rect 948 -3725 982 -3632
rect 1038 -3783 1072 -3632
rect 1126 -3725 1160 -3632
rect 1216 -3802 1250 -3509
rect 1306 -3724 1340 -3200
rect 1394 -3564 1428 -2611
rect 1928 -2885 1962 -2479
rect 2087 -2555 2160 -2554
rect 2087 -2607 2097 -2555
rect 2149 -2607 2160 -2555
rect 1997 -2666 2070 -2665
rect 1997 -2718 2007 -2666
rect 2059 -2718 2070 -2666
rect 2017 -2831 2051 -2718
rect 2105 -2881 2139 -2607
rect 2176 -2666 2249 -2665
rect 2176 -2718 2186 -2666
rect 2238 -2718 2249 -2666
rect 2195 -2831 2229 -2718
rect 2285 -2887 2319 -2479
rect 3183 -2480 3193 -2428
rect 3245 -2480 3256 -2428
rect 2443 -2555 2931 -2554
rect 2443 -2607 2453 -2555
rect 2505 -2606 2931 -2555
rect 2505 -2607 2516 -2606
rect 2353 -2666 2426 -2665
rect 2353 -2718 2363 -2666
rect 2415 -2718 2426 -2666
rect 2373 -2831 2407 -2718
rect 2462 -2885 2496 -2607
rect 1482 -3283 1516 -3199
rect 1572 -3283 1606 -3140
rect 1662 -3283 1696 -3199
rect 1750 -3283 1784 -3140
rect 1840 -3283 1874 -3199
rect 1482 -3302 1874 -3283
rect 1482 -3317 1654 -3302
rect 1644 -3354 1654 -3317
rect 1706 -3317 1874 -3302
rect 1706 -3354 1717 -3317
rect 1552 -3457 1625 -3456
rect 1552 -3509 1562 -3457
rect 1614 -3509 1625 -3457
rect 1909 -3457 1982 -3456
rect 1909 -3509 1919 -3457
rect 1971 -3509 1982 -3457
rect 1374 -3565 1447 -3564
rect 1374 -3617 1384 -3565
rect 1436 -3617 1447 -3565
rect 1394 -3809 1428 -3617
rect 1572 -3784 1606 -3509
rect 1731 -3565 1804 -3564
rect 1731 -3617 1741 -3565
rect 1793 -3617 1804 -3565
rect 1750 -3786 1784 -3617
rect 1929 -3787 1963 -3509
rect 2017 -3724 2051 -3200
rect 2087 -3565 2160 -3564
rect 2087 -3617 2097 -3565
rect 2149 -3617 2160 -3565
rect 2106 -3785 2140 -3617
rect 2196 -3724 2230 -3200
rect 2265 -3457 2338 -3456
rect 2265 -3509 2275 -3457
rect 2327 -3509 2338 -3457
rect 2284 -3785 2318 -3509
rect 2373 -3724 2407 -3200
rect 2462 -3284 2496 -3141
rect 2551 -3284 2585 -3199
rect 2641 -3284 2675 -3141
rect 2462 -3318 2675 -3284
rect 2441 -3565 2514 -3564
rect 2441 -3617 2451 -3565
rect 2503 -3617 2514 -3565
rect 2462 -3786 2496 -3617
rect -1454 -4184 -1420 -4041
rect -1366 -4184 -1332 -4099
rect -1276 -4184 -1242 -4040
rect -1454 -4218 -1242 -4184
rect -1454 -4541 -1242 -4507
rect -1454 -4685 -1420 -4541
rect -1365 -4624 -1331 -4541
rect -1276 -4706 -1242 -4541
rect -1187 -4625 -1153 -4101
rect -1009 -4624 -975 -4100
rect -831 -4192 -797 -4100
rect -653 -4192 -619 -4101
rect -474 -4192 -440 -4101
rect -297 -4192 -263 -4100
rect -851 -4193 -778 -4192
rect -851 -4245 -841 -4193
rect -789 -4245 -778 -4193
rect -672 -4193 -599 -4192
rect -672 -4245 -662 -4193
rect -610 -4245 -599 -4193
rect -493 -4193 -420 -4192
rect -493 -4245 -483 -4193
rect -431 -4245 -420 -4193
rect -316 -4193 -243 -4192
rect -316 -4245 -306 -4193
rect -254 -4245 -243 -4193
rect -831 -4624 -797 -4245
rect -653 -4625 -619 -4245
rect -474 -4625 -440 -4245
rect -297 -4624 -263 -4245
rect -119 -4624 -85 -4100
rect -1277 -5097 -1243 -4939
rect -1297 -5098 -1224 -5097
rect -1297 -5150 -1287 -5098
rect -1235 -5150 -1224 -5098
rect -1656 -5283 -1575 -5278
rect -1876 -5337 -1823 -5285
rect -1875 -6364 -1823 -5337
rect -1656 -5335 -1642 -5283
rect -1590 -5335 -1575 -5283
rect -1656 -5339 -1575 -5335
rect -1454 -5442 -1242 -5408
rect -1454 -5585 -1420 -5442
rect -1363 -5524 -1329 -5442
rect -1276 -5592 -1242 -5442
rect -1187 -5525 -1153 -4995
rect -1097 -5213 -1063 -4938
rect -1115 -5214 -1042 -5213
rect -1115 -5266 -1105 -5214
rect -1053 -5266 -1042 -5214
rect -1009 -5524 -975 -4994
rect -919 -5097 -885 -4937
rect -939 -5098 -866 -5097
rect -939 -5150 -929 -5098
rect -877 -5150 -866 -5098
rect -830 -5524 -796 -4994
rect -741 -5213 -707 -4937
rect -563 -5097 -529 -4940
rect -582 -5098 -509 -5097
rect -582 -5150 -572 -5098
rect -520 -5150 -509 -5098
rect -386 -5213 -352 -4937
rect -208 -5097 -174 -4910
rect -228 -5098 -155 -5097
rect -228 -5150 -218 -5098
rect -166 -5150 -155 -5098
rect -761 -5214 -688 -5213
rect -761 -5266 -751 -5214
rect -699 -5266 -688 -5214
rect -406 -5214 -333 -5213
rect -406 -5266 -396 -5214
rect -344 -5266 -333 -5214
rect -654 -5434 -262 -5400
rect -654 -5523 -620 -5434
rect -563 -5604 -529 -5434
rect -474 -5524 -440 -5434
rect -385 -5612 -351 -5434
rect -296 -5524 -262 -5434
rect -1274 -6364 -1240 -5839
rect -1886 -6365 -1813 -6364
rect -1886 -6417 -1876 -6365
rect -1824 -6417 -1813 -6365
rect -1292 -6365 -1219 -6364
rect -1292 -6417 -1282 -6365
rect -1230 -6417 -1219 -6365
rect -1099 -6479 -1065 -5845
rect -919 -6365 -885 -5833
rect -938 -6417 -928 -6365
rect -876 -6417 -866 -6365
rect -742 -6479 -708 -5839
rect -1120 -6480 -1047 -6479
rect -1120 -6532 -1110 -6480
rect -1058 -6532 -1047 -6480
rect -762 -6480 -689 -6479
rect -762 -6532 -752 -6480
rect -700 -6532 -689 -6480
rect -476 -6493 -442 -5901
rect -208 -6077 -174 -5150
rect -119 -5380 -85 -4994
rect -30 -5213 4 -4938
rect 59 -5091 93 -4992
rect 148 -5091 182 -3952
rect 326 -4304 360 -4040
rect 416 -4192 450 -4094
rect 397 -4193 470 -4192
rect 397 -4245 407 -4193
rect 459 -4245 470 -4193
rect 307 -4305 380 -4304
rect 307 -4357 317 -4305
rect 369 -4357 380 -4305
rect 326 -4706 360 -4357
rect 416 -4624 450 -4245
rect 504 -4412 538 -4040
rect 593 -4192 627 -4101
rect 573 -4193 646 -4192
rect 573 -4245 583 -4193
rect 635 -4245 646 -4193
rect 485 -4413 558 -4412
rect 485 -4465 495 -4413
rect 547 -4465 558 -4413
rect 504 -4703 538 -4465
rect 593 -4625 627 -4245
rect 682 -4304 716 -4040
rect 771 -4192 805 -4100
rect 751 -4193 824 -4192
rect 751 -4245 761 -4193
rect 813 -4245 824 -4193
rect 663 -4305 736 -4304
rect 663 -4357 673 -4305
rect 725 -4357 736 -4305
rect 682 -4687 716 -4357
rect 771 -4624 805 -4245
rect 860 -4412 894 -4040
rect 840 -4413 913 -4412
rect 840 -4465 850 -4413
rect 902 -4465 913 -4413
rect 860 -4716 894 -4465
rect 236 -5091 270 -4999
rect 948 -5091 982 -5000
rect 1039 -5091 1073 -3989
rect 1305 -4624 1339 -4094
rect 1484 -4192 1518 -4094
rect 1661 -4192 1695 -4094
rect 1839 -4192 1873 -4094
rect 2017 -4192 2051 -4094
rect 1464 -4193 1537 -4192
rect 1464 -4245 1474 -4193
rect 1526 -4245 1537 -4193
rect 1642 -4193 1715 -4192
rect 1642 -4245 1652 -4193
rect 1704 -4245 1715 -4193
rect 1820 -4193 1893 -4192
rect 1820 -4245 1830 -4193
rect 1882 -4245 1893 -4193
rect 1998 -4193 2071 -4192
rect 1998 -4245 2008 -4193
rect 2060 -4245 2071 -4193
rect 1484 -4624 1518 -4245
rect 1661 -4624 1695 -4245
rect 1839 -4624 1873 -4245
rect 2017 -4624 2051 -4245
rect 2195 -4625 2229 -4095
rect 2373 -4624 2407 -4094
rect 2463 -4182 2497 -4038
rect 2552 -4182 2586 -4104
rect 2640 -4180 2674 -4020
rect 2640 -4182 2792 -4180
rect 2463 -4214 2792 -4182
rect 2463 -4216 2674 -4214
rect 2528 -4271 2609 -4266
rect 2528 -4323 2542 -4271
rect 2594 -4323 2609 -4271
rect 2528 -4327 2609 -4323
rect 2550 -4506 2584 -4327
rect 2758 -4446 2792 -4214
rect 2736 -4451 2817 -4446
rect 2736 -4503 2750 -4451
rect 2802 -4503 2817 -4451
rect 2462 -4540 2674 -4506
rect 2736 -4507 2817 -4503
rect 2758 -4508 2792 -4507
rect 2462 -4683 2496 -4540
rect 2550 -4623 2584 -4540
rect 2640 -4713 2674 -4540
rect 1128 -5091 1162 -5002
rect 59 -5125 1162 -5091
rect -51 -5214 22 -5213
rect -51 -5266 -41 -5214
rect 11 -5266 22 -5214
rect 306 -5214 379 -5213
rect 306 -5266 316 -5214
rect 368 -5266 379 -5214
rect -138 -5381 -65 -5380
rect -138 -5433 -128 -5381
rect -76 -5433 -65 -5381
rect -119 -5524 -85 -5433
rect -30 -5603 4 -5266
rect 40 -5381 113 -5380
rect 40 -5433 50 -5381
rect 102 -5433 113 -5381
rect 218 -5381 291 -5380
rect 218 -5433 228 -5381
rect 280 -5433 291 -5381
rect 59 -5524 93 -5433
rect 238 -5524 272 -5433
rect 326 -5586 360 -5266
rect 593 -5315 627 -5125
rect 1216 -5213 1250 -4940
rect 840 -5214 913 -5213
rect 840 -5266 850 -5214
rect 902 -5266 913 -5214
rect 1197 -5214 1270 -5213
rect 1197 -5266 1207 -5214
rect 1259 -5266 1270 -5214
rect 415 -5349 804 -5315
rect 415 -5524 449 -5349
rect 505 -5620 539 -5349
rect 592 -5523 626 -5349
rect 681 -5606 715 -5349
rect 770 -5524 804 -5349
rect 860 -5585 894 -5266
rect 1109 -5381 1182 -5380
rect 930 -5382 1003 -5381
rect 930 -5434 940 -5382
rect 992 -5434 1003 -5382
rect 1109 -5433 1119 -5381
rect 1171 -5433 1182 -5381
rect 949 -5524 983 -5434
rect 1128 -5524 1162 -5433
rect 1216 -5623 1250 -5266
rect 1306 -5380 1340 -4994
rect 1394 -5093 1428 -4913
rect 1375 -5094 1448 -5093
rect 1375 -5146 1385 -5094
rect 1437 -5146 1448 -5094
rect 1286 -5381 1359 -5380
rect 1286 -5433 1296 -5381
rect 1348 -5433 1359 -5381
rect 1306 -5524 1340 -5433
rect 149 -6077 183 -5822
rect -208 -6111 183 -6077
rect 237 -6250 271 -5901
rect 217 -6251 290 -6250
rect 217 -6303 227 -6251
rect 279 -6303 290 -6251
rect 594 -6493 628 -5899
rect 951 -6250 985 -5899
rect 1038 -6081 1072 -5808
rect 1394 -6081 1428 -5146
rect 1572 -5213 1606 -4938
rect 1750 -5093 1784 -4938
rect 1730 -5094 1803 -5093
rect 1730 -5146 1740 -5094
rect 1792 -5146 1803 -5094
rect 1927 -5213 1961 -4940
rect 1553 -5214 1626 -5213
rect 1553 -5266 1563 -5214
rect 1615 -5266 1626 -5214
rect 1907 -5214 1980 -5213
rect 1907 -5266 1917 -5214
rect 1969 -5266 1980 -5214
rect 1482 -5433 1874 -5399
rect 1482 -5523 1516 -5433
rect 1573 -5607 1607 -5433
rect 1661 -5523 1695 -5433
rect 1749 -5604 1783 -5433
rect 1840 -5523 1874 -5433
rect 2018 -5523 2052 -4993
rect 2106 -5093 2140 -4939
rect 2086 -5094 2159 -5093
rect 2086 -5146 2096 -5094
rect 2148 -5146 2159 -5094
rect 2195 -5525 2229 -4995
rect 2284 -5213 2318 -4939
rect 2264 -5214 2337 -5213
rect 2264 -5266 2274 -5214
rect 2326 -5266 2337 -5214
rect 2373 -5525 2407 -4995
rect 2462 -5093 2496 -4937
rect 2443 -5094 2516 -5093
rect 2443 -5146 2453 -5094
rect 2505 -5146 2516 -5094
rect 2463 -5442 2674 -5408
rect 2463 -5585 2497 -5442
rect 2550 -5525 2584 -5442
rect 2640 -5587 2674 -5442
rect 1038 -6115 1428 -6081
rect 932 -6251 1005 -6250
rect 932 -6303 942 -6251
rect 994 -6303 1005 -6251
rect 1662 -6493 1696 -5901
rect 1928 -6124 1962 -5839
rect 2106 -6007 2140 -5842
rect 2086 -6008 2159 -6007
rect 2086 -6060 2096 -6008
rect 2148 -6060 2159 -6008
rect 2284 -6124 2318 -5841
rect 2462 -6007 2496 -5839
rect 2442 -6008 2515 -6007
rect 2442 -6060 2452 -6008
rect 2504 -6060 2515 -6008
rect 1908 -6125 1981 -6124
rect 1908 -6177 1918 -6125
rect 1970 -6177 1981 -6125
rect 2265 -6125 2338 -6124
rect 2265 -6177 2275 -6125
rect 2327 -6177 2338 -6125
rect 2879 -6365 2931 -2606
rect 3194 -4805 3246 -2480
rect 3184 -4857 3194 -4805
rect 3246 -4857 3256 -4805
rect 4761 -4857 4771 -4805
rect 4823 -4857 4833 -4805
rect 2869 -6417 2879 -6365
rect 2931 -6417 2941 -6365
rect -476 -6527 1696 -6493
rect -742 -6598 -708 -6532
rect 4771 -6597 4823 -4857
rect 5027 -5007 5100 -5006
rect 5027 -5059 5037 -5007
rect 5089 -5059 5100 -5007
rect 4895 -5213 4968 -5212
rect 4895 -5265 4905 -5213
rect 4957 -5265 4968 -5213
rect 4762 -6598 4835 -6597
rect -763 -6599 -690 -6598
rect -763 -6651 -753 -6599
rect -701 -6651 -690 -6599
rect 4762 -6650 4772 -6598
rect 4824 -6650 4835 -6598
rect -2013 -6715 -1940 -6714
rect -2013 -6767 -2003 -6715
rect -1951 -6767 -1940 -6715
rect 4771 -6891 4823 -6650
rect 4905 -6889 4958 -5265
rect 5037 -6887 5090 -5059
rect 5337 -5527 5390 -2258
rect 6670 -2263 6754 -2257
rect 7034 -2687 7080 -2509
rect 16034 -2687 16080 -2509
rect 6212 -3457 6296 -3451
rect 6212 -3509 6228 -3457
rect 6280 -3509 6296 -3457
rect 6212 -3515 6296 -3509
rect 7034 -3709 7080 -3537
rect 16034 -3709 16080 -3537
rect 7034 -4487 7080 -4309
rect 16034 -4487 16080 -4309
rect 5604 -5213 5688 -5207
rect 5604 -5265 5620 -5213
rect 5672 -5265 5688 -5213
rect 5604 -5271 5688 -5265
rect 7034 -5509 7080 -5337
rect 16034 -5509 16080 -5337
rect 5327 -5528 5400 -5527
rect 5327 -5580 5337 -5528
rect 5389 -5580 5400 -5528
rect 7034 -6287 7080 -6109
rect 16034 -6287 16080 -6109
rect 17826 -6521 17901 -4862
rect 17821 -6527 17905 -6521
rect 17821 -6579 17837 -6527
rect 17889 -6579 17905 -6527
rect 17821 -6585 17905 -6579
rect 5028 -6888 5101 -6887
rect 4896 -6890 4969 -6889
rect 4760 -6892 4833 -6891
rect 4760 -6944 4770 -6892
rect 4822 -6944 4833 -6892
rect 4896 -6942 4906 -6890
rect 4958 -6942 4969 -6890
rect 5028 -6940 5038 -6888
rect 5090 -6940 5101 -6888
rect 7034 -7309 7080 -7137
rect 16034 -7309 16080 -7137
rect -3883 -7697 -3873 -7691
rect -5629 -7731 -3873 -7697
rect -5628 -7875 -5594 -7731
rect -5544 -7824 -5500 -7731
rect -5450 -7875 -5416 -7731
rect -5366 -7830 -5322 -7731
rect -5188 -7830 -5144 -7731
rect -5094 -7876 -5060 -7731
rect -5010 -7830 -4966 -7731
rect -4832 -7830 -4788 -7731
rect -4738 -7876 -4704 -7731
rect -4654 -7830 -4610 -7731
rect -4476 -7830 -4432 -7731
rect -4382 -7876 -4348 -7731
rect -4298 -7830 -4254 -7731
rect -3883 -7743 -3873 -7731
rect -3821 -7743 -3811 -7691
rect -3741 -7790 -3731 -7785
rect -4026 -7824 -3731 -7790
rect -4026 -7880 -3992 -7824
rect -3741 -7837 -3731 -7824
rect -3679 -7837 -3669 -7785
rect -3551 -7840 -3541 -7788
rect -3489 -7840 -3479 -7788
rect -5628 -11756 -5594 -8130
rect -5544 -8340 -5500 -8214
rect -5544 -8890 -5500 -8764
rect -5544 -9440 -5500 -9314
rect -5544 -9990 -5500 -9864
rect -5544 -10540 -5500 -10414
rect -5544 -11090 -5500 -10964
rect -5544 -11655 -5500 -11485
rect -5450 -11799 -5416 -8130
rect -5366 -8340 -5322 -8214
rect -5366 -8890 -5322 -8764
rect -5366 -9440 -5322 -9314
rect -5366 -9990 -5322 -9864
rect -5366 -10540 -5322 -10414
rect -5366 -11090 -5322 -10964
rect -5272 -11174 -5238 -8130
rect -5188 -8340 -5144 -8214
rect -5188 -8890 -5144 -8764
rect -5188 -9440 -5144 -9314
rect -5188 -9990 -5144 -9864
rect -5188 -10540 -5144 -10414
rect -5188 -11090 -5144 -10964
rect -5364 -11655 -5320 -11485
rect -5272 -12119 -5238 -11431
rect -5188 -11656 -5144 -11486
rect -5094 -11830 -5060 -8131
rect -5010 -8341 -4966 -8215
rect -5010 -8890 -4966 -8764
rect -5010 -9440 -4966 -9314
rect -5010 -9990 -4966 -9864
rect -5010 -10540 -4966 -10414
rect -5010 -11090 -4966 -10964
rect -4916 -11174 -4882 -8130
rect -4832 -8340 -4788 -8214
rect -4832 -8890 -4788 -8764
rect -4832 -9440 -4788 -9314
rect -4832 -9990 -4788 -9864
rect -4832 -10540 -4788 -10414
rect -4832 -11090 -4788 -10964
rect -5010 -11655 -4966 -11485
rect -4916 -12119 -4882 -11430
rect -4832 -11657 -4788 -11487
rect -4738 -11788 -4704 -8130
rect -4654 -8340 -4610 -8214
rect -4654 -8890 -4610 -8764
rect -4654 -9440 -4610 -9314
rect -4654 -9990 -4610 -9864
rect -4654 -10540 -4610 -10414
rect -4654 -11090 -4610 -10964
rect -4560 -11174 -4526 -8130
rect -4476 -8340 -4432 -8214
rect -4476 -8890 -4432 -8764
rect -4476 -9440 -4432 -9314
rect -4476 -9990 -4432 -9864
rect -4476 -10540 -4432 -10414
rect -4476 -11090 -4432 -10964
rect -4654 -11657 -4610 -11487
rect -4560 -12119 -4526 -11430
rect -4476 -11656 -4432 -11486
rect -4382 -11804 -4348 -8130
rect -4298 -8340 -4254 -8214
rect -4298 -8890 -4254 -8764
rect -4298 -9440 -4254 -9314
rect -4298 -9990 -4254 -9864
rect -4298 -10540 -4254 -10414
rect -4298 -11090 -4254 -10964
rect -4204 -11174 -4170 -8130
rect -4120 -8340 -4076 -8214
rect -4120 -8890 -4076 -8764
rect -4120 -9440 -4076 -9314
rect -4120 -9990 -4076 -9864
rect -4120 -10540 -4076 -10414
rect -4120 -11090 -4076 -10964
rect -4026 -11174 -3992 -8130
rect -4298 -11656 -4254 -11486
rect -4204 -12119 -4170 -11430
rect -4120 -11656 -4076 -11486
rect -4113 -12119 -4079 -12030
rect -4026 -12119 -3992 -11430
rect -5272 -12153 -3611 -12119
rect -5512 -12272 -5439 -12271
rect -4512 -12272 -4439 -12271
rect -5512 -12324 -5502 -12272
rect -5450 -12324 -5439 -12272
rect -5010 -12273 -4937 -12272
rect -6976 -12513 -6014 -12512
rect -6976 -12565 -6077 -12513
rect -6025 -12565 -6014 -12513
rect -5636 -12513 -5563 -12512
rect -5636 -12565 -5626 -12513
rect -5574 -12565 -5563 -12513
rect -6233 -13063 -6160 -13062
rect -6233 -13115 -6223 -13063
rect -6171 -13115 -6160 -13063
rect -6976 -13853 -6363 -13852
rect -6976 -13905 -6426 -13853
rect -6374 -13905 -6363 -13853
rect -6223 -14055 -6170 -13115
rect -6077 -13745 -6024 -12565
rect -5922 -12628 -5877 -12612
rect -5922 -12700 -5876 -12628
rect -5817 -12668 -5778 -12612
rect -5617 -12662 -5583 -12565
rect -5824 -12700 -5778 -12668
rect -5492 -12700 -5458 -12324
rect -5010 -12325 -5000 -12273
rect -4948 -12325 -4937 -12273
rect -4512 -12324 -4502 -12272
rect -4450 -12324 -4439 -12272
rect -5386 -12389 -5313 -12388
rect -5386 -12441 -5376 -12389
rect -5324 -12441 -5313 -12389
rect -5137 -12389 -5064 -12388
rect -5137 -12441 -5127 -12389
rect -5075 -12441 -5064 -12389
rect -5367 -12668 -5333 -12441
rect -5117 -12668 -5083 -12441
rect -4992 -12700 -4958 -12325
rect -4887 -12513 -4814 -12512
rect -4887 -12565 -4877 -12513
rect -4825 -12565 -4814 -12513
rect -4637 -12513 -4564 -12512
rect -4637 -12565 -4627 -12513
rect -4575 -12565 -4564 -12513
rect -4867 -12668 -4833 -12565
rect -4617 -12668 -4583 -12565
rect -4492 -12700 -4458 -12324
rect -4387 -12389 -4314 -12388
rect -4387 -12441 -4377 -12389
rect -4325 -12441 -4314 -12389
rect -3938 -12390 -3865 -12389
rect -4367 -12668 -4333 -12441
rect -3938 -12442 -3928 -12390
rect -3876 -12442 -3865 -12390
rect -4172 -12700 -4126 -12612
rect -5824 -12740 -5626 -12700
rect -5574 -12740 -5376 -12700
rect -5324 -12740 -5126 -12700
rect -5074 -12740 -4876 -12700
rect -4823 -12740 -4625 -12700
rect -4574 -12740 -4376 -12700
rect -4324 -12740 -4126 -12700
rect -4074 -12712 -4028 -12612
rect -5818 -12940 -5632 -12900
rect -5574 -12940 -5376 -12900
rect -5324 -12940 -5126 -12900
rect -5074 -12940 -4876 -12900
rect -4825 -12940 -4627 -12900
rect -4574 -12940 -4376 -12900
rect -4324 -12940 -4126 -12900
rect -5744 -13062 -5704 -12940
rect -5761 -13063 -5688 -13062
rect -5761 -13115 -5751 -13063
rect -5699 -13115 -5688 -13063
rect -5495 -13380 -5455 -12940
rect -5245 -13189 -5205 -12940
rect -5261 -13190 -5188 -13189
rect -5261 -13242 -5251 -13190
rect -5199 -13242 -5188 -13190
rect -4995 -13380 -4955 -12940
rect -4746 -13062 -4706 -12940
rect -4762 -13063 -4689 -13062
rect -4762 -13115 -4752 -13063
rect -4700 -13115 -4689 -13063
rect -4495 -13380 -4455 -12940
rect -4244 -13189 -4204 -12940
rect -4261 -13190 -4188 -13189
rect -4261 -13242 -4251 -13190
rect -4199 -13242 -4188 -13190
rect -5824 -13420 -5626 -13380
rect -5574 -13420 -5376 -13380
rect -5324 -13420 -5126 -13380
rect -5074 -13420 -4876 -13380
rect -4824 -13420 -4626 -13380
rect -4574 -13420 -4376 -13380
rect -4324 -13420 -4126 -13380
rect -5922 -13708 -5876 -13608
rect -5824 -13620 -5626 -13580
rect -5574 -13620 -5376 -13580
rect -5324 -13620 -5126 -13580
rect -5074 -13620 -4876 -13580
rect -4824 -13620 -4626 -13580
rect -4574 -13620 -4376 -13580
rect -4324 -13620 -4126 -13580
rect -5824 -13708 -5778 -13620
rect -6087 -13746 -6014 -13745
rect -6087 -13798 -6077 -13746
rect -6025 -13798 -6014 -13746
rect -5720 -13957 -5686 -13620
rect -5617 -13852 -5583 -13652
rect -5367 -13745 -5333 -13652
rect -5386 -13746 -5313 -13745
rect -5386 -13798 -5376 -13746
rect -5324 -13798 -5313 -13746
rect -5636 -13853 -5563 -13852
rect -5636 -13905 -5626 -13853
rect -5574 -13905 -5563 -13853
rect -5740 -13958 -5667 -13957
rect -5740 -14010 -5730 -13958
rect -5678 -14010 -5667 -13958
rect -5240 -14055 -5206 -13620
rect -5117 -13745 -5083 -13652
rect -5136 -13746 -5063 -13745
rect -5136 -13798 -5126 -13746
rect -5074 -13798 -5063 -13746
rect -4867 -13852 -4833 -13652
rect -4887 -13853 -4814 -13852
rect -4887 -13905 -4877 -13853
rect -4825 -13905 -4814 -13853
rect -4742 -13957 -4708 -13620
rect -4617 -13852 -4583 -13652
rect -4367 -13745 -4333 -13652
rect -4386 -13746 -4313 -13745
rect -4386 -13798 -4376 -13746
rect -4324 -13798 -4313 -13746
rect -4637 -13853 -4564 -13852
rect -4637 -13905 -4627 -13853
rect -4575 -13905 -4564 -13853
rect -4762 -13958 -4689 -13957
rect -4762 -14010 -4752 -13958
rect -4700 -14010 -4689 -13958
rect -4240 -14055 -4206 -13620
rect -4172 -13708 -4126 -13620
rect -4074 -13708 -4028 -13608
rect -3928 -13852 -3875 -12442
rect -3798 -13190 -3725 -13189
rect -3798 -13242 -3788 -13190
rect -3736 -13242 -3725 -13190
rect -3938 -13853 -3865 -13852
rect -3938 -13905 -3928 -13853
rect -3876 -13905 -3865 -13853
rect -3928 -13906 -3875 -13905
rect -3788 -13957 -3735 -13242
rect -3798 -13958 -3725 -13957
rect -3798 -14010 -3788 -13958
rect -3736 -14010 -3725 -13958
rect -6233 -14056 -6160 -14055
rect -6233 -14108 -6223 -14056
rect -6171 -14108 -6160 -14056
rect -5260 -14056 -5187 -14055
rect -5260 -14108 -5250 -14056
rect -5198 -14108 -5187 -14056
rect -4260 -14056 -4187 -14055
rect -4260 -14108 -4250 -14056
rect -4198 -14108 -4187 -14056
rect -6965 -14260 -4303 -14226
rect -6028 -14394 -5994 -14260
rect -5939 -14350 -5905 -14260
rect -5850 -14394 -5816 -14260
rect -5761 -14350 -5727 -14260
rect -5583 -14350 -5549 -14260
rect -5405 -14350 -5371 -14260
rect -5227 -14350 -5193 -14260
rect -5049 -14350 -5015 -14260
rect -4871 -14350 -4837 -14260
rect -4693 -14350 -4659 -14260
rect -4515 -14350 -4481 -14260
rect -4337 -14350 -4303 -14260
rect -4248 -14260 -4036 -14226
rect -4248 -14394 -4214 -14260
rect -4159 -14344 -4125 -14260
rect -4070 -14394 -4036 -14260
rect -5850 -14795 -5816 -14651
rect -6169 -14796 -6096 -14795
rect -6169 -14848 -6159 -14796
rect -6107 -14848 -6096 -14796
rect -5870 -14796 -5797 -14795
rect -5870 -14848 -5860 -14796
rect -5808 -14848 -5797 -14796
rect -6159 -15482 -6106 -14848
rect -6028 -14959 -5816 -14925
rect -6027 -15093 -5993 -14959
rect -5939 -15050 -5905 -14959
rect -5850 -15094 -5816 -14959
rect -5761 -15010 -5727 -14700
rect -5672 -15094 -5638 -14650
rect -5583 -15035 -5549 -14719
rect -5494 -14901 -5460 -14650
rect -5514 -14902 -5441 -14901
rect -5514 -14954 -5504 -14902
rect -5452 -14954 -5441 -14902
rect -5405 -15033 -5371 -14717
rect -6169 -15483 -6096 -15482
rect -6169 -15535 -6159 -15483
rect -6107 -15535 -6096 -15483
rect -6159 -16193 -6106 -15535
rect -5850 -15588 -5816 -15350
rect -5870 -15589 -5797 -15588
rect -5870 -15641 -5860 -15589
rect -5808 -15641 -5797 -15589
rect -5761 -15717 -5727 -15401
rect -5672 -15803 -5638 -15350
rect -5583 -15724 -5549 -15408
rect -5494 -15481 -5460 -15350
rect -5514 -15482 -5441 -15481
rect -5514 -15534 -5504 -15482
rect -5452 -15534 -5441 -15482
rect -5405 -15731 -5371 -15415
rect -6028 -16185 -5994 -16049
rect -5939 -16185 -5905 -16094
rect -5850 -16185 -5816 -16050
rect -6169 -16194 -6096 -16193
rect -6169 -16246 -6159 -16194
rect -6107 -16246 -6096 -16194
rect -6028 -16219 -5816 -16185
rect -6159 -17007 -6106 -16246
rect -5850 -16294 -5816 -16219
rect -5870 -16295 -5797 -16294
rect -5870 -16347 -5860 -16295
rect -5808 -16347 -5797 -16295
rect -5761 -16426 -5727 -16110
rect -5672 -16494 -5638 -16050
rect -5583 -16428 -5549 -16112
rect -5494 -16193 -5460 -16050
rect -5514 -16194 -5441 -16193
rect -5514 -16246 -5504 -16194
rect -5452 -16246 -5441 -16194
rect -5405 -16427 -5371 -16111
rect -5316 -16494 -5282 -14650
rect -5227 -15032 -5193 -14716
rect -5138 -14795 -5104 -14651
rect -5157 -14796 -5084 -14795
rect -5157 -14848 -5147 -14796
rect -5095 -14848 -5084 -14796
rect -5049 -15032 -5015 -14716
rect -5227 -15729 -5193 -15413
rect -5138 -15589 -5104 -15350
rect -5158 -15590 -5085 -15589
rect -5158 -15642 -5148 -15590
rect -5096 -15642 -5085 -15590
rect -5049 -15730 -5015 -15414
rect -5227 -16427 -5193 -16111
rect -5138 -16294 -5104 -16051
rect -5158 -16295 -5085 -16294
rect -5158 -16347 -5148 -16295
rect -5096 -16347 -5085 -16295
rect -5049 -16427 -5015 -16111
rect -4960 -16494 -4926 -14650
rect -4871 -15031 -4837 -14715
rect -4782 -14901 -4748 -14650
rect -4801 -14902 -4728 -14901
rect -4801 -14954 -4791 -14902
rect -4739 -14954 -4728 -14902
rect -4693 -15030 -4659 -14714
rect -4871 -15730 -4837 -15414
rect -4782 -15481 -4748 -15350
rect -4802 -15482 -4729 -15481
rect -4802 -15534 -4792 -15482
rect -4740 -15534 -4729 -15482
rect -4693 -15729 -4659 -15413
rect -4871 -16427 -4837 -16111
rect -4782 -16193 -4748 -16050
rect -4802 -16194 -4729 -16193
rect -4802 -16246 -4792 -16194
rect -4740 -16246 -4729 -16194
rect -4693 -16427 -4659 -16111
rect -4604 -16494 -4570 -14650
rect -4515 -15030 -4481 -14714
rect -4426 -14795 -4392 -14650
rect -4446 -14796 -4373 -14795
rect -4446 -14848 -4436 -14796
rect -4384 -14848 -4373 -14796
rect -4337 -15028 -4303 -14712
rect -4248 -14925 -4214 -14650
rect -4159 -14750 -4125 -14700
rect -3664 -14901 -3611 -12153
rect -3541 -13137 -3489 -7840
rect 5027 -7851 5100 -7850
rect 4896 -7853 4969 -7852
rect 4761 -7855 4834 -7854
rect 4761 -7907 4771 -7855
rect 4823 -7907 4834 -7855
rect 4896 -7905 4906 -7853
rect 4958 -7905 4969 -7853
rect 5027 -7903 5037 -7851
rect 5089 -7903 5100 -7851
rect 5327 -7851 5400 -7850
rect 5174 -7856 5247 -7855
rect -1392 -7923 -1319 -7922
rect -1035 -7923 -962 -7922
rect -3392 -7934 -3319 -7933
rect -3392 -7986 -3382 -7934
rect -3330 -7986 -3319 -7934
rect -1392 -7975 -1382 -7923
rect -1330 -7975 -1319 -7923
rect -1213 -7924 -1140 -7923
rect -3542 -13189 -3489 -13137
rect -3552 -13190 -3479 -13189
rect -3552 -13242 -3542 -13190
rect -3490 -13242 -3479 -13190
rect -3382 -14055 -3329 -7986
rect -1372 -8080 -1338 -7975
rect -1213 -7976 -1203 -7924
rect -1151 -7976 -1140 -7924
rect -1035 -7975 -1025 -7923
rect -973 -7975 -962 -7923
rect -858 -7923 -785 -7922
rect -858 -7975 -848 -7923
rect -796 -7975 -785 -7923
rect -680 -7923 -607 -7922
rect -680 -7975 -670 -7923
rect -618 -7975 -607 -7923
rect -500 -7923 -427 -7922
rect -500 -7975 -490 -7923
rect -438 -7975 -427 -7923
rect 745 -7923 818 -7922
rect 745 -7975 755 -7923
rect 807 -7975 818 -7923
rect 922 -7923 995 -7922
rect 922 -7975 932 -7923
rect 984 -7975 995 -7923
rect 1102 -7923 1175 -7922
rect 1457 -7923 1530 -7922
rect 1102 -7975 1112 -7923
rect 1164 -7975 1175 -7923
rect 1279 -7924 1352 -7923
rect -1194 -8081 -1160 -7976
rect -1016 -8081 -982 -7975
rect -838 -8081 -804 -7975
rect -660 -8081 -626 -7975
rect -481 -8081 -447 -7975
rect 765 -8082 799 -7975
rect 942 -8081 976 -7975
rect 1121 -8081 1155 -7975
rect 1279 -7976 1289 -7924
rect 1341 -7976 1352 -7924
rect 1457 -7975 1467 -7923
rect 1519 -7975 1530 -7923
rect 1634 -7923 1707 -7922
rect 1634 -7975 1644 -7923
rect 1696 -7975 1707 -7923
rect 2880 -7923 2953 -7922
rect 2880 -7975 2890 -7923
rect 2942 -7975 2953 -7923
rect 3059 -7923 3132 -7922
rect 3059 -7975 3069 -7923
rect 3121 -7975 3132 -7923
rect 3237 -7923 3310 -7922
rect 3237 -7975 3247 -7923
rect 3299 -7975 3310 -7923
rect 3414 -7923 3487 -7922
rect 3768 -7923 3841 -7922
rect 3414 -7975 3424 -7923
rect 3476 -7975 3487 -7923
rect 3593 -7924 3666 -7923
rect 1298 -8082 1332 -7976
rect 1476 -8081 1510 -7975
rect 1654 -8081 1688 -7975
rect 2900 -8081 2934 -7975
rect 3078 -8082 3112 -7975
rect 3256 -8081 3290 -7975
rect 3434 -8081 3468 -7975
rect 3593 -7976 3603 -7924
rect 3655 -7976 3666 -7924
rect 3768 -7975 3778 -7923
rect 3830 -7975 3841 -7923
rect 4198 -7924 4271 -7923
rect 3612 -8081 3646 -7976
rect 3790 -8081 3824 -7975
rect 4198 -7976 4208 -7924
rect 4260 -7976 4271 -7924
rect -2171 -8440 -2137 -8358
rect -1995 -8440 -1961 -8389
rect -2171 -8474 -1961 -8440
rect -1995 -8767 -1961 -8474
rect -1906 -8534 -1872 -8438
rect -1926 -8535 -1853 -8534
rect -1926 -8587 -1916 -8535
rect -1864 -8587 -1853 -8535
rect -1817 -8653 -1783 -8389
rect -1729 -8534 -1695 -8438
rect -1749 -8535 -1676 -8534
rect -1749 -8587 -1739 -8535
rect -1687 -8587 -1676 -8535
rect -1836 -8654 -1763 -8653
rect -1836 -8706 -1826 -8654
rect -1774 -8706 -1763 -8654
rect -2457 -8768 -2384 -8767
rect -2457 -8820 -2447 -8768
rect -2395 -8820 -2384 -8768
rect -2015 -8768 -1942 -8767
rect -2015 -8820 -2005 -8768
rect -1953 -8820 -1942 -8768
rect -2447 -12272 -2394 -8820
rect -2174 -9439 -2140 -9360
rect -1995 -9439 -1961 -8820
rect -2174 -9473 -1961 -9439
rect -2325 -9926 -2252 -9925
rect -2325 -9978 -2315 -9926
rect -2263 -9978 -2252 -9926
rect -2457 -12273 -2384 -12272
rect -2457 -12325 -2447 -12273
rect -2395 -12325 -2384 -12273
rect -3392 -14056 -3319 -14055
rect -3392 -14108 -3382 -14056
rect -3330 -14108 -3319 -14056
rect -3946 -14902 -3611 -14901
rect -4248 -14959 -4036 -14925
rect -3946 -14954 -3936 -14902
rect -3884 -14954 -3611 -14902
rect -4515 -15727 -4481 -15411
rect -4426 -15589 -4392 -15351
rect -4445 -15641 -4435 -15589
rect -4383 -15641 -4373 -15589
rect -4337 -15727 -4303 -15411
rect -4515 -16427 -4481 -16111
rect -4426 -16294 -4392 -16050
rect -4446 -16295 -4373 -16294
rect -4446 -16347 -4436 -16295
rect -4384 -16347 -4373 -16295
rect -4337 -16427 -4303 -16111
rect -4248 -16185 -4214 -14959
rect -4159 -15050 -4125 -14959
rect -4070 -15094 -4036 -14959
rect -3936 -15006 -3883 -14954
rect -3935 -15589 -3883 -15006
rect -3945 -15641 -3935 -15589
rect -3883 -15641 -3873 -15589
rect -4159 -16185 -4125 -16094
rect -4070 -16185 -4036 -16050
rect -4248 -16219 -4036 -16185
rect -4248 -16494 -4214 -16219
rect -3935 -16295 -3883 -15641
rect -2447 -15821 -2394 -12325
rect -2315 -14543 -2262 -9978
rect -1995 -10049 -1961 -9473
rect -1906 -9546 -1872 -9441
rect -1926 -9547 -1853 -9546
rect -1926 -9599 -1916 -9547
rect -1864 -9599 -1853 -9547
rect -1926 -9926 -1853 -9925
rect -1926 -9978 -1916 -9926
rect -1864 -9978 -1853 -9926
rect -2175 -10083 -1961 -10049
rect -1906 -10082 -1872 -9978
rect -2175 -10174 -2141 -10083
rect -1995 -10263 -1961 -10083
rect -1817 -10195 -1783 -8706
rect -1639 -8767 -1605 -8378
rect -1549 -8534 -1515 -8439
rect -1568 -8535 -1495 -8534
rect -1568 -8587 -1558 -8535
rect -1506 -8587 -1495 -8535
rect -1461 -8653 -1427 -8380
rect -1392 -8535 -1319 -8534
rect -1392 -8587 -1382 -8535
rect -1330 -8587 -1319 -8535
rect -1480 -8654 -1407 -8653
rect -1480 -8706 -1470 -8654
rect -1418 -8706 -1407 -8654
rect -1658 -8768 -1585 -8767
rect -1658 -8820 -1648 -8768
rect -1596 -8820 -1585 -8768
rect -1728 -9546 -1694 -9439
rect -1748 -9547 -1675 -9546
rect -1748 -9599 -1738 -9547
rect -1686 -9599 -1675 -9547
rect -1748 -9927 -1675 -9926
rect -1748 -9979 -1738 -9927
rect -1686 -9979 -1675 -9927
rect -1728 -10081 -1694 -9979
rect -1639 -10253 -1605 -8820
rect -1549 -9546 -1515 -9438
rect -1568 -9547 -1495 -9546
rect -1568 -9599 -1558 -9547
rect -1506 -9599 -1495 -9547
rect -1570 -9926 -1497 -9925
rect -1570 -9978 -1560 -9926
rect -1508 -9978 -1497 -9926
rect -1550 -10081 -1516 -9978
rect -1461 -10200 -1427 -8706
rect -1372 -9081 -1338 -8587
rect -1283 -8767 -1249 -8381
rect -1213 -8535 -1140 -8534
rect -1213 -8587 -1203 -8535
rect -1151 -8587 -1140 -8535
rect -1303 -8768 -1230 -8767
rect -1303 -8820 -1293 -8768
rect -1241 -8820 -1230 -8768
rect -1372 -9924 -1338 -9439
rect -1392 -9925 -1319 -9924
rect -1392 -9977 -1382 -9925
rect -1330 -9977 -1319 -9925
rect -1283 -10256 -1249 -8820
rect -1193 -9081 -1159 -8587
rect -1105 -8653 -1071 -8370
rect -1036 -8535 -963 -8534
rect -1036 -8587 -1026 -8535
rect -974 -8587 -963 -8535
rect -1125 -8654 -1052 -8653
rect -1125 -8706 -1115 -8654
rect -1063 -8706 -1052 -8654
rect -1105 -10208 -1071 -8706
rect -1016 -9081 -982 -8587
rect -927 -8767 -893 -8382
rect -858 -8535 -785 -8534
rect -858 -8587 -848 -8535
rect -796 -8587 -785 -8535
rect -946 -8768 -873 -8767
rect -946 -8820 -936 -8768
rect -884 -8820 -873 -8768
rect -927 -10257 -893 -8820
rect -838 -9080 -804 -8587
rect -749 -8653 -715 -8368
rect -680 -8535 -607 -8534
rect -680 -8587 -670 -8535
rect -618 -8587 -607 -8535
rect -768 -8654 -695 -8653
rect -768 -8706 -758 -8654
rect -706 -8706 -695 -8654
rect -749 -10180 -715 -8706
rect -660 -9082 -626 -8587
rect -571 -8766 -537 -8373
rect -501 -8535 -428 -8534
rect -501 -8587 -491 -8535
rect -439 -8587 -428 -8535
rect -590 -8767 -517 -8766
rect -590 -8819 -580 -8767
rect -528 -8819 -517 -8767
rect -571 -10248 -537 -8819
rect -482 -9081 -448 -8587
rect -393 -8653 -359 -8358
rect -304 -8534 -270 -8439
rect -324 -8535 -251 -8534
rect -324 -8587 -314 -8535
rect -262 -8587 -251 -8535
rect -412 -8654 -339 -8653
rect -412 -8706 -402 -8654
rect -350 -8706 -339 -8654
rect -393 -10180 -359 -8706
rect -215 -8767 -181 -8371
rect -126 -8534 -92 -8439
rect -146 -8535 -73 -8534
rect -146 -8587 -136 -8535
rect -84 -8587 -73 -8535
rect -37 -8653 -3 -8353
rect 52 -8534 86 -8438
rect 32 -8535 105 -8534
rect 32 -8587 42 -8535
rect 94 -8587 105 -8535
rect -57 -8654 16 -8653
rect -57 -8706 -47 -8654
rect 5 -8706 16 -8654
rect -235 -8768 -162 -8767
rect -235 -8820 -225 -8768
rect -173 -8820 -162 -8768
rect -303 -9546 -269 -9440
rect -322 -9547 -249 -9546
rect -322 -9599 -312 -9547
rect -260 -9599 -249 -9547
rect -324 -9926 -251 -9925
rect -324 -9978 -314 -9926
rect -262 -9978 -251 -9926
rect -304 -10082 -270 -9978
rect -215 -10246 -181 -8820
rect -126 -9545 -92 -9438
rect -146 -9546 -73 -9545
rect -146 -9598 -136 -9546
rect -84 -9598 -73 -9546
rect -146 -9927 -73 -9926
rect -146 -9979 -136 -9927
rect -84 -9979 -73 -9927
rect -126 -10081 -92 -9979
rect -37 -10184 -3 -8706
rect 141 -8768 175 -8380
rect 230 -8534 264 -8440
rect 211 -8535 284 -8534
rect 211 -8587 221 -8535
rect 273 -8587 284 -8535
rect 319 -8653 353 -8362
rect 408 -8534 442 -8440
rect 388 -8535 461 -8534
rect 388 -8587 398 -8535
rect 450 -8587 461 -8535
rect 300 -8654 373 -8653
rect 300 -8706 310 -8654
rect 362 -8706 373 -8654
rect 122 -8769 195 -8768
rect 122 -8821 132 -8769
rect 184 -8821 195 -8769
rect 52 -9546 86 -9440
rect 32 -9547 105 -9546
rect 32 -9599 42 -9547
rect 94 -9599 105 -9547
rect 33 -9926 106 -9925
rect 33 -9978 43 -9926
rect 95 -9978 106 -9926
rect 52 -10082 86 -9978
rect 141 -10255 175 -8821
rect 231 -9545 265 -9439
rect 212 -9546 285 -9545
rect 212 -9598 222 -9546
rect 274 -9598 285 -9546
rect 210 -9926 283 -9925
rect 210 -9978 220 -9926
rect 272 -9978 283 -9926
rect 230 -10081 264 -9978
rect 319 -10194 353 -8706
rect 497 -8766 531 -8370
rect 586 -8534 620 -8439
rect 567 -8535 640 -8534
rect 567 -8587 577 -8535
rect 629 -8587 640 -8535
rect 675 -8653 709 -8365
rect 744 -8535 817 -8534
rect 744 -8587 754 -8535
rect 806 -8587 817 -8535
rect 656 -8654 729 -8653
rect 656 -8706 666 -8654
rect 718 -8706 729 -8654
rect 479 -8767 552 -8766
rect 479 -8819 489 -8767
rect 541 -8819 552 -8767
rect 408 -9546 442 -9438
rect 389 -9547 462 -9546
rect 389 -9599 399 -9547
rect 451 -9599 462 -9547
rect 388 -9926 461 -9925
rect 388 -9978 398 -9926
rect 450 -9978 461 -9926
rect 408 -10082 442 -9978
rect 497 -10245 531 -8819
rect 587 -9546 621 -9440
rect 567 -9547 640 -9546
rect 567 -9599 577 -9547
rect 629 -9599 640 -9547
rect 566 -9926 639 -9925
rect 566 -9978 576 -9926
rect 628 -9978 639 -9926
rect 586 -10082 620 -9978
rect 675 -10189 709 -8706
rect 764 -9082 798 -8587
rect 853 -8766 887 -8369
rect 922 -8535 995 -8534
rect 922 -8587 932 -8535
rect 984 -8587 995 -8535
rect 833 -8767 906 -8766
rect 833 -8819 843 -8767
rect 895 -8819 906 -8767
rect 853 -9191 887 -8819
rect 942 -9081 976 -8587
rect 1031 -8653 1065 -8366
rect 1101 -8535 1174 -8534
rect 1101 -8587 1111 -8535
rect 1163 -8587 1174 -8535
rect 1012 -8654 1085 -8653
rect 1012 -8706 1022 -8654
rect 1074 -8706 1085 -8654
rect 1031 -10213 1065 -8706
rect 1120 -9081 1154 -8587
rect 1209 -8767 1243 -8364
rect 1279 -8535 1352 -8534
rect 1279 -8587 1289 -8535
rect 1341 -8587 1352 -8535
rect 1191 -8768 1264 -8767
rect 1191 -8820 1201 -8768
rect 1253 -8820 1264 -8768
rect 1209 -10239 1243 -8820
rect 1298 -9081 1332 -8587
rect 1387 -8653 1421 -8365
rect 1456 -8535 1529 -8534
rect 1456 -8587 1466 -8535
rect 1518 -8587 1529 -8535
rect 1367 -8654 1440 -8653
rect 1367 -8706 1377 -8654
rect 1429 -8706 1440 -8654
rect 1387 -10213 1421 -8706
rect 1476 -9081 1510 -8587
rect 1565 -8767 1599 -8372
rect 1634 -8535 1707 -8534
rect 1634 -8587 1644 -8535
rect 1696 -8587 1707 -8535
rect 1546 -8768 1619 -8767
rect 1546 -8820 1556 -8768
rect 1608 -8820 1619 -8768
rect 1565 -10247 1599 -8820
rect 1654 -9081 1688 -8587
rect 1743 -8653 1777 -8363
rect 1832 -8534 1866 -8439
rect 1812 -8535 1885 -8534
rect 1812 -8587 1822 -8535
rect 1874 -8587 1885 -8535
rect 1723 -8654 1796 -8653
rect 1723 -8706 1733 -8654
rect 1785 -8706 1796 -8654
rect 1743 -10181 1777 -8706
rect 1921 -8767 1955 -8372
rect 2010 -8534 2044 -8439
rect 1990 -8535 2063 -8534
rect 1990 -8587 2000 -8535
rect 2052 -8587 2063 -8535
rect 2099 -8653 2133 -8368
rect 2188 -8534 2222 -8439
rect 2168 -8535 2241 -8534
rect 2168 -8587 2178 -8535
rect 2230 -8587 2241 -8535
rect 2080 -8654 2153 -8653
rect 2080 -8706 2090 -8654
rect 2142 -8706 2153 -8654
rect 1901 -8768 1974 -8767
rect 1901 -8820 1911 -8768
rect 1963 -8820 1974 -8768
rect 1832 -10082 1866 -9426
rect 1921 -10247 1955 -8820
rect 2010 -10082 2044 -9426
rect 2099 -10209 2133 -8706
rect 2277 -8767 2311 -8372
rect 2367 -8534 2401 -8439
rect 2347 -8535 2420 -8534
rect 2347 -8587 2357 -8535
rect 2409 -8587 2420 -8535
rect 2455 -8653 2489 -8370
rect 2544 -8534 2578 -8439
rect 2524 -8535 2597 -8534
rect 2524 -8587 2534 -8535
rect 2586 -8587 2597 -8535
rect 2436 -8654 2509 -8653
rect 2436 -8706 2446 -8654
rect 2498 -8706 2509 -8654
rect 2257 -8768 2330 -8767
rect 2257 -8820 2267 -8768
rect 2319 -8820 2330 -8768
rect 2188 -9547 2222 -9426
rect 2168 -9548 2241 -9547
rect 2168 -9600 2178 -9548
rect 2230 -9600 2241 -9548
rect 2188 -10082 2222 -9600
rect 2277 -10247 2311 -8820
rect 2366 -9546 2400 -9440
rect 2347 -9547 2420 -9546
rect 2347 -9599 2357 -9547
rect 2409 -9599 2420 -9547
rect 2346 -9926 2419 -9925
rect 2346 -9978 2356 -9926
rect 2408 -9978 2419 -9926
rect 2366 -10082 2400 -9978
rect 2455 -10186 2489 -8706
rect 2633 -8767 2667 -8375
rect 2722 -8534 2756 -8440
rect 2702 -8535 2775 -8534
rect 2702 -8587 2712 -8535
rect 2764 -8587 2775 -8535
rect 2811 -8653 2845 -8374
rect 2880 -8535 2953 -8534
rect 2880 -8587 2890 -8535
rect 2942 -8587 2953 -8535
rect 2792 -8654 2865 -8653
rect 2792 -8706 2802 -8654
rect 2854 -8706 2865 -8654
rect 2614 -8768 2687 -8767
rect 2614 -8820 2624 -8768
rect 2676 -8820 2687 -8768
rect 2544 -9546 2578 -9441
rect 2524 -9547 2597 -9546
rect 2524 -9599 2534 -9547
rect 2586 -9599 2597 -9547
rect 2524 -9926 2597 -9925
rect 2524 -9978 2534 -9926
rect 2586 -9978 2597 -9926
rect 2544 -10081 2578 -9978
rect 2633 -10250 2667 -8820
rect 2722 -9546 2756 -9441
rect 2703 -9547 2776 -9546
rect 2703 -9599 2713 -9547
rect 2765 -9599 2776 -9547
rect 2702 -9927 2775 -9926
rect 2702 -9979 2712 -9927
rect 2764 -9979 2775 -9927
rect 2722 -10081 2756 -9979
rect 2811 -10205 2845 -8706
rect 2900 -9082 2934 -8587
rect 2989 -8767 3023 -8376
rect 3058 -8535 3131 -8534
rect 3058 -8587 3068 -8535
rect 3120 -8587 3131 -8535
rect 2970 -8768 3043 -8767
rect 2970 -8820 2980 -8768
rect 3032 -8820 3043 -8768
rect 2881 -9926 2954 -9925
rect 2881 -9978 2891 -9926
rect 2943 -9978 2954 -9926
rect 2900 -10080 2934 -9978
rect 2989 -10251 3023 -8820
rect 3078 -9082 3112 -8587
rect 3167 -8653 3201 -8362
rect 3236 -8535 3309 -8534
rect 3236 -8587 3246 -8535
rect 3298 -8587 3309 -8535
rect 3148 -8654 3221 -8653
rect 3148 -8706 3158 -8654
rect 3210 -8706 3221 -8654
rect 3059 -9926 3132 -9925
rect 3059 -9978 3069 -9926
rect 3121 -9978 3132 -9926
rect 3078 -10080 3112 -9978
rect 3167 -10176 3201 -8706
rect 3256 -9081 3290 -8587
rect 3345 -8767 3379 -8374
rect 3414 -8535 3487 -8534
rect 3414 -8587 3424 -8535
rect 3476 -8587 3487 -8535
rect 3326 -8768 3399 -8767
rect 3326 -8820 3336 -8768
rect 3388 -8820 3399 -8768
rect 3256 -9925 3290 -9443
rect 3236 -9926 3309 -9925
rect 3236 -9978 3246 -9926
rect 3298 -9978 3309 -9926
rect 3256 -10081 3290 -9978
rect 3345 -10249 3379 -8820
rect 3434 -9082 3468 -8587
rect 3523 -8653 3557 -8365
rect 3592 -8535 3665 -8534
rect 3592 -8587 3602 -8535
rect 3654 -8587 3665 -8535
rect 3503 -8654 3576 -8653
rect 3503 -8706 3513 -8654
rect 3565 -8706 3576 -8654
rect 3523 -10190 3557 -8706
rect 3612 -9082 3646 -8587
rect 3701 -8767 3735 -8376
rect 3879 -8440 3913 -8365
rect 4056 -8440 4090 -8360
rect 3879 -8474 4090 -8440
rect 3771 -8535 3844 -8534
rect 3771 -8587 3781 -8535
rect 3833 -8587 3844 -8535
rect 3682 -8768 3755 -8767
rect 3682 -8820 3692 -8768
rect 3744 -8820 3755 -8768
rect 3701 -10251 3735 -8820
rect 3790 -9081 3824 -8587
rect 3879 -8653 3913 -8474
rect 3859 -8654 3932 -8653
rect 3859 -8706 3869 -8654
rect 3921 -8706 3932 -8654
rect 3879 -9439 3913 -8706
rect 4056 -9439 4090 -9361
rect 3879 -9473 4090 -9439
rect 3879 -10047 3913 -9473
rect 4208 -9546 4261 -7976
rect 4771 -9262 4823 -7907
rect 4771 -9314 4824 -9262
rect 4761 -9315 4834 -9314
rect 4761 -9367 4771 -9315
rect 4823 -9367 4834 -9315
rect 4198 -9547 4271 -9546
rect 4198 -9599 4208 -9547
rect 4260 -9599 4271 -9547
rect 3879 -10081 4092 -10047
rect 3879 -10205 3913 -10081
rect 4058 -10174 4092 -10081
rect -1837 -10909 -1764 -10908
rect -1837 -10961 -1827 -10909
rect -1775 -10961 -1764 -10909
rect -1480 -10909 -1407 -10908
rect -1480 -10961 -1470 -10909
rect -1418 -10961 -1407 -10909
rect -2172 -11439 -2138 -11345
rect -1995 -11439 -1961 -11189
rect -2172 -11473 -1961 -11439
rect -1995 -11637 -1961 -11473
rect -2014 -11638 -1941 -11637
rect -2014 -11690 -2004 -11638
rect -1952 -11690 -1941 -11638
rect -1995 -12047 -1961 -11690
rect -1905 -11919 -1871 -11445
rect -1925 -11920 -1852 -11919
rect -1925 -11972 -1915 -11920
rect -1863 -11972 -1852 -11920
rect -2176 -12081 -1961 -12047
rect -2176 -12171 -2142 -12081
rect -1995 -12542 -1961 -12081
rect -1905 -12083 -1871 -11972
rect -2015 -12543 -1942 -12542
rect -2015 -12595 -2005 -12543
rect -1953 -12595 -1942 -12543
rect -1995 -13046 -1961 -12595
rect -2174 -13080 -1961 -13046
rect -1906 -13077 -1872 -12439
rect -2174 -13165 -2140 -13080
rect -1995 -13200 -1961 -13080
rect -1818 -13220 -1784 -10961
rect -1728 -11919 -1694 -11447
rect -1639 -11528 -1605 -11374
rect -1659 -11529 -1586 -11528
rect -1659 -11581 -1649 -11529
rect -1597 -11581 -1586 -11529
rect -1549 -11919 -1515 -11447
rect -1748 -11920 -1675 -11919
rect -1748 -11972 -1738 -11920
rect -1686 -11972 -1675 -11920
rect -1569 -11920 -1496 -11919
rect -1569 -11972 -1559 -11920
rect -1507 -11972 -1496 -11920
rect -1728 -12081 -1694 -11972
rect -1549 -12081 -1515 -11972
rect -1728 -13080 -1694 -12442
rect -1639 -12542 -1605 -12386
rect -1659 -12543 -1586 -12542
rect -1659 -12595 -1649 -12543
rect -1597 -12595 -1586 -12543
rect -1549 -13079 -1515 -12441
rect -1461 -13228 -1427 -10961
rect -1372 -11081 -1338 -10438
rect -1193 -11081 -1159 -10432
rect -1124 -10909 -1051 -10908
rect -1124 -10961 -1114 -10909
rect -1062 -10961 -1051 -10909
rect -1372 -11919 -1338 -11448
rect -1283 -11526 -1249 -11373
rect -1284 -11528 -1249 -11526
rect -1303 -11529 -1230 -11528
rect -1303 -11581 -1293 -11529
rect -1241 -11581 -1230 -11529
rect -1391 -11920 -1318 -11919
rect -1391 -11972 -1381 -11920
rect -1329 -11972 -1318 -11920
rect -1372 -12080 -1338 -11972
rect -1372 -13080 -1338 -12442
rect -1284 -12654 -1250 -11581
rect -1194 -11919 -1160 -11448
rect -1213 -11920 -1140 -11919
rect -1213 -11972 -1203 -11920
rect -1151 -11972 -1140 -11920
rect -1194 -12081 -1160 -11972
rect -1304 -12655 -1231 -12654
rect -1304 -12707 -1294 -12655
rect -1242 -12707 -1231 -12655
rect -1194 -13079 -1160 -12441
rect -1105 -13202 -1071 -10961
rect -1016 -11081 -982 -10432
rect -838 -11082 -804 -10433
rect -768 -10909 -695 -10908
rect -768 -10961 -758 -10909
rect -706 -10961 -695 -10909
rect -1016 -11919 -982 -11448
rect -927 -11528 -893 -11367
rect -947 -11529 -874 -11528
rect -947 -11581 -937 -11529
rect -885 -11581 -874 -11529
rect -838 -11919 -804 -11448
rect -1035 -11920 -962 -11919
rect -1035 -11972 -1025 -11920
rect -973 -11972 -962 -11920
rect -858 -11920 -785 -11919
rect -858 -11972 -848 -11920
rect -796 -11972 -785 -11920
rect -1016 -12080 -982 -11972
rect -838 -12081 -804 -11972
rect -1016 -13080 -982 -12442
rect -927 -12783 -893 -12389
rect -947 -12784 -874 -12783
rect -947 -12836 -937 -12784
rect -885 -12836 -874 -12784
rect -927 -13174 -893 -12836
rect -838 -13079 -804 -12441
rect -749 -13222 -715 -10961
rect -659 -11081 -625 -10432
rect -482 -11081 -448 -10432
rect 853 -10438 887 -10368
rect 941 -10438 975 -10431
rect 1031 -10438 1065 -10360
rect 759 -10472 1159 -10438
rect 941 -10908 975 -10472
rect -412 -10909 -339 -10908
rect -412 -10961 -402 -10909
rect -350 -10961 -339 -10909
rect -56 -10909 17 -10908
rect -56 -10961 -46 -10909
rect 6 -10961 17 -10909
rect 299 -10909 372 -10908
rect 299 -10961 309 -10909
rect 361 -10961 372 -10909
rect 655 -10909 728 -10908
rect 655 -10961 665 -10909
rect 717 -10961 728 -10909
rect 921 -10909 994 -10908
rect 921 -10961 931 -10909
rect 983 -10961 994 -10909
rect 1189 -10909 1262 -10908
rect 1189 -10961 1199 -10909
rect 1251 -10961 1262 -10909
rect -660 -11919 -626 -11448
rect -571 -11637 -537 -11388
rect -590 -11638 -517 -11637
rect -590 -11690 -580 -11638
rect -528 -11690 -517 -11638
rect -482 -11919 -448 -11448
rect -680 -11920 -607 -11919
rect -680 -11972 -670 -11920
rect -618 -11972 -607 -11920
rect -502 -11920 -429 -11919
rect -502 -11972 -492 -11920
rect -440 -11972 -429 -11920
rect -660 -12081 -626 -11972
rect -482 -12081 -448 -11972
rect -660 -13081 -626 -12443
rect -571 -12653 -537 -12387
rect -592 -12654 -519 -12653
rect -592 -12706 -582 -12654
rect -530 -12706 -519 -12654
rect -482 -13081 -448 -12443
rect -393 -13207 -359 -10961
rect -304 -11919 -270 -11448
rect -215 -11757 -181 -11385
rect -234 -11758 -161 -11757
rect -234 -11810 -224 -11758
rect -172 -11810 -161 -11758
rect -324 -11920 -251 -11919
rect -324 -11972 -314 -11920
rect -262 -11972 -251 -11920
rect -304 -12080 -270 -11972
rect -304 -13082 -270 -12444
rect -215 -12783 -181 -11810
rect -126 -11919 -92 -11448
rect -146 -11920 -73 -11919
rect -146 -11972 -136 -11920
rect -84 -11972 -73 -11920
rect -126 -12079 -92 -11972
rect -234 -12784 -161 -12783
rect -234 -12836 -224 -12784
rect -172 -12836 -161 -12784
rect -126 -13081 -92 -12443
rect -36 -13199 -2 -10961
rect 52 -11919 86 -11448
rect 141 -11757 175 -11387
rect 121 -11758 194 -11757
rect 121 -11810 131 -11758
rect 183 -11810 194 -11758
rect 141 -11811 175 -11810
rect 230 -11919 264 -11448
rect 32 -11920 105 -11919
rect 32 -11972 42 -11920
rect 94 -11972 105 -11920
rect 210 -11920 283 -11919
rect 210 -11972 220 -11920
rect 272 -11972 283 -11920
rect 52 -12081 86 -11972
rect 230 -12080 264 -11972
rect 52 -13080 86 -12442
rect 141 -12653 175 -12384
rect 120 -12654 193 -12653
rect 120 -12706 130 -12654
rect 182 -12706 193 -12654
rect -1995 -13545 -1961 -13383
rect -2014 -13546 -1941 -13545
rect -2014 -13598 -2004 -13546
rect -1952 -13598 -1941 -13546
rect -1905 -14082 -1871 -13444
rect -1728 -14081 -1694 -13443
rect -1638 -13672 -1604 -13385
rect -1658 -13673 -1585 -13672
rect -1658 -13725 -1648 -13673
rect -1596 -13725 -1585 -13673
rect -1550 -14082 -1516 -13444
rect -1282 -13672 -1248 -13383
rect -927 -13672 -893 -13387
rect -571 -13545 -537 -13385
rect -591 -13546 -518 -13545
rect -591 -13598 -581 -13546
rect -529 -13598 -518 -13546
rect -1301 -13673 -1228 -13672
rect -1301 -13725 -1291 -13673
rect -1239 -13725 -1228 -13673
rect -947 -13673 -874 -13672
rect -947 -13725 -937 -13673
rect -885 -13725 -874 -13673
rect -927 -13726 -893 -13725
rect -304 -14081 -270 -13437
rect -216 -13794 -182 -13386
rect -235 -13795 -162 -13794
rect -235 -13847 -225 -13795
rect -173 -13847 -162 -13795
rect -125 -14082 -91 -13438
rect 52 -14081 86 -13437
rect 141 -13794 175 -12706
rect 230 -13080 264 -12442
rect 319 -13207 353 -10961
rect 408 -11919 442 -11448
rect 497 -11757 531 -11380
rect 477 -11758 550 -11757
rect 477 -11810 487 -11758
rect 539 -11810 550 -11758
rect 389 -11920 462 -11919
rect 389 -11972 399 -11920
rect 451 -11972 462 -11920
rect 408 -12081 442 -11972
rect 408 -13082 442 -12444
rect 496 -12784 530 -11810
rect 586 -11919 620 -11448
rect 567 -11920 640 -11919
rect 567 -11972 577 -11920
rect 629 -11972 640 -11920
rect 586 -12081 620 -11972
rect 476 -12785 549 -12784
rect 476 -12837 486 -12785
rect 538 -12837 549 -12785
rect 587 -13082 621 -12444
rect 675 -13231 709 -10961
rect 941 -11080 975 -10961
rect 853 -11438 887 -11362
rect 942 -11438 976 -11432
rect 1031 -11438 1065 -11357
rect 757 -11472 1159 -11438
rect 764 -12081 798 -12032
rect 942 -12081 976 -11472
rect 1120 -12080 1154 -12032
rect 852 -12438 886 -12353
rect 942 -12438 976 -12432
rect 1031 -12438 1065 -12377
rect 759 -12472 1160 -12438
rect 942 -13048 976 -12472
rect 761 -13082 1160 -13048
rect 852 -13154 886 -13082
rect 1032 -13165 1066 -13082
rect 1209 -13212 1243 -10961
rect 1299 -11081 1333 -10432
rect 1477 -11081 1511 -10432
rect 1546 -10909 1619 -10908
rect 1546 -10961 1556 -10909
rect 1608 -10961 1619 -10909
rect 1298 -11919 1332 -11448
rect 1387 -11528 1421 -11389
rect 1367 -11529 1440 -11528
rect 1367 -11581 1377 -11529
rect 1429 -11581 1440 -11529
rect 1477 -11919 1511 -11448
rect 1278 -11920 1351 -11919
rect 1278 -11972 1288 -11920
rect 1340 -11972 1351 -11920
rect 1458 -11920 1531 -11919
rect 1458 -11972 1468 -11920
rect 1520 -11972 1531 -11920
rect 1298 -12080 1332 -11972
rect 1477 -12081 1511 -11972
rect 1299 -13081 1333 -12443
rect 1388 -12783 1422 -12389
rect 1368 -12784 1441 -12783
rect 1368 -12836 1378 -12784
rect 1430 -12836 1441 -12784
rect 1388 -13187 1422 -12836
rect 1476 -13081 1510 -12443
rect 1566 -13217 1600 -10961
rect 1653 -11080 1687 -10431
rect 1832 -11082 1866 -10433
rect 1903 -10909 1976 -10908
rect 1903 -10961 1913 -10909
rect 1965 -10961 1976 -10909
rect 1654 -11920 1688 -11448
rect 1743 -11528 1777 -11386
rect 1723 -11529 1796 -11528
rect 1723 -11581 1733 -11529
rect 1785 -11581 1796 -11529
rect 1634 -11921 1707 -11920
rect 1634 -11973 1644 -11921
rect 1696 -11973 1707 -11921
rect 1654 -12080 1688 -11973
rect 1655 -13082 1689 -12444
rect 1744 -12654 1778 -11581
rect 1832 -11919 1866 -11448
rect 1813 -11920 1886 -11919
rect 1813 -11972 1823 -11920
rect 1875 -11972 1886 -11920
rect 1832 -12081 1866 -11972
rect 1725 -12655 1798 -12654
rect 1725 -12707 1735 -12655
rect 1787 -12707 1798 -12655
rect 1833 -13081 1867 -12443
rect 1922 -13187 1956 -10961
rect 2010 -11081 2044 -10432
rect 2188 -11081 2222 -10432
rect 2258 -10909 2331 -10908
rect 2258 -10961 2268 -10909
rect 2320 -10961 2331 -10909
rect 2613 -10909 2686 -10908
rect 2613 -10961 2623 -10909
rect 2675 -10961 2686 -10909
rect 2970 -10909 3043 -10908
rect 2970 -10961 2980 -10909
rect 3032 -10961 3043 -10909
rect 3325 -10909 3398 -10908
rect 3325 -10961 3335 -10909
rect 3387 -10961 3398 -10909
rect 2010 -11919 2044 -11448
rect 2099 -11528 2133 -11380
rect 2079 -11529 2152 -11528
rect 2079 -11581 2089 -11529
rect 2141 -11581 2152 -11529
rect 2188 -11919 2222 -11448
rect 1990 -11920 2063 -11919
rect 1990 -11972 2000 -11920
rect 2052 -11972 2063 -11920
rect 2168 -11920 2241 -11919
rect 2168 -11972 2178 -11920
rect 2230 -11972 2241 -11920
rect 2010 -12079 2044 -11972
rect 2188 -12079 2222 -11972
rect 2009 -13079 2043 -12441
rect 2098 -12782 2132 -12375
rect 2078 -12783 2151 -12782
rect 2078 -12835 2088 -12783
rect 2140 -12835 2151 -12783
rect 2098 -13193 2132 -12835
rect 2188 -13079 2222 -12441
rect 2277 -13199 2311 -10961
rect 2366 -11919 2400 -11448
rect 2456 -11637 2490 -11386
rect 2436 -11638 2509 -11637
rect 2436 -11690 2446 -11638
rect 2498 -11690 2509 -11638
rect 2544 -11919 2578 -11448
rect 2347 -11920 2420 -11919
rect 2347 -11972 2357 -11920
rect 2409 -11972 2420 -11920
rect 2524 -11920 2597 -11919
rect 2524 -11972 2534 -11920
rect 2586 -11972 2597 -11920
rect 2366 -12083 2400 -11972
rect 2544 -12081 2578 -11972
rect 2366 -13082 2400 -12444
rect 2455 -12653 2489 -12385
rect 2435 -12654 2508 -12653
rect 2435 -12706 2445 -12654
rect 2497 -12706 2508 -12654
rect 2544 -13082 2578 -12444
rect 2633 -13204 2667 -10961
rect 2722 -11919 2756 -11448
rect 2810 -11757 2844 -11387
rect 2790 -11758 2863 -11757
rect 2790 -11810 2800 -11758
rect 2852 -11810 2863 -11758
rect 2703 -11920 2776 -11919
rect 2703 -11972 2713 -11920
rect 2765 -11972 2776 -11920
rect 2722 -12080 2756 -11972
rect 2722 -13079 2756 -12441
rect 2811 -12782 2845 -11810
rect 2900 -11919 2934 -11448
rect 2880 -11920 2953 -11919
rect 2880 -11972 2890 -11920
rect 2942 -11972 2953 -11920
rect 2900 -12080 2934 -11972
rect 2791 -12783 2864 -12782
rect 2791 -12835 2801 -12783
rect 2853 -12835 2864 -12783
rect 2900 -13082 2934 -12444
rect 2989 -13212 3023 -10961
rect 3078 -11919 3112 -11448
rect 3166 -11757 3200 -11384
rect 3147 -11758 3220 -11757
rect 3147 -11810 3157 -11758
rect 3209 -11810 3220 -11758
rect 3256 -11919 3290 -11448
rect 3058 -11920 3131 -11919
rect 3058 -11972 3068 -11920
rect 3120 -11972 3131 -11920
rect 3237 -11920 3310 -11919
rect 3237 -11972 3247 -11920
rect 3299 -11972 3310 -11920
rect 3078 -12081 3112 -11972
rect 3256 -12080 3290 -11972
rect 3078 -13081 3112 -12443
rect 3167 -12650 3201 -12387
rect 3166 -12652 3201 -12650
rect 3148 -12653 3221 -12652
rect 3148 -12705 3158 -12653
rect 3210 -12705 3221 -12653
rect 123 -13795 196 -13794
rect 123 -13847 133 -13795
rect 185 -13847 196 -13795
rect 230 -14081 264 -13437
rect 408 -14081 442 -13437
rect 496 -13795 530 -13385
rect 477 -13796 550 -13795
rect 477 -13848 487 -13796
rect 539 -13848 550 -13796
rect 587 -14081 621 -13437
rect 942 -14048 976 -13430
rect 1388 -13672 1422 -13380
rect 1743 -13672 1777 -13382
rect 2100 -13672 2134 -13382
rect 1369 -13673 1442 -13672
rect 1369 -13725 1379 -13673
rect 1431 -13725 1442 -13673
rect 1722 -13673 1795 -13672
rect 1722 -13725 1732 -13673
rect 1784 -13725 1795 -13673
rect 2081 -13673 2154 -13672
rect 2081 -13725 2091 -13673
rect 2143 -13725 2154 -13673
rect 762 -14082 1159 -14048
rect 2366 -14081 2400 -13432
rect 2455 -13545 2489 -13388
rect 2436 -13546 2509 -13545
rect 2436 -13598 2446 -13546
rect 2498 -13598 2509 -13546
rect 2544 -14081 2578 -13432
rect 2723 -14082 2757 -13433
rect 2812 -13794 2846 -13379
rect 2792 -13795 2865 -13794
rect 2792 -13847 2802 -13795
rect 2854 -13847 2865 -13795
rect 2901 -14081 2935 -13432
rect 3078 -14082 3112 -13433
rect 3166 -13795 3200 -12705
rect 3256 -13082 3290 -12444
rect 3345 -13223 3379 -10961
rect 3434 -11082 3468 -10433
rect 3613 -11082 3647 -10433
rect 3682 -10909 3755 -10908
rect 3682 -10961 3692 -10909
rect 3744 -10961 3755 -10909
rect 3434 -11919 3468 -11448
rect 3522 -11757 3556 -11369
rect 3503 -11758 3576 -11757
rect 3503 -11810 3513 -11758
rect 3565 -11810 3576 -11758
rect 3612 -11919 3646 -11448
rect 3415 -11920 3488 -11919
rect 3415 -11972 3425 -11920
rect 3477 -11972 3488 -11920
rect 3593 -11920 3666 -11919
rect 3593 -11972 3603 -11920
rect 3655 -11972 3666 -11920
rect 3434 -12081 3468 -11972
rect 3612 -12080 3646 -11972
rect 3434 -13080 3468 -12442
rect 3524 -12542 3558 -12386
rect 3504 -12543 3577 -12542
rect 3504 -12595 3514 -12543
rect 3566 -12595 3577 -12543
rect 3613 -13080 3647 -12442
rect 3701 -13213 3735 -10961
rect 3791 -11081 3825 -10432
rect 3881 -11437 3915 -11232
rect 4056 -11437 4090 -11365
rect 3790 -11919 3824 -11448
rect 3881 -11471 4090 -11437
rect 3881 -11638 3915 -11471
rect 3861 -11639 3934 -11638
rect 3861 -11691 3871 -11639
rect 3923 -11691 3934 -11639
rect 3771 -11920 3844 -11919
rect 3771 -11972 3781 -11920
rect 3833 -11972 3844 -11920
rect 3790 -12079 3824 -11972
rect 3881 -12436 3915 -11691
rect 4058 -12436 4092 -12363
rect 3790 -13080 3824 -12442
rect 3881 -12470 4092 -12436
rect 3881 -12542 3915 -12470
rect 3861 -12543 3934 -12542
rect 3861 -12595 3871 -12543
rect 3923 -12595 3934 -12543
rect 3881 -13047 3915 -12595
rect 3881 -13081 4090 -13047
rect 3881 -13192 3915 -13081
rect 4056 -13165 4090 -13081
rect 3147 -13796 3220 -13795
rect 3147 -13848 3157 -13796
rect 3209 -13848 3220 -13796
rect 3257 -14080 3291 -13431
rect 3523 -13794 3557 -13336
rect 3879 -13545 3913 -13387
rect 3860 -13546 3933 -13545
rect 3860 -13598 3870 -13546
rect 3922 -13598 3933 -13546
rect 3502 -13795 3575 -13794
rect 3502 -13847 3512 -13795
rect 3564 -13847 3575 -13795
rect 3523 -13848 3557 -13847
rect 853 -14160 887 -14082
rect 1032 -14164 1066 -14082
rect -2173 -14441 -2139 -14361
rect -1995 -14441 -1961 -14228
rect -2173 -14475 -1961 -14441
rect -2325 -14544 -2252 -14543
rect -2325 -14596 -2315 -14544
rect -2263 -14596 -2252 -14544
rect -1995 -15045 -1961 -14475
rect -2176 -15079 -1961 -15045
rect -2176 -15163 -2142 -15079
rect -2457 -15822 -2384 -15821
rect -1995 -15822 -1961 -15079
rect -2457 -15874 -2447 -15822
rect -2395 -15874 -2384 -15822
rect -2015 -15823 -1942 -15822
rect -2015 -15875 -2005 -15823
rect -1953 -15875 -1942 -15823
rect -1995 -16050 -1961 -15875
rect -1906 -15933 -1872 -15441
rect -1925 -15934 -1852 -15933
rect -1925 -15986 -1915 -15934
rect -1863 -15986 -1852 -15934
rect -2173 -16084 -1961 -16050
rect -2173 -16156 -2139 -16084
rect -1995 -16132 -1961 -16084
rect -3945 -16347 -3935 -16295
rect -3883 -16347 -3873 -16295
rect -6028 -16886 -5994 -16750
rect -5939 -16886 -5905 -16794
rect -5850 -16886 -5816 -16750
rect -5672 -16886 -5638 -16750
rect -6028 -16920 -5816 -16886
rect -5850 -17007 -5816 -16920
rect -5692 -16887 -5619 -16886
rect -5692 -16939 -5682 -16887
rect -5630 -16939 -5619 -16887
rect -6169 -17008 -6096 -17007
rect -6169 -17060 -6159 -17008
rect -6107 -17060 -6096 -17008
rect -5869 -17008 -5796 -17007
rect -5869 -17060 -5859 -17008
rect -5807 -17060 -5796 -17008
rect -5494 -17118 -5460 -16751
rect -5316 -16886 -5282 -16750
rect -5336 -16887 -5263 -16886
rect -5336 -16939 -5326 -16887
rect -5274 -16939 -5263 -16887
rect -5138 -17007 -5104 -16751
rect -4960 -16886 -4926 -16751
rect -4980 -16887 -4907 -16886
rect -4980 -16939 -4970 -16887
rect -4918 -16939 -4907 -16887
rect -5158 -17008 -5085 -17007
rect -5158 -17060 -5148 -17008
rect -5096 -17060 -5085 -17008
rect -5514 -17119 -5441 -17118
rect -5514 -17171 -5504 -17119
rect -5452 -17171 -5441 -17119
rect -7605 -17251 -7329 -17250
rect -4970 -17251 -4917 -16939
rect -4782 -17118 -4748 -16751
rect -4604 -16886 -4570 -16751
rect -4624 -16887 -4551 -16886
rect -4624 -16939 -4614 -16887
rect -4562 -16939 -4551 -16887
rect -4426 -17007 -4392 -16750
rect -4248 -16886 -4214 -16750
rect -4159 -16886 -4125 -16794
rect -4070 -16886 -4036 -16750
rect -4268 -16887 -4036 -16886
rect -4268 -16939 -4258 -16887
rect -4206 -16939 -4036 -16887
rect -4447 -17008 -4374 -17007
rect -4447 -17060 -4437 -17008
rect -4385 -17060 -4374 -17008
rect -3935 -17118 -3883 -16347
rect -1906 -16542 -1872 -16438
rect -1927 -16543 -1854 -16542
rect -1927 -16595 -1917 -16543
rect -1865 -16595 -1854 -16543
rect -1817 -16665 -1783 -14309
rect -1728 -15933 -1694 -15438
rect -1639 -15822 -1605 -14231
rect -1659 -15823 -1586 -15822
rect -1659 -15875 -1649 -15823
rect -1597 -15875 -1586 -15823
rect -1748 -15934 -1675 -15933
rect -1748 -15986 -1738 -15934
rect -1686 -15986 -1675 -15934
rect -1639 -16135 -1605 -15875
rect -1550 -15933 -1516 -15438
rect -1570 -15934 -1497 -15933
rect -1570 -15986 -1560 -15934
rect -1508 -15986 -1497 -15934
rect -1728 -16542 -1694 -16440
rect -1550 -16541 -1516 -16439
rect -1571 -16542 -1498 -16541
rect -1748 -16543 -1675 -16542
rect -1748 -16595 -1738 -16543
rect -1686 -16595 -1675 -16543
rect -1571 -16594 -1561 -16542
rect -1509 -16594 -1498 -16542
rect -1837 -16666 -1764 -16665
rect -1837 -16718 -1827 -16666
rect -1775 -16718 -1764 -16666
rect -1736 -16666 -1528 -16655
rect -1461 -16666 -1427 -14309
rect -1371 -14543 -1337 -14438
rect -1391 -14544 -1318 -14543
rect -1391 -14596 -1381 -14544
rect -1329 -14596 -1318 -14544
rect -1371 -15076 -1337 -14596
rect -1372 -15933 -1338 -15440
rect -1283 -15822 -1249 -14234
rect -1194 -14543 -1160 -14438
rect -1214 -14544 -1141 -14543
rect -1214 -14596 -1204 -14544
rect -1152 -14596 -1141 -14544
rect -1303 -15823 -1230 -15822
rect -1303 -15875 -1293 -15823
rect -1241 -15875 -1230 -15823
rect -1392 -15934 -1319 -15933
rect -1392 -15986 -1382 -15934
rect -1330 -15986 -1319 -15934
rect -1283 -16138 -1249 -15875
rect -1194 -15933 -1160 -15438
rect -1214 -15934 -1141 -15933
rect -1214 -15986 -1204 -15934
rect -1152 -15986 -1141 -15934
rect -1372 -16543 -1338 -16440
rect -1194 -16542 -1160 -16440
rect -1214 -16543 -1141 -16542
rect -1391 -16544 -1318 -16543
rect -1391 -16596 -1381 -16544
rect -1329 -16596 -1318 -16544
rect -1214 -16595 -1204 -16543
rect -1152 -16595 -1141 -16543
rect -1104 -16665 -1070 -14312
rect -1016 -14543 -982 -14439
rect -1036 -14544 -963 -14543
rect -1036 -14596 -1026 -14544
rect -974 -14596 -963 -14544
rect -1015 -15933 -981 -15439
rect -927 -15822 -893 -14231
rect -838 -14543 -804 -14438
rect -858 -14544 -785 -14543
rect -858 -14596 -848 -14544
rect -796 -14596 -785 -14544
rect -857 -14927 -784 -14926
rect -857 -14979 -847 -14927
rect -795 -14979 -784 -14927
rect -838 -15081 -804 -14979
rect -947 -15823 -874 -15822
rect -947 -15875 -937 -15823
rect -885 -15875 -874 -15823
rect -1035 -15934 -962 -15933
rect -1035 -15986 -1025 -15934
rect -973 -15986 -962 -15934
rect -927 -16135 -893 -15875
rect -857 -15934 -784 -15933
rect -857 -15986 -847 -15934
rect -795 -15986 -784 -15934
rect -838 -16080 -804 -15986
rect -1016 -16542 -982 -16439
rect -1036 -16543 -963 -16542
rect -1036 -16595 -1026 -16543
rect -974 -16595 -963 -16543
rect -749 -16664 -715 -14310
rect -659 -14543 -625 -14440
rect -679 -14544 -606 -14543
rect -679 -14596 -669 -14544
rect -617 -14596 -606 -14544
rect -679 -14927 -606 -14926
rect -679 -14979 -669 -14927
rect -617 -14979 -606 -14927
rect -660 -15081 -626 -14979
rect -571 -15822 -537 -14231
rect -482 -14543 -448 -14439
rect -501 -14544 -428 -14543
rect -501 -14596 -491 -14544
rect -439 -14596 -428 -14544
rect -501 -14927 -428 -14926
rect -501 -14979 -491 -14927
rect -439 -14979 -428 -14927
rect -481 -15081 -447 -14979
rect -591 -15823 -518 -15822
rect -591 -15875 -581 -15823
rect -529 -15875 -518 -15823
rect -680 -15934 -607 -15933
rect -680 -15986 -670 -15934
rect -618 -15986 -607 -15934
rect -660 -16082 -626 -15986
rect -571 -16135 -537 -15875
rect -501 -15934 -428 -15933
rect -501 -15986 -491 -15934
rect -439 -15986 -428 -15934
rect -482 -16081 -448 -15986
rect -769 -16665 -696 -16664
rect -1124 -16666 -1051 -16665
rect -1736 -16718 -1692 -16666
rect -1640 -16718 -1628 -16666
rect -1576 -16718 -1528 -16666
rect -4802 -17119 -4729 -17118
rect -4802 -17171 -4792 -17119
rect -4740 -17171 -4729 -17119
rect -3945 -17170 -3935 -17118
rect -3883 -17170 -3873 -17118
rect -1736 -17251 -1528 -16718
rect -1481 -16667 -1408 -16666
rect -1481 -16719 -1471 -16667
rect -1419 -16719 -1408 -16667
rect -1124 -16718 -1114 -16666
rect -1062 -16718 -1051 -16666
rect -769 -16717 -759 -16665
rect -707 -16717 -696 -16665
rect -658 -16666 -450 -16656
rect -393 -16665 -359 -14306
rect -304 -14927 -270 -14437
rect -324 -14928 -251 -14927
rect -324 -14980 -314 -14928
rect -262 -14980 -251 -14928
rect -304 -15081 -270 -14980
rect -215 -15822 -181 -14230
rect -126 -14926 -92 -14440
rect -147 -14927 -74 -14926
rect -147 -14979 -137 -14927
rect -85 -14979 -74 -14927
rect -126 -15081 -92 -14979
rect -235 -15823 -162 -15822
rect -235 -15875 -225 -15823
rect -173 -15875 -162 -15823
rect -323 -15934 -250 -15933
rect -323 -15986 -313 -15934
rect -261 -15986 -250 -15934
rect -304 -16080 -270 -15986
rect -215 -16134 -181 -15875
rect -146 -15934 -73 -15933
rect -146 -15986 -136 -15934
rect -84 -15986 -73 -15934
rect -126 -16080 -92 -15986
rect -37 -16665 -3 -14312
rect 52 -14926 86 -14445
rect 33 -14927 106 -14926
rect 33 -14979 43 -14927
rect 95 -14979 106 -14927
rect 52 -15081 86 -14979
rect 141 -15821 175 -14231
rect 122 -15822 195 -15821
rect 122 -15874 132 -15822
rect 184 -15874 195 -15822
rect 33 -15934 106 -15933
rect 33 -15986 43 -15934
rect 95 -15986 106 -15934
rect 52 -16080 86 -15986
rect 141 -16135 175 -15874
rect 230 -15933 264 -15439
rect 211 -15934 284 -15933
rect 211 -15986 221 -15934
rect 273 -15986 284 -15934
rect 230 -16542 264 -16438
rect 210 -16543 283 -16542
rect 210 -16595 220 -16543
rect 272 -16595 283 -16543
rect -658 -16718 -617 -16666
rect -565 -16718 -553 -16666
rect -501 -16718 -450 -16666
rect -413 -16666 -340 -16665
rect -413 -16718 -403 -16666
rect -351 -16718 -340 -16666
rect -57 -16666 16 -16665
rect 319 -16666 353 -14307
rect 408 -15933 442 -15439
rect 497 -15822 531 -14231
rect 477 -15823 550 -15822
rect 477 -15875 487 -15823
rect 539 -15875 550 -15823
rect 388 -15934 461 -15933
rect 388 -15986 398 -15934
rect 450 -15986 461 -15934
rect 497 -16135 531 -15875
rect 585 -15933 619 -15439
rect 565 -15934 638 -15933
rect 565 -15986 575 -15934
rect 627 -15986 638 -15934
rect 408 -16542 442 -16439
rect 586 -16542 620 -16439
rect 387 -16543 460 -16542
rect 387 -16595 397 -16543
rect 449 -16595 460 -16543
rect 566 -16543 639 -16542
rect 566 -16595 576 -16543
rect 628 -16595 639 -16543
rect 408 -16666 616 -16649
rect 675 -16665 709 -14307
rect 764 -15933 798 -15438
rect 853 -15822 887 -15340
rect 833 -15823 906 -15822
rect 833 -15875 843 -15823
rect 895 -15875 906 -15823
rect 745 -15934 818 -15933
rect 745 -15986 755 -15934
rect 807 -15986 818 -15934
rect 853 -16136 887 -15875
rect 941 -15933 975 -15439
rect 921 -15934 994 -15933
rect 921 -15986 931 -15934
rect 983 -15986 994 -15934
rect 765 -16542 799 -16438
rect 943 -16542 977 -16439
rect 745 -16543 818 -16542
rect 745 -16595 755 -16543
rect 807 -16595 818 -16543
rect 923 -16543 996 -16542
rect 923 -16595 933 -16543
rect 985 -16595 996 -16543
rect 1031 -16665 1065 -14308
rect 1120 -15933 1154 -15440
rect 1209 -15822 1243 -14231
rect 1298 -14543 1332 -14439
rect 1278 -14544 1351 -14543
rect 1278 -14596 1288 -14544
rect 1340 -14596 1351 -14544
rect 1279 -14928 1352 -14927
rect 1279 -14980 1289 -14928
rect 1341 -14980 1352 -14928
rect 1298 -15081 1332 -14980
rect 1191 -15823 1264 -15822
rect 1191 -15875 1201 -15823
rect 1253 -15875 1264 -15823
rect 1100 -15934 1173 -15933
rect 1100 -15986 1110 -15934
rect 1162 -15986 1173 -15934
rect 1209 -16135 1243 -15875
rect 1279 -15934 1352 -15933
rect 1279 -15986 1289 -15934
rect 1341 -15986 1352 -15934
rect 1298 -16081 1332 -15986
rect 1120 -16542 1154 -16439
rect 1101 -16543 1174 -16542
rect 1101 -16595 1111 -16543
rect 1163 -16595 1174 -16543
rect 1387 -16665 1421 -14307
rect 1477 -14543 1511 -14439
rect 1456 -14544 1529 -14543
rect 1456 -14596 1466 -14544
rect 1518 -14596 1529 -14544
rect 1457 -14927 1530 -14926
rect 1457 -14979 1467 -14927
rect 1519 -14979 1530 -14927
rect 1476 -15081 1510 -14979
rect 1565 -15822 1599 -14231
rect 1654 -14543 1688 -14438
rect 1634 -14544 1707 -14543
rect 1634 -14596 1644 -14544
rect 1696 -14596 1707 -14544
rect 1634 -14927 1707 -14926
rect 1634 -14979 1644 -14927
rect 1696 -14979 1707 -14927
rect 1654 -15082 1688 -14979
rect 1545 -15823 1618 -15822
rect 1545 -15875 1555 -15823
rect 1607 -15875 1618 -15823
rect 1456 -15934 1529 -15933
rect 1456 -15986 1466 -15934
rect 1518 -15986 1529 -15934
rect 1476 -16082 1510 -15986
rect 1565 -16135 1599 -15875
rect 1633 -15934 1706 -15933
rect 1633 -15986 1643 -15934
rect 1695 -15986 1706 -15934
rect 1653 -16081 1687 -15986
rect -57 -16718 -47 -16666
rect 5 -16718 16 -16666
rect 299 -16667 372 -16666
rect -658 -17251 -450 -16718
rect 299 -16719 309 -16667
rect 361 -16719 372 -16667
rect 408 -16718 452 -16666
rect 504 -16718 516 -16666
rect 568 -16718 616 -16666
rect 655 -16666 728 -16665
rect 655 -16718 665 -16666
rect 717 -16718 728 -16666
rect 1011 -16666 1084 -16665
rect 1011 -16718 1021 -16666
rect 1073 -16718 1084 -16666
rect 1367 -16666 1440 -16665
rect 1367 -16718 1377 -16666
rect 1429 -16718 1440 -16666
rect 1488 -16666 1696 -16658
rect 1744 -16665 1778 -14312
rect 1832 -14542 1866 -14438
rect 1813 -14543 1886 -14542
rect 1813 -14595 1823 -14543
rect 1875 -14595 1886 -14543
rect 1812 -14927 1885 -14926
rect 1812 -14979 1822 -14927
rect 1874 -14979 1885 -14927
rect 1833 -15081 1867 -14979
rect 1921 -15822 1955 -14231
rect 2010 -14543 2044 -14438
rect 1990 -14544 2063 -14543
rect 1990 -14596 2000 -14544
rect 2052 -14596 2063 -14544
rect 1989 -14927 2062 -14926
rect 1989 -14979 1999 -14927
rect 2051 -14979 2062 -14927
rect 2010 -15082 2044 -14979
rect 1900 -15823 1973 -15822
rect 1900 -15875 1910 -15823
rect 1962 -15875 1973 -15823
rect 1812 -15934 1885 -15933
rect 1812 -15986 1822 -15934
rect 1874 -15986 1885 -15934
rect 1832 -16080 1866 -15986
rect 1921 -16135 1955 -15875
rect 1990 -15934 2063 -15933
rect 1990 -15986 2000 -15934
rect 2052 -15986 2063 -15934
rect 2010 -16081 2044 -15986
rect 2100 -16664 2134 -14313
rect 2188 -14543 2222 -14439
rect 2168 -14544 2241 -14543
rect 2168 -14596 2178 -14544
rect 2230 -14596 2241 -14544
rect 2170 -14927 2243 -14926
rect 2170 -14979 2180 -14927
rect 2232 -14979 2243 -14927
rect 2189 -15081 2223 -14979
rect 2277 -15822 2311 -14231
rect 2257 -15823 2330 -15822
rect 2257 -15875 2267 -15823
rect 2319 -15875 2330 -15823
rect 2169 -15934 2242 -15933
rect 2169 -15986 2179 -15934
rect 2231 -15986 2242 -15934
rect 2189 -16081 2223 -15986
rect 2277 -16135 2311 -15875
rect 2366 -15933 2400 -15440
rect 2346 -15934 2419 -15933
rect 2346 -15986 2356 -15934
rect 2408 -15986 2419 -15934
rect 2366 -16542 2400 -16439
rect 2346 -16543 2419 -16542
rect 2346 -16595 2356 -16543
rect 2408 -16595 2419 -16543
rect 2080 -16665 2153 -16664
rect 2455 -16665 2489 -14311
rect 2544 -15933 2578 -15440
rect 2633 -15822 2667 -14232
rect 2614 -15823 2687 -15822
rect 2614 -15875 2624 -15823
rect 2676 -15875 2687 -15823
rect 2524 -15934 2597 -15933
rect 2524 -15986 2534 -15934
rect 2586 -15986 2597 -15934
rect 2633 -16136 2667 -15875
rect 2722 -15933 2756 -15440
rect 2702 -15934 2775 -15933
rect 2702 -15986 2712 -15934
rect 2764 -15986 2775 -15934
rect 2544 -16542 2578 -16439
rect 2722 -16541 2756 -16441
rect 2703 -16542 2776 -16541
rect 2524 -16543 2597 -16542
rect 2524 -16595 2534 -16543
rect 2586 -16595 2597 -16543
rect 2703 -16594 2713 -16542
rect 2765 -16594 2776 -16542
rect 1488 -16718 1528 -16666
rect 1580 -16718 1592 -16666
rect 1644 -16718 1696 -16666
rect 1725 -16666 1798 -16665
rect 1725 -16718 1735 -16666
rect 1787 -16718 1798 -16666
rect 2080 -16717 2090 -16665
rect 2142 -16717 2153 -16665
rect 2435 -16666 2508 -16665
rect 2435 -16718 2445 -16666
rect 2497 -16718 2508 -16666
rect 2547 -16666 2755 -16653
rect 2811 -16665 2845 -14310
rect 2900 -15933 2934 -15439
rect 2989 -15822 3023 -14231
rect 2969 -15823 3042 -15822
rect 2969 -15875 2979 -15823
rect 3031 -15875 3042 -15823
rect 2881 -15934 2954 -15933
rect 2881 -15986 2891 -15934
rect 2943 -15986 2954 -15934
rect 2989 -16135 3023 -15875
rect 3078 -15933 3112 -15438
rect 3058 -15934 3131 -15933
rect 3058 -15986 3068 -15934
rect 3120 -15986 3131 -15934
rect 2901 -16542 2935 -16441
rect 3079 -16542 3113 -16439
rect 2881 -16543 2954 -16542
rect 2881 -16595 2891 -16543
rect 2943 -16595 2954 -16543
rect 3060 -16543 3133 -16542
rect 3060 -16595 3070 -16543
rect 3122 -16595 3133 -16543
rect 3167 -16664 3201 -14315
rect 3236 -14545 3309 -14544
rect 3236 -14597 3246 -14545
rect 3298 -14597 3309 -14545
rect 3256 -15080 3290 -14597
rect 3256 -15933 3290 -15439
rect 3345 -15822 3379 -14231
rect 3434 -14543 3468 -14439
rect 3414 -14544 3487 -14543
rect 3414 -14596 3424 -14544
rect 3476 -14596 3487 -14544
rect 3415 -14927 3488 -14926
rect 3415 -14979 3425 -14927
rect 3477 -14979 3488 -14927
rect 3434 -15081 3468 -14979
rect 3325 -15823 3398 -15822
rect 3325 -15875 3335 -15823
rect 3387 -15875 3398 -15823
rect 3237 -15934 3310 -15933
rect 3237 -15986 3247 -15934
rect 3299 -15986 3310 -15934
rect 3345 -16135 3379 -15875
rect 3414 -15934 3487 -15933
rect 3414 -15986 3424 -15934
rect 3476 -15986 3487 -15934
rect 3434 -16081 3468 -15986
rect 3257 -16542 3291 -16440
rect 3239 -16543 3312 -16542
rect 3239 -16595 3249 -16543
rect 3301 -16595 3312 -16543
rect 3147 -16665 3220 -16664
rect 2547 -16718 2592 -16666
rect 2644 -16718 2656 -16666
rect 2708 -16718 2755 -16666
rect 2791 -16666 2864 -16665
rect 2791 -16718 2801 -16666
rect 2853 -16718 2864 -16666
rect 3147 -16717 3157 -16665
rect 3209 -16717 3220 -16665
rect 3524 -16666 3558 -14310
rect 3612 -14543 3646 -14439
rect 3592 -14544 3665 -14543
rect 3592 -14596 3602 -14544
rect 3654 -14596 3665 -14544
rect 3593 -14927 3666 -14926
rect 3593 -14979 3603 -14927
rect 3655 -14979 3666 -14927
rect 3612 -15082 3646 -14979
rect 3701 -15822 3735 -14232
rect 3879 -14439 3913 -14307
rect 4057 -14439 4091 -14357
rect 3791 -14543 3825 -14439
rect 3879 -14473 4091 -14439
rect 3771 -14544 3844 -14543
rect 3771 -14596 3781 -14544
rect 3833 -14596 3844 -14544
rect 3770 -14927 3843 -14926
rect 3770 -14979 3780 -14927
rect 3832 -14979 3843 -14927
rect 3790 -15082 3824 -14979
rect 3879 -15047 3913 -14473
rect 4905 -14545 4958 -7905
rect 5037 -13296 5090 -7903
rect 5174 -7908 5184 -7856
rect 5236 -7908 5247 -7856
rect 5327 -7903 5337 -7851
rect 5389 -7903 5400 -7851
rect 5185 -8635 5237 -7908
rect 5175 -8687 5185 -8635
rect 5237 -8687 5247 -8635
rect 5337 -9925 5390 -7903
rect 11647 -8716 11681 -8715
rect 11044 -8717 11117 -8716
rect 6690 -8760 6815 -8726
rect 6690 -8907 6724 -8760
rect 6781 -8844 6815 -8760
rect 11044 -8769 11054 -8717
rect 11106 -8769 11117 -8717
rect 11335 -8717 11408 -8716
rect 11335 -8769 11345 -8717
rect 11397 -8769 11408 -8717
rect 11628 -8717 11701 -8716
rect 11628 -8769 11638 -8717
rect 11690 -8769 11701 -8717
rect 11922 -8717 11995 -8716
rect 11922 -8769 11932 -8717
rect 11984 -8769 11995 -8717
rect 12212 -8717 12285 -8716
rect 12212 -8769 12222 -8717
rect 12274 -8769 12285 -8717
rect 9004 -8842 9395 -8808
rect 6513 -9201 6547 -9125
rect 6689 -9201 6723 -8954
rect 6513 -9235 6723 -9201
rect 6779 -9314 6813 -9198
rect 6759 -9315 6832 -9314
rect 6759 -9367 6769 -9315
rect 6821 -9367 6832 -9315
rect 6669 -9546 6742 -9545
rect 6669 -9598 6679 -9546
rect 6731 -9598 6742 -9546
rect 5327 -9926 5400 -9925
rect 5327 -9978 5337 -9926
rect 5389 -9978 5400 -9926
rect 6513 -10099 6547 -10017
rect 6690 -10099 6724 -9598
rect 6779 -9740 6813 -9367
rect 6513 -10133 6724 -10099
rect 6690 -10313 6724 -10133
rect 6670 -10314 6743 -10313
rect 6670 -10366 6680 -10314
rect 6732 -10366 6743 -10314
rect 6868 -10467 6902 -9042
rect 6957 -9315 6991 -9197
rect 6937 -9316 7010 -9315
rect 6937 -9368 6947 -9316
rect 6999 -9368 7010 -9316
rect 6957 -9621 6991 -9368
rect 7046 -9621 7080 -9046
rect 7135 -9315 7169 -9198
rect 7116 -9316 7189 -9315
rect 7116 -9368 7126 -9316
rect 7178 -9368 7189 -9316
rect 6957 -9655 7080 -9621
rect 6957 -9743 6991 -9655
rect 6848 -10468 6921 -10467
rect 6848 -10520 6858 -10468
rect 6910 -10520 6921 -10468
rect 6510 -11003 6544 -10910
rect 6688 -11003 6722 -10920
rect 6868 -11003 6902 -10520
rect 6958 -10643 6992 -10097
rect 6510 -11037 6902 -11003
rect 6511 -11900 6545 -11823
rect 6688 -11900 6722 -11819
rect 6868 -11900 6902 -11037
rect 6958 -11544 6992 -10995
rect 7046 -11366 7080 -9655
rect 7135 -9744 7169 -9368
rect 7136 -10643 7170 -10097
rect 7224 -10466 7258 -9049
rect 7313 -9313 7347 -9197
rect 7293 -9314 7366 -9313
rect 7293 -9366 7303 -9314
rect 7355 -9366 7366 -9314
rect 7313 -9743 7347 -9366
rect 7204 -10467 7277 -10466
rect 7204 -10519 7214 -10467
rect 7266 -10519 7277 -10467
rect 7027 -11367 7100 -11366
rect 7027 -11419 7037 -11367
rect 7089 -11419 7100 -11367
rect 7046 -11671 7080 -11419
rect 7135 -11543 7169 -10994
rect 6511 -11934 6902 -11900
rect 6868 -12040 6902 -11934
rect 7224 -12040 7258 -10519
rect 7313 -10644 7347 -10098
rect 7313 -11542 7347 -10993
rect 7402 -11366 7436 -9048
rect 7491 -9313 7525 -9198
rect 7472 -9314 7545 -9313
rect 7472 -9366 7482 -9314
rect 7534 -9366 7545 -9314
rect 7491 -9744 7525 -9366
rect 7492 -10643 7526 -10097
rect 7580 -10466 7614 -9051
rect 7669 -9315 7703 -9198
rect 7649 -9316 7722 -9315
rect 7649 -9368 7659 -9316
rect 7711 -9368 7722 -9316
rect 7669 -9744 7703 -9368
rect 7561 -10467 7634 -10466
rect 7561 -10519 7571 -10467
rect 7623 -10519 7634 -10467
rect 7383 -11367 7456 -11366
rect 7383 -11419 7393 -11367
rect 7445 -11419 7456 -11367
rect 7402 -11673 7436 -11419
rect 7491 -11542 7525 -10993
rect 7580 -12040 7614 -10519
rect 7669 -10644 7703 -10098
rect 7669 -11542 7703 -10993
rect 7758 -11367 7792 -9054
rect 7847 -9314 7881 -9198
rect 7827 -9315 7900 -9314
rect 7827 -9367 7837 -9315
rect 7889 -9367 7900 -9315
rect 7847 -9744 7881 -9367
rect 7847 -10643 7881 -10097
rect 7936 -10466 7970 -9051
rect 8025 -9315 8059 -9198
rect 8005 -9316 8078 -9315
rect 8005 -9368 8015 -9316
rect 8067 -9368 8078 -9316
rect 8025 -9744 8059 -9368
rect 7917 -10467 7990 -10466
rect 7917 -10519 7927 -10467
rect 7979 -10519 7990 -10467
rect 7738 -11368 7811 -11367
rect 7738 -11420 7748 -11368
rect 7800 -11420 7811 -11368
rect 7758 -11679 7792 -11420
rect 7848 -11542 7882 -10993
rect 7936 -12040 7970 -10519
rect 8025 -10643 8059 -10097
rect 8024 -11543 8058 -10994
rect 8113 -11366 8147 -9056
rect 8203 -9314 8237 -9198
rect 8184 -9315 8257 -9314
rect 8184 -9367 8194 -9315
rect 8246 -9367 8257 -9315
rect 8203 -9744 8237 -9367
rect 8203 -10642 8237 -10096
rect 8292 -10467 8326 -9060
rect 8381 -9314 8415 -9198
rect 8361 -9315 8434 -9314
rect 8361 -9367 8371 -9315
rect 8423 -9367 8434 -9315
rect 8381 -9744 8415 -9367
rect 8273 -10468 8346 -10467
rect 8273 -10520 8283 -10468
rect 8335 -10520 8346 -10468
rect 8093 -11367 8166 -11366
rect 8093 -11419 8103 -11367
rect 8155 -11419 8166 -11367
rect 8113 -11681 8147 -11419
rect 8203 -11544 8237 -10995
rect 8292 -12040 8326 -10520
rect 8382 -10644 8416 -10098
rect 8381 -11543 8415 -10994
rect 8470 -11366 8504 -9056
rect 8559 -9314 8593 -9198
rect 8539 -9315 8612 -9314
rect 8539 -9367 8549 -9315
rect 8601 -9367 8612 -9315
rect 8559 -9744 8593 -9367
rect 8559 -10642 8593 -10096
rect 8648 -10466 8682 -9064
rect 8737 -9315 8771 -9198
rect 8717 -9316 8790 -9315
rect 8717 -9368 8727 -9316
rect 8779 -9368 8790 -9316
rect 8737 -9744 8771 -9368
rect 8628 -10467 8701 -10466
rect 8628 -10519 8638 -10467
rect 8690 -10519 8701 -10467
rect 8451 -11367 8524 -11366
rect 8451 -11419 8461 -11367
rect 8513 -11419 8524 -11367
rect 8470 -11681 8504 -11419
rect 8559 -11543 8593 -10994
rect 8648 -12040 8682 -10519
rect 8737 -10644 8771 -10098
rect 8737 -11543 8771 -10994
rect 8826 -11366 8860 -9063
rect 9004 -9068 9038 -8842
rect 9183 -8926 9217 -8842
rect 9361 -8923 9395 -8842
rect 8915 -9314 8949 -9198
rect 8896 -9315 8969 -9314
rect 8896 -9367 8906 -9315
rect 8958 -9367 8969 -9315
rect 8915 -9744 8949 -9367
rect 9004 -9709 9038 -9113
rect 11063 -9145 11097 -8769
rect 11354 -8986 11388 -8769
rect 11647 -8981 11681 -8769
rect 11941 -9011 11975 -8769
rect 12231 -8840 12265 -8769
rect 12231 -8874 12738 -8840
rect 12231 -9013 12265 -8874
rect 12522 -8947 12556 -8874
rect 12704 -8953 12738 -8874
rect 10968 -9152 11097 -9145
rect 10772 -9230 10806 -9156
rect 10950 -9179 11097 -9152
rect 10950 -9230 10984 -9179
rect 10772 -9264 10984 -9230
rect 10861 -9638 10895 -9264
rect 11063 -9387 11097 -9179
rect 11154 -9374 11188 -9259
rect 11134 -9375 11207 -9374
rect 11134 -9387 11144 -9375
rect 11063 -9421 11144 -9387
rect 11134 -9427 11144 -9421
rect 11196 -9427 11207 -9375
rect 11154 -9642 11188 -9427
rect 9004 -9743 9394 -9709
rect 11242 -9716 11276 -9180
rect 11445 -9375 11479 -9252
rect 11426 -9376 11499 -9375
rect 11426 -9428 11436 -9376
rect 11488 -9428 11499 -9376
rect 11445 -9635 11479 -9428
rect 11534 -9706 11568 -9170
rect 11738 -9375 11772 -9256
rect 11718 -9376 11791 -9375
rect 11718 -9428 11728 -9376
rect 11780 -9428 11791 -9376
rect 11738 -9639 11772 -9428
rect 11825 -9711 11859 -9175
rect 12030 -9376 12064 -9251
rect 12010 -9377 12083 -9376
rect 12010 -9429 12020 -9377
rect 12072 -9429 12083 -9377
rect 12030 -9634 12064 -9429
rect 12118 -9704 12152 -9168
rect 12321 -9375 12355 -9252
rect 12302 -9376 12375 -9375
rect 12302 -9428 12312 -9376
rect 12364 -9428 12375 -9376
rect 12321 -9635 12355 -9428
rect 12410 -9718 12444 -9182
rect 12613 -9610 12647 -9228
rect 12525 -9644 12736 -9610
rect 12525 -9737 12559 -9644
rect 12702 -9731 12736 -9644
rect 8915 -10643 8949 -10097
rect 9004 -10467 9038 -9743
rect 9182 -9824 9216 -9743
rect 9360 -9833 9394 -9743
rect 10773 -10001 10807 -9926
rect 10951 -10001 10985 -9912
rect 10773 -10035 10985 -10001
rect 9161 -10315 9234 -10314
rect 9161 -10367 9171 -10315
rect 9223 -10367 9234 -10315
rect 8985 -10468 9058 -10467
rect 8985 -10520 8995 -10468
rect 9047 -10520 9058 -10468
rect 8807 -11367 8880 -11366
rect 8807 -11419 8817 -11367
rect 8869 -11419 8880 -11367
rect 8826 -11688 8860 -11419
rect 8915 -11543 8949 -10994
rect 9004 -11679 9038 -10520
rect 9181 -10614 9215 -10367
rect 10862 -10380 10896 -10035
rect 10772 -10414 10986 -10380
rect 10772 -10485 10806 -10414
rect 10952 -10507 10986 -10414
rect 11063 -10490 11097 -9954
rect 11153 -10400 11187 -10017
rect 11356 -10481 11390 -9941
rect 11446 -10400 11480 -10017
rect 11648 -10486 11682 -9946
rect 11737 -10400 11771 -10017
rect 11940 -10482 11974 -9942
rect 12028 -10399 12062 -10016
rect 12232 -10488 12266 -9948
rect 12320 -10398 12354 -10015
rect 12613 -10413 12647 -9999
rect 9181 -10648 9393 -10614
rect 9181 -10695 9215 -10648
rect 9359 -10726 9393 -10648
rect 9093 -11541 9127 -11005
rect 10772 -11149 10806 -11148
rect 10860 -11149 10894 -10785
rect 10772 -11183 10986 -11149
rect 11152 -11175 11186 -10792
rect 10772 -11253 10806 -11183
rect 10952 -11268 10986 -11183
rect 11244 -11260 11278 -10720
rect 11446 -11171 11480 -10788
rect 11534 -11258 11568 -10718
rect 11737 -11173 11771 -10790
rect 11826 -11260 11860 -10720
rect 12029 -11172 12063 -10789
rect 12118 -11263 12152 -10723
rect 12322 -11171 12356 -10788
rect 12410 -11263 12444 -10723
rect 12525 -10772 12559 -10649
rect 12613 -10772 12647 -10770
rect 12700 -10772 12734 -10681
rect 12525 -10806 12734 -10772
rect 12613 -11184 12647 -10806
rect 9182 -11544 9394 -11510
rect 8912 -11985 8946 -11900
rect 9095 -11985 9129 -11900
rect 9182 -11985 9216 -11544
rect 9360 -11633 9394 -11544
rect 11063 -11674 11097 -11383
rect 11043 -11675 11116 -11674
rect 11356 -11675 11390 -11417
rect 11648 -11674 11682 -11402
rect 11940 -11674 11974 -11405
rect 12233 -11674 12267 -11403
rect 12525 -11541 12559 -11396
rect 12701 -11541 12735 -11460
rect 12525 -11575 12735 -11541
rect 13012 -11674 13085 -11673
rect 11628 -11675 11701 -11674
rect 11043 -11727 11053 -11675
rect 11105 -11727 11116 -11675
rect 11337 -11676 11410 -11675
rect 11337 -11728 11347 -11676
rect 11399 -11728 11410 -11676
rect 11628 -11727 11638 -11675
rect 11690 -11727 11701 -11675
rect 11921 -11675 11994 -11674
rect 11921 -11727 11931 -11675
rect 11983 -11727 11994 -11675
rect 12213 -11675 12286 -11674
rect 12213 -11727 12223 -11675
rect 12275 -11727 12286 -11675
rect 13012 -11726 13022 -11674
rect 13074 -11726 13085 -11674
rect 8912 -12019 9216 -11985
rect 6868 -12074 8682 -12040
rect 5027 -13297 5100 -13296
rect 5027 -13349 5037 -13297
rect 5089 -13349 5100 -13297
rect 5524 -13297 5597 -13296
rect 5524 -13349 5534 -13297
rect 5586 -13349 5597 -13297
rect 5021 -13434 5094 -13433
rect 5021 -13486 5031 -13434
rect 5083 -13486 5094 -13434
rect 4895 -14546 4968 -14545
rect 4895 -14598 4905 -14546
rect 4957 -14598 4968 -14546
rect 4229 -14927 4302 -14926
rect 4229 -14979 4239 -14927
rect 4291 -14979 4302 -14927
rect 3879 -15081 4091 -15047
rect 3682 -15823 3755 -15822
rect 3682 -15875 3692 -15823
rect 3744 -15875 3755 -15823
rect 3593 -15934 3666 -15933
rect 3593 -15986 3603 -15934
rect 3655 -15986 3666 -15934
rect 3612 -16080 3646 -15986
rect 3701 -16136 3735 -15875
rect 3770 -15934 3843 -15933
rect 3770 -15986 3780 -15934
rect 3832 -15986 3843 -15934
rect 3790 -16080 3824 -15986
rect 3879 -16047 3913 -15081
rect 4057 -15169 4091 -15081
rect 4238 -15539 4291 -14979
rect 4228 -15540 4301 -15539
rect 5031 -15540 5084 -13486
rect 5390 -13546 5463 -13545
rect 5390 -13598 5400 -13546
rect 5452 -13598 5463 -13546
rect 5132 -13795 5205 -13794
rect 5132 -13847 5142 -13795
rect 5194 -13847 5205 -13795
rect 5142 -14658 5195 -13847
rect 5133 -14659 5206 -14658
rect 5133 -14711 5143 -14659
rect 5195 -14711 5206 -14659
rect 4228 -15592 4238 -15540
rect 4290 -15592 4301 -15540
rect 5021 -15541 5094 -15540
rect 3879 -16081 4090 -16047
rect 3614 -16666 3822 -16658
rect 3879 -16665 3913 -16081
rect 4056 -16170 4090 -16081
rect 4238 -16542 4291 -15592
rect 5021 -15593 5031 -15541
rect 5083 -15593 5094 -15541
rect 4228 -16543 4301 -16542
rect 4228 -16595 4238 -16543
rect 4290 -16595 4301 -16543
rect 3504 -16667 3577 -16666
rect 408 -17251 616 -16718
rect 1488 -17251 1696 -16718
rect 2547 -17251 2755 -16718
rect 3504 -16719 3514 -16667
rect 3566 -16719 3577 -16667
rect 3614 -16718 3660 -16666
rect 3712 -16718 3724 -16666
rect 3776 -16718 3822 -16666
rect 3858 -16666 3931 -16665
rect 3858 -16718 3868 -16666
rect 3920 -16718 3931 -16666
rect 3614 -17251 3822 -16718
rect 5031 -16782 5084 -15593
rect 5400 -15653 5453 -13598
rect 5534 -13672 5587 -13349
rect 5524 -13673 5597 -13672
rect 5524 -13725 5534 -13673
rect 5586 -13725 5597 -13673
rect 6912 -13922 6946 -12074
rect 8940 -13434 9013 -13433
rect 8940 -13486 8950 -13434
rect 9002 -13486 9013 -13434
rect 9295 -13434 9368 -13433
rect 9295 -13486 9305 -13434
rect 9357 -13486 9368 -13434
rect 8762 -13557 8835 -13556
rect 8762 -13609 8772 -13557
rect 8824 -13609 8835 -13557
rect 8228 -13672 8301 -13671
rect 7516 -13673 7589 -13672
rect 7516 -13725 7526 -13673
rect 7578 -13725 7589 -13673
rect 7872 -13674 7945 -13673
rect 7338 -13797 7411 -13796
rect 7338 -13849 7348 -13797
rect 7400 -13849 7411 -13797
rect 5823 -13923 5896 -13922
rect 5823 -13975 5833 -13923
rect 5885 -13975 5896 -13923
rect 6003 -13923 6076 -13922
rect 6359 -13923 6432 -13922
rect 6715 -13923 6788 -13922
rect 6003 -13975 6013 -13923
rect 6065 -13975 6076 -13923
rect 6180 -13924 6253 -13923
rect 5577 -14082 5790 -14048
rect 5843 -14078 5877 -13975
rect 6022 -14080 6056 -13975
rect 6180 -13976 6190 -13924
rect 6242 -13976 6253 -13924
rect 6359 -13975 6369 -13923
rect 6421 -13975 6432 -13923
rect 6537 -13924 6610 -13923
rect 6200 -14080 6234 -13976
rect 6378 -14080 6412 -13975
rect 6537 -13976 6547 -13924
rect 6599 -13976 6610 -13924
rect 6715 -13975 6725 -13923
rect 6777 -13975 6788 -13923
rect 6892 -13923 6965 -13922
rect 6892 -13975 6902 -13923
rect 6954 -13975 6965 -13923
rect 6556 -14080 6590 -13976
rect 6734 -14081 6768 -13975
rect 6912 -14079 6946 -13975
rect 7103 -14082 7297 -14048
rect 5577 -14164 5611 -14082
rect 5756 -14545 5790 -14082
rect 7179 -14161 7213 -14082
rect 5736 -14546 5809 -14545
rect 5736 -14598 5746 -14546
rect 5798 -14598 5809 -14546
rect 5575 -15081 5789 -15047
rect 5843 -15075 5877 -14442
rect 5933 -14658 5967 -14388
rect 5914 -14659 5987 -14658
rect 5914 -14711 5924 -14659
rect 5976 -14711 5987 -14659
rect 6022 -15080 6056 -14447
rect 6111 -14545 6145 -14392
rect 6091 -14546 6164 -14545
rect 6091 -14598 6101 -14546
rect 6153 -14598 6164 -14546
rect 6200 -15079 6234 -14446
rect 6289 -14658 6323 -14387
rect 6269 -14659 6342 -14658
rect 6269 -14711 6279 -14659
rect 6331 -14711 6342 -14659
rect 6378 -15081 6412 -14448
rect 6468 -14545 6502 -14388
rect 6449 -14546 6522 -14545
rect 6449 -14598 6459 -14546
rect 6511 -14598 6522 -14546
rect 6557 -15081 6591 -14448
rect 6645 -14658 6679 -14387
rect 6823 -14545 6857 -14387
rect 6803 -14546 6876 -14545
rect 6803 -14598 6813 -14546
rect 6865 -14598 6876 -14546
rect 7000 -14658 7034 -14397
rect 6626 -14659 6699 -14658
rect 6626 -14711 6636 -14659
rect 6688 -14711 6699 -14659
rect 6981 -14659 7054 -14658
rect 6981 -14711 6991 -14659
rect 7043 -14711 7054 -14659
rect 7179 -14749 7213 -14387
rect 6822 -14783 7213 -14749
rect 5575 -15172 5609 -15081
rect 5755 -15539 5789 -15081
rect 5735 -15540 5808 -15539
rect 5735 -15592 5745 -15540
rect 5797 -15592 5808 -15540
rect 5390 -15654 5463 -15653
rect 5390 -15706 5400 -15654
rect 5452 -15706 5463 -15654
rect 5400 -16667 5453 -15706
rect 5737 -15751 5810 -15750
rect 5737 -15803 5747 -15751
rect 5799 -15803 5810 -15751
rect 5576 -16438 5610 -16353
rect 5756 -16438 5790 -15803
rect 5844 -16081 5878 -15448
rect 5933 -15652 5967 -15376
rect 5913 -15653 5986 -15652
rect 5913 -15705 5923 -15653
rect 5975 -15705 5986 -15653
rect 5911 -15949 5984 -15948
rect 5911 -16001 5921 -15949
rect 5973 -16001 5984 -15949
rect 5931 -16133 5965 -16001
rect 6022 -16082 6056 -15449
rect 6111 -15539 6145 -15380
rect 6091 -15540 6164 -15539
rect 6091 -15592 6101 -15540
rect 6153 -15592 6164 -15540
rect 6091 -15750 6164 -15749
rect 6091 -15802 6101 -15750
rect 6153 -15802 6164 -15750
rect 6112 -16136 6146 -15802
rect 6201 -16082 6235 -15449
rect 6289 -15652 6323 -15364
rect 6269 -15653 6342 -15652
rect 6269 -15705 6279 -15653
rect 6331 -15705 6342 -15653
rect 6269 -15949 6342 -15948
rect 6269 -16001 6279 -15949
rect 6331 -16001 6342 -15949
rect 6288 -16137 6322 -16001
rect 6379 -16081 6413 -15448
rect 6468 -15539 6502 -15375
rect 6448 -15540 6521 -15539
rect 6448 -15592 6458 -15540
rect 6510 -15592 6521 -15540
rect 6446 -15751 6519 -15750
rect 6446 -15803 6456 -15751
rect 6508 -15803 6519 -15751
rect 6467 -16137 6501 -15803
rect 6556 -16081 6590 -15448
rect 6645 -15652 6679 -15357
rect 6822 -15368 6856 -14783
rect 7357 -14824 7391 -13849
rect 7427 -13923 7500 -13922
rect 7427 -13975 7437 -13923
rect 7489 -13975 7500 -13923
rect 7446 -14081 7480 -13975
rect 6983 -14825 7056 -14824
rect 6983 -14877 6993 -14825
rect 7045 -14877 7056 -14825
rect 7337 -14825 7410 -14824
rect 7337 -14877 7347 -14825
rect 7399 -14877 7410 -14825
rect 6822 -15438 6857 -15368
rect 6748 -15472 6942 -15438
rect 6625 -15653 6698 -15652
rect 6625 -15705 6635 -15653
rect 6687 -15705 6698 -15653
rect 6703 -15752 6776 -15751
rect 6703 -15804 6713 -15752
rect 6765 -15804 6776 -15752
rect 6624 -15949 6697 -15948
rect 6624 -16001 6634 -15949
rect 6686 -16001 6697 -15949
rect 6734 -15956 6768 -15804
rect 6822 -15851 6856 -15472
rect 6803 -15852 6876 -15851
rect 6803 -15904 6813 -15852
rect 6865 -15904 6876 -15852
rect 7002 -15951 7036 -14877
rect 7070 -14924 7143 -14923
rect 7070 -14976 7080 -14924
rect 7132 -14976 7143 -14924
rect 7250 -14925 7323 -14924
rect 7090 -15080 7124 -14976
rect 7250 -14977 7260 -14925
rect 7312 -14977 7323 -14925
rect 7269 -15080 7303 -14977
rect 7357 -15182 7391 -14877
rect 7447 -14923 7481 -14448
rect 7429 -14924 7502 -14923
rect 7429 -14976 7439 -14924
rect 7491 -14976 7502 -14924
rect 7447 -15081 7481 -14976
rect 7535 -15163 7569 -13725
rect 7872 -13726 7882 -13674
rect 7934 -13726 7945 -13674
rect 8228 -13724 8238 -13672
rect 8290 -13724 8301 -13672
rect 7694 -13796 7767 -13795
rect 7694 -13848 7704 -13796
rect 7756 -13848 7767 -13796
rect 7605 -13923 7678 -13922
rect 7605 -13975 7615 -13923
rect 7667 -13975 7678 -13923
rect 7624 -14080 7658 -13975
rect 7713 -14130 7747 -13848
rect 7783 -13924 7856 -13923
rect 7783 -13976 7793 -13924
rect 7845 -13976 7856 -13924
rect 7802 -14081 7836 -13976
rect 7892 -14124 7926 -13726
rect 8051 -13797 8124 -13796
rect 8051 -13849 8061 -13797
rect 8113 -13849 8124 -13797
rect 7960 -13923 8033 -13922
rect 7960 -13975 7970 -13923
rect 8022 -13975 8033 -13923
rect 7980 -14081 8014 -13975
rect 8069 -14134 8103 -13849
rect 8138 -13923 8211 -13922
rect 8138 -13975 8148 -13923
rect 8200 -13975 8211 -13923
rect 8158 -14081 8192 -13975
rect 8248 -14137 8282 -13724
rect 8405 -13797 8478 -13796
rect 8405 -13849 8415 -13797
rect 8467 -13849 8478 -13797
rect 8316 -13923 8389 -13922
rect 8316 -13975 8326 -13923
rect 8378 -13975 8389 -13923
rect 8336 -14080 8370 -13975
rect 8425 -14142 8459 -13849
rect 8529 -14082 8723 -14048
rect 8603 -14165 8637 -14082
rect 8781 -14129 8815 -13609
rect 8851 -13923 8924 -13922
rect 8851 -13975 8861 -13923
rect 8913 -13975 8924 -13923
rect 8871 -14081 8905 -13975
rect 8960 -14131 8994 -13486
rect 9117 -13557 9190 -13556
rect 9117 -13609 9127 -13557
rect 9179 -13609 9190 -13557
rect 9028 -13923 9101 -13922
rect 9028 -13975 9038 -13923
rect 9090 -13975 9101 -13923
rect 9048 -14081 9082 -13975
rect 9137 -14134 9171 -13609
rect 9207 -13923 9280 -13922
rect 9207 -13975 9217 -13923
rect 9269 -13975 9280 -13923
rect 9227 -14081 9261 -13975
rect 9315 -14130 9349 -13486
rect 9473 -13557 9546 -13556
rect 9473 -13609 9483 -13557
rect 9535 -13609 9546 -13557
rect 9384 -13923 9457 -13922
rect 9384 -13975 9394 -13923
rect 9446 -13975 9457 -13923
rect 9404 -14081 9438 -13975
rect 9493 -14132 9527 -13609
rect 11432 -13673 11505 -13672
rect 11432 -13725 11442 -13673
rect 11494 -13725 11505 -13673
rect 11788 -13673 11861 -13672
rect 12499 -13673 12572 -13672
rect 11788 -13725 11798 -13673
rect 11850 -13725 11861 -13673
rect 12142 -13674 12215 -13673
rect 11254 -13797 11327 -13796
rect 11254 -13849 11264 -13797
rect 11316 -13849 11327 -13797
rect 10098 -13923 10171 -13922
rect 10630 -13923 10703 -13922
rect 9919 -13924 9992 -13923
rect 9919 -13976 9929 -13924
rect 9981 -13976 9992 -13924
rect 10098 -13975 10108 -13923
rect 10160 -13975 10171 -13923
rect 10274 -13924 10347 -13923
rect 9594 -14082 9788 -14048
rect 9938 -14081 9972 -13976
rect 10117 -14082 10151 -13975
rect 10274 -13976 10284 -13924
rect 10336 -13976 10347 -13924
rect 10452 -13924 10525 -13923
rect 10452 -13976 10462 -13924
rect 10514 -13976 10525 -13924
rect 10630 -13975 10640 -13923
rect 10692 -13975 10703 -13923
rect 10809 -13924 10882 -13923
rect 10294 -14082 10328 -13976
rect 10472 -14081 10506 -13976
rect 10650 -14081 10684 -13975
rect 10809 -13976 10819 -13924
rect 10871 -13976 10882 -13924
rect 10828 -14081 10862 -13976
rect 11018 -14082 11212 -14048
rect 9671 -14159 9705 -14082
rect 11095 -14158 11129 -14082
rect 7625 -15081 7659 -14448
rect 7694 -14826 7767 -14825
rect 7694 -14878 7704 -14826
rect 7756 -14878 7767 -14826
rect 7714 -15135 7748 -14878
rect 7802 -15081 7836 -14448
rect 8226 -14546 8299 -14545
rect 8226 -14598 8236 -14546
rect 8288 -14598 8299 -14546
rect 8050 -14822 8123 -14821
rect 8050 -14874 8060 -14822
rect 8112 -14874 8123 -14822
rect 7179 -15750 7213 -15384
rect 7159 -15751 7232 -15750
rect 7159 -15803 7169 -15751
rect 7221 -15803 7232 -15751
rect 7159 -15853 7232 -15852
rect 7159 -15905 7169 -15853
rect 7221 -15905 7232 -15853
rect 6984 -15952 7057 -15951
rect 6734 -15990 6858 -15956
rect 6644 -16145 6678 -16001
rect 6824 -16163 6858 -15990
rect 6984 -16004 6994 -15952
rect 7046 -16004 7057 -15952
rect 7002 -16273 7036 -16004
rect 7178 -16438 7212 -15905
rect 7447 -16080 7481 -15447
rect 7536 -15749 7570 -15382
rect 7516 -15750 7589 -15749
rect 7516 -15802 7526 -15750
rect 7578 -15802 7589 -15750
rect 7516 -15954 7589 -15953
rect 7516 -16006 7526 -15954
rect 7578 -16006 7589 -15954
rect 7535 -16147 7569 -16006
rect 7624 -16081 7658 -15448
rect 7803 -16081 7837 -15448
rect 7891 -15749 7925 -15369
rect 8069 -15438 8103 -14874
rect 8000 -15472 8194 -15438
rect 7872 -15750 7945 -15749
rect 7872 -15802 7882 -15750
rect 7934 -15802 7945 -15750
rect 8069 -15851 8103 -15472
rect 8050 -15852 8123 -15851
rect 8050 -15904 8060 -15852
rect 8112 -15904 8123 -15852
rect 8247 -15952 8281 -14598
rect 8336 -14923 8370 -14448
rect 8407 -14658 8480 -14657
rect 8407 -14710 8417 -14658
rect 8469 -14710 8480 -14658
rect 8317 -14924 8390 -14923
rect 8317 -14976 8327 -14924
rect 8379 -14976 8390 -14924
rect 8336 -15081 8370 -14976
rect 7871 -15953 7944 -15952
rect 7871 -16005 7881 -15953
rect 7933 -16005 7944 -15953
rect 8227 -15953 8300 -15952
rect 8227 -16005 8237 -15953
rect 8289 -16005 8300 -15953
rect 7891 -16167 7925 -16005
rect 8247 -16221 8281 -16005
rect 8336 -16080 8370 -15447
rect 5576 -16472 5790 -16438
rect 6557 -16544 6591 -16441
rect 6735 -16544 6769 -16440
rect 6538 -16545 6611 -16544
rect 6538 -16597 6548 -16545
rect 6600 -16597 6611 -16545
rect 6716 -16545 6789 -16544
rect 6912 -16545 6946 -16442
rect 7101 -16472 7295 -16438
rect 6716 -16597 6726 -16545
rect 6778 -16597 6789 -16545
rect 6893 -16546 6966 -16545
rect 6893 -16598 6903 -16546
rect 6955 -16598 6966 -16546
rect 5389 -16668 5462 -16667
rect 5389 -16720 5399 -16668
rect 5451 -16720 5462 -16668
rect 5021 -16783 5094 -16782
rect 5021 -16835 5031 -16783
rect 5083 -16835 5094 -16783
rect 7357 -16890 7391 -16342
rect 7713 -16890 7747 -16345
rect 7980 -16545 8014 -16453
rect 7960 -16546 8033 -16545
rect 7960 -16598 7970 -16546
rect 8022 -16598 8033 -16546
rect 8069 -16890 8103 -16382
rect 8158 -16544 8192 -16445
rect 8139 -16545 8212 -16544
rect 8139 -16597 8149 -16545
rect 8201 -16597 8212 -16545
rect 8426 -16890 8460 -14710
rect 8514 -14806 8548 -14438
rect 8585 -14546 8658 -14545
rect 8585 -14598 8595 -14546
rect 8647 -14598 8658 -14546
rect 8494 -14807 8567 -14806
rect 8494 -14859 8504 -14807
rect 8556 -14859 8567 -14807
rect 8514 -14871 8548 -14859
rect 8495 -14925 8568 -14924
rect 8495 -14977 8505 -14925
rect 8557 -14977 8568 -14925
rect 8514 -15080 8548 -14977
rect 8604 -15136 8638 -14598
rect 8762 -14659 8835 -14658
rect 8762 -14711 8772 -14659
rect 8824 -14711 8835 -14659
rect 8692 -14924 8726 -14923
rect 8673 -14925 8746 -14924
rect 8673 -14977 8683 -14925
rect 8735 -14977 8746 -14925
rect 8692 -15080 8726 -14977
rect 8781 -15148 8815 -14711
rect 8870 -15081 8904 -14448
rect 8940 -14547 9013 -14546
rect 8940 -14599 8950 -14547
rect 9002 -14599 9013 -14547
rect 8960 -15139 8994 -14599
rect 9048 -15081 9082 -14448
rect 9117 -14660 9190 -14659
rect 9117 -14712 9127 -14660
rect 9179 -14712 9190 -14660
rect 9137 -15140 9171 -14712
rect 9226 -15081 9260 -14448
rect 9294 -14546 9367 -14545
rect 9294 -14598 9304 -14546
rect 9356 -14598 9367 -14546
rect 9314 -15144 9348 -14598
rect 9404 -15081 9438 -14448
rect 9651 -14546 9724 -14545
rect 9651 -14598 9661 -14546
rect 9713 -14598 9724 -14546
rect 9473 -14659 9546 -14658
rect 9473 -14711 9483 -14659
rect 9535 -14711 9546 -14659
rect 9493 -15135 9527 -14711
rect 9562 -14924 9635 -14923
rect 9562 -14976 9572 -14924
rect 9624 -14976 9635 -14924
rect 9582 -15077 9616 -14976
rect 9671 -15139 9705 -14598
rect 9763 -14806 9797 -14453
rect 9848 -14659 9882 -14383
rect 9827 -14660 9900 -14659
rect 9827 -14712 9837 -14660
rect 9889 -14712 9900 -14660
rect 9743 -14807 9816 -14806
rect 9743 -14859 9753 -14807
rect 9805 -14859 9816 -14807
rect 9763 -14871 9797 -14859
rect 9740 -14924 9813 -14923
rect 9740 -14976 9750 -14924
rect 9802 -14976 9813 -14924
rect 9760 -15078 9794 -14976
rect 9848 -15200 9882 -14712
rect 9939 -14923 9973 -14449
rect 10026 -14545 10060 -14384
rect 10006 -14546 10079 -14545
rect 10006 -14598 10016 -14546
rect 10068 -14598 10079 -14546
rect 9919 -14924 9992 -14923
rect 9919 -14976 9929 -14924
rect 9981 -14976 9992 -14924
rect 9939 -15082 9973 -14976
rect 10026 -15216 10060 -14598
rect 10205 -14658 10239 -14385
rect 10383 -14546 10417 -14385
rect 10363 -14547 10436 -14546
rect 10363 -14599 10373 -14547
rect 10425 -14599 10436 -14547
rect 10186 -14659 10259 -14658
rect 10186 -14711 10196 -14659
rect 10248 -14711 10259 -14659
rect 10185 -14823 10258 -14822
rect 10185 -14875 10195 -14823
rect 10247 -14875 10258 -14823
rect 10205 -15438 10239 -14875
rect 10472 -15081 10506 -14448
rect 10560 -14658 10594 -14383
rect 10540 -14659 10613 -14658
rect 10540 -14711 10550 -14659
rect 10602 -14711 10613 -14659
rect 10542 -14816 10615 -14815
rect 10542 -14868 10552 -14816
rect 10604 -14868 10615 -14816
rect 10561 -15136 10595 -14868
rect 10650 -15081 10684 -14448
rect 10738 -14545 10772 -14383
rect 10719 -14546 10792 -14545
rect 10719 -14598 10729 -14546
rect 10781 -14598 10792 -14546
rect 10828 -14923 10862 -14448
rect 10917 -14658 10951 -14387
rect 11096 -14658 11130 -14334
rect 10898 -14659 10971 -14658
rect 10898 -14711 10908 -14659
rect 10960 -14711 10971 -14659
rect 11077 -14659 11150 -14658
rect 11077 -14711 11087 -14659
rect 11139 -14711 11150 -14659
rect 10898 -14814 10971 -14813
rect 10898 -14866 10908 -14814
rect 10960 -14866 10971 -14814
rect 11273 -14815 11307 -13849
rect 11343 -13923 11416 -13922
rect 11343 -13975 11353 -13923
rect 11405 -13975 11416 -13923
rect 11362 -14081 11396 -13975
rect 11452 -14133 11486 -13725
rect 11610 -13798 11683 -13797
rect 11610 -13850 11620 -13798
rect 11672 -13850 11683 -13798
rect 11520 -13923 11593 -13922
rect 11520 -13975 11530 -13923
rect 11582 -13975 11593 -13923
rect 11540 -14080 11574 -13975
rect 11630 -14135 11664 -13850
rect 11699 -13923 11772 -13922
rect 11699 -13975 11709 -13923
rect 11761 -13975 11772 -13923
rect 11719 -14081 11753 -13975
rect 11807 -14133 11841 -13725
rect 12142 -13726 12152 -13674
rect 12204 -13726 12215 -13674
rect 12499 -13725 12509 -13673
rect 12561 -13725 12572 -13673
rect 11967 -13797 12040 -13796
rect 11967 -13849 11977 -13797
rect 12029 -13849 12040 -13797
rect 11876 -13924 11949 -13923
rect 11876 -13976 11886 -13924
rect 11938 -13976 11949 -13924
rect 11895 -14080 11929 -13976
rect 11986 -14131 12020 -13849
rect 12054 -13923 12127 -13922
rect 12054 -13975 12064 -13923
rect 12116 -13975 12127 -13923
rect 12073 -14082 12107 -13975
rect 12162 -14137 12196 -13726
rect 12324 -13797 12397 -13796
rect 12324 -13849 12334 -13797
rect 12386 -13849 12397 -13797
rect 12232 -13924 12305 -13923
rect 12232 -13976 12242 -13924
rect 12294 -13976 12305 -13924
rect 12252 -14081 12286 -13976
rect 12342 -14133 12376 -13849
rect 12410 -13923 12483 -13922
rect 12410 -13975 12420 -13923
rect 12472 -13975 12483 -13923
rect 12430 -14081 12464 -13975
rect 12519 -14048 12553 -13725
rect 12519 -14082 12731 -14048
rect 12519 -14134 12553 -14082
rect 12697 -14154 12731 -14082
rect 11430 -14657 11503 -14656
rect 11430 -14709 11440 -14657
rect 11492 -14709 11503 -14657
rect 11254 -14816 11327 -14815
rect 10809 -14924 10882 -14923
rect 10809 -14976 10819 -14924
rect 10871 -14976 10882 -14924
rect 10828 -15081 10862 -14976
rect 8583 -15853 8656 -15852
rect 8583 -15905 8593 -15853
rect 8645 -15905 8656 -15853
rect 8603 -16438 8637 -15905
rect 8870 -16080 8904 -15447
rect 9049 -16081 9083 -15448
rect 9226 -16080 9260 -15447
rect 9404 -16080 9438 -15447
rect 9653 -15853 9726 -15852
rect 9653 -15905 9663 -15853
rect 9715 -15905 9726 -15853
rect 8519 -16472 8713 -16438
rect 8781 -16666 8815 -16386
rect 8761 -16667 8834 -16666
rect 8761 -16719 8771 -16667
rect 8823 -16719 8834 -16667
rect 8960 -16782 8994 -16389
rect 9138 -16666 9172 -16383
rect 9118 -16667 9191 -16666
rect 9118 -16719 9128 -16667
rect 9180 -16719 9191 -16667
rect 9315 -16782 9349 -16393
rect 9493 -16666 9527 -16380
rect 9672 -16438 9706 -15905
rect 9939 -16081 9973 -15448
rect 10122 -15472 10316 -15438
rect 10205 -15852 10239 -15472
rect 10383 -15751 10417 -15349
rect 10363 -15752 10436 -15751
rect 10363 -15804 10373 -15752
rect 10425 -15804 10436 -15752
rect 10184 -15853 10257 -15852
rect 10184 -15905 10194 -15853
rect 10246 -15905 10257 -15853
rect 10472 -16080 10506 -15447
rect 10650 -16080 10684 -15447
rect 10739 -15750 10773 -15359
rect 10720 -15751 10793 -15750
rect 10720 -15803 10730 -15751
rect 10782 -15803 10793 -15751
rect 10739 -16238 10773 -15803
rect 10828 -16080 10862 -15447
rect 10916 -16215 10950 -14866
rect 11254 -14868 11264 -14816
rect 11316 -14868 11327 -14816
rect 10986 -14924 11059 -14923
rect 10986 -14976 10996 -14924
rect 11048 -14976 11059 -14924
rect 11165 -14924 11238 -14923
rect 11165 -14976 11175 -14924
rect 11227 -14976 11238 -14924
rect 11006 -15061 11040 -14976
rect 11184 -15063 11218 -14976
rect 11273 -15189 11307 -14868
rect 11095 -15750 11129 -15348
rect 11451 -15438 11485 -14709
rect 11717 -15078 11751 -14439
rect 11897 -15079 11931 -14440
rect 12075 -15079 12109 -14440
rect 12253 -15081 12287 -14442
rect 12430 -15081 12464 -14442
rect 12520 -15083 12730 -15049
rect 11390 -15472 11584 -15438
rect 11076 -15751 11149 -15750
rect 11076 -15803 11086 -15751
rect 11138 -15803 11149 -15751
rect 11451 -15841 11485 -15472
rect 11629 -15652 11663 -15392
rect 11609 -15653 11682 -15652
rect 11609 -15705 11619 -15653
rect 11671 -15705 11682 -15653
rect 11629 -15706 11663 -15705
rect 11430 -15842 11503 -15841
rect 11074 -15853 11147 -15852
rect 11074 -15905 11084 -15853
rect 11136 -15905 11147 -15853
rect 11430 -15894 11440 -15842
rect 11492 -15894 11503 -15842
rect 11451 -15902 11485 -15894
rect 9595 -16472 9789 -16438
rect 9474 -16667 9547 -16666
rect 9474 -16719 9484 -16667
rect 9536 -16719 9547 -16667
rect 8940 -16783 9013 -16782
rect 8940 -16835 8950 -16783
rect 9002 -16835 9013 -16783
rect 9295 -16783 9368 -16782
rect 9295 -16835 9305 -16783
rect 9357 -16835 9368 -16783
rect 7337 -16891 7410 -16890
rect 7337 -16943 7347 -16891
rect 7399 -16943 7410 -16891
rect 7694 -16891 7767 -16890
rect 7694 -16943 7704 -16891
rect 7756 -16943 7767 -16891
rect 8050 -16891 8123 -16890
rect 8050 -16943 8060 -16891
rect 8112 -16943 8123 -16891
rect 8406 -16891 8479 -16890
rect 8406 -16943 8416 -16891
rect 8468 -16943 8479 -16891
rect 9672 -17251 9706 -16472
rect 9848 -16666 9882 -16349
rect 9938 -16544 9972 -16458
rect 9919 -16545 9992 -16544
rect 9919 -16597 9929 -16545
rect 9981 -16597 9992 -16545
rect 9828 -16667 9901 -16666
rect 9828 -16719 9838 -16667
rect 9890 -16719 9901 -16667
rect 10028 -16781 10062 -16383
rect 10117 -16545 10151 -16456
rect 10097 -16546 10170 -16545
rect 10097 -16598 10107 -16546
rect 10159 -16598 10170 -16546
rect 10205 -16665 10239 -16334
rect 10296 -16545 10330 -16458
rect 10277 -16546 10350 -16545
rect 10277 -16598 10287 -16546
rect 10339 -16598 10350 -16546
rect 10185 -16666 10258 -16665
rect 10185 -16718 10195 -16666
rect 10247 -16718 10258 -16666
rect 10383 -16781 10417 -16377
rect 10561 -16665 10595 -16352
rect 10540 -16666 10613 -16665
rect 10540 -16718 10550 -16666
rect 10602 -16718 10613 -16666
rect 10739 -16779 10773 -16359
rect 10917 -16665 10951 -16377
rect 11094 -16437 11128 -15905
rect 11431 -15953 11504 -15952
rect 11431 -16005 11441 -15953
rect 11493 -16005 11504 -15953
rect 11451 -16138 11485 -16005
rect 11718 -16081 11752 -15448
rect 11808 -15540 11842 -15394
rect 11788 -15541 11861 -15540
rect 11788 -15593 11798 -15541
rect 11850 -15593 11861 -15541
rect 11787 -15953 11860 -15952
rect 11787 -16005 11797 -15953
rect 11849 -16005 11860 -15953
rect 11806 -16136 11840 -16005
rect 11897 -16081 11931 -15448
rect 11985 -15652 12019 -15387
rect 11965 -15653 12038 -15652
rect 11965 -15705 11975 -15653
rect 12027 -15705 12038 -15653
rect 12074 -16080 12108 -15447
rect 12165 -15539 12199 -15372
rect 12145 -15540 12218 -15539
rect 12145 -15592 12155 -15540
rect 12207 -15592 12218 -15540
rect 12144 -15953 12217 -15952
rect 12144 -16005 12154 -15953
rect 12206 -16005 12217 -15953
rect 12163 -16136 12197 -16005
rect 12252 -16081 12286 -15448
rect 12342 -15652 12376 -15386
rect 12322 -15653 12395 -15652
rect 12322 -15705 12332 -15653
rect 12384 -15705 12395 -15653
rect 12431 -16081 12465 -15448
rect 12520 -15539 12554 -15083
rect 12696 -15154 12730 -15083
rect 12501 -15540 12574 -15539
rect 12501 -15592 12511 -15540
rect 12563 -15592 12574 -15540
rect 12501 -15953 12574 -15952
rect 12501 -16005 12511 -15953
rect 12563 -16005 12574 -15953
rect 11019 -16471 11213 -16437
rect 10897 -16666 10970 -16665
rect 10897 -16718 10907 -16666
rect 10959 -16718 10970 -16666
rect 10721 -16780 10794 -16779
rect 10007 -16782 10080 -16781
rect 10007 -16834 10017 -16782
rect 10069 -16834 10080 -16782
rect 10364 -16782 10437 -16781
rect 10364 -16834 10374 -16782
rect 10426 -16834 10437 -16782
rect 10721 -16832 10731 -16780
rect 10783 -16832 10794 -16780
rect 11273 -16890 11307 -16340
rect 11362 -16545 11396 -16455
rect 11342 -16546 11415 -16545
rect 11540 -16546 11574 -16453
rect 11342 -16598 11352 -16546
rect 11404 -16598 11415 -16546
rect 11520 -16547 11593 -16546
rect 11520 -16599 11530 -16547
rect 11582 -16599 11593 -16547
rect 11630 -16890 11664 -16362
rect 11718 -16545 11752 -16457
rect 11699 -16546 11772 -16545
rect 11699 -16598 11709 -16546
rect 11761 -16598 11772 -16546
rect 11985 -16889 12019 -16353
rect 12340 -16889 12374 -16380
rect 12520 -16440 12554 -16005
rect 12698 -16440 12732 -16356
rect 12520 -16474 12732 -16440
rect 11965 -16890 12038 -16889
rect 11253 -16891 11326 -16890
rect 11253 -16943 11263 -16891
rect 11315 -16943 11326 -16891
rect 11610 -16891 11683 -16890
rect 11610 -16943 11620 -16891
rect 11672 -16943 11683 -16891
rect 11965 -16942 11975 -16890
rect 12027 -16942 12038 -16890
rect 12321 -16890 12394 -16889
rect 12321 -16942 12331 -16890
rect 12383 -16942 12394 -16890
rect 13022 -17251 13075 -11726
rect 18337 -13421 18412 -6747
rect 18327 -13433 18422 -13421
rect 18327 -13485 18348 -13433
rect 18400 -13485 18422 -13433
rect 18327 -13496 18422 -13485
rect 18337 -13506 18412 -13496
rect -7605 -17492 13720 -17251
rect -7605 -17526 -7319 -17492
rect -7285 -17526 -7247 -17492
rect -7213 -17526 -7175 -17492
rect -7141 -17526 -7103 -17492
rect -7069 -17526 -7031 -17492
rect -6997 -17526 -6959 -17492
rect -6925 -17526 -6887 -17492
rect -6853 -17526 -6815 -17492
rect -6781 -17526 -6743 -17492
rect -6709 -17526 -6671 -17492
rect -6637 -17526 -6599 -17492
rect -6565 -17526 -6527 -17492
rect -6493 -17526 -6455 -17492
rect -6421 -17526 -6383 -17492
rect -6349 -17526 -6311 -17492
rect -6277 -17526 -6239 -17492
rect -6205 -17526 -6167 -17492
rect -6133 -17526 -6095 -17492
rect -6061 -17526 -6023 -17492
rect -5989 -17526 -5951 -17492
rect -5917 -17526 -5879 -17492
rect -5845 -17526 -5807 -17492
rect -5773 -17526 -5735 -17492
rect -5701 -17526 -5663 -17492
rect -5629 -17526 -5591 -17492
rect -5557 -17526 -5519 -17492
rect -5485 -17526 -5447 -17492
rect -5413 -17526 -5375 -17492
rect -5341 -17526 -5303 -17492
rect -5269 -17526 -5231 -17492
rect -5197 -17526 -5159 -17492
rect -5125 -17526 -5087 -17492
rect -5053 -17526 -5015 -17492
rect -4981 -17526 -4943 -17492
rect -4909 -17526 -4871 -17492
rect -4837 -17526 -4799 -17492
rect -4765 -17526 -4727 -17492
rect -4693 -17526 -4655 -17492
rect -4621 -17526 -4583 -17492
rect -4549 -17526 -4511 -17492
rect -4477 -17526 -4439 -17492
rect -4405 -17526 -4367 -17492
rect -4333 -17526 -4295 -17492
rect -4261 -17526 -4223 -17492
rect -4189 -17526 -4151 -17492
rect -4117 -17526 -4079 -17492
rect -4045 -17526 -4007 -17492
rect -3973 -17526 -3935 -17492
rect -3901 -17526 -3863 -17492
rect -3829 -17526 -3791 -17492
rect -3757 -17526 -3719 -17492
rect -3685 -17526 -3647 -17492
rect -3613 -17526 -3575 -17492
rect -3541 -17526 -3503 -17492
rect -3469 -17526 -3431 -17492
rect -3397 -17526 -3359 -17492
rect -3325 -17526 -3287 -17492
rect -3253 -17526 -3215 -17492
rect -3181 -17526 -3143 -17492
rect -3109 -17526 -3071 -17492
rect -3037 -17526 -2999 -17492
rect -2965 -17526 -2927 -17492
rect -2893 -17526 -2855 -17492
rect -2821 -17526 -2783 -17492
rect -2749 -17526 -2711 -17492
rect -2677 -17526 -2639 -17492
rect -2605 -17526 -2567 -17492
rect -2533 -17526 -2495 -17492
rect -2461 -17526 -2423 -17492
rect -2389 -17526 -2351 -17492
rect -2317 -17526 -2279 -17492
rect -2245 -17526 -2207 -17492
rect -2173 -17526 -2135 -17492
rect -2101 -17526 -2063 -17492
rect -2029 -17526 -1991 -17492
rect -1957 -17526 -1919 -17492
rect -1885 -17526 -1847 -17492
rect -1813 -17526 -1775 -17492
rect -1741 -17526 -1703 -17492
rect -1669 -17526 -1631 -17492
rect -1597 -17526 -1559 -17492
rect -1525 -17526 -1487 -17492
rect -1453 -17526 -1415 -17492
rect -1381 -17526 -1343 -17492
rect -1309 -17526 -1271 -17492
rect -1237 -17526 -1199 -17492
rect -1165 -17526 -1127 -17492
rect -1093 -17526 -1055 -17492
rect -1021 -17526 -983 -17492
rect -949 -17526 -911 -17492
rect -877 -17526 -839 -17492
rect -805 -17526 -767 -17492
rect -733 -17526 -695 -17492
rect -661 -17526 -623 -17492
rect -589 -17526 -551 -17492
rect -517 -17526 -479 -17492
rect -445 -17526 -407 -17492
rect -373 -17526 -335 -17492
rect -301 -17526 -263 -17492
rect -229 -17526 -191 -17492
rect -157 -17526 -119 -17492
rect -85 -17526 -47 -17492
rect -13 -17526 25 -17492
rect 59 -17526 97 -17492
rect 131 -17526 169 -17492
rect 203 -17526 241 -17492
rect 275 -17526 313 -17492
rect 347 -17526 385 -17492
rect 419 -17526 457 -17492
rect 491 -17526 529 -17492
rect 563 -17526 601 -17492
rect 635 -17526 673 -17492
rect 707 -17526 745 -17492
rect 779 -17526 817 -17492
rect 851 -17526 889 -17492
rect 923 -17526 961 -17492
rect 995 -17526 1033 -17492
rect 1067 -17526 1105 -17492
rect 1139 -17526 1177 -17492
rect 1211 -17526 1249 -17492
rect 1283 -17526 1321 -17492
rect 1355 -17526 1393 -17492
rect 1427 -17526 1465 -17492
rect 1499 -17526 1537 -17492
rect 1571 -17526 1609 -17492
rect 1643 -17526 1681 -17492
rect 1715 -17526 1753 -17492
rect 1787 -17526 1825 -17492
rect 1859 -17526 1897 -17492
rect 1931 -17526 1969 -17492
rect 2003 -17526 2041 -17492
rect 2075 -17526 2113 -17492
rect 2147 -17526 2185 -17492
rect 2219 -17526 2257 -17492
rect 2291 -17526 2329 -17492
rect 2363 -17526 2401 -17492
rect 2435 -17526 2473 -17492
rect 2507 -17526 2545 -17492
rect 2579 -17526 2617 -17492
rect 2651 -17526 2689 -17492
rect 2723 -17526 2761 -17492
rect 2795 -17526 2833 -17492
rect 2867 -17526 2905 -17492
rect 2939 -17526 2977 -17492
rect 3011 -17526 3049 -17492
rect 3083 -17526 3121 -17492
rect 3155 -17526 3193 -17492
rect 3227 -17526 3265 -17492
rect 3299 -17526 3337 -17492
rect 3371 -17526 3409 -17492
rect 3443 -17526 3481 -17492
rect 3515 -17526 3553 -17492
rect 3587 -17526 3625 -17492
rect 3659 -17526 3697 -17492
rect 3731 -17526 3769 -17492
rect 3803 -17526 3841 -17492
rect 3875 -17526 3913 -17492
rect 3947 -17526 3985 -17492
rect 4019 -17526 4057 -17492
rect 4091 -17526 4129 -17492
rect 4163 -17526 4201 -17492
rect 4235 -17526 4273 -17492
rect 4307 -17526 4345 -17492
rect 4379 -17526 4417 -17492
rect 4451 -17526 4489 -17492
rect 4523 -17526 4561 -17492
rect 4595 -17526 4633 -17492
rect 4667 -17526 4705 -17492
rect 4739 -17526 4777 -17492
rect 4811 -17526 4849 -17492
rect 4883 -17526 4921 -17492
rect 4955 -17526 4993 -17492
rect 5027 -17526 5065 -17492
rect 5099 -17526 5137 -17492
rect 5171 -17526 5209 -17492
rect 5243 -17526 5281 -17492
rect 5315 -17526 5353 -17492
rect 5387 -17526 5425 -17492
rect 5459 -17526 5497 -17492
rect 5531 -17526 5569 -17492
rect 5603 -17526 5641 -17492
rect 5675 -17526 5713 -17492
rect 5747 -17526 5785 -17492
rect 5819 -17526 5857 -17492
rect 5891 -17526 5929 -17492
rect 5963 -17526 6001 -17492
rect 6035 -17526 6073 -17492
rect 6107 -17526 6145 -17492
rect 6179 -17526 6217 -17492
rect 6251 -17526 6289 -17492
rect 6323 -17526 6361 -17492
rect 6395 -17526 6433 -17492
rect 6467 -17526 6505 -17492
rect 6539 -17526 6577 -17492
rect 6611 -17526 6649 -17492
rect 6683 -17526 6721 -17492
rect 6755 -17526 6793 -17492
rect 6827 -17526 6865 -17492
rect 6899 -17526 6937 -17492
rect 6971 -17526 7009 -17492
rect 7043 -17526 7081 -17492
rect 7115 -17526 7153 -17492
rect 7187 -17526 7225 -17492
rect 7259 -17526 7297 -17492
rect 7331 -17526 7369 -17492
rect 7403 -17526 7441 -17492
rect 7475 -17526 7513 -17492
rect 7547 -17526 7585 -17492
rect 7619 -17526 7657 -17492
rect 7691 -17526 7729 -17492
rect 7763 -17526 7801 -17492
rect 7835 -17526 7873 -17492
rect 7907 -17526 7945 -17492
rect 7979 -17526 8017 -17492
rect 8051 -17526 8089 -17492
rect 8123 -17526 8161 -17492
rect 8195 -17526 8233 -17492
rect 8267 -17526 8305 -17492
rect 8339 -17526 8377 -17492
rect 8411 -17526 8449 -17492
rect 8483 -17526 8521 -17492
rect 8555 -17526 8593 -17492
rect 8627 -17526 8665 -17492
rect 8699 -17526 8737 -17492
rect 8771 -17526 8809 -17492
rect 8843 -17526 8881 -17492
rect 8915 -17526 8953 -17492
rect 8987 -17526 9025 -17492
rect 9059 -17526 9097 -17492
rect 9131 -17526 9169 -17492
rect 9203 -17526 9241 -17492
rect 9275 -17526 9313 -17492
rect 9347 -17526 9385 -17492
rect 9419 -17526 9457 -17492
rect 9491 -17526 9529 -17492
rect 9563 -17526 9601 -17492
rect 9635 -17526 9673 -17492
rect 9707 -17526 9745 -17492
rect 9779 -17526 9817 -17492
rect 9851 -17526 9889 -17492
rect 9923 -17526 9961 -17492
rect 9995 -17526 10033 -17492
rect 10067 -17526 10105 -17492
rect 10139 -17526 10177 -17492
rect 10211 -17526 10249 -17492
rect 10283 -17526 10321 -17492
rect 10355 -17526 10393 -17492
rect 10427 -17526 10465 -17492
rect 10499 -17526 10537 -17492
rect 10571 -17526 10609 -17492
rect 10643 -17526 10681 -17492
rect 10715 -17526 10753 -17492
rect 10787 -17526 10825 -17492
rect 10859 -17526 10897 -17492
rect 10931 -17526 10969 -17492
rect 11003 -17526 11041 -17492
rect 11075 -17526 11113 -17492
rect 11147 -17526 11185 -17492
rect 11219 -17526 11257 -17492
rect 11291 -17526 11329 -17492
rect 11363 -17526 11401 -17492
rect 11435 -17526 11473 -17492
rect 11507 -17526 11545 -17492
rect 11579 -17526 11617 -17492
rect 11651 -17526 11689 -17492
rect 11723 -17526 11761 -17492
rect 11795 -17526 11833 -17492
rect 11867 -17526 11905 -17492
rect 11939 -17526 11977 -17492
rect 12011 -17526 12049 -17492
rect 12083 -17526 12121 -17492
rect 12155 -17526 12193 -17492
rect 12227 -17526 12265 -17492
rect 12299 -17526 12337 -17492
rect 12371 -17526 12409 -17492
rect 12443 -17526 12481 -17492
rect 12515 -17526 12553 -17492
rect 12587 -17526 12625 -17492
rect 12659 -17526 12697 -17492
rect 12731 -17526 12769 -17492
rect 12803 -17526 12841 -17492
rect 12875 -17526 12913 -17492
rect 12947 -17526 12985 -17492
rect 13019 -17526 13057 -17492
rect 13091 -17526 13129 -17492
rect 13163 -17526 13201 -17492
rect 13235 -17526 13273 -17492
rect 13307 -17526 13345 -17492
rect 13379 -17526 13720 -17492
rect -7605 -17527 13720 -17526
rect -7605 -17587 13719 -17527
<< via1 >>
rect -5867 -1963 -5815 -1911
rect -5689 -1963 -5637 -1911
rect -5510 -1963 -5458 -1911
rect -5333 -1963 -5281 -1911
rect -5155 -1963 -5103 -1911
rect -4976 -1963 -4924 -1911
rect -4799 -1963 -4747 -1911
rect -4621 -1963 -4569 -1911
rect -4443 -1963 -4391 -1911
rect -4265 -1963 -4213 -1911
rect -4086 -1963 -4034 -1911
rect -3909 -1963 -3857 -1911
rect -1109 -1963 -1057 -1911
rect -6498 -2582 -6446 -2530
rect -6625 -3454 -6573 -3402
rect -6044 -2833 -5992 -2781
rect -6134 -3454 -6082 -3402
rect -6498 -3693 -6446 -3641
rect -6498 -4324 -6446 -4272
rect -6134 -4443 -6082 -4391
rect -6498 -5194 -6446 -5142
rect -6625 -5375 -6573 -5323
rect -6134 -5285 -6082 -5233
rect -5777 -2583 -5725 -2531
rect -5866 -2833 -5814 -2781
rect -5777 -3569 -5725 -3517
rect -5778 -4324 -5726 -4272
rect -5777 -5468 -5725 -5416
rect -5421 -2721 -5369 -2669
rect -5422 -3693 -5370 -3641
rect -5422 -4559 -5370 -4507
rect -5422 -5194 -5370 -5142
rect -5066 -2583 -5014 -2531
rect -5066 -3454 -5014 -3402
rect -5066 -4443 -5014 -4391
rect -5066 -5286 -5014 -5234
rect -4710 -2721 -4658 -2669
rect -4710 -3454 -4658 -3402
rect -4709 -4443 -4657 -4391
rect -4710 -5375 -4658 -5323
rect -4354 -2583 -4302 -2531
rect -4353 -3693 -4301 -3641
rect -4353 -4559 -4301 -4507
rect -4353 -5194 -4301 -5142
rect -3998 -2721 -3946 -2669
rect -1109 -2478 -1057 -2426
rect -752 -2478 -700 -2426
rect -3908 -2833 -3856 -2781
rect -3998 -3569 -3946 -3517
rect -3998 -4324 -3946 -4272
rect -3997 -5468 -3945 -5416
rect -2624 -2611 -2572 -2559
rect -1285 -2611 -1233 -2559
rect -3298 -2721 -3246 -2669
rect -3731 -2833 -3679 -2781
rect -3642 -3454 -3590 -3402
rect -3131 -3454 -3079 -3402
rect -3298 -3569 -3246 -3517
rect -3642 -4443 -3590 -4391
rect -3298 -4559 -3246 -4507
rect -3642 -5372 -3590 -5320
rect -3130 -5286 -3078 -5234
rect -1197 -2718 -1145 -2666
rect -930 -2611 -878 -2559
rect -1019 -2718 -967 -2666
rect -841 -2718 -789 -2666
rect -129 -2718 -77 -2666
rect 50 -2718 102 -2666
rect 227 -2718 279 -2666
rect 5337 -2258 5389 -2206
rect 6686 -2257 6738 -2205
rect 1919 -2479 1971 -2427
rect 2275 -2479 2327 -2427
rect 940 -2718 992 -2666
rect 1117 -2718 1169 -2666
rect 1295 -2718 1347 -2666
rect -1641 -3506 -1589 -3454
rect -2004 -4465 -1952 -4413
rect -2624 -5377 -2572 -5325
rect -3298 -5469 -3246 -5417
rect -5956 -6069 -5904 -6017
rect -5601 -6069 -5549 -6017
rect -5778 -6184 -5726 -6132
rect -5244 -6069 -5192 -6017
rect -5065 -6184 -5013 -6132
rect -6498 -6301 -6446 -6249
rect -5421 -6301 -5369 -6249
rect -4888 -6069 -4836 -6017
rect -4710 -6301 -4658 -6249
rect -4532 -6069 -4480 -6017
rect -4175 -6069 -4123 -6017
rect -4354 -6184 -4302 -6132
rect -3820 -6069 -3768 -6017
rect -2624 -6060 -2572 -6008
rect -3298 -6184 -3246 -6132
rect -3998 -6300 -3946 -6248
rect -4786 -6431 -4734 -6379
rect -1876 -5285 -1824 -5233
rect -1286 -3624 -1234 -3572
rect -1108 -3509 -1056 -3457
rect -929 -3624 -877 -3572
rect -484 -3354 -432 -3302
rect -750 -3509 -698 -3457
rect -396 -3509 -344 -3457
rect -573 -3624 -521 -3572
rect -217 -3624 -165 -3572
rect 583 -3354 635 -3302
rect -39 -3509 13 -3457
rect 317 -3509 369 -3457
rect 850 -3509 902 -3457
rect 1206 -3509 1258 -3457
rect 2097 -2607 2149 -2555
rect 2007 -2718 2059 -2666
rect 2186 -2718 2238 -2666
rect 3193 -2480 3245 -2428
rect 2453 -2607 2505 -2555
rect 2363 -2718 2415 -2666
rect 1654 -3354 1706 -3302
rect 1562 -3509 1614 -3457
rect 1919 -3509 1971 -3457
rect 1384 -3617 1436 -3565
rect 1741 -3617 1793 -3565
rect 2097 -3617 2149 -3565
rect 2275 -3509 2327 -3457
rect 2451 -3617 2503 -3565
rect -841 -4245 -789 -4193
rect -662 -4245 -610 -4193
rect -483 -4245 -431 -4193
rect -306 -4245 -254 -4193
rect -1287 -5150 -1235 -5098
rect -1642 -5335 -1590 -5283
rect -1105 -5266 -1053 -5214
rect -929 -5150 -877 -5098
rect -572 -5150 -520 -5098
rect -218 -5150 -166 -5098
rect -751 -5266 -699 -5214
rect -396 -5266 -344 -5214
rect -1876 -6417 -1824 -6365
rect -1282 -6417 -1230 -6365
rect -928 -6417 -876 -6365
rect -1110 -6532 -1058 -6480
rect -752 -6532 -700 -6480
rect 407 -4245 459 -4193
rect 317 -4357 369 -4305
rect 583 -4245 635 -4193
rect 495 -4465 547 -4413
rect 761 -4245 813 -4193
rect 673 -4357 725 -4305
rect 850 -4465 902 -4413
rect 1474 -4245 1526 -4193
rect 1652 -4245 1704 -4193
rect 1830 -4245 1882 -4193
rect 2008 -4245 2060 -4193
rect 2542 -4323 2594 -4271
rect 2750 -4503 2802 -4451
rect -41 -5266 11 -5214
rect 316 -5266 368 -5214
rect -128 -5433 -76 -5381
rect 50 -5433 102 -5381
rect 228 -5433 280 -5381
rect 850 -5266 902 -5214
rect 1207 -5266 1259 -5214
rect 940 -5434 992 -5382
rect 1119 -5433 1171 -5381
rect 1385 -5146 1437 -5094
rect 1296 -5433 1348 -5381
rect 227 -6303 279 -6251
rect 1740 -5146 1792 -5094
rect 1563 -5266 1615 -5214
rect 1917 -5266 1969 -5214
rect 2096 -5146 2148 -5094
rect 2274 -5266 2326 -5214
rect 2453 -5146 2505 -5094
rect 942 -6303 994 -6251
rect 2096 -6060 2148 -6008
rect 2452 -6060 2504 -6008
rect 1918 -6177 1970 -6125
rect 2275 -6177 2327 -6125
rect 3194 -4857 3246 -4805
rect 4771 -4857 4823 -4805
rect 2879 -6417 2931 -6365
rect 5037 -5059 5089 -5007
rect 4905 -5265 4957 -5213
rect -753 -6651 -701 -6599
rect 4772 -6650 4824 -6598
rect -2003 -6767 -1951 -6715
rect 6228 -3509 6280 -3457
rect 5620 -5265 5672 -5213
rect 5337 -5580 5389 -5528
rect 17837 -6579 17889 -6527
rect 4770 -6944 4822 -6892
rect 4906 -6942 4958 -6890
rect 5038 -6940 5090 -6888
rect -3873 -7743 -3821 -7691
rect -3731 -7837 -3679 -7785
rect -3541 -7840 -3489 -7788
rect -5502 -12324 -5450 -12272
rect -6077 -12565 -6025 -12513
rect -5626 -12565 -5574 -12513
rect -6223 -13115 -6171 -13063
rect -6426 -13905 -6374 -13853
rect -5000 -12325 -4948 -12273
rect -4502 -12324 -4450 -12272
rect -5376 -12441 -5324 -12389
rect -5127 -12441 -5075 -12389
rect -4877 -12565 -4825 -12513
rect -4627 -12565 -4575 -12513
rect -4377 -12441 -4325 -12389
rect -3928 -12442 -3876 -12390
rect -5751 -13115 -5699 -13063
rect -5251 -13242 -5199 -13190
rect -4752 -13115 -4700 -13063
rect -4251 -13242 -4199 -13190
rect -6077 -13798 -6025 -13746
rect -5376 -13798 -5324 -13746
rect -5626 -13905 -5574 -13853
rect -5730 -14010 -5678 -13958
rect -5126 -13798 -5074 -13746
rect -4877 -13905 -4825 -13853
rect -4376 -13798 -4324 -13746
rect -4627 -13905 -4575 -13853
rect -4752 -14010 -4700 -13958
rect -3788 -13242 -3736 -13190
rect -3928 -13905 -3876 -13853
rect -3788 -14010 -3736 -13958
rect -6223 -14108 -6171 -14056
rect -5250 -14108 -5198 -14056
rect -4250 -14108 -4198 -14056
rect -6159 -14848 -6107 -14796
rect -5860 -14848 -5808 -14796
rect -5504 -14954 -5452 -14902
rect -6159 -15535 -6107 -15483
rect -5860 -15641 -5808 -15589
rect -5504 -15534 -5452 -15482
rect -6159 -16246 -6107 -16194
rect -5860 -16347 -5808 -16295
rect -5504 -16246 -5452 -16194
rect -5147 -14848 -5095 -14796
rect -5148 -15642 -5096 -15590
rect -5148 -16347 -5096 -16295
rect -4791 -14954 -4739 -14902
rect -4792 -15534 -4740 -15482
rect -4792 -16246 -4740 -16194
rect -4436 -14848 -4384 -14796
rect 4771 -7907 4823 -7855
rect 4906 -7905 4958 -7853
rect 5037 -7903 5089 -7851
rect -3382 -7986 -3330 -7934
rect -1382 -7975 -1330 -7923
rect -3542 -13242 -3490 -13190
rect -1203 -7976 -1151 -7924
rect -1025 -7975 -973 -7923
rect -848 -7975 -796 -7923
rect -670 -7975 -618 -7923
rect -490 -7975 -438 -7923
rect 755 -7975 807 -7923
rect 932 -7975 984 -7923
rect 1112 -7975 1164 -7923
rect 1289 -7976 1341 -7924
rect 1467 -7975 1519 -7923
rect 1644 -7975 1696 -7923
rect 2890 -7975 2942 -7923
rect 3069 -7975 3121 -7923
rect 3247 -7975 3299 -7923
rect 3424 -7975 3476 -7923
rect 3603 -7976 3655 -7924
rect 3778 -7975 3830 -7923
rect 4208 -7976 4260 -7924
rect -1916 -8587 -1864 -8535
rect -1739 -8587 -1687 -8535
rect -1826 -8706 -1774 -8654
rect -2447 -8820 -2395 -8768
rect -2005 -8820 -1953 -8768
rect -2315 -9978 -2263 -9926
rect -2447 -12325 -2395 -12273
rect -3382 -14108 -3330 -14056
rect -3936 -14954 -3884 -14902
rect -4435 -15641 -4383 -15589
rect -4436 -16347 -4384 -16295
rect -3935 -15641 -3883 -15589
rect -1916 -9599 -1864 -9547
rect -1916 -9978 -1864 -9926
rect -1558 -8587 -1506 -8535
rect -1382 -8587 -1330 -8535
rect -1470 -8706 -1418 -8654
rect -1648 -8820 -1596 -8768
rect -1738 -9599 -1686 -9547
rect -1738 -9979 -1686 -9927
rect -1558 -9599 -1506 -9547
rect -1560 -9978 -1508 -9926
rect -1203 -8587 -1151 -8535
rect -1293 -8820 -1241 -8768
rect -1382 -9977 -1330 -9925
rect -1026 -8587 -974 -8535
rect -1115 -8706 -1063 -8654
rect -848 -8587 -796 -8535
rect -936 -8820 -884 -8768
rect -670 -8587 -618 -8535
rect -758 -8706 -706 -8654
rect -491 -8587 -439 -8535
rect -580 -8819 -528 -8767
rect -314 -8587 -262 -8535
rect -402 -8706 -350 -8654
rect -136 -8587 -84 -8535
rect 42 -8587 94 -8535
rect -47 -8706 5 -8654
rect -225 -8820 -173 -8768
rect -312 -9599 -260 -9547
rect -314 -9978 -262 -9926
rect -136 -9598 -84 -9546
rect -136 -9979 -84 -9927
rect 221 -8587 273 -8535
rect 398 -8587 450 -8535
rect 310 -8706 362 -8654
rect 132 -8821 184 -8769
rect 42 -9599 94 -9547
rect 43 -9978 95 -9926
rect 222 -9598 274 -9546
rect 220 -9978 272 -9926
rect 577 -8587 629 -8535
rect 754 -8587 806 -8535
rect 666 -8706 718 -8654
rect 489 -8819 541 -8767
rect 399 -9599 451 -9547
rect 398 -9978 450 -9926
rect 577 -9599 629 -9547
rect 576 -9978 628 -9926
rect 932 -8587 984 -8535
rect 843 -8819 895 -8767
rect 1111 -8587 1163 -8535
rect 1022 -8706 1074 -8654
rect 1289 -8587 1341 -8535
rect 1201 -8820 1253 -8768
rect 1466 -8587 1518 -8535
rect 1377 -8706 1429 -8654
rect 1644 -8587 1696 -8535
rect 1556 -8820 1608 -8768
rect 1822 -8587 1874 -8535
rect 1733 -8706 1785 -8654
rect 2000 -8587 2052 -8535
rect 2178 -8587 2230 -8535
rect 2090 -8706 2142 -8654
rect 1911 -8820 1963 -8768
rect 2357 -8587 2409 -8535
rect 2534 -8587 2586 -8535
rect 2446 -8706 2498 -8654
rect 2267 -8820 2319 -8768
rect 2178 -9600 2230 -9548
rect 2357 -9599 2409 -9547
rect 2356 -9978 2408 -9926
rect 2712 -8587 2764 -8535
rect 2890 -8587 2942 -8535
rect 2802 -8706 2854 -8654
rect 2624 -8820 2676 -8768
rect 2534 -9599 2586 -9547
rect 2534 -9978 2586 -9926
rect 2713 -9599 2765 -9547
rect 2712 -9979 2764 -9927
rect 3068 -8587 3120 -8535
rect 2980 -8820 3032 -8768
rect 2891 -9978 2943 -9926
rect 3246 -8587 3298 -8535
rect 3158 -8706 3210 -8654
rect 3069 -9978 3121 -9926
rect 3424 -8587 3476 -8535
rect 3336 -8820 3388 -8768
rect 3246 -9978 3298 -9926
rect 3602 -8587 3654 -8535
rect 3513 -8706 3565 -8654
rect 3781 -8587 3833 -8535
rect 3692 -8820 3744 -8768
rect 3869 -8706 3921 -8654
rect 4771 -9367 4823 -9315
rect 4208 -9599 4260 -9547
rect -1827 -10961 -1775 -10909
rect -1470 -10961 -1418 -10909
rect -2004 -11690 -1952 -11638
rect -1915 -11972 -1863 -11920
rect -2005 -12595 -1953 -12543
rect -1649 -11581 -1597 -11529
rect -1738 -11972 -1686 -11920
rect -1559 -11972 -1507 -11920
rect -1649 -12595 -1597 -12543
rect -1114 -10961 -1062 -10909
rect -1293 -11581 -1241 -11529
rect -1381 -11972 -1329 -11920
rect -1203 -11972 -1151 -11920
rect -1294 -12707 -1242 -12655
rect -758 -10961 -706 -10909
rect -937 -11581 -885 -11529
rect -1025 -11972 -973 -11920
rect -848 -11972 -796 -11920
rect -937 -12836 -885 -12784
rect -402 -10961 -350 -10909
rect -46 -10961 6 -10909
rect 309 -10961 361 -10909
rect 665 -10961 717 -10909
rect 931 -10961 983 -10909
rect 1199 -10961 1251 -10909
rect -580 -11690 -528 -11638
rect -670 -11972 -618 -11920
rect -492 -11972 -440 -11920
rect -582 -12706 -530 -12654
rect -224 -11810 -172 -11758
rect -314 -11972 -262 -11920
rect -136 -11972 -84 -11920
rect -224 -12836 -172 -12784
rect 131 -11810 183 -11758
rect 42 -11972 94 -11920
rect 220 -11972 272 -11920
rect 130 -12706 182 -12654
rect -2004 -13598 -1952 -13546
rect -1648 -13725 -1596 -13673
rect -581 -13598 -529 -13546
rect -1291 -13725 -1239 -13673
rect -937 -13725 -885 -13673
rect -225 -13847 -173 -13795
rect 487 -11810 539 -11758
rect 399 -11972 451 -11920
rect 577 -11972 629 -11920
rect 486 -12837 538 -12785
rect 1556 -10961 1608 -10909
rect 1377 -11581 1429 -11529
rect 1288 -11972 1340 -11920
rect 1468 -11972 1520 -11920
rect 1378 -12836 1430 -12784
rect 1913 -10961 1965 -10909
rect 1733 -11581 1785 -11529
rect 1644 -11973 1696 -11921
rect 1823 -11972 1875 -11920
rect 1735 -12707 1787 -12655
rect 2268 -10961 2320 -10909
rect 2623 -10961 2675 -10909
rect 2980 -10961 3032 -10909
rect 3335 -10961 3387 -10909
rect 2089 -11581 2141 -11529
rect 2000 -11972 2052 -11920
rect 2178 -11972 2230 -11920
rect 2088 -12835 2140 -12783
rect 2446 -11690 2498 -11638
rect 2357 -11972 2409 -11920
rect 2534 -11972 2586 -11920
rect 2445 -12706 2497 -12654
rect 2800 -11810 2852 -11758
rect 2713 -11972 2765 -11920
rect 2890 -11972 2942 -11920
rect 2801 -12835 2853 -12783
rect 3157 -11810 3209 -11758
rect 3068 -11972 3120 -11920
rect 3247 -11972 3299 -11920
rect 3158 -12705 3210 -12653
rect 133 -13847 185 -13795
rect 487 -13848 539 -13796
rect 1379 -13725 1431 -13673
rect 1732 -13725 1784 -13673
rect 2091 -13725 2143 -13673
rect 2446 -13598 2498 -13546
rect 2802 -13847 2854 -13795
rect 3692 -10961 3744 -10909
rect 3513 -11810 3565 -11758
rect 3425 -11972 3477 -11920
rect 3603 -11972 3655 -11920
rect 3514 -12595 3566 -12543
rect 3871 -11691 3923 -11639
rect 3781 -11972 3833 -11920
rect 3871 -12595 3923 -12543
rect 3157 -13848 3209 -13796
rect 3870 -13598 3922 -13546
rect 3512 -13847 3564 -13795
rect -2315 -14596 -2263 -14544
rect -2447 -15874 -2395 -15822
rect -2005 -15875 -1953 -15823
rect -1915 -15986 -1863 -15934
rect -3935 -16347 -3883 -16295
rect -5682 -16939 -5630 -16887
rect -6159 -17060 -6107 -17008
rect -5859 -17060 -5807 -17008
rect -5326 -16939 -5274 -16887
rect -4970 -16939 -4918 -16887
rect -5148 -17060 -5096 -17008
rect -5504 -17171 -5452 -17119
rect -4614 -16939 -4562 -16887
rect -4258 -16939 -4206 -16887
rect -4437 -17060 -4385 -17008
rect -1917 -16595 -1865 -16543
rect -1649 -15875 -1597 -15823
rect -1738 -15986 -1686 -15934
rect -1560 -15986 -1508 -15934
rect -1738 -16595 -1686 -16543
rect -1561 -16594 -1509 -16542
rect -1827 -16718 -1775 -16666
rect -1381 -14596 -1329 -14544
rect -1204 -14596 -1152 -14544
rect -1293 -15875 -1241 -15823
rect -1382 -15986 -1330 -15934
rect -1204 -15986 -1152 -15934
rect -1381 -16596 -1329 -16544
rect -1204 -16595 -1152 -16543
rect -1026 -14596 -974 -14544
rect -848 -14596 -796 -14544
rect -847 -14979 -795 -14927
rect -937 -15875 -885 -15823
rect -1025 -15986 -973 -15934
rect -847 -15986 -795 -15934
rect -1026 -16595 -974 -16543
rect -669 -14596 -617 -14544
rect -669 -14979 -617 -14927
rect -491 -14596 -439 -14544
rect -491 -14979 -439 -14927
rect -581 -15875 -529 -15823
rect -670 -15986 -618 -15934
rect -491 -15986 -439 -15934
rect -1692 -16718 -1640 -16666
rect -1628 -16718 -1576 -16666
rect -4792 -17171 -4740 -17119
rect -3935 -17170 -3883 -17118
rect -1471 -16719 -1419 -16667
rect -1114 -16718 -1062 -16666
rect -759 -16717 -707 -16665
rect -314 -14980 -262 -14928
rect -137 -14979 -85 -14927
rect -225 -15875 -173 -15823
rect -313 -15986 -261 -15934
rect -136 -15986 -84 -15934
rect 43 -14979 95 -14927
rect 132 -15874 184 -15822
rect 43 -15986 95 -15934
rect 221 -15986 273 -15934
rect 220 -16595 272 -16543
rect -617 -16718 -565 -16666
rect -553 -16718 -501 -16666
rect -403 -16718 -351 -16666
rect 487 -15875 539 -15823
rect 398 -15986 450 -15934
rect 575 -15986 627 -15934
rect 397 -16595 449 -16543
rect 576 -16595 628 -16543
rect 843 -15875 895 -15823
rect 755 -15986 807 -15934
rect 931 -15986 983 -15934
rect 755 -16595 807 -16543
rect 933 -16595 985 -16543
rect 1288 -14596 1340 -14544
rect 1289 -14980 1341 -14928
rect 1201 -15875 1253 -15823
rect 1110 -15986 1162 -15934
rect 1289 -15986 1341 -15934
rect 1111 -16595 1163 -16543
rect 1466 -14596 1518 -14544
rect 1467 -14979 1519 -14927
rect 1644 -14596 1696 -14544
rect 1644 -14979 1696 -14927
rect 1555 -15875 1607 -15823
rect 1466 -15986 1518 -15934
rect 1643 -15986 1695 -15934
rect -47 -16718 5 -16666
rect 309 -16719 361 -16667
rect 452 -16718 504 -16666
rect 516 -16718 568 -16666
rect 665 -16718 717 -16666
rect 1021 -16718 1073 -16666
rect 1377 -16718 1429 -16666
rect 1823 -14595 1875 -14543
rect 1822 -14979 1874 -14927
rect 2000 -14596 2052 -14544
rect 1999 -14979 2051 -14927
rect 1910 -15875 1962 -15823
rect 1822 -15986 1874 -15934
rect 2000 -15986 2052 -15934
rect 2178 -14596 2230 -14544
rect 2180 -14979 2232 -14927
rect 2267 -15875 2319 -15823
rect 2179 -15986 2231 -15934
rect 2356 -15986 2408 -15934
rect 2356 -16595 2408 -16543
rect 2624 -15875 2676 -15823
rect 2534 -15986 2586 -15934
rect 2712 -15986 2764 -15934
rect 2534 -16595 2586 -16543
rect 2713 -16594 2765 -16542
rect 1528 -16718 1580 -16666
rect 1592 -16718 1644 -16666
rect 1735 -16718 1787 -16666
rect 2090 -16717 2142 -16665
rect 2445 -16718 2497 -16666
rect 2979 -15875 3031 -15823
rect 2891 -15986 2943 -15934
rect 3068 -15986 3120 -15934
rect 2891 -16595 2943 -16543
rect 3070 -16595 3122 -16543
rect 3246 -14597 3298 -14545
rect 3424 -14596 3476 -14544
rect 3425 -14979 3477 -14927
rect 3335 -15875 3387 -15823
rect 3247 -15986 3299 -15934
rect 3424 -15986 3476 -15934
rect 3249 -16595 3301 -16543
rect 2592 -16718 2644 -16666
rect 2656 -16718 2708 -16666
rect 2801 -16718 2853 -16666
rect 3157 -16717 3209 -16665
rect 3602 -14596 3654 -14544
rect 3603 -14979 3655 -14927
rect 3781 -14596 3833 -14544
rect 3780 -14979 3832 -14927
rect 5184 -7908 5236 -7856
rect 5337 -7903 5389 -7851
rect 5185 -8687 5237 -8635
rect 11054 -8769 11106 -8717
rect 11345 -8769 11397 -8717
rect 11638 -8769 11690 -8717
rect 11932 -8769 11984 -8717
rect 12222 -8769 12274 -8717
rect 6769 -9367 6821 -9315
rect 6679 -9598 6731 -9546
rect 5337 -9978 5389 -9926
rect 6680 -10366 6732 -10314
rect 6947 -9368 6999 -9316
rect 7126 -9368 7178 -9316
rect 6858 -10520 6910 -10468
rect 7303 -9366 7355 -9314
rect 7214 -10519 7266 -10467
rect 7037 -11419 7089 -11367
rect 7482 -9366 7534 -9314
rect 7659 -9368 7711 -9316
rect 7571 -10519 7623 -10467
rect 7393 -11419 7445 -11367
rect 7837 -9367 7889 -9315
rect 8015 -9368 8067 -9316
rect 7927 -10519 7979 -10467
rect 7748 -11420 7800 -11368
rect 8194 -9367 8246 -9315
rect 8371 -9367 8423 -9315
rect 8283 -10520 8335 -10468
rect 8103 -11419 8155 -11367
rect 8549 -9367 8601 -9315
rect 8727 -9368 8779 -9316
rect 8638 -10519 8690 -10467
rect 8461 -11419 8513 -11367
rect 8906 -9367 8958 -9315
rect 11144 -9427 11196 -9375
rect 11436 -9428 11488 -9376
rect 11728 -9428 11780 -9376
rect 12020 -9429 12072 -9377
rect 12312 -9428 12364 -9376
rect 9171 -10367 9223 -10315
rect 8995 -10520 9047 -10468
rect 8817 -11419 8869 -11367
rect 11053 -11727 11105 -11675
rect 11347 -11728 11399 -11676
rect 11638 -11727 11690 -11675
rect 11931 -11727 11983 -11675
rect 12223 -11727 12275 -11675
rect 13022 -11726 13074 -11674
rect 5037 -13349 5089 -13297
rect 5534 -13349 5586 -13297
rect 5031 -13486 5083 -13434
rect 4905 -14598 4957 -14546
rect 4239 -14979 4291 -14927
rect 3692 -15875 3744 -15823
rect 3603 -15986 3655 -15934
rect 3780 -15986 3832 -15934
rect 5400 -13598 5452 -13546
rect 5142 -13847 5194 -13795
rect 5143 -14711 5195 -14659
rect 4238 -15592 4290 -15540
rect 5031 -15593 5083 -15541
rect 4238 -16595 4290 -16543
rect 3514 -16719 3566 -16667
rect 3660 -16718 3712 -16666
rect 3724 -16718 3776 -16666
rect 3868 -16718 3920 -16666
rect 5534 -13725 5586 -13673
rect 8950 -13486 9002 -13434
rect 9305 -13486 9357 -13434
rect 8772 -13609 8824 -13557
rect 7526 -13725 7578 -13673
rect 7348 -13849 7400 -13797
rect 5833 -13975 5885 -13923
rect 6013 -13975 6065 -13923
rect 6190 -13976 6242 -13924
rect 6369 -13975 6421 -13923
rect 6547 -13976 6599 -13924
rect 6725 -13975 6777 -13923
rect 6902 -13975 6954 -13923
rect 5746 -14598 5798 -14546
rect 5924 -14711 5976 -14659
rect 6101 -14598 6153 -14546
rect 6279 -14711 6331 -14659
rect 6459 -14598 6511 -14546
rect 6813 -14598 6865 -14546
rect 6636 -14711 6688 -14659
rect 6991 -14711 7043 -14659
rect 5745 -15592 5797 -15540
rect 5400 -15706 5452 -15654
rect 5747 -15803 5799 -15751
rect 5923 -15705 5975 -15653
rect 5921 -16001 5973 -15949
rect 6101 -15592 6153 -15540
rect 6101 -15802 6153 -15750
rect 6279 -15705 6331 -15653
rect 6279 -16001 6331 -15949
rect 6458 -15592 6510 -15540
rect 6456 -15803 6508 -15751
rect 7437 -13975 7489 -13923
rect 6993 -14877 7045 -14825
rect 7347 -14877 7399 -14825
rect 6635 -15705 6687 -15653
rect 6713 -15804 6765 -15752
rect 6634 -16001 6686 -15949
rect 6813 -15904 6865 -15852
rect 7080 -14976 7132 -14924
rect 7260 -14977 7312 -14925
rect 7439 -14976 7491 -14924
rect 7882 -13726 7934 -13674
rect 8238 -13724 8290 -13672
rect 7704 -13848 7756 -13796
rect 7615 -13975 7667 -13923
rect 7793 -13976 7845 -13924
rect 8061 -13849 8113 -13797
rect 7970 -13975 8022 -13923
rect 8148 -13975 8200 -13923
rect 8415 -13849 8467 -13797
rect 8326 -13975 8378 -13923
rect 8861 -13975 8913 -13923
rect 9127 -13609 9179 -13557
rect 9038 -13975 9090 -13923
rect 9217 -13975 9269 -13923
rect 9483 -13609 9535 -13557
rect 9394 -13975 9446 -13923
rect 11442 -13725 11494 -13673
rect 11798 -13725 11850 -13673
rect 11264 -13849 11316 -13797
rect 9929 -13976 9981 -13924
rect 10108 -13975 10160 -13923
rect 10284 -13976 10336 -13924
rect 10462 -13976 10514 -13924
rect 10640 -13975 10692 -13923
rect 10819 -13976 10871 -13924
rect 7704 -14878 7756 -14826
rect 8236 -14598 8288 -14546
rect 8060 -14874 8112 -14822
rect 7169 -15803 7221 -15751
rect 7169 -15905 7221 -15853
rect 6994 -16004 7046 -15952
rect 7526 -15802 7578 -15750
rect 7526 -16006 7578 -15954
rect 7882 -15802 7934 -15750
rect 8060 -15904 8112 -15852
rect 8417 -14710 8469 -14658
rect 8327 -14976 8379 -14924
rect 7881 -16005 7933 -15953
rect 8237 -16005 8289 -15953
rect 6548 -16597 6600 -16545
rect 6726 -16597 6778 -16545
rect 6903 -16598 6955 -16546
rect 5399 -16720 5451 -16668
rect 5031 -16835 5083 -16783
rect 7970 -16598 8022 -16546
rect 8149 -16597 8201 -16545
rect 8595 -14598 8647 -14546
rect 8504 -14859 8556 -14807
rect 8505 -14977 8557 -14925
rect 8772 -14711 8824 -14659
rect 8683 -14977 8735 -14925
rect 8950 -14599 9002 -14547
rect 9127 -14712 9179 -14660
rect 9304 -14598 9356 -14546
rect 9661 -14598 9713 -14546
rect 9483 -14711 9535 -14659
rect 9572 -14976 9624 -14924
rect 9837 -14712 9889 -14660
rect 9753 -14859 9805 -14807
rect 9750 -14976 9802 -14924
rect 10016 -14598 10068 -14546
rect 9929 -14976 9981 -14924
rect 10373 -14599 10425 -14547
rect 10196 -14711 10248 -14659
rect 10195 -14875 10247 -14823
rect 10550 -14711 10602 -14659
rect 10552 -14868 10604 -14816
rect 10729 -14598 10781 -14546
rect 10908 -14711 10960 -14659
rect 11087 -14711 11139 -14659
rect 10908 -14866 10960 -14814
rect 11353 -13975 11405 -13923
rect 11620 -13850 11672 -13798
rect 11530 -13975 11582 -13923
rect 11709 -13975 11761 -13923
rect 12152 -13726 12204 -13674
rect 12509 -13725 12561 -13673
rect 11977 -13849 12029 -13797
rect 11886 -13976 11938 -13924
rect 12064 -13975 12116 -13923
rect 12334 -13849 12386 -13797
rect 12242 -13976 12294 -13924
rect 12420 -13975 12472 -13923
rect 11440 -14709 11492 -14657
rect 10819 -14976 10871 -14924
rect 8593 -15905 8645 -15853
rect 9663 -15905 9715 -15853
rect 8771 -16719 8823 -16667
rect 9128 -16719 9180 -16667
rect 10373 -15804 10425 -15752
rect 10194 -15905 10246 -15853
rect 10730 -15803 10782 -15751
rect 11264 -14868 11316 -14816
rect 10996 -14976 11048 -14924
rect 11175 -14976 11227 -14924
rect 11086 -15803 11138 -15751
rect 11619 -15705 11671 -15653
rect 11084 -15905 11136 -15853
rect 11440 -15894 11492 -15842
rect 9484 -16719 9536 -16667
rect 8950 -16835 9002 -16783
rect 9305 -16835 9357 -16783
rect 7347 -16943 7399 -16891
rect 7704 -16943 7756 -16891
rect 8060 -16943 8112 -16891
rect 8416 -16943 8468 -16891
rect 9929 -16597 9981 -16545
rect 9838 -16719 9890 -16667
rect 10107 -16598 10159 -16546
rect 10287 -16598 10339 -16546
rect 10195 -16718 10247 -16666
rect 10550 -16718 10602 -16666
rect 11441 -16005 11493 -15953
rect 11798 -15593 11850 -15541
rect 11797 -16005 11849 -15953
rect 11975 -15705 12027 -15653
rect 12155 -15592 12207 -15540
rect 12154 -16005 12206 -15953
rect 12332 -15705 12384 -15653
rect 12511 -15592 12563 -15540
rect 12511 -16005 12563 -15953
rect 10907 -16718 10959 -16666
rect 10017 -16834 10069 -16782
rect 10374 -16834 10426 -16782
rect 10731 -16832 10783 -16780
rect 11352 -16598 11404 -16546
rect 11530 -16599 11582 -16547
rect 11709 -16598 11761 -16546
rect 11263 -16943 11315 -16891
rect 11620 -16943 11672 -16891
rect 11975 -16942 12027 -16890
rect 12331 -16942 12383 -16890
rect 18348 -13485 18400 -13433
<< metal2 >>
rect -5867 -1910 -5814 -1900
rect -5689 -1910 -5636 -1900
rect -5510 -1910 -5457 -1900
rect -5333 -1910 -5280 -1900
rect -5155 -1910 -5102 -1900
rect -4976 -1910 -4923 -1900
rect -4799 -1910 -4746 -1900
rect -4621 -1910 -4568 -1900
rect -4443 -1910 -4390 -1900
rect -4265 -1910 -4212 -1900
rect -4086 -1910 -4033 -1900
rect -3909 -1910 -3856 -1900
rect -1109 -1910 -1056 -1900
rect -5867 -1911 -1056 -1910
rect -5815 -1963 -5689 -1911
rect -5637 -1963 -5510 -1911
rect -5458 -1963 -5333 -1911
rect -5281 -1963 -5155 -1911
rect -5103 -1963 -4976 -1911
rect -4924 -1963 -4799 -1911
rect -4747 -1963 -4621 -1911
rect -4569 -1963 -4443 -1911
rect -4391 -1963 -4265 -1911
rect -4213 -1963 -4086 -1911
rect -4034 -1963 -3909 -1911
rect -3857 -1963 -1109 -1911
rect -1057 -1963 -1056 -1911
rect -5867 -1973 -5814 -1963
rect -5689 -1973 -5636 -1963
rect -5510 -1973 -5457 -1963
rect -5333 -1973 -5280 -1963
rect -5155 -1973 -5102 -1963
rect -4976 -1973 -4923 -1963
rect -4799 -1973 -4746 -1963
rect -4621 -1973 -4568 -1963
rect -4443 -1973 -4390 -1963
rect -4265 -1973 -4212 -1963
rect -4086 -1973 -4033 -1963
rect -3909 -1973 -3856 -1963
rect -1109 -1973 -1056 -1963
rect 5337 -2205 5390 -2195
rect 6680 -2205 6744 -2189
rect 5337 -2206 6686 -2205
rect 5389 -2257 6686 -2206
rect 6738 -2257 6748 -2205
rect 5389 -2258 6748 -2257
rect 5337 -2268 5390 -2258
rect 6680 -2273 6744 -2258
rect -1109 -2425 -1056 -2415
rect -752 -2425 -699 -2415
rect -1109 -2426 -699 -2425
rect -1057 -2478 -752 -2426
rect -700 -2478 -699 -2426
rect -1109 -2488 -1056 -2478
rect -752 -2488 -699 -2478
rect 1919 -2426 1972 -2416
rect 2275 -2426 2328 -2416
rect 3193 -2426 3246 -2417
rect 1919 -2427 3246 -2426
rect 1971 -2479 2275 -2427
rect 2327 -2428 3246 -2427
rect 2327 -2479 3193 -2428
rect 1919 -2489 1972 -2479
rect 2275 -2489 2328 -2479
rect 3245 -2480 3246 -2428
rect 3193 -2490 3246 -2480
rect -6498 -2529 -6445 -2519
rect -5777 -2529 -5724 -2520
rect -6498 -2530 -5724 -2529
rect -5066 -2530 -5013 -2520
rect -4354 -2530 -4301 -2520
rect -6446 -2531 -4301 -2530
rect -6446 -2582 -5777 -2531
rect -6498 -2592 -6445 -2582
rect -5725 -2583 -5066 -2531
rect -5014 -2583 -4354 -2531
rect -4302 -2583 -4301 -2531
rect -5777 -2593 -5724 -2583
rect -5066 -2593 -5013 -2583
rect -4354 -2593 -4301 -2583
rect -2624 -2558 -2571 -2548
rect -1285 -2558 -1232 -2548
rect -930 -2558 -877 -2548
rect -2624 -2559 -877 -2558
rect -2572 -2611 -1285 -2559
rect -1233 -2611 -930 -2559
rect -878 -2611 -877 -2559
rect -2624 -2621 -2571 -2611
rect -1285 -2621 -1232 -2611
rect -930 -2621 -877 -2611
rect 2097 -2554 2150 -2544
rect 2453 -2554 2506 -2544
rect 2097 -2555 2506 -2554
rect 2149 -2607 2453 -2555
rect 2505 -2607 2506 -2555
rect 2097 -2617 2150 -2607
rect 2453 -2617 2506 -2607
rect -5421 -2668 -5368 -2658
rect -4710 -2668 -4657 -2658
rect -3998 -2668 -3945 -2658
rect -3298 -2668 -3245 -2658
rect -5421 -2669 -3245 -2668
rect -5369 -2721 -4710 -2669
rect -4658 -2721 -3998 -2669
rect -3946 -2721 -3298 -2669
rect -3246 -2721 -3245 -2669
rect -5421 -2731 -5368 -2721
rect -4710 -2731 -4657 -2721
rect -3998 -2731 -3945 -2721
rect -3298 -2731 -3245 -2721
rect -1197 -2665 -1144 -2655
rect -1019 -2665 -966 -2655
rect -841 -2665 -788 -2655
rect -129 -2665 -76 -2655
rect 50 -2665 103 -2655
rect 227 -2665 280 -2655
rect 940 -2665 993 -2655
rect 1117 -2665 1170 -2655
rect 1295 -2665 1348 -2655
rect 2007 -2665 2060 -2655
rect 2186 -2665 2239 -2655
rect 2363 -2665 2416 -2655
rect -1197 -2666 2416 -2665
rect -1145 -2718 -1019 -2666
rect -967 -2718 -841 -2666
rect -789 -2718 -129 -2666
rect -77 -2718 50 -2666
rect 102 -2718 227 -2666
rect 279 -2718 940 -2666
rect 992 -2718 1117 -2666
rect 1169 -2718 1295 -2666
rect 1347 -2718 2007 -2666
rect 2059 -2718 2186 -2666
rect 2238 -2718 2363 -2666
rect 2415 -2718 2416 -2666
rect -1197 -2728 -1144 -2718
rect -1019 -2728 -966 -2718
rect -841 -2728 -788 -2718
rect -129 -2728 -76 -2718
rect 50 -2728 103 -2718
rect 227 -2728 280 -2718
rect 940 -2728 993 -2718
rect 1117 -2728 1170 -2718
rect 1295 -2728 1348 -2718
rect 2007 -2728 2060 -2718
rect 2186 -2728 2239 -2718
rect 2363 -2728 2416 -2718
rect -6044 -2780 -5991 -2770
rect -5866 -2780 -5813 -2770
rect -6044 -2781 -5813 -2780
rect -5992 -2833 -5866 -2781
rect -5814 -2833 -5813 -2781
rect -6044 -2843 -5991 -2833
rect -5866 -2843 -5813 -2833
rect -3908 -2780 -3855 -2770
rect -3731 -2780 -3678 -2770
rect -3908 -2781 -3678 -2780
rect -3856 -2833 -3731 -2781
rect -3679 -2833 -3678 -2781
rect -3908 -2843 -3855 -2833
rect -3731 -2843 -3678 -2833
rect -484 -3301 -431 -3291
rect 583 -3301 636 -3291
rect 1654 -3301 1707 -3291
rect -484 -3302 1707 -3301
rect -432 -3354 583 -3302
rect 635 -3354 1654 -3302
rect 1706 -3354 1707 -3302
rect -484 -3364 -431 -3354
rect 583 -3364 636 -3354
rect 1654 -3364 1707 -3354
rect -6625 -3401 -6572 -3391
rect -6134 -3401 -6081 -3391
rect -5066 -3401 -5013 -3391
rect -6625 -3402 -5013 -3401
rect -6573 -3454 -6134 -3402
rect -6082 -3454 -5066 -3402
rect -5014 -3454 -5013 -3402
rect -6625 -3464 -6572 -3454
rect -6134 -3464 -6081 -3454
rect -5066 -3464 -5013 -3454
rect -4710 -3401 -4657 -3391
rect -3642 -3401 -3589 -3391
rect -3131 -3401 -3078 -3391
rect -4710 -3402 -3078 -3401
rect -4658 -3454 -3642 -3402
rect -3590 -3454 -3131 -3402
rect -3079 -3454 -3078 -3402
rect -4710 -3464 -4657 -3454
rect -3642 -3464 -3589 -3454
rect -3131 -3464 -3078 -3454
rect -1645 -3454 -1584 -3439
rect -1645 -3506 -1641 -3454
rect -1589 -3456 -1584 -3454
rect -1108 -3456 -1055 -3446
rect -750 -3456 -697 -3446
rect -396 -3456 -343 -3446
rect -39 -3456 14 -3446
rect 317 -3456 370 -3446
rect -1589 -3457 370 -3456
rect -1589 -3506 -1108 -3457
rect -5777 -3516 -5724 -3506
rect -3998 -3516 -3945 -3506
rect -3298 -3516 -3245 -3506
rect -5777 -3517 -3245 -3516
rect -5725 -3569 -3998 -3517
rect -3946 -3569 -3298 -3517
rect -3246 -3569 -3245 -3517
rect -1645 -3509 -1108 -3506
rect -1056 -3509 -750 -3457
rect -698 -3509 -396 -3457
rect -344 -3509 -39 -3457
rect 13 -3509 317 -3457
rect 369 -3509 370 -3457
rect -1645 -3520 -1584 -3509
rect -1108 -3519 -1055 -3509
rect -750 -3519 -697 -3509
rect -396 -3519 -343 -3509
rect -39 -3519 14 -3509
rect 317 -3519 370 -3509
rect 850 -3456 903 -3446
rect 1206 -3456 1259 -3446
rect 1562 -3456 1615 -3446
rect 1919 -3456 1972 -3446
rect 2275 -3456 2328 -3446
rect 3019 -3455 3080 -3442
rect 3019 -3456 3021 -3455
rect 850 -3457 3021 -3456
rect 902 -3509 1206 -3457
rect 1258 -3509 1562 -3457
rect 1614 -3509 1919 -3457
rect 1971 -3509 2275 -3457
rect 2327 -3509 3021 -3457
rect 850 -3519 903 -3509
rect 1206 -3519 1259 -3509
rect 1562 -3519 1615 -3509
rect 1919 -3519 1972 -3509
rect 2275 -3519 2328 -3509
rect 3019 -3511 3021 -3509
rect 3077 -3456 3080 -3455
rect 6222 -3456 6286 -3441
rect 3077 -3457 6297 -3456
rect 3077 -3509 6228 -3457
rect 6280 -3509 6297 -3457
rect 3077 -3511 3080 -3509
rect 3019 -3523 3080 -3511
rect 6222 -3525 6286 -3509
rect -5777 -3579 -5724 -3569
rect -3998 -3579 -3945 -3569
rect -3298 -3579 -3245 -3569
rect -1286 -3571 -1233 -3561
rect -929 -3571 -876 -3561
rect -573 -3571 -520 -3561
rect -217 -3571 -164 -3561
rect -1702 -3572 -164 -3571
rect -1702 -3624 -1286 -3572
rect -1234 -3624 -929 -3572
rect -877 -3624 -573 -3572
rect -521 -3624 -217 -3572
rect -165 -3624 -164 -3572
rect -6498 -3640 -6445 -3630
rect -5422 -3640 -5369 -3630
rect -4353 -3640 -4300 -3630
rect -1702 -3640 -1649 -3624
rect -1286 -3634 -1233 -3624
rect -929 -3634 -876 -3624
rect -573 -3634 -520 -3624
rect -217 -3634 -164 -3624
rect 1384 -3564 1437 -3554
rect 1741 -3564 1794 -3554
rect 2097 -3564 2150 -3554
rect 2451 -3564 2504 -3554
rect 1384 -3565 2504 -3564
rect 1436 -3617 1741 -3565
rect 1793 -3617 2097 -3565
rect 2149 -3617 2451 -3565
rect 2503 -3617 2504 -3565
rect 1384 -3627 1437 -3617
rect 1741 -3627 1794 -3617
rect 2097 -3627 2150 -3617
rect 2451 -3627 2504 -3617
rect -6498 -3641 -1649 -3640
rect -6446 -3693 -5422 -3641
rect -5370 -3693 -4353 -3641
rect -4301 -3693 -1649 -3641
rect -6498 -3703 -6445 -3693
rect -5422 -3703 -5369 -3693
rect -4353 -3703 -4300 -3693
rect -2546 -3931 -2485 -3693
rect -2546 -3987 -2544 -3931
rect -2488 -3987 -2485 -3931
rect -2546 -3999 -2485 -3987
rect -841 -4192 -788 -4182
rect -662 -4192 -609 -4182
rect -483 -4192 -430 -4182
rect -306 -4192 -253 -4182
rect 407 -4192 460 -4182
rect 583 -4192 636 -4182
rect 761 -4192 814 -4182
rect 1474 -4192 1527 -4182
rect 1652 -4192 1705 -4182
rect 1830 -4192 1883 -4182
rect 2008 -4192 2061 -4182
rect -841 -4193 2061 -4192
rect -789 -4245 -662 -4193
rect -610 -4245 -483 -4193
rect -431 -4245 -306 -4193
rect -254 -4245 407 -4193
rect 459 -4245 583 -4193
rect 635 -4245 761 -4193
rect 813 -4245 1474 -4193
rect 1526 -4245 1652 -4193
rect 1704 -4245 1830 -4193
rect 1882 -4245 2008 -4193
rect 2060 -4245 2061 -4193
rect -841 -4255 -788 -4245
rect -662 -4255 -609 -4245
rect -483 -4255 -430 -4245
rect -306 -4255 -253 -4245
rect 407 -4255 460 -4245
rect 583 -4255 636 -4245
rect 761 -4255 814 -4245
rect 1474 -4255 1527 -4245
rect 1652 -4255 1705 -4245
rect 1830 -4255 1883 -4245
rect 2008 -4255 2061 -4245
rect -6498 -4271 -6445 -4261
rect -5778 -4271 -5725 -4261
rect -3998 -4271 -3945 -4261
rect -6498 -4272 -3945 -4271
rect -6446 -4324 -5778 -4272
rect -5726 -4324 -3998 -4272
rect -3946 -4324 -3945 -4272
rect 2538 -4269 2599 -4256
rect 317 -4304 370 -4294
rect 673 -4304 726 -4294
rect -6498 -4334 -6445 -4324
rect -5778 -4334 -5725 -4324
rect -3998 -4334 -3945 -4324
rect -2357 -4305 726 -4304
rect -2357 -4357 317 -4305
rect 369 -4357 673 -4305
rect 725 -4357 726 -4305
rect 2538 -4325 2540 -4269
rect 2596 -4325 2599 -4269
rect 2538 -4337 2599 -4325
rect -6134 -4390 -6081 -4380
rect -5066 -4390 -5013 -4380
rect -4709 -4390 -4656 -4380
rect -3642 -4390 -3589 -4380
rect -2357 -4390 -2304 -4357
rect 317 -4367 370 -4357
rect 673 -4367 726 -4357
rect -6134 -4391 -2304 -4390
rect -6082 -4443 -5066 -4391
rect -5014 -4443 -4709 -4391
rect -4657 -4443 -3642 -4391
rect -3590 -4443 -2304 -4391
rect -2004 -4412 -1951 -4402
rect 495 -4412 548 -4402
rect 850 -4412 903 -4402
rect -2004 -4413 903 -4412
rect -6134 -4453 -6081 -4443
rect -5066 -4453 -5013 -4443
rect -4709 -4453 -4656 -4443
rect -3642 -4453 -3589 -4443
rect -1952 -4465 495 -4413
rect 547 -4465 850 -4413
rect 902 -4465 903 -4413
rect -2004 -4475 -1951 -4465
rect 495 -4475 548 -4465
rect 850 -4475 903 -4465
rect 2746 -4449 2807 -4436
rect -5422 -4506 -5369 -4496
rect -4353 -4506 -4300 -4496
rect -3298 -4506 -3245 -4496
rect -2385 -4506 -2324 -4495
rect -5422 -4507 -2324 -4506
rect -5370 -4559 -4353 -4507
rect -4301 -4559 -3298 -4507
rect -3246 -4508 -2324 -4507
rect -3246 -4559 -2383 -4508
rect -5422 -4569 -5369 -4559
rect -4353 -4569 -4300 -4559
rect -3298 -4569 -3245 -4559
rect -2385 -4564 -2383 -4559
rect -2327 -4564 -2324 -4508
rect 2746 -4505 2748 -4449
rect 2804 -4505 2807 -4449
rect 2746 -4517 2807 -4505
rect -2385 -4576 -2324 -4564
rect 3194 -4805 3246 -4795
rect 4771 -4805 4823 -4795
rect 3246 -4857 4771 -4805
rect 3194 -4867 3246 -4857
rect 4771 -4867 4823 -4857
rect 3021 -5005 3082 -4992
rect 3021 -5061 3023 -5005
rect 3079 -5007 3082 -5005
rect 5037 -5006 5090 -4996
rect 4985 -5007 5090 -5006
rect 3079 -5059 5037 -5007
rect 5089 -5059 5090 -5007
rect 3079 -5061 3082 -5059
rect 3021 -5073 3082 -5061
rect 5037 -5069 5090 -5059
rect -2385 -5096 -2324 -5083
rect -6498 -5142 -6445 -5131
rect -6446 -5147 -6445 -5142
rect -5422 -5142 -5369 -5131
rect -6446 -5187 -5422 -5147
rect -6446 -5194 -6445 -5187
rect -6498 -5204 -6445 -5194
rect -5370 -5148 -5369 -5142
rect -4353 -5142 -4300 -5131
rect -5370 -5188 -4353 -5148
rect -5370 -5194 -5369 -5188
rect -5422 -5204 -5369 -5194
rect -4301 -5194 -4300 -5142
rect -2385 -5152 -2383 -5096
rect -2327 -5097 -2324 -5096
rect -1287 -5097 -1234 -5087
rect -929 -5097 -876 -5087
rect -572 -5097 -519 -5087
rect -218 -5097 -165 -5087
rect -2327 -5098 -165 -5097
rect -2327 -5150 -1287 -5098
rect -1235 -5150 -929 -5098
rect -877 -5150 -572 -5098
rect -520 -5150 -218 -5098
rect -166 -5150 -165 -5098
rect 1385 -5093 1438 -5083
rect 1740 -5093 1793 -5083
rect 2096 -5093 2149 -5083
rect 2453 -5093 2506 -5083
rect 1385 -5094 2506 -5093
rect -2327 -5152 -2324 -5150
rect -2385 -5164 -2324 -5152
rect -1287 -5160 -1234 -5150
rect -929 -5160 -876 -5150
rect -572 -5160 -519 -5150
rect -218 -5160 -165 -5150
rect 311 -5151 372 -5138
rect -4353 -5204 -4300 -5194
rect -1105 -5213 -1052 -5203
rect -751 -5213 -698 -5203
rect -396 -5213 -343 -5203
rect -41 -5213 12 -5203
rect 311 -5207 313 -5151
rect 369 -5207 372 -5151
rect 1437 -5146 1740 -5094
rect 1792 -5146 2096 -5094
rect 2148 -5146 2453 -5094
rect 2505 -5146 2506 -5094
rect 1385 -5156 1438 -5146
rect 1740 -5156 1793 -5146
rect 2096 -5156 2149 -5146
rect 2453 -5156 2506 -5146
rect 311 -5213 372 -5207
rect -1105 -5214 372 -5213
rect -6134 -5233 -6081 -5222
rect -6082 -5239 -6081 -5233
rect -5066 -5234 -5013 -5223
rect -6082 -5279 -5066 -5239
rect -6082 -5285 -6081 -5279
rect -6134 -5295 -6081 -5285
rect -5014 -5239 -5013 -5234
rect -3130 -5234 -3077 -5223
rect -5014 -5279 -3130 -5239
rect -5014 -5286 -5013 -5279
rect -5066 -5296 -5013 -5286
rect -3078 -5239 -3077 -5234
rect -1876 -5233 -1823 -5222
rect -3078 -5279 -1876 -5239
rect -3078 -5286 -3077 -5279
rect -3130 -5296 -3077 -5286
rect -1824 -5285 -1823 -5233
rect -1053 -5266 -751 -5214
rect -699 -5266 -396 -5214
rect -344 -5266 -41 -5214
rect 11 -5266 316 -5214
rect 368 -5219 372 -5214
rect 846 -5213 903 -5203
rect 1207 -5213 1260 -5203
rect 1563 -5213 1616 -5203
rect 1917 -5213 1970 -5203
rect 2274 -5213 2327 -5203
rect 4905 -5213 4958 -5202
rect 5614 -5213 5678 -5197
rect 846 -5214 4905 -5213
rect 368 -5266 369 -5219
rect -1876 -5295 -1823 -5285
rect -1646 -5281 -1585 -5268
rect -1105 -5276 -1052 -5266
rect -751 -5276 -698 -5266
rect -396 -5276 -343 -5266
rect -41 -5276 12 -5266
rect 316 -5276 369 -5266
rect 846 -5266 850 -5214
rect 902 -5266 1207 -5214
rect 1259 -5266 1563 -5214
rect 1615 -5266 1917 -5214
rect 1969 -5266 2274 -5214
rect 2326 -5265 4905 -5214
rect 4957 -5265 5620 -5213
rect 5672 -5265 5685 -5213
rect 2326 -5266 5685 -5265
rect -6625 -5323 -6572 -5312
rect -6573 -5329 -6572 -5323
rect -4710 -5323 -4657 -5312
rect -6573 -5369 -4710 -5329
rect -6573 -5375 -6572 -5369
rect -6625 -5385 -6572 -5375
rect -4658 -5329 -4657 -5323
rect -3642 -5320 -3589 -5309
rect -4658 -5369 -3642 -5329
rect -4658 -5375 -4657 -5369
rect -4710 -5385 -4657 -5375
rect -3590 -5329 -3589 -5320
rect -2624 -5325 -2571 -5314
rect -3590 -5369 -2624 -5329
rect -3590 -5372 -3589 -5369
rect -3642 -5382 -3589 -5372
rect -2572 -5377 -2571 -5325
rect -1646 -5337 -1644 -5281
rect -1588 -5337 -1585 -5281
rect -1646 -5349 -1585 -5337
rect 846 -5281 907 -5266
rect 1207 -5276 1260 -5266
rect 1563 -5276 1616 -5266
rect 1917 -5276 1970 -5266
rect 2274 -5276 2327 -5266
rect 4905 -5275 4958 -5266
rect 5614 -5281 5678 -5266
rect 846 -5337 848 -5281
rect 904 -5337 907 -5281
rect 846 -5349 907 -5337
rect -2624 -5387 -2571 -5377
rect -128 -5380 -75 -5370
rect 50 -5380 103 -5370
rect 228 -5380 281 -5370
rect 940 -5380 993 -5371
rect 1119 -5380 1172 -5370
rect 1296 -5380 1349 -5370
rect -128 -5381 1349 -5380
rect -5777 -5416 -5724 -5405
rect -5725 -5422 -5724 -5416
rect -3997 -5416 -3944 -5405
rect -5725 -5462 -3997 -5422
rect -5725 -5468 -5724 -5462
rect -5777 -5478 -5724 -5468
rect -3945 -5422 -3944 -5416
rect -3298 -5417 -3245 -5406
rect -3945 -5462 -3298 -5422
rect -3945 -5468 -3944 -5462
rect -3997 -5478 -3944 -5468
rect -3246 -5469 -3245 -5417
rect -76 -5433 50 -5381
rect 102 -5433 228 -5381
rect 280 -5382 1119 -5381
rect 280 -5433 940 -5382
rect -128 -5443 -75 -5433
rect 50 -5443 103 -5433
rect 228 -5443 281 -5433
rect 992 -5433 1119 -5382
rect 1171 -5433 1296 -5381
rect 1348 -5433 1349 -5381
rect 992 -5434 993 -5433
rect 940 -5444 993 -5434
rect 1119 -5443 1172 -5433
rect 1296 -5443 1349 -5433
rect -3298 -5479 -3245 -5469
rect 5337 -5528 5390 -5517
rect 5389 -5580 5390 -5528
rect -5956 -6016 -5903 -6006
rect -5601 -6016 -5548 -6006
rect -5244 -6016 -5191 -6006
rect -4888 -6016 -4835 -6006
rect -4532 -6016 -4479 -6006
rect -4175 -6016 -4122 -6006
rect -3820 -6016 -3767 -6006
rect -5956 -6017 -3767 -6016
rect -5904 -6069 -5601 -6017
rect -5549 -6069 -5244 -6017
rect -5192 -6069 -4888 -6017
rect -4836 -6069 -4532 -6017
rect -4480 -6069 -4175 -6017
rect -4123 -6069 -3820 -6017
rect -3768 -6069 -3767 -6017
rect -5956 -6079 -5903 -6069
rect -5601 -6079 -5548 -6069
rect -5244 -6079 -5191 -6069
rect -4888 -6079 -4835 -6069
rect -4532 -6079 -4479 -6069
rect -4175 -6079 -4122 -6069
rect -3820 -6079 -3767 -6069
rect -2624 -6007 -2571 -5997
rect 2096 -6007 2149 -5997
rect 2452 -6007 2505 -5997
rect -2624 -6008 2505 -6007
rect -2572 -6060 2096 -6008
rect 2148 -6060 2452 -6008
rect 2504 -6060 2505 -6008
rect -2624 -6070 -2571 -6060
rect 2096 -6070 2149 -6060
rect 2452 -6070 2505 -6060
rect -5778 -6131 -5725 -6121
rect -5065 -6131 -5012 -6121
rect -4354 -6131 -4301 -6121
rect -3298 -6131 -3245 -6121
rect 1918 -6124 1971 -6114
rect 2275 -6124 2328 -6114
rect -2821 -6125 2328 -6124
rect -5778 -6132 -3245 -6131
rect -5726 -6184 -5065 -6132
rect -5013 -6184 -4354 -6132
rect -4302 -6184 -3298 -6132
rect -3246 -6184 -3245 -6132
rect -5778 -6194 -5725 -6184
rect -5065 -6194 -5012 -6184
rect -4354 -6194 -4301 -6184
rect -3298 -6194 -3245 -6184
rect -2856 -6177 1918 -6125
rect 1970 -6177 2275 -6125
rect 2327 -6177 2328 -6125
rect -6498 -6248 -6445 -6238
rect -5421 -6248 -5368 -6238
rect -4710 -6248 -4657 -6238
rect -3998 -6248 -3945 -6237
rect -6498 -6249 -3998 -6248
rect -6446 -6301 -5421 -6249
rect -5369 -6301 -4710 -6249
rect -4658 -6300 -3998 -6249
rect -3946 -6300 -3945 -6248
rect -4658 -6301 -3945 -6300
rect -6498 -6311 -6445 -6301
rect -5421 -6311 -5368 -6301
rect -4710 -6311 -4657 -6301
rect -3998 -6310 -3945 -6301
rect -4786 -6379 -4733 -6368
rect -4734 -6408 -4733 -6379
rect -2856 -6401 -2803 -6177
rect 1918 -6187 1971 -6177
rect 2275 -6187 2328 -6177
rect -3874 -6408 -2803 -6401
rect -4734 -6431 -2803 -6408
rect -4786 -6454 -2803 -6431
rect -2702 -6250 -2649 -6249
rect 227 -6250 280 -6240
rect 942 -6250 995 -6240
rect -2702 -6251 995 -6250
rect -2702 -6303 227 -6251
rect 279 -6303 942 -6251
rect 994 -6303 995 -6251
rect -4786 -6461 -3820 -6454
rect -3874 -7691 -3821 -6461
rect -2702 -6542 -2649 -6303
rect 227 -6313 280 -6303
rect 942 -6313 995 -6303
rect -1876 -6364 -1823 -6354
rect -1282 -6364 -1229 -6354
rect -1876 -6365 -1177 -6364
rect -928 -6365 -876 -6355
rect 2879 -6365 2931 -6355
rect -1824 -6417 -1282 -6365
rect -1230 -6417 -928 -6365
rect -876 -6417 2879 -6365
rect -1876 -6427 -1823 -6417
rect -1282 -6427 -1229 -6417
rect -928 -6427 -876 -6417
rect 2879 -6427 2931 -6417
rect -1110 -6479 -1057 -6469
rect -752 -6479 -699 -6469
rect -1110 -6480 -699 -6479
rect -1058 -6532 -752 -6480
rect -700 -6532 -699 -6480
rect -1110 -6542 -1057 -6532
rect -752 -6542 -699 -6532
rect -3874 -7743 -3873 -7691
rect -3873 -7753 -3821 -7743
rect -3731 -6595 -2649 -6542
rect -3731 -7785 -3678 -6595
rect -753 -6598 -700 -6588
rect 4772 -6598 4825 -6587
rect -753 -6599 4772 -6598
rect -701 -6650 4772 -6599
rect 4824 -6650 4825 -6598
rect -701 -6651 4825 -6650
rect -753 -6661 -700 -6651
rect 4772 -6660 4825 -6651
rect -2003 -6714 -1950 -6704
rect -2003 -6715 5237 -6714
rect -1951 -6767 5237 -6715
rect -2003 -6777 -1950 -6767
rect -3545 -6809 -3484 -6796
rect -3545 -6865 -3543 -6809
rect -3487 -6865 -3484 -6809
rect -3545 -6877 -3484 -6865
rect -3679 -7837 -3678 -7785
rect -3541 -7788 -3489 -6877
rect 4770 -6892 4823 -6881
rect 4822 -6944 4823 -6892
rect -3386 -6982 -3325 -6969
rect -3386 -7038 -3384 -6982
rect -3328 -7038 -3325 -6982
rect 4770 -6996 4823 -6944
rect 4906 -6890 4959 -6879
rect 4958 -6942 4959 -6890
rect 4906 -6994 4959 -6942
rect -3386 -7050 -3325 -7038
rect -3731 -7847 -3679 -7837
rect -3541 -7850 -3489 -7840
rect -3382 -7934 -3329 -7050
rect 4771 -7844 4823 -6996
rect 4907 -7842 4959 -6994
rect 5038 -6888 5091 -6877
rect 5090 -6940 5091 -6888
rect 5038 -7840 5091 -6940
rect 4771 -7855 4824 -7844
rect 4823 -7907 4824 -7855
rect -3330 -7986 -3329 -7934
rect -1382 -7922 -1329 -7912
rect -1203 -7922 -1150 -7913
rect -1025 -7922 -972 -7912
rect -848 -7922 -795 -7912
rect -670 -7922 -617 -7912
rect -490 -7922 -437 -7912
rect 755 -7922 808 -7912
rect 932 -7922 985 -7912
rect 1112 -7922 1165 -7912
rect 1289 -7922 1342 -7913
rect 1467 -7922 1520 -7912
rect 1644 -7922 1697 -7912
rect 2890 -7922 2943 -7912
rect 3069 -7922 3122 -7912
rect 3247 -7922 3300 -7912
rect 3424 -7922 3477 -7912
rect 3603 -7922 3656 -7913
rect 3778 -7922 3831 -7912
rect -1382 -7923 3831 -7922
rect 4208 -7923 4261 -7913
rect 4771 -7917 4824 -7907
rect 4906 -7853 4959 -7842
rect 4958 -7905 4959 -7853
rect 4906 -7915 4959 -7905
rect 5037 -7851 5091 -7840
rect 5089 -7898 5091 -7851
rect 5184 -7856 5237 -6767
rect 5089 -7903 5090 -7898
rect 5037 -7913 5090 -7903
rect 5236 -7908 5237 -7856
rect 5184 -7918 5237 -7908
rect 5337 -7851 5390 -5580
rect 5389 -7903 5390 -7851
rect 5337 -7913 5390 -7903
rect 17831 -6527 17895 -6511
rect 17831 -6579 17837 -6527
rect 17889 -6579 17895 -6527
rect -1330 -7924 -1025 -7923
rect -1330 -7975 -1203 -7924
rect -1382 -7985 -1329 -7975
rect -1151 -7975 -1025 -7924
rect -973 -7975 -848 -7923
rect -796 -7975 -670 -7923
rect -618 -7975 -490 -7923
rect -438 -7975 755 -7923
rect 807 -7975 932 -7923
rect 984 -7975 1112 -7923
rect 1164 -7924 1467 -7923
rect 1164 -7975 1289 -7924
rect -1151 -7976 -1150 -7975
rect -1203 -7986 -1150 -7976
rect -1025 -7985 -972 -7975
rect -848 -7985 -795 -7975
rect -670 -7985 -617 -7975
rect -490 -7985 -437 -7975
rect 755 -7985 808 -7975
rect 932 -7985 985 -7975
rect 1112 -7985 1165 -7975
rect 1341 -7975 1467 -7924
rect 1519 -7975 1644 -7923
rect 1696 -7975 2890 -7923
rect 2942 -7975 3069 -7923
rect 3121 -7975 3247 -7923
rect 3299 -7975 3424 -7923
rect 3476 -7924 3778 -7923
rect 3476 -7975 3603 -7924
rect 1341 -7976 1342 -7975
rect 1289 -7986 1342 -7976
rect 1467 -7985 1520 -7975
rect 1644 -7985 1697 -7975
rect 2890 -7985 2943 -7975
rect 3069 -7985 3122 -7975
rect 3247 -7985 3300 -7975
rect 3424 -7985 3477 -7975
rect 3655 -7975 3778 -7924
rect 3830 -7924 4261 -7923
rect 3830 -7975 4208 -7924
rect 3655 -7976 3656 -7975
rect 3603 -7986 3656 -7976
rect 3778 -7976 4208 -7975
rect 4260 -7976 4261 -7924
rect 3778 -7985 3831 -7976
rect 4208 -7986 4261 -7976
rect -3382 -7996 -3329 -7986
rect -1916 -8534 -1863 -8524
rect -1739 -8534 -1686 -8524
rect -1558 -8534 -1505 -8524
rect -1382 -8534 -1329 -8524
rect -1203 -8534 -1150 -8524
rect -1026 -8534 -973 -8524
rect -848 -8534 -795 -8524
rect -670 -8534 -617 -8524
rect -491 -8534 -438 -8524
rect -314 -8534 -261 -8524
rect -136 -8534 -83 -8524
rect 42 -8534 95 -8524
rect 221 -8534 274 -8524
rect 398 -8534 451 -8524
rect 577 -8534 630 -8524
rect 754 -8534 807 -8524
rect 932 -8534 985 -8524
rect 1111 -8534 1164 -8524
rect 1289 -8534 1342 -8524
rect 1466 -8534 1519 -8524
rect 1644 -8534 1697 -8524
rect 1822 -8534 1875 -8524
rect 2000 -8534 2053 -8524
rect 2178 -8534 2231 -8524
rect 2357 -8534 2410 -8524
rect 2534 -8534 2587 -8524
rect 2712 -8534 2765 -8524
rect 2890 -8534 2943 -8524
rect 3068 -8534 3121 -8524
rect 3246 -8534 3299 -8524
rect 3424 -8534 3477 -8524
rect 3602 -8534 3655 -8524
rect 3781 -8534 3834 -8524
rect -1916 -8535 3834 -8534
rect -1864 -8587 -1739 -8535
rect -1687 -8587 -1558 -8535
rect -1506 -8587 -1382 -8535
rect -1330 -8587 -1203 -8535
rect -1151 -8587 -1026 -8535
rect -974 -8587 -848 -8535
rect -796 -8587 -670 -8535
rect -618 -8587 -491 -8535
rect -439 -8587 -314 -8535
rect -262 -8587 -136 -8535
rect -84 -8587 42 -8535
rect 94 -8587 221 -8535
rect 273 -8587 398 -8535
rect 450 -8587 577 -8535
rect 629 -8587 754 -8535
rect 806 -8587 932 -8535
rect 984 -8587 1111 -8535
rect 1163 -8587 1289 -8535
rect 1341 -8587 1466 -8535
rect 1518 -8587 1644 -8535
rect 1696 -8587 1822 -8535
rect 1874 -8587 2000 -8535
rect 2052 -8587 2178 -8535
rect 2230 -8587 2357 -8535
rect 2409 -8587 2534 -8535
rect 2586 -8587 2712 -8535
rect 2764 -8587 2890 -8535
rect 2942 -8587 3068 -8535
rect 3120 -8587 3246 -8535
rect 3298 -8587 3424 -8535
rect 3476 -8587 3602 -8535
rect 3654 -8587 3781 -8535
rect 3833 -8587 3834 -8535
rect -1916 -8597 -1863 -8587
rect -1739 -8597 -1686 -8587
rect -1558 -8597 -1505 -8587
rect -1382 -8597 -1329 -8587
rect -1203 -8597 -1150 -8587
rect -1026 -8597 -973 -8587
rect -848 -8597 -795 -8587
rect -670 -8597 -617 -8587
rect -491 -8597 -438 -8587
rect -314 -8597 -261 -8587
rect -136 -8597 -83 -8587
rect 42 -8597 95 -8587
rect 221 -8597 274 -8587
rect 398 -8597 451 -8587
rect 577 -8597 630 -8587
rect 754 -8597 807 -8587
rect 932 -8597 985 -8587
rect 1111 -8597 1164 -8587
rect 1289 -8597 1342 -8587
rect 1466 -8597 1519 -8587
rect 1644 -8597 1697 -8587
rect 1822 -8597 1875 -8587
rect 2000 -8597 2053 -8587
rect 2178 -8597 2231 -8587
rect 2357 -8597 2410 -8587
rect 2534 -8597 2587 -8587
rect 2712 -8597 2765 -8587
rect 2890 -8597 2943 -8587
rect 3068 -8597 3121 -8587
rect 3246 -8597 3299 -8587
rect 3424 -8597 3477 -8587
rect 3602 -8597 3655 -8587
rect 3781 -8597 3834 -8587
rect 5185 -8633 5237 -8625
rect 5185 -8635 10564 -8633
rect -1826 -8653 -1773 -8643
rect -1470 -8653 -1417 -8643
rect -1115 -8653 -1062 -8643
rect -758 -8653 -705 -8643
rect -402 -8653 -349 -8643
rect -47 -8653 6 -8643
rect 310 -8653 363 -8643
rect 666 -8653 719 -8643
rect 1022 -8653 1075 -8643
rect 1377 -8653 1430 -8643
rect 1733 -8653 1786 -8643
rect 2090 -8653 2143 -8643
rect 2446 -8653 2499 -8643
rect 2802 -8653 2855 -8643
rect 3158 -8653 3211 -8643
rect 3513 -8653 3566 -8643
rect 3869 -8653 3922 -8643
rect -1826 -8654 3922 -8653
rect -1774 -8706 -1470 -8654
rect -1418 -8706 -1115 -8654
rect -1063 -8706 -758 -8654
rect -706 -8706 -402 -8654
rect -350 -8706 -47 -8654
rect 5 -8706 310 -8654
rect 362 -8706 666 -8654
rect 718 -8706 1022 -8654
rect 1074 -8706 1377 -8654
rect 1429 -8706 1733 -8654
rect 1785 -8706 2090 -8654
rect 2142 -8706 2446 -8654
rect 2498 -8706 2802 -8654
rect 2854 -8706 3158 -8654
rect 3210 -8706 3513 -8654
rect 3565 -8706 3869 -8654
rect 3921 -8706 3922 -8654
rect 5237 -8685 10564 -8635
rect 5185 -8697 5237 -8687
rect -1826 -8716 -1773 -8706
rect -1470 -8716 -1417 -8706
rect -1115 -8716 -1062 -8706
rect -758 -8716 -705 -8706
rect -402 -8716 -349 -8706
rect -47 -8716 6 -8706
rect 310 -8716 363 -8706
rect 666 -8716 719 -8706
rect 1022 -8716 1075 -8706
rect 1377 -8716 1430 -8706
rect 1733 -8716 1786 -8706
rect 2090 -8716 2143 -8706
rect 2446 -8716 2499 -8706
rect 2802 -8716 2855 -8706
rect 3158 -8716 3211 -8706
rect 3513 -8716 3566 -8706
rect 3869 -8716 3922 -8706
rect 10512 -8716 10564 -8685
rect 11054 -8716 11107 -8706
rect 11345 -8716 11398 -8706
rect 11638 -8716 11691 -8706
rect 11932 -8716 11985 -8706
rect 12222 -8716 12275 -8706
rect 17831 -8716 17895 -6579
rect 10512 -8717 17895 -8716
rect -2447 -8767 -2394 -8757
rect -2005 -8767 -1952 -8757
rect -1648 -8767 -1595 -8757
rect -1293 -8767 -1240 -8757
rect -936 -8767 -883 -8757
rect -580 -8767 -527 -8756
rect -225 -8767 -172 -8757
rect 132 -8767 185 -8758
rect 489 -8767 542 -8756
rect 843 -8767 896 -8756
rect 1201 -8767 1254 -8757
rect 1556 -8767 1609 -8757
rect 1911 -8767 1964 -8757
rect 2267 -8767 2320 -8757
rect 2624 -8767 2677 -8757
rect 2980 -8767 3033 -8757
rect 3336 -8767 3389 -8757
rect 3692 -8767 3745 -8757
rect -2447 -8768 -580 -8767
rect -2395 -8820 -2005 -8768
rect -1953 -8820 -1648 -8768
rect -1596 -8820 -1293 -8768
rect -1241 -8820 -936 -8768
rect -884 -8819 -580 -8768
rect -528 -8768 489 -8767
rect -528 -8819 -225 -8768
rect -884 -8820 -225 -8819
rect -173 -8769 489 -8768
rect -173 -8820 132 -8769
rect -2447 -8830 -2394 -8820
rect -2005 -8830 -1952 -8820
rect -1648 -8830 -1595 -8820
rect -1293 -8830 -1240 -8820
rect -936 -8830 -883 -8820
rect -580 -8829 -527 -8820
rect -225 -8830 -172 -8820
rect 184 -8819 489 -8769
rect 541 -8819 843 -8767
rect 895 -8768 3745 -8767
rect 10512 -8768 11054 -8717
rect 895 -8819 1201 -8768
rect 184 -8820 1201 -8819
rect 1253 -8820 1556 -8768
rect 1608 -8820 1911 -8768
rect 1963 -8820 2267 -8768
rect 2319 -8820 2624 -8768
rect 2676 -8820 2980 -8768
rect 3032 -8820 3336 -8768
rect 3388 -8820 3692 -8768
rect 3744 -8820 3745 -8768
rect 10584 -8769 11054 -8768
rect 11106 -8769 11345 -8717
rect 11397 -8769 11638 -8717
rect 11690 -8769 11932 -8717
rect 11984 -8769 12222 -8717
rect 12274 -8769 17895 -8717
rect 11054 -8779 11107 -8769
rect 11345 -8779 11398 -8769
rect 11638 -8779 11691 -8769
rect 11932 -8779 11985 -8769
rect 12222 -8779 12275 -8769
rect 184 -8821 185 -8820
rect 132 -8831 185 -8821
rect 489 -8829 542 -8820
rect 843 -8829 896 -8820
rect 1201 -8830 1254 -8820
rect 1556 -8830 1609 -8820
rect 1911 -8830 1964 -8820
rect 2267 -8830 2320 -8820
rect 2624 -8830 2677 -8820
rect 2980 -8830 3033 -8820
rect 3336 -8830 3389 -8820
rect 3692 -8830 3745 -8820
rect 4771 -9314 4824 -9304
rect 6769 -9314 6822 -9304
rect 6947 -9314 7000 -9305
rect 7126 -9314 7179 -9305
rect 7303 -9314 7356 -9303
rect 7482 -9314 7535 -9303
rect 7659 -9314 7712 -9305
rect 7837 -9314 7890 -9304
rect 8015 -9314 8068 -9305
rect 8194 -9314 8247 -9304
rect 8371 -9314 8424 -9304
rect 8549 -9314 8602 -9304
rect 8727 -9314 8780 -9305
rect 8906 -9314 8959 -9304
rect 4771 -9315 7303 -9314
rect 4823 -9367 6769 -9315
rect 6821 -9316 7303 -9315
rect 6821 -9367 6947 -9316
rect 4771 -9377 4824 -9367
rect 6769 -9377 6822 -9367
rect 6999 -9367 7126 -9316
rect 6999 -9368 7000 -9367
rect 6947 -9378 7000 -9368
rect 7178 -9366 7303 -9316
rect 7355 -9366 7482 -9314
rect 7534 -9315 8959 -9314
rect 7534 -9316 7837 -9315
rect 7534 -9366 7659 -9316
rect 7178 -9367 7659 -9366
rect 7178 -9368 7179 -9367
rect 7126 -9378 7179 -9368
rect 7303 -9376 7356 -9367
rect 7482 -9376 7535 -9367
rect 7711 -9367 7837 -9316
rect 7889 -9316 8194 -9315
rect 7889 -9367 8015 -9316
rect 7711 -9368 7712 -9367
rect 7659 -9378 7712 -9368
rect 7837 -9377 7890 -9367
rect 8067 -9367 8194 -9316
rect 8246 -9367 8371 -9315
rect 8423 -9367 8549 -9315
rect 8601 -9316 8906 -9315
rect 8601 -9367 8727 -9316
rect 8067 -9368 8068 -9367
rect 8015 -9378 8068 -9368
rect 8194 -9377 8247 -9367
rect 8371 -9377 8424 -9367
rect 8549 -9377 8602 -9367
rect 8779 -9367 8906 -9316
rect 8958 -9367 8959 -9315
rect 8779 -9368 8780 -9367
rect 8727 -9378 8780 -9368
rect 8906 -9377 8959 -9367
rect 11144 -9375 11197 -9364
rect 11436 -9375 11489 -9365
rect 11728 -9375 11781 -9365
rect 12020 -9375 12073 -9366
rect 12312 -9375 12365 -9365
rect 11196 -9376 12365 -9375
rect 11196 -9427 11436 -9376
rect 11144 -9428 11436 -9427
rect 11488 -9428 11728 -9376
rect 11780 -9377 12312 -9376
rect 11780 -9428 12020 -9377
rect 11144 -9437 11197 -9428
rect 11436 -9438 11489 -9428
rect 11728 -9438 11781 -9428
rect 12072 -9428 12312 -9377
rect 12364 -9428 12365 -9376
rect 12072 -9429 12073 -9428
rect 12020 -9439 12073 -9429
rect 12312 -9438 12365 -9428
rect -1916 -9546 -1863 -9536
rect -1738 -9546 -1685 -9536
rect -1558 -9546 -1505 -9536
rect -312 -9546 -259 -9536
rect -136 -9546 -83 -9535
rect 42 -9546 95 -9536
rect 222 -9546 275 -9535
rect 399 -9546 452 -9536
rect 577 -9546 630 -9536
rect 2178 -9546 2231 -9537
rect 2357 -9546 2410 -9536
rect 2534 -9546 2587 -9536
rect 2713 -9546 2766 -9536
rect 4208 -9546 4261 -9536
rect 6679 -9546 6732 -9535
rect -1916 -9547 -136 -9546
rect -1864 -9599 -1738 -9547
rect -1686 -9599 -1558 -9547
rect -1506 -9599 -312 -9547
rect -260 -9598 -136 -9547
rect -84 -9547 222 -9546
rect -84 -9598 42 -9547
rect -260 -9599 42 -9598
rect 94 -9598 222 -9547
rect 274 -9547 6679 -9546
rect 274 -9598 399 -9547
rect 94 -9599 399 -9598
rect 451 -9599 577 -9547
rect 629 -9548 2357 -9547
rect 629 -9599 2178 -9548
rect -1916 -9609 -1863 -9599
rect -1738 -9609 -1685 -9599
rect -1558 -9609 -1505 -9599
rect -312 -9609 -259 -9599
rect -136 -9608 -83 -9599
rect 42 -9609 95 -9599
rect 222 -9608 275 -9599
rect 399 -9609 452 -9599
rect 577 -9609 630 -9599
rect 2230 -9599 2357 -9548
rect 2409 -9599 2534 -9547
rect 2586 -9599 2713 -9547
rect 2765 -9599 4208 -9547
rect 4260 -9598 6679 -9547
rect 6731 -9598 6732 -9546
rect 4260 -9599 6732 -9598
rect 2230 -9600 2231 -9599
rect 2178 -9610 2231 -9600
rect 2357 -9609 2410 -9599
rect 2534 -9609 2587 -9599
rect 2713 -9609 2766 -9599
rect 4208 -9609 4261 -9599
rect 6679 -9608 6732 -9599
rect -2315 -9925 -2262 -9915
rect -1916 -9925 -1863 -9915
rect -1738 -9925 -1685 -9916
rect -1560 -9925 -1507 -9915
rect -1382 -9925 -1329 -9914
rect -314 -9925 -261 -9915
rect -136 -9925 -83 -9916
rect 43 -9925 96 -9915
rect 220 -9925 273 -9915
rect 398 -9925 451 -9915
rect 576 -9925 629 -9915
rect 2356 -9925 2409 -9915
rect 2534 -9925 2587 -9915
rect 2712 -9925 2765 -9916
rect 2891 -9925 2944 -9915
rect 3069 -9925 3122 -9915
rect 3246 -9925 3299 -9915
rect 5337 -9925 5390 -9915
rect -2315 -9926 -1382 -9925
rect -2263 -9978 -1916 -9926
rect -1864 -9927 -1560 -9926
rect -1864 -9978 -1738 -9927
rect -2315 -9988 -2262 -9978
rect -1916 -9988 -1863 -9978
rect -1686 -9978 -1560 -9927
rect -1508 -9977 -1382 -9926
rect -1330 -9926 5390 -9925
rect -1330 -9977 -314 -9926
rect -1508 -9978 -314 -9977
rect -262 -9927 43 -9926
rect -262 -9978 -136 -9927
rect -1686 -9979 -1685 -9978
rect -1738 -9989 -1685 -9979
rect -1560 -9988 -1507 -9978
rect -1382 -9987 -1329 -9978
rect -314 -9988 -261 -9978
rect -84 -9978 43 -9927
rect 95 -9978 220 -9926
rect 272 -9978 398 -9926
rect 450 -9978 576 -9926
rect 628 -9978 2356 -9926
rect 2408 -9978 2534 -9926
rect 2586 -9927 2891 -9926
rect 2586 -9978 2712 -9927
rect -84 -9979 -83 -9978
rect -136 -9989 -83 -9979
rect 43 -9988 96 -9978
rect 220 -9988 273 -9978
rect 398 -9988 451 -9978
rect 576 -9988 629 -9978
rect 2356 -9988 2409 -9978
rect 2534 -9988 2587 -9978
rect 2764 -9978 2891 -9927
rect 2943 -9978 3069 -9926
rect 3121 -9978 3246 -9926
rect 3298 -9978 5337 -9926
rect 5389 -9978 5390 -9926
rect 2764 -9979 2765 -9978
rect 2712 -9989 2765 -9979
rect 2891 -9988 2944 -9978
rect 3069 -9988 3122 -9978
rect 3246 -9988 3299 -9978
rect 5337 -9988 5390 -9978
rect 6680 -10313 6733 -10303
rect 9171 -10313 9224 -10304
rect 6680 -10314 9224 -10313
rect 6732 -10315 9224 -10314
rect 6732 -10366 9171 -10315
rect 6680 -10376 6733 -10366
rect 9223 -10367 9224 -10315
rect 9171 -10377 9224 -10367
rect 6858 -10466 6911 -10457
rect 7214 -10466 7267 -10456
rect 7571 -10466 7624 -10456
rect 7927 -10466 7980 -10456
rect 8283 -10466 8336 -10457
rect 8638 -10466 8691 -10456
rect 8995 -10466 9048 -10457
rect 6858 -10467 9048 -10466
rect 6858 -10468 7214 -10467
rect 6910 -10519 7214 -10468
rect 7266 -10519 7571 -10467
rect 7623 -10519 7927 -10467
rect 7979 -10468 8638 -10467
rect 7979 -10519 8283 -10468
rect 6910 -10520 6911 -10519
rect 6858 -10530 6911 -10520
rect 7214 -10529 7267 -10519
rect 7571 -10529 7624 -10519
rect 7927 -10529 7980 -10519
rect 8335 -10519 8638 -10468
rect 8690 -10468 9048 -10467
rect 8690 -10519 8995 -10468
rect 8335 -10520 8336 -10519
rect 8283 -10530 8336 -10520
rect 8638 -10529 8691 -10519
rect 9047 -10520 9048 -10468
rect 8995 -10530 9048 -10520
rect -1827 -10908 -1774 -10898
rect -1470 -10908 -1417 -10898
rect -1114 -10908 -1061 -10898
rect -758 -10908 -705 -10898
rect -402 -10908 -349 -10898
rect -46 -10908 7 -10898
rect 309 -10908 362 -10898
rect 665 -10908 718 -10898
rect 931 -10908 984 -10898
rect 1199 -10908 1252 -10898
rect 1556 -10908 1609 -10898
rect 1913 -10908 1966 -10898
rect 2268 -10908 2321 -10898
rect 2623 -10908 2676 -10898
rect 2980 -10908 3033 -10898
rect 3335 -10908 3388 -10898
rect 3692 -10908 3745 -10898
rect -1827 -10909 3745 -10908
rect -1775 -10961 -1470 -10909
rect -1418 -10961 -1114 -10909
rect -1062 -10961 -758 -10909
rect -706 -10961 -402 -10909
rect -350 -10961 -46 -10909
rect 6 -10961 309 -10909
rect 361 -10961 665 -10909
rect 717 -10961 931 -10909
rect 983 -10961 1199 -10909
rect 1251 -10961 1556 -10909
rect 1608 -10961 1913 -10909
rect 1965 -10961 2268 -10909
rect 2320 -10961 2623 -10909
rect 2675 -10961 2980 -10909
rect 3032 -10961 3335 -10909
rect 3387 -10961 3692 -10909
rect 3744 -10961 3745 -10909
rect -1827 -10971 -1774 -10961
rect -1470 -10971 -1417 -10961
rect -1114 -10971 -1061 -10961
rect -758 -10971 -705 -10961
rect -402 -10971 -349 -10961
rect -46 -10971 7 -10961
rect 309 -10971 362 -10961
rect 665 -10971 718 -10961
rect 931 -10971 984 -10961
rect 1199 -10971 1252 -10961
rect 1556 -10971 1609 -10961
rect 1913 -10971 1966 -10961
rect 2268 -10971 2321 -10961
rect 2623 -10971 2676 -10961
rect 2980 -10971 3033 -10961
rect 3335 -10971 3388 -10961
rect 3692 -10971 3745 -10961
rect 7037 -11366 7090 -11356
rect 7393 -11366 7446 -11356
rect 7748 -11366 7801 -11357
rect 8103 -11366 8156 -11356
rect 8461 -11366 8514 -11356
rect 8817 -11366 8870 -11356
rect 7037 -11367 8870 -11366
rect 7089 -11419 7393 -11367
rect 7445 -11368 8103 -11367
rect 7445 -11419 7748 -11368
rect 7037 -11429 7090 -11419
rect 7393 -11429 7446 -11419
rect 7800 -11419 8103 -11368
rect 8155 -11419 8461 -11367
rect 8513 -11419 8817 -11367
rect 8869 -11419 8870 -11367
rect 7800 -11420 7801 -11419
rect 7748 -11430 7801 -11420
rect 8103 -11429 8156 -11419
rect 8461 -11429 8514 -11419
rect 8817 -11429 8870 -11419
rect -1649 -11528 -1596 -11518
rect -1293 -11528 -1240 -11518
rect -937 -11528 -884 -11518
rect 1377 -11528 1430 -11518
rect 1733 -11528 1786 -11518
rect 2089 -11528 2142 -11518
rect -1649 -11529 2142 -11528
rect -1597 -11581 -1293 -11529
rect -1241 -11581 -937 -11529
rect -885 -11581 1377 -11529
rect 1429 -11581 1733 -11529
rect 1785 -11581 2089 -11529
rect 2141 -11581 2142 -11529
rect -1649 -11591 -1596 -11581
rect -1293 -11591 -1240 -11581
rect -937 -11591 -884 -11581
rect 1377 -11591 1430 -11581
rect 1733 -11591 1786 -11581
rect 2089 -11591 2142 -11581
rect -2004 -11637 -1951 -11627
rect -580 -11637 -527 -11627
rect 2446 -11637 2499 -11627
rect 3871 -11637 3924 -11628
rect -2004 -11638 3924 -11637
rect -1952 -11690 -580 -11638
rect -528 -11690 2446 -11638
rect 2498 -11639 3924 -11638
rect 2498 -11690 3871 -11639
rect -2004 -11700 -1951 -11690
rect -580 -11700 -527 -11690
rect 2446 -11700 2499 -11690
rect 3923 -11691 3924 -11639
rect 3871 -11701 3924 -11691
rect 11053 -11674 11106 -11664
rect 11347 -11674 11400 -11665
rect 11638 -11674 11691 -11664
rect 11931 -11674 11984 -11664
rect 12223 -11674 12276 -11664
rect 13022 -11674 13075 -11663
rect 11053 -11675 13022 -11674
rect 11105 -11676 11638 -11675
rect 11105 -11727 11347 -11676
rect 11053 -11737 11106 -11727
rect 11399 -11727 11638 -11676
rect 11690 -11727 11931 -11675
rect 11983 -11727 12223 -11675
rect 12275 -11726 13022 -11675
rect 13074 -11726 13075 -11674
rect 12275 -11727 13075 -11726
rect 11399 -11728 11400 -11727
rect 11347 -11738 11400 -11728
rect 11638 -11737 11691 -11727
rect 11931 -11737 11984 -11727
rect 12223 -11737 12276 -11727
rect 13022 -11736 13075 -11727
rect -224 -11757 -171 -11747
rect 131 -11757 184 -11747
rect 487 -11757 540 -11747
rect 2800 -11757 2853 -11747
rect 3157 -11757 3210 -11747
rect 3513 -11757 3566 -11747
rect -224 -11758 3566 -11757
rect -172 -11810 131 -11758
rect 183 -11810 487 -11758
rect 539 -11810 2800 -11758
rect 2852 -11810 3157 -11758
rect 3209 -11810 3513 -11758
rect 3565 -11810 3566 -11758
rect -224 -11820 -171 -11810
rect 131 -11820 184 -11810
rect 487 -11820 540 -11810
rect 2800 -11820 2853 -11810
rect 3157 -11820 3210 -11810
rect 3513 -11820 3566 -11810
rect -1915 -11919 -1862 -11909
rect -1738 -11919 -1685 -11909
rect -1559 -11919 -1506 -11909
rect -1381 -11919 -1328 -11909
rect -1203 -11919 -1150 -11909
rect -1025 -11919 -972 -11909
rect -848 -11919 -795 -11909
rect -670 -11919 -617 -11909
rect -492 -11919 -439 -11909
rect -314 -11919 -261 -11909
rect -136 -11919 -83 -11909
rect 42 -11919 95 -11909
rect 220 -11919 273 -11909
rect 399 -11919 452 -11909
rect 577 -11919 630 -11909
rect 1288 -11919 1341 -11909
rect 1468 -11919 1521 -11909
rect 1644 -11919 1697 -11910
rect 1823 -11919 1876 -11909
rect 2000 -11919 2053 -11909
rect 2178 -11919 2231 -11909
rect 2357 -11919 2410 -11909
rect 2534 -11919 2587 -11909
rect 2713 -11919 2766 -11909
rect 2890 -11919 2943 -11909
rect 3068 -11919 3121 -11909
rect 3247 -11919 3300 -11909
rect 3425 -11919 3478 -11909
rect 3603 -11919 3656 -11909
rect 3781 -11919 3834 -11909
rect -1915 -11920 3834 -11919
rect -1863 -11972 -1738 -11920
rect -1686 -11972 -1559 -11920
rect -1507 -11972 -1381 -11920
rect -1329 -11972 -1203 -11920
rect -1151 -11972 -1025 -11920
rect -973 -11972 -848 -11920
rect -796 -11972 -670 -11920
rect -618 -11972 -492 -11920
rect -440 -11972 -314 -11920
rect -262 -11972 -136 -11920
rect -84 -11972 42 -11920
rect 94 -11972 220 -11920
rect 272 -11972 399 -11920
rect 451 -11972 577 -11920
rect 629 -11972 1288 -11920
rect 1340 -11972 1468 -11920
rect 1520 -11921 1823 -11920
rect 1520 -11972 1644 -11921
rect -1915 -11982 -1862 -11972
rect -1738 -11982 -1685 -11972
rect -1559 -11982 -1506 -11972
rect -1381 -11982 -1328 -11972
rect -1203 -11982 -1150 -11972
rect -1025 -11982 -972 -11972
rect -848 -11982 -795 -11972
rect -670 -11982 -617 -11972
rect -492 -11982 -439 -11972
rect -314 -11982 -261 -11972
rect -136 -11982 -83 -11972
rect 42 -11982 95 -11972
rect 220 -11982 273 -11972
rect 399 -11982 452 -11972
rect 577 -11982 630 -11972
rect 1288 -11982 1341 -11972
rect 1468 -11982 1521 -11972
rect 1696 -11972 1823 -11921
rect 1875 -11972 2000 -11920
rect 2052 -11972 2178 -11920
rect 2230 -11972 2357 -11920
rect 2409 -11972 2534 -11920
rect 2586 -11972 2713 -11920
rect 2765 -11972 2890 -11920
rect 2942 -11972 3068 -11920
rect 3120 -11972 3247 -11920
rect 3299 -11972 3425 -11920
rect 3477 -11972 3603 -11920
rect 3655 -11972 3781 -11920
rect 3833 -11972 3834 -11920
rect 1696 -11973 1697 -11972
rect 1644 -11983 1697 -11973
rect 1823 -11982 1876 -11972
rect 2000 -11982 2053 -11972
rect 2178 -11982 2231 -11972
rect 2357 -11982 2410 -11972
rect 2534 -11982 2587 -11972
rect 2713 -11982 2766 -11972
rect 2890 -11982 2943 -11972
rect 3068 -11982 3121 -11972
rect 3247 -11982 3300 -11972
rect 3425 -11982 3478 -11972
rect 3603 -11982 3656 -11972
rect 3781 -11982 3834 -11972
rect -5502 -12271 -5449 -12261
rect -5000 -12271 -4947 -12262
rect -4502 -12271 -4449 -12261
rect -5502 -12272 -4449 -12271
rect -2447 -12272 -2394 -12262
rect -5450 -12273 -4502 -12272
rect -5450 -12324 -5000 -12273
rect -5502 -12334 -5449 -12324
rect -4948 -12324 -4502 -12273
rect -4450 -12273 -2394 -12272
rect -4450 -12324 -2447 -12273
rect -4948 -12325 -4947 -12324
rect -5000 -12335 -4947 -12325
rect -4502 -12325 -2447 -12324
rect -2395 -12325 -2394 -12273
rect -4502 -12334 -4449 -12325
rect -2447 -12335 -2394 -12325
rect -5376 -12388 -5323 -12378
rect -5127 -12388 -5074 -12378
rect -4377 -12388 -4324 -12378
rect -3928 -12388 -3875 -12379
rect -5376 -12389 -3875 -12388
rect -5324 -12441 -5127 -12389
rect -5075 -12441 -4377 -12389
rect -4325 -12390 -3875 -12389
rect -4325 -12441 -3928 -12390
rect -5376 -12451 -5323 -12441
rect -5127 -12451 -5074 -12441
rect -4377 -12451 -4324 -12441
rect -3876 -12442 -3875 -12390
rect -3928 -12452 -3875 -12442
rect -6077 -12512 -6024 -12502
rect -5626 -12512 -5573 -12502
rect -4877 -12512 -4824 -12502
rect -4627 -12512 -4574 -12502
rect -6077 -12513 -4574 -12512
rect -6025 -12565 -5626 -12513
rect -5574 -12565 -4877 -12513
rect -4825 -12565 -4627 -12513
rect -4575 -12565 -4574 -12513
rect -6077 -12575 -6024 -12565
rect -5626 -12575 -5573 -12565
rect -4877 -12575 -4824 -12565
rect -4627 -12575 -4574 -12565
rect -2005 -12542 -1952 -12532
rect -1649 -12542 -1596 -12532
rect 3514 -12542 3567 -12532
rect 3871 -12542 3924 -12532
rect -2005 -12543 -1284 -12542
rect -1953 -12595 -1649 -12543
rect -1597 -12544 -1284 -12543
rect -1250 -12543 3924 -12542
rect -1250 -12544 3514 -12543
rect -1597 -12595 3514 -12544
rect 3566 -12595 3871 -12543
rect 3923 -12595 3924 -12543
rect -2005 -12605 -1952 -12595
rect -1649 -12605 -1596 -12595
rect 3514 -12605 3567 -12595
rect 3871 -12605 3924 -12595
rect -1294 -12653 -1241 -12644
rect -582 -12653 -529 -12643
rect 130 -12653 183 -12643
rect 1735 -12653 1788 -12644
rect 2445 -12653 2498 -12643
rect 3158 -12653 3211 -12642
rect -1294 -12654 3158 -12653
rect -1294 -12655 -582 -12654
rect -1242 -12706 -582 -12655
rect -530 -12706 130 -12654
rect 182 -12655 2445 -12654
rect 182 -12706 1735 -12655
rect -1242 -12707 -1241 -12706
rect -1294 -12717 -1241 -12707
rect -582 -12716 -529 -12706
rect 130 -12716 183 -12706
rect 1787 -12706 2445 -12655
rect 2497 -12705 3158 -12654
rect 3210 -12705 3211 -12653
rect 2497 -12706 3211 -12705
rect 1787 -12707 1788 -12706
rect 1735 -12717 1788 -12707
rect 2445 -12716 2498 -12706
rect 3158 -12715 3211 -12706
rect -937 -12783 -884 -12773
rect -224 -12783 -171 -12773
rect 486 -12783 539 -12774
rect 1378 -12783 1431 -12773
rect 2088 -12783 2141 -12772
rect 2801 -12783 2854 -12772
rect -937 -12784 2088 -12783
rect -885 -12836 -224 -12784
rect -172 -12785 1378 -12784
rect -172 -12836 486 -12785
rect -937 -12846 -884 -12836
rect -224 -12846 -171 -12836
rect 538 -12836 1378 -12785
rect 1430 -12835 2088 -12784
rect 2140 -12835 2801 -12783
rect 2853 -12835 2854 -12783
rect 1430 -12836 2854 -12835
rect 538 -12837 539 -12836
rect 486 -12847 539 -12837
rect 1378 -12846 1431 -12836
rect 2088 -12845 2141 -12836
rect 2801 -12845 2854 -12836
rect -6223 -13062 -6170 -13052
rect -5751 -13062 -5698 -13052
rect -4752 -13062 -4699 -13052
rect -6223 -13063 -4699 -13062
rect -6171 -13115 -5751 -13063
rect -5699 -13115 -4752 -13063
rect -4700 -13115 -4699 -13063
rect -6223 -13125 -6170 -13115
rect -5751 -13125 -5698 -13115
rect -4752 -13125 -4699 -13115
rect -5251 -13189 -5198 -13179
rect -4251 -13189 -4198 -13179
rect -3788 -13189 -3735 -13179
rect -3542 -13189 -3489 -13179
rect -5251 -13190 -3489 -13189
rect -5199 -13242 -4251 -13190
rect -4199 -13242 -3788 -13190
rect -3736 -13242 -3542 -13190
rect -3490 -13242 -3489 -13190
rect -5251 -13252 -5198 -13242
rect -4251 -13252 -4198 -13242
rect -3788 -13252 -3735 -13242
rect -3542 -13252 -3489 -13242
rect 5037 -13296 5090 -13286
rect 5534 -13296 5587 -13286
rect 5037 -13297 5587 -13296
rect 5089 -13349 5534 -13297
rect 5586 -13349 5587 -13297
rect 5037 -13359 5090 -13349
rect 5534 -13359 5587 -13349
rect 5031 -13433 5084 -13423
rect 8950 -13433 9003 -13423
rect 9305 -13433 9358 -13423
rect 18337 -13433 18412 -13411
rect 5031 -13434 18348 -13433
rect 5083 -13486 8950 -13434
rect 9002 -13486 9305 -13434
rect 9357 -13485 18348 -13434
rect 18400 -13485 18422 -13433
rect 9357 -13486 18422 -13485
rect 5031 -13496 5084 -13486
rect 8950 -13496 9003 -13486
rect 9305 -13496 9358 -13486
rect 18337 -13506 18412 -13486
rect -2004 -13545 -1951 -13535
rect -581 -13545 -528 -13535
rect 2446 -13545 2499 -13535
rect 3870 -13545 3923 -13535
rect 5400 -13545 5453 -13535
rect -2004 -13546 8828 -13545
rect -1952 -13598 -581 -13546
rect -529 -13598 2446 -13546
rect 2498 -13598 3870 -13546
rect 3922 -13598 5400 -13546
rect 5452 -13556 8828 -13546
rect 9127 -13556 9180 -13546
rect 9483 -13556 9536 -13546
rect 5452 -13557 9536 -13556
rect 5452 -13598 8772 -13557
rect -2004 -13608 -1951 -13598
rect -581 -13608 -528 -13598
rect 2446 -13608 2499 -13598
rect 3870 -13608 3923 -13598
rect 5400 -13608 5453 -13598
rect 8824 -13609 9127 -13557
rect 9179 -13609 9483 -13557
rect 9535 -13609 9536 -13557
rect 8772 -13619 8825 -13609
rect 9127 -13619 9180 -13609
rect 9483 -13619 9536 -13609
rect -1648 -13672 -1595 -13662
rect -1291 -13672 -1238 -13662
rect -937 -13672 -884 -13662
rect 1379 -13672 1432 -13662
rect 1732 -13672 1785 -13662
rect 2091 -13672 2144 -13662
rect 5534 -13672 5587 -13662
rect 7526 -13672 7579 -13662
rect 7882 -13672 7935 -13663
rect 8238 -13672 8291 -13661
rect 11442 -13672 11495 -13662
rect 11798 -13672 11851 -13662
rect 12152 -13672 12205 -13663
rect 12509 -13672 12562 -13662
rect -1648 -13673 5323 -13672
rect -1596 -13725 -1291 -13673
rect -1239 -13725 -937 -13673
rect -885 -13725 1379 -13673
rect 1431 -13725 1732 -13673
rect 1784 -13725 2091 -13673
rect 2143 -13725 5323 -13673
rect -1648 -13735 -1595 -13725
rect -1291 -13735 -1238 -13725
rect -937 -13735 -884 -13725
rect 1379 -13735 1432 -13725
rect 1732 -13735 1785 -13725
rect 2091 -13735 2144 -13725
rect -6077 -13745 -6024 -13735
rect -5376 -13745 -5323 -13735
rect -5126 -13745 -5073 -13735
rect -4376 -13745 -4323 -13735
rect -6077 -13746 -4323 -13745
rect -6025 -13798 -5376 -13746
rect -5324 -13798 -5126 -13746
rect -5074 -13798 -4376 -13746
rect -4324 -13798 -4323 -13746
rect -6077 -13808 -6024 -13798
rect -5376 -13808 -5323 -13798
rect -5126 -13808 -5073 -13798
rect -4376 -13808 -4323 -13798
rect -225 -13794 -172 -13784
rect 133 -13794 186 -13784
rect 487 -13794 540 -13785
rect 2802 -13794 2855 -13784
rect 3157 -13794 3210 -13785
rect 3512 -13794 3565 -13784
rect 5142 -13794 5195 -13784
rect -225 -13795 5195 -13794
rect -6426 -13852 -6373 -13842
rect -5626 -13852 -5573 -13842
rect -4877 -13852 -4824 -13842
rect -4627 -13852 -4574 -13842
rect -3928 -13852 -3875 -13842
rect -6426 -13853 -3875 -13852
rect -6374 -13905 -5626 -13853
rect -5574 -13905 -4877 -13853
rect -4825 -13905 -4627 -13853
rect -4575 -13905 -3928 -13853
rect -3876 -13905 -3875 -13853
rect -173 -13847 133 -13795
rect 185 -13796 2802 -13795
rect 185 -13847 487 -13796
rect -225 -13857 -172 -13847
rect 133 -13857 186 -13847
rect 539 -13847 2802 -13796
rect 2854 -13796 3512 -13795
rect 2854 -13847 3157 -13796
rect 539 -13848 540 -13847
rect 487 -13858 540 -13848
rect 2802 -13857 2855 -13847
rect 3209 -13847 3512 -13796
rect 3564 -13847 5142 -13795
rect 5194 -13847 5195 -13795
rect 3209 -13848 3210 -13847
rect 3157 -13858 3210 -13848
rect 3512 -13857 3565 -13847
rect 5142 -13857 5195 -13847
rect 5270 -13796 5323 -13725
rect 5534 -13673 8238 -13672
rect 5586 -13725 7526 -13673
rect 7578 -13674 8238 -13673
rect 7578 -13725 7882 -13674
rect 5534 -13735 5587 -13725
rect 7526 -13735 7579 -13725
rect 7934 -13724 8238 -13674
rect 8290 -13673 12562 -13672
rect 8290 -13724 11442 -13673
rect 7934 -13725 11442 -13724
rect 11494 -13725 11798 -13673
rect 11850 -13674 12509 -13673
rect 11850 -13725 12152 -13674
rect 7934 -13726 7935 -13725
rect 7882 -13736 7935 -13726
rect 8238 -13734 8291 -13725
rect 11442 -13735 11495 -13725
rect 11798 -13735 11851 -13725
rect 12204 -13725 12509 -13674
rect 12561 -13725 12562 -13673
rect 12204 -13726 12205 -13725
rect 12152 -13736 12205 -13726
rect 12509 -13735 12562 -13725
rect 7348 -13796 7401 -13786
rect 7704 -13796 7757 -13785
rect 8061 -13796 8114 -13786
rect 8415 -13796 8468 -13786
rect 11264 -13796 11317 -13786
rect 11620 -13796 11673 -13787
rect 11977 -13796 12030 -13786
rect 12334 -13796 12387 -13786
rect 5270 -13797 7704 -13796
rect 5270 -13849 7348 -13797
rect 7400 -13848 7704 -13797
rect 7756 -13797 12387 -13796
rect 7756 -13848 8061 -13797
rect 7400 -13849 8061 -13848
rect 8113 -13849 8415 -13797
rect 8467 -13849 11264 -13797
rect 11316 -13798 11977 -13797
rect 11316 -13849 11620 -13798
rect 7348 -13859 7401 -13849
rect 7704 -13858 7757 -13849
rect 8061 -13859 8114 -13849
rect 8415 -13859 8468 -13849
rect 11264 -13859 11317 -13849
rect 11672 -13849 11977 -13798
rect 12029 -13849 12334 -13797
rect 12386 -13849 12387 -13797
rect 11672 -13850 11673 -13849
rect 11620 -13860 11673 -13850
rect 11977 -13859 12030 -13849
rect 12334 -13859 12387 -13849
rect -6426 -13915 -6373 -13905
rect -5626 -13915 -5573 -13905
rect -4877 -13915 -4824 -13905
rect -4627 -13915 -4574 -13905
rect -3928 -13915 -3875 -13905
rect 5833 -13922 5886 -13912
rect 6013 -13922 6066 -13912
rect 6190 -13922 6243 -13913
rect 6369 -13922 6422 -13912
rect 6547 -13922 6600 -13913
rect 6725 -13922 6778 -13912
rect 6902 -13922 6955 -13912
rect 7437 -13922 7490 -13912
rect 7615 -13922 7668 -13912
rect 7793 -13922 7846 -13913
rect 7970 -13922 8023 -13912
rect 8148 -13922 8201 -13912
rect 8326 -13922 8379 -13912
rect 8861 -13922 8914 -13912
rect 9038 -13922 9091 -13912
rect 9217 -13922 9270 -13912
rect 9394 -13922 9447 -13912
rect 9929 -13922 9982 -13913
rect 10108 -13922 10161 -13912
rect 10284 -13922 10337 -13913
rect 10462 -13922 10515 -13913
rect 10640 -13922 10693 -13912
rect 10819 -13922 10872 -13913
rect 11353 -13922 11406 -13912
rect 11530 -13922 11583 -13912
rect 11709 -13922 11762 -13912
rect 11886 -13922 11939 -13913
rect 12064 -13922 12117 -13912
rect 12242 -13922 12295 -13913
rect 12420 -13922 12473 -13912
rect 5833 -13923 12473 -13922
rect -5730 -13957 -5677 -13947
rect -4752 -13957 -4699 -13947
rect -3788 -13957 -3735 -13947
rect -5730 -13958 -3735 -13957
rect -5678 -14010 -4752 -13958
rect -4700 -14010 -3788 -13958
rect -3736 -14010 -3735 -13958
rect 5885 -13975 6013 -13923
rect 6065 -13924 6369 -13923
rect 6065 -13975 6190 -13924
rect 5833 -13985 5886 -13975
rect 6013 -13985 6066 -13975
rect 6242 -13975 6369 -13924
rect 6421 -13924 6725 -13923
rect 6421 -13975 6547 -13924
rect 6242 -13976 6243 -13975
rect 6190 -13986 6243 -13976
rect 6369 -13985 6422 -13975
rect 6599 -13975 6725 -13924
rect 6777 -13975 6902 -13923
rect 6954 -13975 7437 -13923
rect 7489 -13975 7615 -13923
rect 7667 -13924 7970 -13923
rect 7667 -13975 7793 -13924
rect 6599 -13976 6600 -13975
rect 6547 -13986 6600 -13976
rect 6725 -13985 6778 -13975
rect 6902 -13985 6955 -13975
rect 7437 -13985 7490 -13975
rect 7615 -13985 7668 -13975
rect 7845 -13975 7970 -13924
rect 8022 -13975 8148 -13923
rect 8200 -13975 8326 -13923
rect 8378 -13975 8861 -13923
rect 8913 -13975 9038 -13923
rect 9090 -13975 9217 -13923
rect 9269 -13975 9394 -13923
rect 9446 -13924 10108 -13923
rect 9446 -13975 9929 -13924
rect 7845 -13976 7846 -13975
rect 7793 -13986 7846 -13976
rect 7970 -13985 8023 -13975
rect 8148 -13985 8201 -13975
rect 8326 -13985 8379 -13975
rect 8861 -13985 8914 -13975
rect 9038 -13985 9091 -13975
rect 9217 -13985 9270 -13975
rect 9394 -13985 9447 -13975
rect 9981 -13975 10108 -13924
rect 10160 -13924 10640 -13923
rect 10160 -13975 10284 -13924
rect 9981 -13976 9982 -13975
rect 9929 -13986 9982 -13976
rect 10108 -13985 10161 -13975
rect 10336 -13975 10462 -13924
rect 10336 -13976 10337 -13975
rect 10284 -13986 10337 -13976
rect 10514 -13975 10640 -13924
rect 10692 -13924 11353 -13923
rect 10692 -13975 10819 -13924
rect 10514 -13976 10515 -13975
rect 10462 -13986 10515 -13976
rect 10640 -13985 10693 -13975
rect 10871 -13975 11353 -13924
rect 11405 -13975 11530 -13923
rect 11582 -13975 11709 -13923
rect 11761 -13924 12064 -13923
rect 11761 -13975 11886 -13924
rect 10871 -13976 10872 -13975
rect 10819 -13986 10872 -13976
rect 11353 -13985 11406 -13975
rect 11530 -13985 11583 -13975
rect 11709 -13985 11762 -13975
rect 11938 -13975 12064 -13924
rect 12116 -13924 12420 -13923
rect 12116 -13975 12242 -13924
rect 11938 -13976 11939 -13975
rect 11886 -13986 11939 -13976
rect 12064 -13985 12117 -13975
rect 12294 -13975 12420 -13924
rect 12472 -13975 12473 -13923
rect 12294 -13976 12295 -13975
rect 12242 -13986 12295 -13976
rect 12420 -13985 12473 -13975
rect -5730 -14020 -5677 -14010
rect -4752 -14020 -4699 -14010
rect -3788 -14020 -3735 -14010
rect -6223 -14055 -6170 -14045
rect -5250 -14055 -5197 -14045
rect -4250 -14055 -4197 -14045
rect -3382 -14055 -3329 -14045
rect -6223 -14056 -3329 -14055
rect -6171 -14108 -5250 -14056
rect -5198 -14108 -4250 -14056
rect -4198 -14108 -3382 -14056
rect -3330 -14108 -3329 -14056
rect -6223 -14118 -6170 -14108
rect -5250 -14118 -5197 -14108
rect -4250 -14118 -4197 -14108
rect -3382 -14118 -3329 -14108
rect -2315 -14543 -2262 -14533
rect -1381 -14543 -1328 -14533
rect -1204 -14543 -1151 -14533
rect -1026 -14543 -973 -14533
rect -848 -14543 -795 -14533
rect -669 -14543 -616 -14533
rect -491 -14543 -438 -14533
rect 1288 -14543 1341 -14533
rect 1466 -14543 1519 -14533
rect 1644 -14543 1697 -14533
rect 1823 -14543 1876 -14532
rect 2000 -14543 2053 -14533
rect 2178 -14543 2231 -14533
rect 3246 -14543 3299 -14534
rect 3424 -14543 3477 -14533
rect 3602 -14543 3655 -14533
rect 3781 -14543 3834 -14533
rect -2315 -14544 1823 -14543
rect -2263 -14596 -1381 -14544
rect -1329 -14596 -1204 -14544
rect -1152 -14596 -1026 -14544
rect -974 -14596 -848 -14544
rect -796 -14596 -669 -14544
rect -617 -14596 -491 -14544
rect -439 -14596 1288 -14544
rect 1340 -14596 1466 -14544
rect 1518 -14596 1644 -14544
rect 1696 -14595 1823 -14544
rect 1875 -14544 3834 -14543
rect 1875 -14595 2000 -14544
rect 1696 -14596 2000 -14595
rect 2052 -14596 2178 -14544
rect 2230 -14545 3424 -14544
rect 2230 -14596 3246 -14545
rect -2315 -14606 -2262 -14596
rect -1381 -14606 -1328 -14596
rect -1204 -14606 -1151 -14596
rect -1026 -14606 -973 -14596
rect -848 -14606 -795 -14596
rect -669 -14606 -616 -14596
rect -491 -14606 -438 -14596
rect 1288 -14606 1341 -14596
rect 1466 -14606 1519 -14596
rect 1644 -14606 1697 -14596
rect 1823 -14605 1876 -14596
rect 2000 -14606 2053 -14596
rect 2178 -14606 2231 -14596
rect 3298 -14596 3424 -14545
rect 3476 -14596 3602 -14544
rect 3654 -14596 3781 -14544
rect 3833 -14596 3834 -14544
rect 3298 -14597 3299 -14596
rect 3246 -14607 3299 -14597
rect 3424 -14606 3477 -14596
rect 3602 -14606 3655 -14596
rect 3781 -14606 3834 -14596
rect 4905 -14545 4958 -14535
rect 5746 -14545 5799 -14535
rect 6101 -14545 6154 -14535
rect 6459 -14545 6512 -14535
rect 6813 -14545 6866 -14535
rect 8236 -14545 8289 -14535
rect 8595 -14545 8648 -14535
rect 8950 -14545 9003 -14536
rect 9304 -14545 9357 -14535
rect 9661 -14545 9714 -14535
rect 10016 -14545 10069 -14535
rect 10373 -14545 10426 -14536
rect 10729 -14545 10782 -14535
rect 4905 -14546 10782 -14545
rect 4957 -14598 5746 -14546
rect 5798 -14598 6101 -14546
rect 6153 -14598 6459 -14546
rect 6511 -14598 6813 -14546
rect 6865 -14598 8236 -14546
rect 8288 -14598 8595 -14546
rect 8647 -14547 9304 -14546
rect 8647 -14598 8950 -14547
rect 4905 -14608 4958 -14598
rect 5746 -14608 5799 -14598
rect 6101 -14608 6154 -14598
rect 6459 -14608 6512 -14598
rect 6813 -14608 6866 -14598
rect 8236 -14608 8289 -14598
rect 8595 -14608 8648 -14598
rect 9002 -14598 9304 -14547
rect 9356 -14598 9661 -14546
rect 9713 -14598 10016 -14546
rect 10068 -14547 10729 -14546
rect 10068 -14598 10373 -14547
rect 9002 -14599 9003 -14598
rect 8950 -14609 9003 -14599
rect 9304 -14608 9357 -14598
rect 9661 -14608 9714 -14598
rect 10016 -14608 10069 -14598
rect 10425 -14598 10729 -14547
rect 10781 -14598 10782 -14546
rect 10425 -14599 10426 -14598
rect 10373 -14609 10426 -14599
rect 10729 -14608 10782 -14598
rect 5143 -14658 5196 -14648
rect 5924 -14658 5977 -14648
rect 6279 -14658 6332 -14648
rect 6636 -14658 6689 -14648
rect 6991 -14658 7044 -14648
rect 8417 -14658 8470 -14647
rect 8772 -14658 8825 -14648
rect 9127 -14658 9180 -14649
rect 9483 -14658 9536 -14648
rect 9837 -14658 9890 -14649
rect 10196 -14658 10249 -14648
rect 10550 -14658 10603 -14648
rect 10908 -14658 10961 -14648
rect 5143 -14659 8417 -14658
rect 5195 -14711 5924 -14659
rect 5976 -14711 6279 -14659
rect 6331 -14711 6636 -14659
rect 6688 -14711 6991 -14659
rect 7043 -14710 8417 -14659
rect 8469 -14659 10961 -14658
rect 8469 -14710 8772 -14659
rect 7043 -14711 8772 -14710
rect 8824 -14660 9483 -14659
rect 8824 -14711 9127 -14660
rect 5143 -14721 5196 -14711
rect 5924 -14721 5977 -14711
rect 6279 -14721 6332 -14711
rect 6636 -14721 6689 -14711
rect 6991 -14721 7044 -14711
rect 8417 -14720 8470 -14711
rect 8772 -14721 8825 -14711
rect 9179 -14711 9483 -14660
rect 9535 -14660 10196 -14659
rect 9535 -14711 9837 -14660
rect 9179 -14712 9180 -14711
rect 9127 -14722 9180 -14712
rect 9483 -14721 9536 -14711
rect 9889 -14711 10196 -14660
rect 10248 -14711 10550 -14659
rect 10602 -14711 10908 -14659
rect 10960 -14711 10961 -14659
rect 9889 -14712 9890 -14711
rect 9837 -14722 9890 -14712
rect 10196 -14721 10249 -14711
rect 10550 -14721 10603 -14711
rect 10908 -14721 10961 -14711
rect 11087 -14656 11140 -14648
rect 11440 -14656 11493 -14646
rect 11087 -14657 11493 -14656
rect 11087 -14659 11440 -14657
rect 11139 -14708 11440 -14659
rect 11139 -14709 11192 -14708
rect 11492 -14709 11493 -14657
rect 11139 -14711 11140 -14709
rect 11087 -14721 11140 -14711
rect 11440 -14719 11493 -14709
rect -6159 -14795 -6106 -14785
rect -5860 -14795 -5807 -14785
rect -5147 -14795 -5094 -14785
rect -4436 -14795 -4383 -14785
rect -6159 -14796 -4383 -14795
rect -6107 -14848 -5860 -14796
rect -5808 -14848 -5147 -14796
rect -5095 -14848 -4436 -14796
rect -4384 -14848 -4383 -14796
rect 8504 -14807 8557 -14796
rect -6159 -14858 -6106 -14848
rect -5860 -14858 -5807 -14848
rect -5147 -14858 -5094 -14848
rect -4436 -14858 -4383 -14848
rect 6993 -14824 7046 -14814
rect 7347 -14824 7400 -14814
rect 7704 -14824 7757 -14815
rect 6993 -14825 7757 -14824
rect 7045 -14877 7347 -14825
rect 7399 -14826 7757 -14825
rect 7399 -14877 7704 -14826
rect 6993 -14887 7046 -14877
rect 7347 -14887 7400 -14877
rect 7756 -14878 7757 -14826
rect 7704 -14888 7757 -14878
rect 8060 -14821 8113 -14811
rect 8060 -14822 8504 -14821
rect 8112 -14859 8504 -14822
rect 8556 -14821 8557 -14807
rect 9753 -14807 9806 -14796
rect 8556 -14859 9753 -14821
rect 9805 -14821 9806 -14807
rect 10195 -14821 10248 -14812
rect 9805 -14823 10248 -14821
rect 9805 -14859 10195 -14823
rect 8112 -14874 10195 -14859
rect 8060 -14884 8113 -14874
rect 10247 -14875 10248 -14823
rect 10195 -14885 10248 -14875
rect 10552 -14814 10605 -14805
rect 10908 -14813 10961 -14803
rect 10908 -14814 11013 -14813
rect 11264 -14814 11317 -14805
rect 10552 -14816 10908 -14814
rect 10604 -14866 10908 -14816
rect 10960 -14816 11317 -14814
rect 10960 -14866 11264 -14816
rect 10604 -14868 10605 -14866
rect 10552 -14878 10605 -14868
rect 10908 -14876 10961 -14866
rect 11316 -14868 11317 -14816
rect 11264 -14878 11317 -14868
rect -5504 -14901 -5451 -14891
rect -4791 -14901 -4738 -14891
rect -3936 -14901 -3883 -14891
rect -5504 -14902 -3883 -14901
rect -5452 -14954 -4791 -14902
rect -4739 -14954 -3936 -14902
rect -3884 -14954 -3883 -14902
rect -5504 -14964 -5451 -14954
rect -4791 -14964 -4738 -14954
rect -3936 -14964 -3883 -14954
rect -847 -14926 -794 -14916
rect -669 -14926 -616 -14916
rect -491 -14926 -438 -14916
rect -314 -14926 -261 -14917
rect -137 -14926 -84 -14916
rect 43 -14926 96 -14916
rect 1289 -14926 1342 -14917
rect 1467 -14926 1520 -14916
rect 1644 -14926 1697 -14916
rect 1822 -14926 1875 -14916
rect 1999 -14926 2052 -14916
rect 2180 -14926 2233 -14916
rect 3425 -14926 3478 -14916
rect 3603 -14926 3656 -14916
rect 3780 -14926 3833 -14916
rect 4239 -14926 4292 -14916
rect -847 -14927 4292 -14926
rect -795 -14979 -669 -14927
rect -617 -14979 -491 -14927
rect -439 -14928 -137 -14927
rect -439 -14979 -314 -14928
rect -847 -14989 -794 -14979
rect -669 -14989 -616 -14979
rect -491 -14989 -438 -14979
rect -262 -14979 -137 -14928
rect -85 -14979 43 -14927
rect 95 -14928 1467 -14927
rect 95 -14979 1289 -14928
rect -262 -14980 -261 -14979
rect -314 -14990 -261 -14980
rect -137 -14989 -84 -14979
rect 43 -14989 96 -14979
rect 1341 -14979 1467 -14928
rect 1519 -14979 1644 -14927
rect 1696 -14979 1822 -14927
rect 1874 -14979 1999 -14927
rect 2051 -14979 2180 -14927
rect 2232 -14979 3425 -14927
rect 3477 -14979 3603 -14927
rect 3655 -14979 3780 -14927
rect 3832 -14979 4239 -14927
rect 4291 -14979 4292 -14927
rect 1341 -14980 1342 -14979
rect 1289 -14990 1342 -14980
rect 1467 -14989 1520 -14979
rect 1644 -14989 1697 -14979
rect 1822 -14989 1875 -14979
rect 1999 -14989 2052 -14979
rect 2180 -14989 2233 -14979
rect 3425 -14989 3478 -14979
rect 3603 -14989 3656 -14979
rect 3780 -14989 3833 -14979
rect 4239 -14989 4292 -14979
rect 7080 -14923 7133 -14913
rect 7260 -14923 7313 -14914
rect 7439 -14923 7492 -14913
rect 8327 -14923 8380 -14913
rect 8505 -14923 8558 -14914
rect 8683 -14923 8736 -14914
rect 9572 -14923 9625 -14913
rect 9750 -14923 9803 -14913
rect 9929 -14923 9982 -14913
rect 10819 -14923 10872 -14913
rect 10996 -14923 11049 -14913
rect 11175 -14923 11228 -14913
rect 7080 -14924 11228 -14923
rect 7132 -14925 7439 -14924
rect 7132 -14976 7260 -14925
rect 7080 -14986 7133 -14976
rect 7312 -14976 7439 -14925
rect 7491 -14976 8327 -14924
rect 8379 -14925 9572 -14924
rect 8379 -14976 8505 -14925
rect 7312 -14977 7313 -14976
rect 7260 -14987 7313 -14977
rect 7439 -14986 7492 -14976
rect 8327 -14986 8380 -14976
rect 8557 -14976 8683 -14925
rect 8557 -14977 8558 -14976
rect 8505 -14987 8558 -14977
rect 8735 -14976 9572 -14925
rect 9624 -14976 9750 -14924
rect 9802 -14976 9929 -14924
rect 9981 -14976 10819 -14924
rect 10871 -14976 10996 -14924
rect 11048 -14976 11175 -14924
rect 11227 -14976 11228 -14924
rect 8735 -14977 8736 -14976
rect 8683 -14987 8736 -14977
rect 9572 -14986 9625 -14976
rect 9750 -14986 9803 -14976
rect 9929 -14986 9982 -14976
rect 10819 -14986 10872 -14976
rect 10996 -14986 11049 -14976
rect 11175 -14986 11228 -14976
rect -6159 -15481 -6106 -15472
rect -5504 -15481 -5451 -15471
rect -4792 -15481 -4739 -15471
rect -6159 -15482 -4739 -15481
rect -6159 -15483 -5504 -15482
rect -6107 -15534 -5504 -15483
rect -5452 -15534 -4792 -15482
rect -4740 -15534 -4739 -15482
rect -6107 -15535 -6106 -15534
rect -6159 -15545 -6106 -15535
rect -5504 -15544 -5451 -15534
rect -4792 -15544 -4739 -15534
rect 4238 -15539 4291 -15529
rect 5031 -15539 5084 -15530
rect 5745 -15539 5798 -15529
rect 6101 -15539 6154 -15529
rect 6458 -15539 6511 -15529
rect 11798 -15539 11851 -15530
rect 12155 -15539 12208 -15529
rect 12511 -15539 12564 -15529
rect 4238 -15540 12564 -15539
rect -5860 -15589 -5807 -15578
rect -5148 -15589 -5095 -15579
rect -4435 -15589 -4383 -15579
rect -3935 -15589 -3883 -15579
rect -5808 -15590 -4435 -15589
rect -5808 -15641 -5148 -15590
rect -5860 -15651 -5807 -15641
rect -5096 -15641 -4435 -15590
rect -4383 -15641 -3935 -15589
rect 4290 -15541 5745 -15540
rect 4290 -15592 5031 -15541
rect 4238 -15602 4291 -15592
rect 5083 -15592 5745 -15541
rect 5797 -15592 6101 -15540
rect 6153 -15592 6458 -15540
rect 6510 -15541 12155 -15540
rect 6510 -15592 11798 -15541
rect 5083 -15593 5084 -15592
rect 5031 -15603 5084 -15593
rect 5745 -15602 5798 -15592
rect 6101 -15602 6154 -15592
rect 6458 -15602 6511 -15592
rect 11850 -15592 12155 -15541
rect 12207 -15592 12511 -15540
rect 12563 -15592 12564 -15540
rect 11850 -15593 11851 -15592
rect 11798 -15603 11851 -15593
rect 12155 -15602 12208 -15592
rect 12511 -15602 12564 -15592
rect -5096 -15642 -5095 -15641
rect -5148 -15652 -5095 -15642
rect -4435 -15651 -4383 -15641
rect -3935 -15651 -3883 -15641
rect 5400 -15652 5453 -15643
rect 5923 -15652 5976 -15642
rect 6279 -15652 6332 -15642
rect 6635 -15652 6688 -15642
rect 11619 -15652 11672 -15642
rect 11975 -15652 12028 -15642
rect 12332 -15652 12385 -15642
rect 5400 -15653 12385 -15652
rect 5400 -15654 5923 -15653
rect 5452 -15705 5923 -15654
rect 5975 -15705 6279 -15653
rect 6331 -15705 6635 -15653
rect 6687 -15705 11619 -15653
rect 11671 -15705 11975 -15653
rect 12027 -15705 12332 -15653
rect 12384 -15705 12385 -15653
rect 5452 -15706 5453 -15705
rect 5400 -15716 5453 -15706
rect 5923 -15715 5976 -15705
rect 6279 -15715 6332 -15705
rect 6635 -15715 6688 -15705
rect 11619 -15715 11672 -15705
rect 11975 -15715 12028 -15705
rect 12332 -15715 12385 -15705
rect 5747 -15750 5800 -15740
rect 6101 -15750 6154 -15739
rect 6456 -15750 6509 -15740
rect 6713 -15750 6766 -15741
rect 7169 -15750 7222 -15740
rect 7526 -15750 7579 -15739
rect 7882 -15750 7935 -15739
rect 10373 -15750 10426 -15741
rect 10730 -15750 10783 -15740
rect 11086 -15750 11139 -15740
rect 5747 -15751 6101 -15750
rect 5799 -15802 6101 -15751
rect 6153 -15751 7526 -15750
rect 6153 -15802 6456 -15751
rect 5799 -15803 6456 -15802
rect 6508 -15752 7169 -15751
rect 6508 -15803 6713 -15752
rect -2447 -15821 -2394 -15811
rect -2005 -15821 -1952 -15812
rect -2447 -15822 -1952 -15821
rect -1649 -15822 -1596 -15812
rect -1293 -15822 -1240 -15812
rect -937 -15822 -884 -15812
rect -581 -15822 -528 -15812
rect -225 -15822 -172 -15812
rect 132 -15822 185 -15811
rect 487 -15822 540 -15812
rect 843 -15822 896 -15812
rect 1201 -15822 1254 -15812
rect 1555 -15822 1608 -15812
rect 1910 -15822 1963 -15812
rect 2267 -15822 2320 -15812
rect 2624 -15822 2677 -15812
rect 2979 -15822 3032 -15812
rect 3335 -15822 3388 -15812
rect 3692 -15822 3745 -15812
rect 5747 -15813 5800 -15803
rect 6101 -15812 6154 -15803
rect 6456 -15813 6509 -15803
rect 6765 -15803 7169 -15752
rect 7221 -15802 7526 -15751
rect 7578 -15802 7882 -15750
rect 7934 -15751 11139 -15750
rect 7934 -15752 10730 -15751
rect 7934 -15802 10373 -15752
rect 7221 -15803 10373 -15802
rect 6765 -15804 6766 -15803
rect 6713 -15814 6766 -15804
rect 7169 -15813 7222 -15803
rect 7526 -15812 7579 -15803
rect 7882 -15812 7935 -15803
rect 10425 -15803 10730 -15752
rect 10782 -15803 11086 -15751
rect 11138 -15803 11139 -15751
rect 10425 -15804 10426 -15803
rect 10373 -15814 10426 -15804
rect 10730 -15813 10783 -15803
rect 11086 -15813 11139 -15803
rect -2395 -15823 132 -15822
rect -2395 -15874 -2005 -15823
rect -2447 -15884 -2394 -15874
rect -1953 -15875 -1649 -15823
rect -1597 -15875 -1293 -15823
rect -1241 -15875 -937 -15823
rect -885 -15875 -581 -15823
rect -529 -15875 -225 -15823
rect -173 -15874 132 -15823
rect 184 -15823 3745 -15822
rect 184 -15874 487 -15823
rect -173 -15875 487 -15874
rect 539 -15875 843 -15823
rect 895 -15875 1201 -15823
rect 1253 -15875 1555 -15823
rect 1607 -15875 1910 -15823
rect 1962 -15875 2267 -15823
rect 2319 -15875 2624 -15823
rect 2676 -15875 2979 -15823
rect 3031 -15875 3335 -15823
rect 3387 -15875 3692 -15823
rect 3744 -15875 3745 -15823
rect -2005 -15885 -1952 -15875
rect -1649 -15885 -1596 -15875
rect -1293 -15885 -1240 -15875
rect -937 -15885 -884 -15875
rect -581 -15885 -528 -15875
rect -225 -15885 -172 -15875
rect 132 -15884 185 -15875
rect 487 -15885 540 -15875
rect 843 -15885 896 -15875
rect 1201 -15885 1254 -15875
rect 1555 -15885 1608 -15875
rect 1910 -15885 1963 -15875
rect 2267 -15885 2320 -15875
rect 2624 -15885 2677 -15875
rect 2979 -15885 3032 -15875
rect 3335 -15885 3388 -15875
rect 3692 -15885 3745 -15875
rect 6813 -15851 6866 -15841
rect 7169 -15851 7222 -15842
rect 8060 -15851 8113 -15841
rect 11440 -15842 11493 -15831
rect 8593 -15851 8646 -15842
rect 9663 -15851 9716 -15842
rect 10194 -15851 10247 -15842
rect 11084 -15851 11137 -15842
rect 6813 -15852 11440 -15851
rect 6865 -15853 8060 -15852
rect 6865 -15904 7169 -15853
rect 6813 -15914 6866 -15904
rect 7221 -15904 8060 -15853
rect 8112 -15853 11440 -15852
rect 8112 -15904 8593 -15853
rect 7221 -15905 7222 -15904
rect 7169 -15915 7222 -15905
rect 8060 -15914 8113 -15904
rect 8645 -15904 9663 -15853
rect 8645 -15905 8646 -15904
rect 8593 -15915 8646 -15905
rect 9715 -15904 10194 -15853
rect 9715 -15905 9716 -15904
rect 9663 -15915 9716 -15905
rect 10246 -15904 11084 -15853
rect 10246 -15905 10247 -15904
rect 10194 -15915 10247 -15905
rect 11136 -15894 11440 -15853
rect 11492 -15894 11493 -15842
rect 11136 -15904 11493 -15894
rect 11136 -15905 11137 -15904
rect 11084 -15915 11137 -15905
rect -1915 -15933 -1862 -15923
rect -1738 -15933 -1685 -15923
rect -1560 -15933 -1507 -15923
rect -1382 -15933 -1329 -15923
rect -1204 -15933 -1151 -15923
rect -1025 -15933 -972 -15923
rect -847 -15933 -794 -15923
rect -670 -15933 -617 -15923
rect -491 -15933 -438 -15923
rect -313 -15933 -260 -15923
rect -136 -15933 -83 -15923
rect 43 -15933 96 -15923
rect 221 -15933 274 -15923
rect 398 -15933 451 -15923
rect 575 -15933 628 -15923
rect 755 -15933 808 -15923
rect 931 -15933 984 -15923
rect 1110 -15933 1163 -15923
rect 1289 -15933 1342 -15923
rect 1466 -15933 1519 -15923
rect 1643 -15933 1696 -15923
rect 1822 -15933 1875 -15923
rect 2000 -15933 2053 -15923
rect 2179 -15933 2232 -15923
rect 2356 -15933 2409 -15923
rect 2534 -15933 2587 -15923
rect 2712 -15933 2765 -15923
rect 2891 -15933 2944 -15923
rect 3068 -15933 3121 -15923
rect 3247 -15933 3300 -15923
rect 3424 -15933 3477 -15923
rect 3603 -15933 3656 -15923
rect 3780 -15933 3833 -15923
rect -1915 -15934 3833 -15933
rect -1863 -15986 -1738 -15934
rect -1686 -15986 -1560 -15934
rect -1508 -15986 -1382 -15934
rect -1330 -15986 -1204 -15934
rect -1152 -15986 -1025 -15934
rect -973 -15986 -847 -15934
rect -795 -15986 -670 -15934
rect -618 -15986 -491 -15934
rect -439 -15986 -313 -15934
rect -261 -15986 -136 -15934
rect -84 -15986 43 -15934
rect 95 -15986 221 -15934
rect 273 -15986 398 -15934
rect 450 -15986 575 -15934
rect 627 -15986 755 -15934
rect 807 -15986 931 -15934
rect 983 -15986 1110 -15934
rect 1162 -15986 1289 -15934
rect 1341 -15986 1466 -15934
rect 1518 -15986 1643 -15934
rect 1695 -15986 1822 -15934
rect 1874 -15986 2000 -15934
rect 2052 -15986 2179 -15934
rect 2231 -15986 2356 -15934
rect 2408 -15986 2534 -15934
rect 2586 -15986 2712 -15934
rect 2764 -15986 2891 -15934
rect 2943 -15986 3068 -15934
rect 3120 -15986 3247 -15934
rect 3299 -15986 3424 -15934
rect 3476 -15986 3603 -15934
rect 3655 -15986 3780 -15934
rect 3832 -15986 3833 -15934
rect -1915 -15996 -1862 -15986
rect -1738 -15996 -1685 -15986
rect -1560 -15996 -1507 -15986
rect -1382 -15996 -1329 -15986
rect -1204 -15996 -1151 -15986
rect -1025 -15996 -972 -15986
rect -847 -15996 -794 -15986
rect -670 -15996 -617 -15986
rect -491 -15996 -438 -15986
rect -313 -15996 -260 -15986
rect -136 -15996 -83 -15986
rect 43 -15996 96 -15986
rect 221 -15996 274 -15986
rect 398 -15996 451 -15986
rect 575 -15996 628 -15986
rect 755 -15996 808 -15986
rect 931 -15996 984 -15986
rect 1110 -15996 1163 -15986
rect 1289 -15996 1342 -15986
rect 1466 -15996 1519 -15986
rect 1643 -15996 1696 -15986
rect 1822 -15996 1875 -15986
rect 2000 -15996 2053 -15986
rect 2179 -15996 2232 -15986
rect 2356 -15996 2409 -15986
rect 2534 -15996 2587 -15986
rect 2712 -15996 2765 -15986
rect 2891 -15996 2944 -15986
rect 3068 -15996 3121 -15986
rect 3247 -15996 3300 -15986
rect 3424 -15996 3477 -15986
rect 3603 -15996 3656 -15986
rect 3780 -15996 3833 -15986
rect 5921 -15947 5974 -15938
rect 6279 -15947 6332 -15938
rect 6634 -15947 6687 -15938
rect 6994 -15947 7047 -15941
rect 5921 -15949 7047 -15947
rect 5973 -16000 6279 -15949
rect 5973 -16001 5974 -16000
rect 5921 -16011 5974 -16001
rect 6331 -16000 6634 -15949
rect 6331 -16001 6332 -16000
rect 6279 -16011 6332 -16001
rect 6686 -15952 7047 -15949
rect 6686 -16000 6994 -15952
rect 6686 -16001 6687 -16000
rect 6634 -16011 6687 -16001
rect 7046 -16004 7047 -15952
rect 6994 -16014 7047 -16004
rect 7526 -15952 7579 -15943
rect 7881 -15952 7934 -15942
rect 8237 -15952 8290 -15942
rect 11441 -15952 11494 -15942
rect 11797 -15952 11850 -15942
rect 12154 -15952 12207 -15942
rect 12511 -15952 12564 -15942
rect 7526 -15953 12564 -15952
rect 7526 -15954 7881 -15953
rect 7578 -16005 7881 -15954
rect 7933 -16005 8237 -15953
rect 8289 -16005 11441 -15953
rect 11493 -16005 11797 -15953
rect 11849 -16005 12154 -15953
rect 12206 -16005 12511 -15953
rect 12563 -16005 12564 -15953
rect 7578 -16006 7579 -16005
rect 7526 -16016 7579 -16006
rect 7881 -16015 7934 -16005
rect 8237 -16015 8290 -16005
rect 11441 -16015 11494 -16005
rect 11797 -16015 11850 -16005
rect 12154 -16015 12207 -16005
rect 12511 -16015 12564 -16005
rect -6159 -16193 -6106 -16183
rect -5504 -16193 -5451 -16183
rect -4792 -16193 -4739 -16183
rect -6159 -16194 -4739 -16193
rect -6107 -16246 -5504 -16194
rect -5452 -16246 -4792 -16194
rect -4740 -16246 -4739 -16194
rect -6159 -16256 -6106 -16246
rect -5504 -16256 -5451 -16246
rect -4792 -16256 -4739 -16246
rect -5860 -16294 -5807 -16284
rect -5148 -16294 -5095 -16284
rect -4436 -16294 -4383 -16284
rect -3935 -16294 -3883 -16285
rect -5860 -16295 -3883 -16294
rect -5808 -16347 -5148 -16295
rect -5096 -16346 -4436 -16295
rect -5096 -16347 -5095 -16346
rect -5860 -16357 -5807 -16347
rect -5148 -16357 -5095 -16347
rect -4384 -16346 -3935 -16295
rect -4384 -16347 -4383 -16346
rect -4436 -16357 -4383 -16347
rect -3935 -16357 -3883 -16347
rect -1917 -16542 -1864 -16532
rect -1738 -16542 -1685 -16532
rect -1561 -16542 -1508 -16531
rect -1381 -16542 -1328 -16533
rect -1204 -16542 -1151 -16532
rect -1026 -16542 -973 -16532
rect 220 -16542 273 -16532
rect 397 -16542 450 -16532
rect 576 -16542 629 -16532
rect 755 -16542 808 -16532
rect 933 -16542 986 -16532
rect 1111 -16542 1164 -16532
rect 2356 -16542 2409 -16532
rect 2534 -16542 2587 -16532
rect 2713 -16542 2766 -16531
rect 2891 -16542 2944 -16532
rect 3070 -16542 3123 -16532
rect 3249 -16542 3302 -16532
rect 4238 -16542 4291 -16532
rect -1917 -16543 -1561 -16542
rect -1865 -16595 -1738 -16543
rect -1686 -16594 -1561 -16543
rect -1509 -16543 2713 -16542
rect -1509 -16544 -1204 -16543
rect -1509 -16594 -1381 -16544
rect -1686 -16595 -1381 -16594
rect -1917 -16605 -1864 -16595
rect -1738 -16605 -1685 -16595
rect -1561 -16604 -1508 -16595
rect -1329 -16595 -1204 -16544
rect -1152 -16595 -1026 -16543
rect -974 -16595 220 -16543
rect 272 -16595 397 -16543
rect 449 -16595 576 -16543
rect 628 -16595 755 -16543
rect 807 -16595 933 -16543
rect 985 -16595 1111 -16543
rect 1163 -16595 2356 -16543
rect 2408 -16595 2534 -16543
rect 2586 -16594 2713 -16543
rect 2765 -16543 4291 -16542
rect 2765 -16594 2891 -16543
rect 2586 -16595 2891 -16594
rect 2943 -16595 3070 -16543
rect 3122 -16595 3249 -16543
rect 3301 -16595 4238 -16543
rect 4290 -16595 4291 -16543
rect -1329 -16596 -1328 -16595
rect -1381 -16606 -1328 -16596
rect -1204 -16605 -1151 -16595
rect -1026 -16605 -973 -16595
rect 220 -16605 273 -16595
rect 397 -16605 450 -16595
rect 576 -16605 629 -16595
rect 755 -16605 808 -16595
rect 933 -16605 986 -16595
rect 1111 -16605 1164 -16595
rect 2356 -16605 2409 -16595
rect 2534 -16605 2587 -16595
rect 2713 -16604 2766 -16595
rect 2891 -16605 2944 -16595
rect 3070 -16605 3123 -16595
rect 3249 -16605 3302 -16595
rect 4238 -16605 4291 -16595
rect 6548 -16545 6601 -16534
rect 6726 -16545 6779 -16534
rect 6903 -16545 6956 -16535
rect 7970 -16545 8023 -16535
rect 8149 -16545 8202 -16534
rect 9929 -16545 9982 -16534
rect 10107 -16545 10160 -16535
rect 10287 -16545 10340 -16535
rect 11352 -16545 11405 -16535
rect 11530 -16545 11583 -16536
rect 11709 -16545 11762 -16535
rect 6600 -16597 6726 -16545
rect 6778 -16546 8149 -16545
rect 6778 -16597 6903 -16546
rect 6548 -16598 6903 -16597
rect 6955 -16598 7970 -16546
rect 8022 -16597 8149 -16546
rect 8201 -16597 9929 -16545
rect 9981 -16546 11762 -16545
rect 9981 -16597 10107 -16546
rect 8022 -16598 10107 -16597
rect 10159 -16598 10287 -16546
rect 10339 -16598 11352 -16546
rect 11404 -16547 11709 -16546
rect 11404 -16598 11530 -16547
rect 6548 -16607 6601 -16598
rect 6726 -16607 6779 -16598
rect 6903 -16608 6956 -16598
rect 7970 -16608 8023 -16598
rect 8149 -16607 8202 -16598
rect 9929 -16607 9982 -16598
rect 10107 -16608 10160 -16598
rect 10287 -16608 10340 -16598
rect 11352 -16608 11405 -16598
rect 11582 -16598 11709 -16547
rect 11761 -16598 11762 -16546
rect 11582 -16599 11583 -16598
rect 11530 -16609 11583 -16599
rect 11709 -16608 11762 -16598
rect -1827 -16665 -1774 -16655
rect -1720 -16665 -1548 -16655
rect -1471 -16665 -1418 -16656
rect -1114 -16665 -1061 -16655
rect -759 -16665 -706 -16654
rect -646 -16665 -471 -16655
rect -403 -16665 -350 -16655
rect -47 -16665 6 -16655
rect 309 -16665 362 -16656
rect 426 -16665 595 -16655
rect 665 -16665 718 -16655
rect 1021 -16665 1074 -16655
rect 1377 -16665 1430 -16655
rect 1501 -16665 1671 -16655
rect 1735 -16665 1788 -16655
rect 2090 -16665 2143 -16654
rect 2445 -16665 2498 -16655
rect 2568 -16665 2732 -16655
rect 2801 -16665 2854 -16655
rect 3157 -16665 3210 -16654
rect 3514 -16665 3567 -16656
rect 3633 -16665 3804 -16655
rect 3868 -16665 3921 -16655
rect -1827 -16666 -759 -16665
rect -1775 -16718 -1692 -16666
rect -1640 -16718 -1628 -16666
rect -1576 -16667 -1114 -16666
rect -1576 -16718 -1471 -16667
rect -1827 -16728 -1774 -16718
rect -1720 -16728 -1548 -16718
rect -1419 -16718 -1114 -16667
rect -1062 -16717 -759 -16666
rect -707 -16666 2090 -16665
rect -707 -16717 -617 -16666
rect -1062 -16718 -617 -16717
rect -565 -16718 -553 -16666
rect -501 -16718 -403 -16666
rect -351 -16718 -47 -16666
rect 5 -16667 452 -16666
rect 5 -16718 309 -16667
rect -1419 -16719 -1418 -16718
rect -1471 -16729 -1418 -16719
rect -1114 -16728 -1061 -16718
rect -759 -16727 -706 -16718
rect -646 -16728 -471 -16718
rect -403 -16728 -350 -16718
rect -47 -16728 6 -16718
rect 361 -16718 452 -16667
rect 504 -16718 516 -16666
rect 568 -16718 665 -16666
rect 717 -16718 1021 -16666
rect 1073 -16718 1377 -16666
rect 1429 -16718 1528 -16666
rect 1580 -16718 1592 -16666
rect 1644 -16718 1735 -16666
rect 1787 -16717 2090 -16666
rect 2142 -16666 3157 -16665
rect 2142 -16717 2445 -16666
rect 1787 -16718 2445 -16717
rect 2497 -16718 2592 -16666
rect 2644 -16718 2656 -16666
rect 2708 -16718 2801 -16666
rect 2853 -16717 3157 -16666
rect 3209 -16666 3921 -16665
rect 3209 -16667 3660 -16666
rect 3209 -16717 3514 -16667
rect 2853 -16718 3514 -16717
rect 361 -16719 362 -16718
rect 309 -16729 362 -16719
rect 426 -16728 595 -16718
rect 665 -16728 718 -16718
rect 1021 -16728 1074 -16718
rect 1377 -16728 1430 -16718
rect 1501 -16728 1671 -16718
rect 1735 -16728 1788 -16718
rect 2090 -16727 2143 -16718
rect 2445 -16728 2498 -16718
rect 2568 -16728 2732 -16718
rect 2801 -16728 2854 -16718
rect 3157 -16727 3210 -16718
rect 3566 -16718 3660 -16667
rect 3712 -16718 3724 -16666
rect 3776 -16718 3868 -16666
rect 3920 -16718 3921 -16666
rect 3566 -16719 3567 -16718
rect 3514 -16729 3567 -16719
rect 3633 -16728 3804 -16718
rect 3868 -16728 3921 -16718
rect 5399 -16666 5452 -16657
rect 8771 -16666 8824 -16656
rect 9128 -16666 9181 -16656
rect 9484 -16666 9537 -16656
rect 5399 -16667 9537 -16666
rect 5399 -16668 8771 -16667
rect 5451 -16719 8771 -16668
rect 8823 -16719 9128 -16667
rect 9180 -16719 9484 -16667
rect 9536 -16719 9537 -16667
rect 5451 -16720 5452 -16719
rect 5399 -16730 5452 -16720
rect 8771 -16729 8824 -16719
rect 9128 -16729 9181 -16719
rect 9484 -16729 9537 -16719
rect 9838 -16665 9891 -16656
rect 10195 -16665 10248 -16655
rect 10550 -16665 10603 -16655
rect 10907 -16665 10960 -16655
rect 9838 -16666 10960 -16665
rect 9838 -16667 10195 -16666
rect 9890 -16718 10195 -16667
rect 10247 -16718 10550 -16666
rect 10602 -16718 10907 -16666
rect 10959 -16718 10960 -16666
rect 9890 -16719 9891 -16718
rect 9838 -16729 9891 -16719
rect 10195 -16728 10248 -16718
rect 10550 -16728 10603 -16718
rect 10907 -16728 10960 -16718
rect 5031 -16782 5084 -16772
rect 8950 -16782 9003 -16772
rect 9305 -16782 9358 -16772
rect 5031 -16783 9358 -16782
rect 5083 -16835 8950 -16783
rect 9002 -16835 9305 -16783
rect 9357 -16835 9358 -16783
rect 5031 -16845 5084 -16835
rect 8950 -16845 9003 -16835
rect 9305 -16845 9358 -16835
rect 10017 -16780 10070 -16771
rect 10374 -16780 10427 -16771
rect 10731 -16780 10784 -16769
rect 10017 -16782 10731 -16780
rect 10069 -16833 10374 -16782
rect 10069 -16834 10070 -16833
rect 10017 -16844 10070 -16834
rect 10426 -16832 10731 -16782
rect 10783 -16832 10784 -16780
rect 10426 -16833 10784 -16832
rect 10426 -16834 10427 -16833
rect 10374 -16844 10427 -16834
rect 10731 -16842 10784 -16833
rect -5682 -16886 -5629 -16876
rect -5326 -16886 -5273 -16876
rect -4970 -16886 -4917 -16876
rect -4614 -16886 -4561 -16876
rect -4258 -16886 -4205 -16876
rect -5682 -16887 -4205 -16886
rect -5630 -16939 -5326 -16887
rect -5274 -16939 -4970 -16887
rect -4918 -16939 -4614 -16887
rect -4562 -16939 -4258 -16887
rect -4206 -16939 -4205 -16887
rect -5682 -16949 -5629 -16939
rect -5326 -16949 -5273 -16939
rect -4970 -16949 -4917 -16939
rect -4614 -16949 -4561 -16939
rect -4258 -16949 -4205 -16939
rect 7347 -16890 7400 -16880
rect 7704 -16890 7757 -16880
rect 8060 -16890 8113 -16880
rect 8416 -16890 8469 -16880
rect 11263 -16890 11316 -16880
rect 11620 -16890 11673 -16880
rect 11975 -16890 12028 -16879
rect 12331 -16890 12384 -16879
rect 7347 -16891 11975 -16890
rect 7399 -16943 7704 -16891
rect 7756 -16943 8060 -16891
rect 8112 -16943 8416 -16891
rect 8468 -16943 11263 -16891
rect 11315 -16943 11620 -16891
rect 11672 -16942 11975 -16891
rect 12027 -16942 12331 -16890
rect 12383 -16942 12384 -16890
rect 11672 -16943 12384 -16942
rect 7347 -16953 7400 -16943
rect 7704 -16953 7757 -16943
rect 8060 -16953 8113 -16943
rect 8416 -16953 8469 -16943
rect 11263 -16953 11316 -16943
rect 11620 -16953 11673 -16943
rect 11975 -16952 12028 -16943
rect 12331 -16952 12384 -16943
rect -6159 -17007 -6106 -16997
rect -5859 -17007 -5806 -16997
rect -5148 -17007 -5095 -16997
rect -4437 -17007 -4384 -16997
rect -6159 -17008 -4384 -17007
rect -6107 -17060 -5859 -17008
rect -5807 -17060 -5148 -17008
rect -5096 -17060 -4437 -17008
rect -4385 -17060 -4384 -17008
rect -6159 -17070 -6106 -17060
rect -5859 -17070 -5806 -17060
rect -5148 -17070 -5095 -17060
rect -4437 -17070 -4384 -17060
rect -5504 -17118 -5451 -17108
rect -4792 -17118 -4739 -17108
rect -3935 -17118 -3883 -17108
rect -5504 -17119 -3935 -17118
rect -5452 -17170 -4792 -17119
rect -5452 -17171 -5451 -17170
rect -5504 -17181 -5451 -17171
rect -4740 -17170 -3935 -17119
rect -4740 -17171 -4739 -17170
rect -4792 -17181 -4739 -17171
rect -3935 -17180 -3883 -17170
<< via2 >>
rect 3021 -3511 3077 -3455
rect -2544 -3987 -2488 -3931
rect 2540 -4271 2596 -4269
rect 2540 -4323 2542 -4271
rect 2542 -4323 2594 -4271
rect 2594 -4323 2596 -4271
rect 2540 -4325 2596 -4323
rect -2383 -4564 -2327 -4508
rect 2748 -4451 2804 -4449
rect 2748 -4503 2750 -4451
rect 2750 -4503 2802 -4451
rect 2802 -4503 2804 -4451
rect 2748 -4505 2804 -4503
rect 3023 -5061 3079 -5005
rect -2383 -5152 -2327 -5096
rect 313 -5207 369 -5151
rect -1644 -5283 -1588 -5281
rect -1644 -5335 -1642 -5283
rect -1642 -5335 -1590 -5283
rect -1590 -5335 -1588 -5283
rect -1644 -5337 -1588 -5335
rect 848 -5337 904 -5281
rect -3543 -6865 -3487 -6809
rect -3384 -7038 -3328 -6982
<< metal3 >>
rect 6451 929 6515 2665
rect 6704 121 6768 1857
rect 17697 122 17761 1858
rect 17950 929 18014 2665
rect 3009 -3455 3090 -3447
rect 3009 -3511 3021 -3455
rect 3077 -3511 3090 -3455
rect 3009 -3518 3090 -3511
rect -2556 -3931 -2475 -3923
rect -2556 -3987 -2544 -3931
rect -2488 -3987 -2475 -3931
rect -2556 -3994 -2475 -3987
rect -2546 -4266 -2485 -3994
rect 2528 -4266 2609 -4261
rect -2546 -4269 2609 -4266
rect -2546 -4325 2540 -4269
rect 2596 -4325 2609 -4269
rect -2546 -4327 2609 -4325
rect -2546 -6637 -2485 -4327
rect 2528 -4332 2609 -4327
rect 2736 -4446 2817 -4441
rect -2385 -4449 2817 -4446
rect -2385 -4500 2748 -4449
rect -2395 -4505 2748 -4500
rect 2804 -4505 2817 -4449
rect -2395 -4507 2817 -4505
rect -2395 -4508 -2314 -4507
rect -2395 -4564 -2383 -4508
rect -2327 -4564 -2314 -4508
rect 2736 -4512 2817 -4507
rect -2395 -4571 -2314 -4564
rect -2385 -5088 -2324 -4571
rect 3021 -4997 3082 -3518
rect 3011 -5005 3092 -4997
rect 3011 -5061 3023 -5005
rect 3079 -5061 3092 -5005
rect 3011 -5068 3092 -5061
rect -2395 -5096 -2314 -5088
rect -2395 -5152 -2383 -5096
rect -2327 -5152 -2314 -5096
rect -2395 -5159 -2314 -5152
rect 301 -5147 382 -5143
rect 3021 -5147 3082 -5068
rect 301 -5151 3082 -5147
rect -3545 -6698 -2485 -6637
rect -3545 -6801 -3484 -6698
rect -2385 -6786 -2324 -5159
rect 301 -5207 313 -5151
rect 369 -5207 3082 -5151
rect 301 -5208 3082 -5207
rect 301 -5214 382 -5208
rect -1656 -5278 -1575 -5273
rect 836 -5278 917 -5273
rect -1656 -5281 917 -5278
rect -1656 -5337 -1644 -5281
rect -1588 -5337 848 -5281
rect 904 -5337 917 -5281
rect -1656 -5339 917 -5337
rect -1656 -5344 -1575 -5339
rect 836 -5344 917 -5339
rect 6451 -6271 6515 -4535
rect 6704 -5279 6768 -3543
rect -3555 -6809 -3474 -6801
rect -3555 -6865 -3543 -6809
rect -3487 -6865 -3474 -6809
rect -3555 -6872 -3474 -6865
rect -3386 -6847 -2324 -6786
rect -3386 -6974 -3325 -6847
rect -3396 -6982 -3315 -6974
rect -3396 -7038 -3384 -6982
rect -3328 -7038 -3315 -6982
rect -3396 -7045 -3315 -7038
rect 17697 -7078 17761 -5342
rect 17950 -6271 18014 -4535
use sc_cmfb  sc_cmfb_0
timestamp 1654583101
transform 1 0 9102 0 1 -5469
box -3494 -1840 9310 8360
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_0
timestamp 1654583101
transform 1 0 7953 0 1 -9022
box -1479 -228 1479 228
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_1
timestamp 1654583101
transform 1 0 7953 0 1 -9922
box -1479 -228 1479 228
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_2
timestamp 1654583101
transform 1 0 7953 0 1 -10822
box -1479 -228 1479 228
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_3
timestamp 1654583101
transform 1 0 7953 0 1 -11722
box -1479 -228 1479 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_0
timestamp 1654583101
transform 1 0 -5032 0 1 -14522
box -1034 -228 1034 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_1
timestamp 1654583101
transform 1 0 -5032 0 1 -15222
box -1034 -228 1034 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_2
timestamp 1654583101
transform 1 0 -5032 0 1 -15922
box -1034 -228 1034 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_3
timestamp 1654583101
transform 1 0 -5032 0 1 -16622
box -1034 -228 1034 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_0
timestamp 1654583101
transform 1 0 959 0 1 -8260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_1
timestamp 1654583101
transform 1 0 959 0 1 -9260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_2
timestamp 1654583101
transform 1 0 959 0 1 -10260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_3
timestamp 1654583101
transform 1 0 959 0 1 -11260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_4
timestamp 1654583101
transform 1 0 959 0 1 -12260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_5
timestamp 1654583101
transform 1 0 959 0 1 -13260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_6
timestamp 1654583101
transform 1 0 959 0 1 -14260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_7
timestamp 1654583101
transform 1 0 959 0 1 -15260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_8
timestamp 1654583101
transform 1 0 959 0 1 -16260
box -3170 -228 3170 228
use sky130_fd_pr__nfet_01v8_DD  sky130_fd_pr__nfet_01v8_DD_0
timestamp 1654583101
transform 1 0 9154 0 1 -14260
box -3615 -228 3615 228
use sky130_fd_pr__nfet_01v8_DD  sky130_fd_pr__nfet_01v8_DD_1
timestamp 1654583101
transform 1 0 9154 0 1 -15260
box -3615 -228 3615 228
use sky130_fd_pr__nfet_01v8_DD  sky130_fd_pr__nfet_01v8_DD_2
timestamp 1654583101
transform 1 0 9154 0 1 -16260
box -3615 -228 3615 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_0
timestamp 1654583101
transform 1 0 11754 0 1 -9052
box -1020 -228 1020 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_1
timestamp 1654583101
transform 1 0 11754 0 1 -9822
box -1020 -228 1020 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_2
timestamp 1654583101
transform 1 0 11754 0 1 -10592
box -1020 -228 1020 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_3
timestamp 1654583101
transform 1 0 11754 0 1 -11362
box -1020 -228 1020 228
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_0
timestamp 1654583101
transform 1 0 -5850 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_1
timestamp 1654583101
transform 1 0 -5600 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_2
timestamp 1654583101
transform 1 0 -5350 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_3
timestamp 1654583101
transform 1 0 -5100 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_4
timestamp 1654583101
transform 1 0 -4850 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_5
timestamp 1654583101
transform 1 0 -4600 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_6
timestamp 1654583101
transform 1 0 -4350 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_7
timestamp 1654583101
transform 1 0 -4100 0 1 -12820
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_8
timestamp 1654583101
transform 1 0 -5850 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_9
timestamp 1654583101
transform 1 0 -5600 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_10
timestamp 1654583101
transform 1 0 -5350 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_11
timestamp 1654583101
transform 1 0 -5100 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_12
timestamp 1654583101
transform 1 0 -4850 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_13
timestamp 1654583101
transform 1 0 -4600 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_14
timestamp 1654583101
transform 1 0 -4350 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_15
timestamp 1654583101
transform 1 0 -4100 0 1 -13500
box -104 -208 104 208
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_0
timestamp 1654583101
transform 1 0 -4810 0 1 -8002
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_1
timestamp 1654583101
transform 1 0 -4810 0 1 -8552
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_2
timestamp 1654583101
transform 1 0 -4810 0 1 -9102
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_3
timestamp 1654583101
transform 1 0 -4810 0 1 -9652
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_4
timestamp 1654583101
transform 1 0 -4810 0 1 -10202
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_5
timestamp 1654583101
transform 1 0 -4810 0 1 -10752
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_6
timestamp 1654583101
transform 1 0 -4810 0 1 -11302
box -856 -228 856 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_7
timestamp 1654583101
transform 1 0 -4810 0 1 -11852
box -856 -228 856 228
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_0
timestamp 1654583101
transform 1 0 610 0 1 -5712
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_1
timestamp 1654583101
transform 1 0 610 0 1 -4812
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_2
timestamp 1654583101
transform 1 0 610 0 1 -3912
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_3
timestamp 1654583101
transform 1 0 610 0 1 -3012
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_0
timestamp 1654583101
transform 1 0 -4861 0 1 -5740
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_1
timestamp 1654583101
transform 1 0 -4861 0 1 -4870
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_2
timestamp 1654583101
transform 1 0 -4861 0 1 -4000
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_3
timestamp 1654583101
transform 1 0 -4861 0 1 -3130
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_4
timestamp 1654583101
transform 1 0 -4861 0 1 -2260
box -1489 -241 1489 241
<< labels >>
flabel metal1 s -6950 -12541 -6950 -12541 1 FreeSans 1500 0 0 0 ip
port 1 nsew
flabel metal1 s -6952 -13880 -6952 -13880 1 FreeSans 1500 0 0 0 in
port 2 nsew
flabel metal3 s 6735 -5207 6735 -5207 1 FreeSans 500 0 0 0 p1
port 3 nsew
flabel metal3 s 17727 -7023 17727 -7023 1 FreeSans 500 0 0 0 p1
port 3 nsew
flabel metal3 s 6486 -6211 6486 -6211 1 FreeSans 500 0 0 0 p1_b
port 4 nsew
flabel metal3 s 17984 -6236 17984 -6236 1 FreeSans 500 0 0 0 p1_b
port 4 nsew
flabel metal3 s 6738 1807 6738 1807 1 FreeSans 500 0 0 0 p2
port 5 nsew
flabel metal3 s 17730 1821 17730 1821 1 FreeSans 500 0 0 0 p2
port 5 nsew
flabel metal3 s 6479 2585 6479 2585 1 FreeSans 500 0 0 0 p2_b
port 6 nsew
flabel metal3 s 17980 2631 17980 2631 1 FreeSans 500 0 0 0 p2_b
port 6 nsew
flabel metal2 s 3431 -5243 3431 -5243 1 FreeSans 1500 0 0 0 op
port 7 nsew
flabel metal2 s 3147 -3484 3147 -3484 1 FreeSans 1500 0 0 0 on
port 8 nsew
flabel metal1 s -6957 -14245 -6957 -14245 1 FreeSans 1500 0 0 0 i_bias
port 9 nsew
flabel metal2 s 17862 -8732 17862 -8732 1 FreeSans 1000 0 0 0 cm
port 10 nsew
flabel metal1 s 4262 -15741 4262 -15741 1 FreeSans 1500 0 0 0 bias_a
port 11 nsew
flabel metal1 s -4277 -7715 -4277 -7715 1 FreeSans 1500 0 0 0 bias_b
port 12 nsew
flabel metal1 s -3636 -12323 -3636 -12323 1 FreeSans 1500 0 0 0 bias_c
port 13 nsew
flabel metal1 s 6929 -13167 6929 -13167 1 FreeSans 1500 0 0 0 bias_d
port 14 nsew
flabel metal2 s 5049 -9956 5049 -9956 1 FreeSans 1500 0 0 0 cmc
port 15 nsew
flabel metal1 s -7420 -1403 -7420 -1403 1 FreeSans 1500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7057 2874 7057 2874 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7058 -739 7058 -739 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7058 -2537 7058 -2537 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7051 -4329 7051 -4329 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 16057 -6136 16057 -6136 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 16057 -2529 16057 -2529 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 16057 1070 16057 1070 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 16057 2870 16057 2870 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7058 1058 7058 1058 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7058 -6144 7058 -6144 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 16056 -4338 16056 -4338 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 16056 -738 16056 -738 1 FreeSans 500 0 0 0 VDD
port 16 nsew
flabel metal1 s 7057 1707 7057 1707 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 7058 -83 7058 -83 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 7058 -1885 7058 -1885 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 7054 -5489 7054 -5489 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 7054 -7288 7054 -7288 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 16056 -7290 16056 -7290 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 16055 -5482 16055 -5482 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 16055 -1886 16055 -1886 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 16057 -86 16057 -86 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 16057 1716 16057 1716 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 7058 -3672 7058 -3672 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 16056 -3678 16056 -3678 1 FreeSans 500 0 0 0 VSS
port 17 nsew
flabel metal1 s 1056 -17349 1056 -17349 1 FreeSans 2000 0 0 0 VSS
port 17 nsew
<< end >>
