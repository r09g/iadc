magic
tech sky130A
magscale 1 2
timestamp 1653212313
<< metal1 >>
rect -6877 -1963 -6867 -1910
rect -6814 -1963 -6804 -1910
rect -6699 -1963 -6689 -1910
rect -6636 -1963 -6626 -1910
rect -6520 -1963 -6510 -1910
rect -6457 -1963 -6447 -1910
rect -6343 -1963 -6333 -1910
rect -6280 -1963 -6270 -1910
rect -6165 -1963 -6155 -1910
rect -6102 -1963 -6092 -1910
rect -5986 -1963 -5976 -1910
rect -5923 -1963 -5913 -1910
rect -5809 -1963 -5799 -1910
rect -5746 -1963 -5736 -1910
rect -5631 -1963 -5621 -1910
rect -5568 -1963 -5558 -1910
rect -5453 -1963 -5443 -1910
rect -5390 -1963 -5380 -1910
rect -5275 -1963 -5265 -1910
rect -5212 -1963 -5202 -1910
rect -5096 -1963 -5086 -1910
rect -5033 -1963 -5023 -1910
rect -4919 -1963 -4909 -1910
rect -4856 -1963 -4846 -1910
rect -6857 -2079 -6823 -1963
rect -6679 -2079 -6645 -1963
rect -6501 -2079 -6467 -1963
rect -6322 -2079 -6288 -1963
rect -6145 -2079 -6111 -1963
rect -5967 -2079 -5933 -1963
rect -5789 -2079 -5755 -1963
rect -5611 -2079 -5577 -1963
rect -5433 -2079 -5399 -1963
rect -5255 -2079 -5221 -1963
rect -5077 -2079 -5043 -1963
rect -4898 -2079 -4864 -1963
rect -7508 -2582 -7498 -2529
rect -7445 -2582 -7435 -2529
rect -7635 -3454 -7625 -3401
rect -7572 -3454 -7562 -3401
rect -7625 -5322 -7572 -3454
rect -7498 -3640 -7445 -2582
rect -7054 -2833 -7044 -2780
rect -6991 -2833 -6981 -2780
rect -7035 -2949 -7001 -2833
rect -7124 -3401 -7090 -3259
rect -7144 -3454 -7134 -3401
rect -7081 -3454 -7071 -3401
rect -7508 -3693 -7498 -3640
rect -7445 -3693 -7435 -3640
rect -7498 -4271 -7445 -3693
rect -7035 -3819 -7001 -3311
rect -7508 -4324 -7498 -4271
rect -7445 -4324 -7435 -4271
rect -7498 -5141 -7445 -4324
rect -7124 -4390 -7090 -4128
rect -7144 -4443 -7134 -4390
rect -7081 -4443 -7071 -4390
rect -7035 -4689 -7001 -4181
rect -7508 -5194 -7498 -5141
rect -7445 -5194 -7435 -5141
rect -7635 -5375 -7625 -5322
rect -7572 -5375 -7562 -5322
rect -7498 -6248 -7445 -5194
rect -7124 -5232 -7090 -4998
rect -7144 -5285 -7134 -5232
rect -7081 -5285 -7071 -5232
rect -6946 -5612 -6912 -2388
rect -6856 -2780 -6822 -2447
rect -6768 -2530 -6734 -2389
rect -6787 -2583 -6777 -2530
rect -6724 -2583 -6714 -2530
rect -6876 -2833 -6866 -2780
rect -6813 -2833 -6803 -2780
rect -6856 -2943 -6822 -2833
rect -6679 -2949 -6645 -2447
rect -6857 -3819 -6823 -3311
rect -6768 -3516 -6734 -3258
rect -6787 -3569 -6777 -3516
rect -6724 -3569 -6714 -3516
rect -6679 -3819 -6645 -3311
rect -6857 -4689 -6823 -4181
rect -6768 -4271 -6734 -4128
rect -6788 -4324 -6778 -4271
rect -6725 -4324 -6715 -4271
rect -6679 -4689 -6645 -4181
rect -6857 -5559 -6823 -5051
rect -6768 -5415 -6734 -4999
rect -6787 -5468 -6777 -5415
rect -6724 -5468 -6714 -5415
rect -6679 -5559 -6645 -5051
rect -6590 -5612 -6556 -2388
rect -6501 -2949 -6467 -2441
rect -6412 -2668 -6378 -2388
rect -6431 -2721 -6421 -2668
rect -6368 -2721 -6358 -2668
rect -6323 -2949 -6289 -2441
rect -6501 -3819 -6467 -3311
rect -6412 -3640 -6378 -3258
rect -6432 -3693 -6422 -3640
rect -6369 -3693 -6359 -3640
rect -6323 -3819 -6289 -3311
rect -6501 -4689 -6467 -4181
rect -6412 -4506 -6378 -4128
rect -6432 -4559 -6422 -4506
rect -6369 -4559 -6359 -4506
rect -6323 -4689 -6289 -4181
rect -6501 -5559 -6467 -5051
rect -6412 -5141 -6378 -4998
rect -6432 -5194 -6422 -5141
rect -6369 -5194 -6359 -5141
rect -6323 -5559 -6289 -5051
rect -6234 -5612 -6200 -2388
rect -6145 -2949 -6111 -2441
rect -6056 -2530 -6022 -2388
rect -6076 -2583 -6066 -2530
rect -6013 -2583 -6003 -2530
rect -5967 -2949 -5933 -2441
rect -6145 -3819 -6111 -3311
rect -6056 -3401 -6022 -3259
rect -6076 -3454 -6066 -3401
rect -6013 -3454 -6003 -3401
rect -5967 -3819 -5933 -3311
rect -6145 -4689 -6111 -4181
rect -6056 -4390 -6022 -4127
rect -6076 -4443 -6066 -4390
rect -6013 -4443 -6003 -4390
rect -5967 -4689 -5933 -4181
rect -6145 -5559 -6111 -5051
rect -6056 -5233 -6022 -4998
rect -6076 -5286 -6066 -5233
rect -6013 -5286 -6003 -5233
rect -5967 -5559 -5933 -5051
rect -5878 -5612 -5844 -2388
rect -5789 -2949 -5755 -2441
rect -5700 -2668 -5666 -2388
rect -5720 -2721 -5710 -2668
rect -5657 -2721 -5647 -2668
rect -5611 -2949 -5577 -2441
rect -5789 -3819 -5755 -3311
rect -5700 -3401 -5666 -3258
rect -5720 -3454 -5710 -3401
rect -5657 -3454 -5647 -3401
rect -5611 -3819 -5577 -3311
rect -5789 -4689 -5755 -4181
rect -5700 -4390 -5666 -4128
rect -5719 -4443 -5709 -4390
rect -5656 -4443 -5646 -4390
rect -5611 -4689 -5577 -4181
rect -5789 -5559 -5755 -5051
rect -5700 -5322 -5666 -4998
rect -5720 -5375 -5710 -5322
rect -5657 -5375 -5647 -5322
rect -5611 -5559 -5577 -5051
rect -5522 -5612 -5488 -2388
rect -5433 -2949 -5399 -2441
rect -5344 -2530 -5310 -2388
rect -5364 -2583 -5354 -2530
rect -5301 -2583 -5291 -2530
rect -5255 -2949 -5221 -2441
rect -5433 -3819 -5399 -3311
rect -5344 -3640 -5310 -3258
rect -5363 -3693 -5353 -3640
rect -5300 -3693 -5290 -3640
rect -5254 -3819 -5220 -3311
rect -5433 -4689 -5399 -4181
rect -5344 -4506 -5310 -4128
rect -5363 -4559 -5353 -4506
rect -5300 -4559 -5290 -4506
rect -5255 -4689 -5221 -4181
rect -5433 -5559 -5399 -5051
rect -5344 -5141 -5310 -4998
rect -5363 -5194 -5353 -5141
rect -5300 -5194 -5290 -5141
rect -5255 -5559 -5221 -5051
rect -5166 -5612 -5132 -2388
rect -5077 -2949 -5043 -2441
rect -4988 -2668 -4954 -2388
rect -5008 -2721 -4998 -2668
rect -4945 -2721 -4935 -2668
rect -4899 -2780 -4865 -2441
rect -4918 -2833 -4908 -2780
rect -4855 -2833 -4845 -2780
rect -4899 -2949 -4865 -2833
rect -5077 -3819 -5043 -3311
rect -4988 -3516 -4954 -3258
rect -5008 -3569 -4998 -3516
rect -4945 -3569 -4935 -3516
rect -4899 -3819 -4865 -3311
rect -5077 -4689 -5043 -4181
rect -4988 -4271 -4954 -4128
rect -5008 -4324 -4998 -4271
rect -4945 -4324 -4935 -4271
rect -4899 -4689 -4865 -4181
rect -5077 -5559 -5043 -5051
rect -4988 -5415 -4954 -4998
rect -5007 -5468 -4997 -5415
rect -4944 -5468 -4934 -5415
rect -4899 -5559 -4865 -5051
rect -4810 -5612 -4776 -2388
rect -4308 -2721 -4298 -2668
rect -4245 -2721 -4235 -2668
rect -4741 -2833 -4731 -2780
rect -4678 -2833 -4668 -2780
rect -4721 -2949 -4687 -2833
rect -4721 -3819 -4687 -3311
rect -4632 -3401 -4598 -3258
rect -4652 -3454 -4642 -3401
rect -4589 -3454 -4579 -3401
rect -4298 -3516 -4245 -2721
rect -4141 -3454 -4131 -3401
rect -4078 -3454 -4068 -3401
rect -4308 -3569 -4298 -3516
rect -4245 -3569 -4235 -3516
rect -4721 -4689 -4687 -4181
rect -4632 -4390 -4598 -4128
rect -4652 -4443 -4642 -4390
rect -4589 -4443 -4579 -4390
rect -4298 -4506 -4245 -3569
rect -4308 -4559 -4298 -4506
rect -4245 -4559 -4235 -4506
rect -4632 -5319 -4598 -4999
rect -4652 -5372 -4642 -5319
rect -4589 -5372 -4579 -5319
rect -4298 -5416 -4245 -4559
rect -4130 -5233 -4077 -3454
rect -4140 -5286 -4130 -5233
rect -4077 -5286 -4067 -5233
rect -4308 -5469 -4298 -5416
rect -4245 -5469 -4235 -5416
rect -6946 -6016 -6912 -5869
rect -6966 -6069 -6956 -6016
rect -6903 -6069 -6893 -6016
rect -6768 -6131 -6734 -5868
rect -6590 -6016 -6556 -5868
rect -6611 -6069 -6601 -6016
rect -6548 -6069 -6538 -6016
rect -6788 -6184 -6778 -6131
rect -6725 -6184 -6715 -6131
rect -6412 -6248 -6378 -5868
rect -6234 -6016 -6200 -5868
rect -6254 -6069 -6244 -6016
rect -6191 -6069 -6181 -6016
rect -6056 -6131 -6022 -5869
rect -5878 -6016 -5844 -5868
rect -5898 -6069 -5888 -6016
rect -5835 -6069 -5825 -6016
rect -6075 -6184 -6065 -6131
rect -6012 -6184 -6002 -6131
rect -5700 -6248 -5666 -5868
rect -5522 -6016 -5488 -5868
rect -5542 -6069 -5532 -6016
rect -5479 -6069 -5469 -6016
rect -5344 -6131 -5310 -5868
rect -5166 -6016 -5132 -5868
rect -5185 -6069 -5175 -6016
rect -5122 -6069 -5112 -6016
rect -5364 -6184 -5354 -6131
rect -5301 -6184 -5291 -6131
rect -4988 -6247 -4954 -5868
rect -4810 -6016 -4776 -5868
rect -4830 -6069 -4820 -6016
rect -4767 -6069 -4757 -6016
rect -4298 -6131 -4245 -5469
rect -4308 -6184 -4298 -6131
rect -4245 -6184 -4235 -6131
rect -7508 -6301 -7498 -6248
rect -7445 -6301 -7435 -6248
rect -6431 -6301 -6421 -6248
rect -6368 -6301 -6358 -6248
rect -5720 -6301 -5710 -6248
rect -5657 -6301 -5647 -6248
rect -5008 -6300 -4998 -6247
rect -4945 -6300 -4935 -6247
rect -4988 -6301 -4954 -6300
rect -3864 -7147 -3830 -6757
rect -5628 -7181 -3830 -7147
rect -5628 -7325 -5594 -7181
rect -5544 -7274 -5500 -7181
rect -5450 -7325 -5416 -7181
rect -5366 -7280 -5322 -7181
rect -5188 -7280 -5144 -7181
rect -5094 -7326 -5060 -7181
rect -5010 -7280 -4966 -7181
rect -4832 -7280 -4788 -7181
rect -4738 -7326 -4704 -7181
rect -4654 -7280 -4610 -7181
rect -4476 -7280 -4432 -7181
rect -4382 -7326 -4348 -7181
rect -4298 -7280 -4254 -7181
rect -3717 -7240 -3683 -6753
rect -4026 -7274 -3683 -7240
rect -4026 -7330 -3992 -7274
rect -7466 -7698 -7422 -7664
rect -5628 -10624 -5594 -7580
rect -5544 -7790 -5500 -7664
rect -5544 -8340 -5500 -8214
rect -5544 -8890 -5500 -8764
rect -5544 -9440 -5500 -9314
rect -5544 -9990 -5500 -9864
rect -5544 -10540 -5500 -10414
rect -5450 -10624 -5416 -7580
rect -5366 -7790 -5322 -7664
rect -5366 -8340 -5322 -8214
rect -5366 -8890 -5322 -8764
rect -5366 -9440 -5322 -9314
rect -5366 -9990 -5322 -9864
rect -5366 -10540 -5322 -10414
rect -5272 -10624 -5238 -7580
rect -5188 -7790 -5144 -7664
rect -5188 -8340 -5144 -8214
rect -5188 -8890 -5144 -8764
rect -5188 -9440 -5144 -9314
rect -5188 -9990 -5144 -9864
rect -5188 -10540 -5144 -10414
rect -5094 -10624 -5060 -7581
rect -5010 -7791 -4966 -7665
rect -5010 -8340 -4966 -8214
rect -5010 -8890 -4966 -8764
rect -5010 -9440 -4966 -9314
rect -5010 -9990 -4966 -9864
rect -5010 -10540 -4966 -10414
rect -4916 -10624 -4882 -7580
rect -4832 -7790 -4788 -7664
rect -4832 -8340 -4788 -8214
rect -4832 -8890 -4788 -8764
rect -4832 -9440 -4788 -9314
rect -4832 -9990 -4788 -9864
rect -4832 -10540 -4788 -10414
rect -4738 -10624 -4704 -7580
rect -4654 -7790 -4610 -7664
rect -4654 -8340 -4610 -8214
rect -4654 -8890 -4610 -8764
rect -4654 -9440 -4610 -9314
rect -4654 -9990 -4610 -9864
rect -4654 -10540 -4610 -10414
rect -4560 -10624 -4526 -7580
rect -4476 -7790 -4432 -7664
rect -4476 -8340 -4432 -8214
rect -4476 -8890 -4432 -8764
rect -4476 -9440 -4432 -9314
rect -4476 -9990 -4432 -9864
rect -4476 -10540 -4432 -10414
rect -4382 -10624 -4348 -7580
rect -4298 -7790 -4254 -7664
rect -4298 -8340 -4254 -8214
rect -4298 -8890 -4254 -8764
rect -4298 -9440 -4254 -9314
rect -4298 -9990 -4254 -9864
rect -4298 -10540 -4254 -10414
rect -4204 -10624 -4170 -7580
rect -4120 -7790 -4076 -7664
rect -4120 -8340 -4076 -8214
rect -4120 -8890 -4076 -8764
rect -4120 -9440 -4076 -9314
rect -4120 -9990 -4076 -9864
rect -4120 -10540 -4076 -10414
rect -4026 -10624 -3992 -7580
rect -5272 -11020 -5238 -10881
rect -4916 -11020 -4882 -10880
rect -4560 -11020 -4526 -10880
rect -4204 -11020 -4170 -10880
rect -4120 -11020 -4076 -10964
rect -4026 -11020 -3992 -10880
rect -5272 -11054 -3611 -11020
rect -5512 -11224 -5502 -11171
rect -5449 -11224 -5439 -11171
rect -6976 -11465 -6077 -11412
rect -6024 -11465 -6014 -11412
rect -5636 -11465 -5626 -11412
rect -5573 -11465 -5563 -11412
rect -6233 -12015 -6223 -11962
rect -6170 -12015 -6160 -11962
rect -6976 -12805 -6426 -12752
rect -6373 -12805 -6363 -12752
rect -6223 -12955 -6170 -12015
rect -6077 -12645 -6024 -11465
rect -5922 -11528 -5877 -11512
rect -5922 -11600 -5876 -11528
rect -5817 -11568 -5778 -11512
rect -5617 -11562 -5583 -11465
rect -5824 -11600 -5778 -11568
rect -5492 -11600 -5458 -11224
rect -5010 -11225 -5000 -11172
rect -4947 -11225 -4937 -11172
rect -4512 -11224 -4502 -11171
rect -4449 -11224 -4439 -11171
rect -5386 -11341 -5376 -11288
rect -5323 -11341 -5313 -11288
rect -5137 -11341 -5127 -11288
rect -5074 -11341 -5064 -11288
rect -5367 -11568 -5333 -11341
rect -5117 -11568 -5083 -11341
rect -4992 -11600 -4958 -11225
rect -4887 -11465 -4877 -11412
rect -4824 -11465 -4814 -11412
rect -4637 -11465 -4627 -11412
rect -4574 -11465 -4564 -11412
rect -4867 -11568 -4833 -11465
rect -4617 -11568 -4583 -11465
rect -4492 -11600 -4458 -11224
rect -4387 -11341 -4377 -11288
rect -4324 -11341 -4314 -11288
rect -4367 -11568 -4333 -11341
rect -3938 -11342 -3928 -11289
rect -3875 -11342 -3865 -11289
rect -4172 -11600 -4126 -11512
rect -5824 -11640 -5626 -11600
rect -5574 -11640 -5376 -11600
rect -5324 -11640 -5126 -11600
rect -5074 -11640 -4876 -11600
rect -4823 -11640 -4625 -11600
rect -4574 -11640 -4376 -11600
rect -4324 -11640 -4126 -11600
rect -4074 -11612 -4028 -11512
rect -5818 -11840 -5632 -11800
rect -5574 -11840 -5376 -11800
rect -5324 -11840 -5126 -11800
rect -5074 -11840 -4876 -11800
rect -4825 -11840 -4627 -11800
rect -4574 -11840 -4376 -11800
rect -4324 -11840 -4126 -11800
rect -5744 -11962 -5704 -11840
rect -5761 -12015 -5751 -11962
rect -5698 -12015 -5688 -11962
rect -5495 -12280 -5455 -11840
rect -5245 -12089 -5205 -11840
rect -5261 -12142 -5251 -12089
rect -5198 -12142 -5188 -12089
rect -4995 -12280 -4955 -11840
rect -4746 -11962 -4706 -11840
rect -4762 -12015 -4752 -11962
rect -4699 -12015 -4689 -11962
rect -4495 -12280 -4455 -11840
rect -4244 -12089 -4204 -11840
rect -4261 -12142 -4251 -12089
rect -4198 -12142 -4188 -12089
rect -5824 -12320 -5626 -12280
rect -5574 -12320 -5376 -12280
rect -5324 -12320 -5126 -12280
rect -5074 -12320 -4876 -12280
rect -4824 -12320 -4626 -12280
rect -4574 -12320 -4376 -12280
rect -4324 -12320 -4126 -12280
rect -5922 -12608 -5876 -12508
rect -5824 -12520 -5626 -12480
rect -5574 -12520 -5376 -12480
rect -5324 -12520 -5126 -12480
rect -5074 -12520 -4876 -12480
rect -4824 -12520 -4626 -12480
rect -4574 -12520 -4376 -12480
rect -4324 -12520 -4126 -12480
rect -5824 -12608 -5778 -12520
rect -6087 -12698 -6077 -12645
rect -6024 -12698 -6014 -12645
rect -5720 -12857 -5686 -12520
rect -5617 -12752 -5583 -12552
rect -5367 -12645 -5333 -12552
rect -5386 -12698 -5376 -12645
rect -5323 -12698 -5313 -12645
rect -5636 -12805 -5626 -12752
rect -5573 -12805 -5563 -12752
rect -5740 -12910 -5730 -12857
rect -5677 -12910 -5667 -12857
rect -5240 -12955 -5206 -12520
rect -5117 -12645 -5083 -12552
rect -5136 -12698 -5126 -12645
rect -5073 -12698 -5063 -12645
rect -4867 -12752 -4833 -12552
rect -4887 -12805 -4877 -12752
rect -4824 -12805 -4814 -12752
rect -4742 -12857 -4708 -12520
rect -4617 -12752 -4583 -12552
rect -4367 -12645 -4333 -12552
rect -4386 -12698 -4376 -12645
rect -4323 -12698 -4313 -12645
rect -4637 -12805 -4627 -12752
rect -4574 -12805 -4564 -12752
rect -4762 -12910 -4752 -12857
rect -4699 -12910 -4689 -12857
rect -4240 -12955 -4206 -12520
rect -4172 -12608 -4126 -12520
rect -4074 -12608 -4028 -12508
rect -3928 -12752 -3875 -11342
rect -3798 -12142 -3788 -12089
rect -3735 -12142 -3725 -12089
rect -3938 -12805 -3928 -12752
rect -3875 -12805 -3865 -12752
rect -3928 -12806 -3875 -12805
rect -3788 -12857 -3735 -12142
rect -3798 -12910 -3788 -12857
rect -3735 -12910 -3725 -12857
rect -6233 -13008 -6223 -12955
rect -6170 -13008 -6160 -12955
rect -5260 -13008 -5250 -12955
rect -5197 -13008 -5187 -12955
rect -4260 -13008 -4250 -12955
rect -4197 -13008 -4187 -12955
rect -6965 -13160 -4303 -13126
rect -6028 -13294 -5994 -13160
rect -5939 -13250 -5905 -13160
rect -5850 -13294 -5816 -13160
rect -5761 -13250 -5727 -13160
rect -5583 -13250 -5549 -13160
rect -5405 -13250 -5371 -13160
rect -5227 -13250 -5193 -13160
rect -5049 -13250 -5015 -13160
rect -4871 -13250 -4837 -13160
rect -4693 -13250 -4659 -13160
rect -4515 -13250 -4481 -13160
rect -4337 -13250 -4303 -13160
rect -4248 -13160 -4036 -13126
rect -4248 -13294 -4214 -13160
rect -4159 -13244 -4125 -13160
rect -4070 -13294 -4036 -13160
rect -5850 -13695 -5816 -13551
rect -6169 -13748 -6159 -13695
rect -6106 -13748 -6096 -13695
rect -5870 -13748 -5860 -13695
rect -5807 -13748 -5797 -13695
rect -6159 -14382 -6106 -13748
rect -6028 -13859 -5816 -13825
rect -6027 -13993 -5993 -13859
rect -5939 -13950 -5905 -13859
rect -5850 -13994 -5816 -13859
rect -5761 -13910 -5727 -13600
rect -5672 -13994 -5638 -13550
rect -5583 -13935 -5549 -13619
rect -5494 -13801 -5460 -13550
rect -5514 -13854 -5504 -13801
rect -5451 -13854 -5441 -13801
rect -5405 -13933 -5371 -13617
rect -6169 -14435 -6159 -14382
rect -6106 -14435 -6096 -14382
rect -6159 -15093 -6106 -14435
rect -5850 -14488 -5816 -14250
rect -5870 -14541 -5860 -14488
rect -5807 -14541 -5797 -14488
rect -5761 -14617 -5727 -14301
rect -5672 -14703 -5638 -14250
rect -5583 -14624 -5549 -14308
rect -5494 -14381 -5460 -14250
rect -5514 -14434 -5504 -14381
rect -5451 -14434 -5441 -14381
rect -5405 -14631 -5371 -14315
rect -6028 -15085 -5994 -14949
rect -5939 -15085 -5905 -14994
rect -5850 -15085 -5816 -14950
rect -6169 -15146 -6159 -15093
rect -6106 -15146 -6096 -15093
rect -6028 -15119 -5816 -15085
rect -6159 -15907 -6106 -15146
rect -5850 -15194 -5816 -15119
rect -5870 -15247 -5860 -15194
rect -5807 -15247 -5797 -15194
rect -5761 -15326 -5727 -15010
rect -5672 -15394 -5638 -14950
rect -5583 -15328 -5549 -15012
rect -5494 -15093 -5460 -14950
rect -5514 -15146 -5504 -15093
rect -5451 -15146 -5441 -15093
rect -5405 -15327 -5371 -15011
rect -5316 -15394 -5282 -13550
rect -5227 -13932 -5193 -13616
rect -5138 -13695 -5104 -13551
rect -5157 -13748 -5147 -13695
rect -5094 -13748 -5084 -13695
rect -5049 -13932 -5015 -13616
rect -5227 -14629 -5193 -14313
rect -5138 -14489 -5104 -14250
rect -5158 -14542 -5148 -14489
rect -5095 -14542 -5085 -14489
rect -5049 -14630 -5015 -14314
rect -5227 -15327 -5193 -15011
rect -5138 -15194 -5104 -14951
rect -5158 -15247 -5148 -15194
rect -5095 -15247 -5085 -15194
rect -5049 -15327 -5015 -15011
rect -4960 -15394 -4926 -13550
rect -4871 -13931 -4837 -13615
rect -4782 -13801 -4748 -13550
rect -4801 -13854 -4791 -13801
rect -4738 -13854 -4728 -13801
rect -4693 -13930 -4659 -13614
rect -4871 -14630 -4837 -14314
rect -4782 -14381 -4748 -14250
rect -4802 -14434 -4792 -14381
rect -4739 -14434 -4729 -14381
rect -4693 -14629 -4659 -14313
rect -4871 -15327 -4837 -15011
rect -4782 -15093 -4748 -14950
rect -4802 -15146 -4792 -15093
rect -4739 -15146 -4729 -15093
rect -4693 -15327 -4659 -15011
rect -4604 -15394 -4570 -13550
rect -4515 -13930 -4481 -13614
rect -4426 -13695 -4392 -13550
rect -4446 -13748 -4436 -13695
rect -4383 -13748 -4373 -13695
rect -4337 -13928 -4303 -13612
rect -4248 -13825 -4214 -13550
rect -4159 -13650 -4125 -13600
rect -3664 -13801 -3611 -11054
rect -4248 -13859 -4036 -13825
rect -3946 -13854 -3936 -13801
rect -3883 -13854 -3611 -13801
rect -4515 -14627 -4481 -14311
rect -4426 -14489 -4392 -14251
rect -4445 -14541 -4435 -14489
rect -4383 -14541 -4373 -14489
rect -4337 -14627 -4303 -14311
rect -4515 -15327 -4481 -15011
rect -4426 -15194 -4392 -14950
rect -4446 -15247 -4436 -15194
rect -4383 -15247 -4373 -15194
rect -4337 -15327 -4303 -15011
rect -4248 -15085 -4214 -13859
rect -4159 -13950 -4125 -13859
rect -4070 -13994 -4036 -13859
rect -3936 -13906 -3883 -13854
rect -3935 -14489 -3883 -13906
rect -3945 -14541 -3935 -14489
rect -3883 -14541 -3873 -14489
rect -4159 -15085 -4125 -14994
rect -4070 -15085 -4036 -14950
rect -4248 -15119 -4036 -15085
rect -4248 -15394 -4214 -15119
rect -3935 -15195 -3883 -14541
rect -3945 -15247 -3935 -15195
rect -3883 -15247 -3873 -15195
rect -6028 -15786 -5994 -15650
rect -5939 -15786 -5905 -15694
rect -5850 -15786 -5816 -15650
rect -5672 -15786 -5638 -15650
rect -6028 -15820 -5816 -15786
rect -5850 -15907 -5816 -15820
rect -5692 -15839 -5682 -15786
rect -5629 -15839 -5619 -15786
rect -6169 -15960 -6159 -15907
rect -6106 -15960 -6096 -15907
rect -5869 -15960 -5859 -15907
rect -5806 -15960 -5796 -15907
rect -5494 -16018 -5460 -15651
rect -5316 -15786 -5282 -15650
rect -5336 -15839 -5326 -15786
rect -5273 -15839 -5263 -15786
rect -5138 -15907 -5104 -15651
rect -4960 -15786 -4926 -15651
rect -4980 -15839 -4970 -15786
rect -4917 -15839 -4907 -15786
rect -5158 -15960 -5148 -15907
rect -5095 -15960 -5085 -15907
rect -5514 -16071 -5504 -16018
rect -5451 -16071 -5441 -16018
rect -4970 -16449 -4917 -15839
rect -4782 -16018 -4748 -15651
rect -4604 -15786 -4570 -15651
rect -4624 -15839 -4614 -15786
rect -4561 -15839 -4551 -15786
rect -4426 -15907 -4392 -15650
rect -4248 -15786 -4214 -15650
rect -4159 -15786 -4125 -15694
rect -4070 -15786 -4036 -15650
rect -4268 -15839 -4258 -15786
rect -4205 -15839 -4036 -15786
rect -4447 -15960 -4437 -15907
rect -4384 -15960 -4374 -15907
rect -3935 -16018 -3883 -15247
rect -4802 -16071 -4792 -16018
rect -4739 -16071 -4729 -16018
rect -3945 -16070 -3935 -16018
rect -3883 -16070 -3873 -16018
<< via1 >>
rect -6867 -1963 -6814 -1910
rect -6689 -1963 -6636 -1910
rect -6510 -1963 -6457 -1910
rect -6333 -1963 -6280 -1910
rect -6155 -1963 -6102 -1910
rect -5976 -1963 -5923 -1910
rect -5799 -1963 -5746 -1910
rect -5621 -1963 -5568 -1910
rect -5443 -1963 -5390 -1910
rect -5265 -1963 -5212 -1910
rect -5086 -1963 -5033 -1910
rect -4909 -1963 -4856 -1910
rect -7498 -2582 -7445 -2529
rect -7625 -3454 -7572 -3401
rect -7044 -2833 -6991 -2780
rect -7134 -3454 -7081 -3401
rect -7498 -3693 -7445 -3640
rect -7498 -4324 -7445 -4271
rect -7134 -4443 -7081 -4390
rect -7498 -5194 -7445 -5141
rect -7625 -5375 -7572 -5322
rect -7134 -5285 -7081 -5232
rect -6777 -2583 -6724 -2530
rect -6866 -2833 -6813 -2780
rect -6777 -3569 -6724 -3516
rect -6778 -4324 -6725 -4271
rect -6777 -5468 -6724 -5415
rect -6421 -2721 -6368 -2668
rect -6422 -3693 -6369 -3640
rect -6422 -4559 -6369 -4506
rect -6422 -5194 -6369 -5141
rect -6066 -2583 -6013 -2530
rect -6066 -3454 -6013 -3401
rect -6066 -4443 -6013 -4390
rect -6066 -5286 -6013 -5233
rect -5710 -2721 -5657 -2668
rect -5710 -3454 -5657 -3401
rect -5709 -4443 -5656 -4390
rect -5710 -5375 -5657 -5322
rect -5354 -2583 -5301 -2530
rect -5353 -3693 -5300 -3640
rect -5353 -4559 -5300 -4506
rect -5353 -5194 -5300 -5141
rect -4998 -2721 -4945 -2668
rect -4908 -2833 -4855 -2780
rect -4998 -3569 -4945 -3516
rect -4998 -4324 -4945 -4271
rect -4997 -5468 -4944 -5415
rect -4298 -2721 -4245 -2668
rect -4731 -2833 -4678 -2780
rect -4642 -3454 -4589 -3401
rect -4131 -3454 -4078 -3401
rect -4298 -3569 -4245 -3516
rect -4642 -4443 -4589 -4390
rect -4298 -4559 -4245 -4506
rect -4642 -5372 -4589 -5319
rect -4130 -5286 -4077 -5233
rect -4298 -5469 -4245 -5416
rect -6956 -6069 -6903 -6016
rect -6601 -6069 -6548 -6016
rect -6778 -6184 -6725 -6131
rect -6244 -6069 -6191 -6016
rect -5888 -6069 -5835 -6016
rect -6065 -6184 -6012 -6131
rect -5532 -6069 -5479 -6016
rect -5175 -6069 -5122 -6016
rect -5354 -6184 -5301 -6131
rect -4820 -6069 -4767 -6016
rect -4298 -6184 -4245 -6131
rect -7498 -6301 -7445 -6248
rect -6421 -6301 -6368 -6248
rect -5710 -6301 -5657 -6248
rect -4998 -6300 -4945 -6247
rect -5502 -11224 -5449 -11171
rect -6077 -11465 -6024 -11412
rect -5626 -11465 -5573 -11412
rect -6223 -12015 -6170 -11962
rect -6426 -12805 -6373 -12752
rect -5000 -11225 -4947 -11172
rect -4502 -11224 -4449 -11171
rect -5376 -11341 -5323 -11288
rect -5127 -11341 -5074 -11288
rect -4877 -11465 -4824 -11412
rect -4627 -11465 -4574 -11412
rect -4377 -11341 -4324 -11288
rect -3928 -11342 -3875 -11289
rect -5751 -12015 -5698 -11962
rect -5251 -12142 -5198 -12089
rect -4752 -12015 -4699 -11962
rect -4251 -12142 -4198 -12089
rect -6077 -12698 -6024 -12645
rect -5376 -12698 -5323 -12645
rect -5626 -12805 -5573 -12752
rect -5730 -12910 -5677 -12857
rect -5126 -12698 -5073 -12645
rect -4877 -12805 -4824 -12752
rect -4376 -12698 -4323 -12645
rect -4627 -12805 -4574 -12752
rect -4752 -12910 -4699 -12857
rect -3788 -12142 -3735 -12089
rect -3928 -12805 -3875 -12752
rect -3788 -12910 -3735 -12857
rect -6223 -13008 -6170 -12955
rect -5250 -13008 -5197 -12955
rect -4250 -13008 -4197 -12955
rect -6159 -13748 -6106 -13695
rect -5860 -13748 -5807 -13695
rect -5504 -13854 -5451 -13801
rect -6159 -14435 -6106 -14382
rect -5860 -14541 -5807 -14488
rect -5504 -14434 -5451 -14381
rect -6159 -15146 -6106 -15093
rect -5860 -15247 -5807 -15194
rect -5504 -15146 -5451 -15093
rect -5147 -13748 -5094 -13695
rect -5148 -14542 -5095 -14489
rect -5148 -15247 -5095 -15194
rect -4791 -13854 -4738 -13801
rect -4792 -14434 -4739 -14381
rect -4792 -15146 -4739 -15093
rect -4436 -13748 -4383 -13695
rect -3936 -13854 -3883 -13801
rect -4435 -14541 -4383 -14489
rect -4436 -15247 -4383 -15194
rect -3935 -14541 -3883 -14489
rect -3935 -15247 -3883 -15195
rect -5682 -15839 -5629 -15786
rect -6159 -15960 -6106 -15907
rect -5859 -15960 -5806 -15907
rect -5326 -15839 -5273 -15786
rect -4970 -15839 -4917 -15786
rect -5148 -15960 -5095 -15907
rect -5504 -16071 -5451 -16018
rect -4614 -15839 -4561 -15786
rect -4258 -15839 -4205 -15786
rect -4437 -15960 -4384 -15907
rect -4792 -16071 -4739 -16018
rect -3935 -16070 -3883 -16018
<< metal2 >>
rect -6867 -1910 -6814 -1900
rect -6689 -1910 -6636 -1900
rect -6510 -1910 -6457 -1900
rect -6333 -1910 -6280 -1900
rect -6155 -1910 -6102 -1900
rect -5976 -1910 -5923 -1900
rect -5799 -1910 -5746 -1900
rect -5621 -1910 -5568 -1900
rect -5443 -1910 -5390 -1900
rect -5265 -1910 -5212 -1900
rect -5086 -1910 -5033 -1900
rect -4909 -1910 -4856 -1900
rect -6814 -1963 -6689 -1910
rect -6636 -1963 -6510 -1910
rect -6457 -1963 -6333 -1910
rect -6280 -1963 -6155 -1910
rect -6102 -1963 -5976 -1910
rect -5923 -1963 -5799 -1910
rect -5746 -1963 -5621 -1910
rect -5568 -1963 -5443 -1910
rect -5390 -1963 -5265 -1910
rect -5212 -1963 -5086 -1910
rect -5033 -1963 -4909 -1910
rect -6867 -1973 -6814 -1963
rect -6689 -1973 -6636 -1963
rect -6510 -1973 -6457 -1963
rect -6333 -1973 -6280 -1963
rect -6155 -1973 -6102 -1963
rect -5976 -1973 -5923 -1963
rect -5799 -1973 -5746 -1963
rect -5621 -1973 -5568 -1963
rect -5443 -1973 -5390 -1963
rect -5265 -1973 -5212 -1963
rect -5086 -1973 -5033 -1963
rect -4909 -1973 -4856 -1963
rect -7498 -2529 -7445 -2519
rect -6777 -2529 -6724 -2520
rect -7445 -2530 -6724 -2529
rect -6066 -2530 -6013 -2520
rect -5354 -2530 -5301 -2520
rect -7445 -2582 -6777 -2530
rect -7498 -2592 -7445 -2582
rect -6724 -2583 -6066 -2530
rect -6013 -2583 -5354 -2530
rect -6777 -2593 -6724 -2583
rect -6066 -2593 -6013 -2583
rect -5354 -2593 -5301 -2583
rect -6421 -2668 -6368 -2658
rect -5710 -2668 -5657 -2658
rect -4998 -2668 -4945 -2658
rect -4298 -2668 -4245 -2658
rect -6368 -2721 -5710 -2668
rect -5657 -2721 -4998 -2668
rect -4945 -2721 -4298 -2668
rect -6421 -2731 -6368 -2721
rect -5710 -2731 -5657 -2721
rect -4998 -2731 -4945 -2721
rect -4298 -2731 -4245 -2721
rect -7044 -2780 -6991 -2770
rect -6866 -2780 -6813 -2770
rect -6991 -2833 -6866 -2780
rect -7044 -2843 -6991 -2833
rect -6866 -2843 -6813 -2833
rect -4908 -2780 -4855 -2770
rect -4731 -2780 -4678 -2770
rect -4855 -2833 -4731 -2780
rect -4908 -2843 -4855 -2833
rect -4731 -2843 -4678 -2833
rect -7625 -3401 -7572 -3391
rect -7134 -3401 -7081 -3391
rect -6066 -3401 -6013 -3391
rect -7572 -3454 -7134 -3401
rect -7081 -3454 -6066 -3401
rect -7625 -3464 -7572 -3454
rect -7134 -3464 -7081 -3454
rect -6066 -3464 -6013 -3454
rect -5710 -3401 -5657 -3391
rect -4642 -3401 -4589 -3391
rect -4131 -3401 -4078 -3391
rect -5657 -3454 -4642 -3401
rect -4589 -3454 -4131 -3401
rect -5710 -3464 -5657 -3454
rect -4642 -3464 -4589 -3454
rect -4131 -3464 -4078 -3454
rect -6777 -3516 -6724 -3506
rect -4998 -3516 -4945 -3506
rect -4298 -3516 -4245 -3506
rect -6724 -3569 -4998 -3516
rect -4945 -3569 -4298 -3516
rect -6777 -3579 -6724 -3569
rect -4998 -3579 -4945 -3569
rect -4298 -3579 -4245 -3569
rect -7498 -3640 -7445 -3630
rect -6422 -3640 -6369 -3630
rect -5353 -3640 -5300 -3630
rect -7445 -3693 -6422 -3640
rect -6369 -3693 -5353 -3640
rect -7498 -3703 -7445 -3693
rect -6422 -3703 -6369 -3693
rect -5353 -3703 -5300 -3693
rect -7498 -4271 -7445 -4261
rect -6778 -4271 -6725 -4261
rect -4998 -4271 -4945 -4261
rect -7445 -4324 -6778 -4271
rect -6725 -4324 -4998 -4271
rect -7498 -4334 -7445 -4324
rect -6778 -4334 -6725 -4324
rect -4998 -4334 -4945 -4324
rect -7134 -4390 -7081 -4380
rect -6066 -4390 -6013 -4380
rect -5709 -4390 -5656 -4380
rect -4642 -4390 -4589 -4380
rect -7081 -4443 -6066 -4390
rect -6013 -4443 -5709 -4390
rect -5656 -4443 -4642 -4390
rect -4589 -4443 -3312 -4390
rect -7134 -4453 -7081 -4443
rect -6066 -4453 -6013 -4443
rect -5709 -4453 -5656 -4443
rect -4642 -4453 -4589 -4443
rect -6422 -4506 -6369 -4496
rect -5353 -4506 -5300 -4496
rect -4298 -4506 -4245 -4496
rect -6369 -4559 -5353 -4506
rect -5300 -4559 -4298 -4506
rect -6422 -4569 -6369 -4559
rect -5353 -4569 -5300 -4559
rect -4298 -4569 -4245 -4559
rect -7498 -5141 -7445 -5131
rect -6422 -5141 -6369 -5131
rect -7445 -5187 -6422 -5147
rect -7498 -5204 -7445 -5194
rect -5353 -5141 -5300 -5131
rect -6369 -5188 -5353 -5148
rect -6422 -5204 -6369 -5194
rect -5353 -5204 -5300 -5194
rect -7134 -5232 -7081 -5222
rect -6066 -5233 -6013 -5223
rect -7081 -5279 -6066 -5239
rect -7134 -5295 -7081 -5285
rect -4130 -5233 -4077 -5223
rect -6013 -5279 -4130 -5239
rect -6066 -5296 -6013 -5286
rect -4130 -5296 -4077 -5286
rect -7625 -5322 -7572 -5312
rect -5710 -5322 -5657 -5312
rect -7572 -5369 -5710 -5329
rect -7625 -5385 -7572 -5375
rect -4642 -5319 -4589 -5309
rect -5657 -5369 -4642 -5329
rect -5710 -5385 -5657 -5375
rect -4642 -5382 -4589 -5372
rect -6777 -5415 -6724 -5405
rect -4997 -5415 -4944 -5405
rect -6724 -5462 -4997 -5422
rect -6777 -5478 -6724 -5468
rect -4298 -5416 -4245 -5406
rect -4944 -5462 -4298 -5422
rect -4997 -5478 -4944 -5468
rect -4298 -5479 -4245 -5469
rect -6956 -6016 -6903 -6006
rect -6601 -6016 -6548 -6006
rect -6244 -6016 -6191 -6006
rect -5888 -6016 -5835 -6006
rect -5532 -6016 -5479 -6006
rect -5175 -6016 -5122 -6006
rect -4820 -6016 -4767 -6006
rect -6903 -6069 -6601 -6016
rect -6548 -6069 -6244 -6016
rect -6191 -6069 -5888 -6016
rect -5835 -6069 -5532 -6016
rect -5479 -6069 -5175 -6016
rect -5122 -6069 -4820 -6016
rect -6956 -6079 -6903 -6069
rect -6601 -6079 -6548 -6069
rect -6244 -6079 -6191 -6069
rect -5888 -6079 -5835 -6069
rect -5532 -6079 -5479 -6069
rect -5175 -6079 -5122 -6069
rect -4820 -6079 -4767 -6069
rect -6778 -6131 -6725 -6121
rect -6065 -6131 -6012 -6121
rect -5354 -6131 -5301 -6121
rect -4298 -6131 -4245 -6121
rect -6725 -6184 -6065 -6131
rect -6012 -6184 -5354 -6131
rect -5301 -6184 -4298 -6131
rect -6778 -6194 -6725 -6184
rect -6065 -6194 -6012 -6184
rect -5354 -6194 -5301 -6184
rect -4298 -6194 -4245 -6184
rect -7498 -6248 -7445 -6238
rect -6421 -6248 -6368 -6238
rect -5710 -6248 -5657 -6238
rect -4998 -6247 -4945 -6237
rect -7445 -6301 -6421 -6248
rect -6368 -6301 -5710 -6248
rect -5657 -6300 -4998 -6248
rect -5657 -6301 -4945 -6300
rect -7498 -6311 -7445 -6301
rect -6421 -6311 -6368 -6301
rect -5710 -6311 -5657 -6301
rect -4998 -6310 -4945 -6301
rect -5502 -11171 -5449 -11161
rect -5000 -11171 -4947 -11162
rect -4502 -11171 -4449 -11161
rect -5449 -11172 -4502 -11171
rect -5449 -11224 -5000 -11172
rect -5502 -11234 -5449 -11224
rect -4947 -11224 -4502 -11172
rect -5000 -11235 -4947 -11225
rect -4502 -11234 -4449 -11224
rect -5376 -11288 -5323 -11278
rect -5127 -11288 -5074 -11278
rect -4377 -11288 -4324 -11278
rect -3928 -11288 -3875 -11279
rect -5323 -11341 -5127 -11288
rect -5074 -11341 -4377 -11288
rect -4324 -11289 -3875 -11288
rect -4324 -11341 -3928 -11289
rect -5376 -11351 -5323 -11341
rect -5127 -11351 -5074 -11341
rect -4377 -11351 -4324 -11341
rect -3928 -11352 -3875 -11342
rect -6077 -11412 -6024 -11402
rect -5626 -11412 -5573 -11402
rect -4877 -11412 -4824 -11402
rect -4627 -11412 -4574 -11402
rect -6024 -11465 -5626 -11412
rect -5573 -11465 -4877 -11412
rect -4824 -11465 -4627 -11412
rect -6077 -11475 -6024 -11465
rect -5626 -11475 -5573 -11465
rect -4877 -11475 -4824 -11465
rect -4627 -11475 -4574 -11465
rect -6223 -11962 -6170 -11952
rect -5751 -11962 -5698 -11952
rect -4752 -11962 -4699 -11952
rect -6170 -12015 -5751 -11962
rect -5698 -12015 -4752 -11962
rect -6223 -12025 -6170 -12015
rect -5751 -12025 -5698 -12015
rect -4752 -12025 -4699 -12015
rect -5251 -12089 -5198 -12079
rect -4251 -12089 -4198 -12079
rect -3788 -12089 -3735 -12079
rect -3542 -12089 -3489 -6756
rect -5198 -12142 -4251 -12089
rect -4198 -12142 -3788 -12089
rect -3735 -12142 -3489 -12089
rect -5251 -12152 -5198 -12142
rect -4251 -12152 -4198 -12142
rect -3788 -12152 -3735 -12142
rect -6077 -12645 -6024 -12635
rect -5376 -12645 -5323 -12635
rect -5126 -12645 -5073 -12635
rect -4376 -12645 -4323 -12635
rect -6024 -12698 -5376 -12645
rect -5323 -12698 -5126 -12645
rect -5073 -12698 -4376 -12645
rect -6077 -12708 -6024 -12698
rect -5376 -12708 -5323 -12698
rect -5126 -12708 -5073 -12698
rect -4376 -12708 -4323 -12698
rect -6426 -12752 -6373 -12742
rect -5626 -12752 -5573 -12742
rect -4877 -12752 -4824 -12742
rect -4627 -12752 -4574 -12742
rect -3928 -12752 -3875 -12742
rect -6373 -12805 -5626 -12752
rect -5573 -12805 -4877 -12752
rect -4824 -12805 -4627 -12752
rect -4574 -12805 -3928 -12752
rect -6426 -12815 -6373 -12805
rect -5626 -12815 -5573 -12805
rect -4877 -12815 -4824 -12805
rect -4627 -12815 -4574 -12805
rect -3928 -12815 -3875 -12805
rect -5730 -12857 -5677 -12847
rect -4752 -12857 -4699 -12847
rect -3788 -12857 -3735 -12847
rect -5677 -12910 -4752 -12857
rect -4699 -12910 -3788 -12857
rect -5730 -12920 -5677 -12910
rect -4752 -12920 -4699 -12910
rect -3788 -12920 -3735 -12910
rect -6223 -12955 -6170 -12945
rect -5250 -12955 -5197 -12945
rect -4250 -12955 -4197 -12945
rect -3432 -12955 -3379 -6747
rect -6170 -13008 -5250 -12955
rect -5197 -13008 -4250 -12955
rect -4197 -13008 -3379 -12955
rect -6223 -13018 -6170 -13008
rect -5250 -13018 -5197 -13008
rect -4250 -13018 -4197 -13008
rect -6159 -13695 -6106 -13685
rect -5860 -13695 -5807 -13685
rect -5147 -13695 -5094 -13685
rect -4436 -13695 -4383 -13685
rect -6106 -13748 -5860 -13695
rect -5807 -13748 -5147 -13695
rect -5094 -13748 -4436 -13695
rect -6159 -13758 -6106 -13748
rect -5860 -13758 -5807 -13748
rect -5147 -13758 -5094 -13748
rect -4436 -13758 -4383 -13748
rect -5504 -13801 -5451 -13791
rect -4791 -13801 -4738 -13791
rect -3936 -13801 -3883 -13791
rect -5451 -13854 -4791 -13801
rect -4738 -13854 -3936 -13801
rect -5504 -13864 -5451 -13854
rect -4791 -13864 -4738 -13854
rect -3936 -13864 -3883 -13854
rect -6159 -14381 -6106 -14372
rect -5504 -14381 -5451 -14371
rect -4792 -14381 -4739 -14371
rect -6159 -14382 -5504 -14381
rect -6106 -14434 -5504 -14382
rect -5451 -14434 -4792 -14381
rect -6159 -14445 -6106 -14435
rect -5504 -14444 -5451 -14434
rect -4792 -14444 -4739 -14434
rect -5860 -14488 -5807 -14478
rect -5148 -14489 -5095 -14479
rect -4435 -14489 -4383 -14479
rect -3935 -14489 -3883 -14479
rect -5807 -14541 -5148 -14489
rect -5860 -14551 -5807 -14541
rect -5095 -14541 -4435 -14489
rect -4383 -14541 -3935 -14489
rect -5148 -14552 -5095 -14542
rect -4435 -14551 -4383 -14541
rect -3935 -14551 -3883 -14541
rect -6159 -15093 -6106 -15083
rect -5504 -15093 -5451 -15083
rect -4792 -15093 -4739 -15083
rect -6106 -15146 -5504 -15093
rect -5451 -15146 -4792 -15093
rect -6159 -15156 -6106 -15146
rect -5504 -15156 -5451 -15146
rect -4792 -15156 -4739 -15146
rect -5860 -15194 -5807 -15184
rect -5148 -15194 -5095 -15184
rect -4436 -15194 -4383 -15184
rect -3935 -15194 -3883 -15185
rect -5807 -15247 -5148 -15194
rect -5095 -15246 -4436 -15194
rect -5860 -15257 -5807 -15247
rect -5148 -15257 -5095 -15247
rect -4383 -15195 -3883 -15194
rect -4383 -15246 -3935 -15195
rect -4436 -15257 -4383 -15247
rect -3935 -15257 -3883 -15247
rect -5682 -15786 -5629 -15776
rect -5326 -15786 -5273 -15776
rect -4970 -15786 -4917 -15776
rect -4614 -15786 -4561 -15776
rect -4258 -15786 -4205 -15776
rect -5629 -15839 -5326 -15786
rect -5273 -15839 -4970 -15786
rect -4917 -15839 -4614 -15786
rect -4561 -15839 -4258 -15786
rect -5682 -15849 -5629 -15839
rect -5326 -15849 -5273 -15839
rect -4970 -15849 -4917 -15839
rect -4614 -15849 -4561 -15839
rect -4258 -15849 -4205 -15839
rect -6159 -15907 -6106 -15897
rect -5859 -15907 -5806 -15897
rect -5148 -15907 -5095 -15897
rect -4437 -15907 -4384 -15897
rect -6106 -15960 -5859 -15907
rect -5806 -15960 -5148 -15907
rect -5095 -15960 -4437 -15907
rect -6159 -15970 -6106 -15960
rect -5859 -15970 -5806 -15960
rect -5148 -15970 -5095 -15960
rect -4437 -15970 -4384 -15960
rect -5504 -16018 -5451 -16008
rect -4792 -16018 -4739 -16008
rect -3935 -16018 -3883 -16008
rect -5451 -16070 -4792 -16018
rect -5504 -16081 -5451 -16071
rect -4739 -16070 -3935 -16018
rect -4792 -16081 -4739 -16071
rect -3935 -16080 -3883 -16070
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_0
timestamp 1653033955
transform 1 0 -5032 0 1 -13422
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_1
timestamp 1653033955
transform 1 0 -5032 0 1 -14122
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_2
timestamp 1653033955
transform 1 0 -5032 0 1 -14822
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_3
timestamp 1653033955
transform 1 0 -5032 0 1 -15522
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_HU75T7  sky130_fd_pr__nfet_01v8_HU75T7_0
timestamp 1653034865
transform 1 0 -7088 0 1 -7452
box -652 -228 652 228
use sky130_fd_pr__nfet_01v8_HU75T7  sky130_fd_pr__nfet_01v8_HU75T7_1
timestamp 1653034865
transform 1 0 -7088 0 1 -8222
box -652 -228 652 228
use sky130_fd_pr__nfet_01v8_HU75T7  sky130_fd_pr__nfet_01v8_HU75T7_2
timestamp 1653034865
transform 1 0 -7088 0 1 -8992
box -652 -228 652 228
use sky130_fd_pr__nfet_01v8_HU75T7  sky130_fd_pr__nfet_01v8_HU75T7_3
timestamp 1653034865
transform 1 0 -7088 0 1 -9762
box -652 -228 652 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_0
timestamp 1653030110
transform 1 0 9 0 1 -7460
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_1
timestamp 1653030110
transform 1 0 9 0 1 -8135
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_2
timestamp 1653030110
transform 1 0 9 0 1 -8810
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_3
timestamp 1653030110
transform 1 0 9 0 1 -9485
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_4
timestamp 1653030110
transform 1 0 9 0 1 -10160
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_5
timestamp 1653030110
transform 1 0 9 0 1 -10835
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_6
timestamp 1653030110
transform 1 0 9 0 1 -11510
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_7
timestamp 1653030110
transform 1 0 9 0 1 -12185
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_8
timestamp 1653030110
transform 1 0 9 0 1 -12860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_9
timestamp 1653030110
transform 1 0 9 0 1 -13535
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_10
timestamp 1653030110
transform 1 0 9 0 1 -14210
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_11
timestamp 1653030110
transform 1 0 9 0 1 -14885
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_12
timestamp 1653030110
transform 1 0 9 0 1 -15560
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_0
timestamp 1653028559
transform 1 0 -5850 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_1
timestamp 1653028559
transform 1 0 -5850 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_2
timestamp 1653028559
transform 1 0 -5600 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_3
timestamp 1653028559
transform 1 0 -5350 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_4
timestamp 1653028559
transform 1 0 -5100 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_5
timestamp 1653028559
transform 1 0 -4850 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_6
timestamp 1653028559
transform 1 0 -4600 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_7
timestamp 1653028559
transform 1 0 -4350 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_8
timestamp 1653028559
transform 1 0 -4100 0 1 -12400
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_9
timestamp 1653028559
transform 1 0 -5600 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_10
timestamp 1653028559
transform 1 0 -5350 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_11
timestamp 1653028559
transform 1 0 -5100 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_12
timestamp 1653028559
transform 1 0 -4850 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_13
timestamp 1653028559
transform 1 0 -4600 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_14
timestamp 1653028559
transform 1 0 -4350 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_15
timestamp 1653028559
transform 1 0 -4100 0 1 -11720
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_0
timestamp 1653032550
transform 1 0 -4810 0 1 -7452
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_1
timestamp 1653032550
transform 1 0 -4810 0 1 -8002
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_2
timestamp 1653032550
transform 1 0 -4810 0 1 -8552
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_3
timestamp 1653032550
transform 1 0 -4810 0 1 -9102
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_4
timestamp 1653032550
transform 1 0 -4810 0 1 -9652
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_5
timestamp 1653032550
transform 1 0 -4810 0 1 -10202
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_6
timestamp 1653032550
transform 1 0 -4810 0 1 -10752
box -830 -228 830 228
use sky130_fd_pr__pfet_01v8_ESNDBA  sky130_fd_pr__pfet_01v8_ESNDBA_0
timestamp 1653026387
transform 1 0 -924 0 1 -3012
box -1578 -240 1578 240
use sky130_fd_pr__pfet_01v8_ESNDBA  sky130_fd_pr__pfet_01v8_ESNDBA_1
timestamp 1653026387
transform 1 0 -924 0 1 -3912
box -1578 -240 1578 240
use sky130_fd_pr__pfet_01v8_ESNDBA  sky130_fd_pr__pfet_01v8_ESNDBA_2
timestamp 1653026387
transform 1 0 -924 0 1 -4812
box -1578 -240 1578 240
use sky130_fd_pr__pfet_01v8_ESNDBA  sky130_fd_pr__pfet_01v8_ESNDBA_3
timestamp 1653026387
transform 1 0 -924 0 1 -5712
box -1578 -240 1578 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_0
timestamp 1653025074
transform 1 0 -5861 0 1 -2260
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_1
timestamp 1653025074
transform 1 0 -5861 0 1 -3130
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_2
timestamp 1653025074
transform 1 0 -5861 0 1 -4000
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_3
timestamp 1653025074
transform 1 0 -5861 0 1 -4870
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_4
timestamp 1653025074
transform 1 0 -5861 0 1 -5740
box -1489 -240 1489 240
<< labels >>
flabel metal1 -6957 -13145 -6957 -13145 1 FreeSans 1200 0 0 0 i_bias
flabel metal1 -4277 -7165 -4277 -7165 1 FreeSans 1200 0 0 0 bias_b
flabel metal1 -3636 -11223 -3636 -11223 1 FreeSans 1200 0 0 0 bias_c
flabel metal1 -6950 -11441 -6950 -11441 1 FreeSans 1200 0 0 0 ip
flabel metal1 -6952 -12780 -6952 -12780 1 FreeSans 1200 0 0 0 in
<< end >>
