magic
tech sky130A
timestamp 1654517900
<< nmos >>
rect -697 -70 -637 70
rect -608 -70 -548 70
rect -519 -70 -459 70
rect -430 -70 -370 70
rect -341 -70 -281 70
rect -252 -70 -192 70
rect -163 -70 -103 70
rect -74 -70 -14 70
rect 14 -70 74 70
rect 103 -70 163 70
rect 192 -70 252 70
rect 281 -70 341 70
rect 370 -70 430 70
rect 459 -70 519 70
rect 548 -70 608 70
rect 637 -70 697 70
<< ndiff >>
rect -726 64 -697 70
rect -726 -64 -720 64
rect -703 -64 -697 64
rect -726 -70 -697 -64
rect -637 64 -608 70
rect -637 -64 -631 64
rect -614 -64 -608 64
rect -637 -70 -608 -64
rect -548 64 -519 70
rect -548 -64 -542 64
rect -525 -64 -519 64
rect -548 -70 -519 -64
rect -459 64 -430 70
rect -459 -64 -453 64
rect -436 -64 -430 64
rect -459 -70 -430 -64
rect -370 64 -341 70
rect -370 -64 -364 64
rect -347 -64 -341 64
rect -370 -70 -341 -64
rect -281 64 -252 70
rect -281 -64 -275 64
rect -258 -64 -252 64
rect -281 -70 -252 -64
rect -192 64 -163 70
rect -192 -64 -186 64
rect -169 -64 -163 64
rect -192 -70 -163 -64
rect -103 64 -74 70
rect -103 -64 -97 64
rect -80 -64 -74 64
rect -103 -70 -74 -64
rect -14 64 14 70
rect -14 -64 -8 64
rect 8 -64 14 64
rect -14 -70 14 -64
rect 74 64 103 70
rect 74 -64 80 64
rect 97 -64 103 64
rect 74 -70 103 -64
rect 163 64 192 70
rect 163 -64 169 64
rect 186 -64 192 64
rect 163 -70 192 -64
rect 252 64 281 70
rect 252 -64 258 64
rect 275 -64 281 64
rect 252 -70 281 -64
rect 341 64 370 70
rect 341 -64 347 64
rect 364 -64 370 64
rect 341 -70 370 -64
rect 430 64 459 70
rect 430 -64 436 64
rect 453 -64 459 64
rect 430 -70 459 -64
rect 519 64 548 70
rect 519 -64 525 64
rect 542 -64 548 64
rect 519 -70 548 -64
rect 608 64 637 70
rect 608 -64 614 64
rect 631 -64 637 64
rect 608 -70 637 -64
rect 697 64 726 70
rect 697 -64 703 64
rect 720 -64 726 64
rect 697 -70 726 -64
<< ndiffc >>
rect -720 -64 -703 64
rect -631 -64 -614 64
rect -542 -64 -525 64
rect -453 -64 -436 64
rect -364 -64 -347 64
rect -275 -64 -258 64
rect -186 -64 -169 64
rect -97 -64 -80 64
rect -8 -64 8 64
rect 80 -64 97 64
rect 169 -64 186 64
rect 258 -64 275 64
rect 347 -64 364 64
rect 436 -64 453 64
rect 525 -64 542 64
rect 614 -64 631 64
rect 703 -64 720 64
<< poly >>
rect -686 106 -648 114
rect -686 97 -678 106
rect -697 89 -678 97
rect -656 97 -648 106
rect -597 106 -559 114
rect -597 97 -589 106
rect -656 89 -637 97
rect -697 70 -637 89
rect -608 89 -589 97
rect -567 97 -559 106
rect -508 106 -470 114
rect -508 97 -500 106
rect -567 89 -548 97
rect -608 70 -548 89
rect -519 89 -500 97
rect -478 97 -470 106
rect -419 106 -381 114
rect -419 97 -411 106
rect -478 89 -459 97
rect -519 70 -459 89
rect -430 89 -411 97
rect -389 97 -381 106
rect -330 106 -292 114
rect -330 97 -322 106
rect -389 89 -370 97
rect -430 70 -370 89
rect -341 89 -322 97
rect -300 97 -292 106
rect -241 106 -203 114
rect -241 97 -233 106
rect -300 89 -281 97
rect -341 70 -281 89
rect -252 89 -233 97
rect -211 97 -203 106
rect -152 106 -114 114
rect -152 97 -144 106
rect -211 89 -192 97
rect -252 70 -192 89
rect -163 89 -144 97
rect -122 97 -114 106
rect -63 106 -25 114
rect -63 97 -55 106
rect -122 89 -103 97
rect -163 70 -103 89
rect -74 89 -55 97
rect -33 97 -25 106
rect 25 106 63 114
rect 25 97 33 106
rect -33 89 -14 97
rect -74 70 -14 89
rect 14 89 33 97
rect 55 97 63 106
rect 114 106 152 114
rect 114 97 122 106
rect 55 89 74 97
rect 14 70 74 89
rect 103 89 122 97
rect 144 97 152 106
rect 203 106 241 114
rect 203 97 211 106
rect 144 89 163 97
rect 103 70 163 89
rect 192 89 211 97
rect 233 97 241 106
rect 292 106 330 114
rect 292 97 300 106
rect 233 89 252 97
rect 192 70 252 89
rect 281 89 300 97
rect 322 97 330 106
rect 381 106 419 114
rect 381 97 389 106
rect 322 89 341 97
rect 281 70 341 89
rect 370 89 389 97
rect 411 97 419 106
rect 470 106 508 114
rect 470 97 478 106
rect 411 89 430 97
rect 370 70 430 89
rect 459 89 478 97
rect 500 97 508 106
rect 559 106 597 114
rect 559 97 567 106
rect 500 89 519 97
rect 459 70 519 89
rect 548 89 567 97
rect 589 97 597 106
rect 648 106 686 114
rect 648 97 656 106
rect 589 89 608 97
rect 548 70 608 89
rect 637 89 656 97
rect 678 97 686 106
rect 678 89 697 97
rect 637 70 697 89
rect -697 -89 -637 -70
rect -697 -97 -678 -89
rect -686 -106 -678 -97
rect -656 -97 -637 -89
rect -608 -89 -548 -70
rect -608 -97 -589 -89
rect -656 -106 -648 -97
rect -686 -114 -648 -106
rect -597 -106 -589 -97
rect -567 -97 -548 -89
rect -519 -89 -459 -70
rect -519 -97 -500 -89
rect -567 -106 -559 -97
rect -597 -114 -559 -106
rect -508 -106 -500 -97
rect -478 -97 -459 -89
rect -430 -89 -370 -70
rect -430 -97 -411 -89
rect -478 -106 -470 -97
rect -508 -114 -470 -106
rect -419 -106 -411 -97
rect -389 -97 -370 -89
rect -341 -89 -281 -70
rect -341 -97 -322 -89
rect -389 -106 -381 -97
rect -419 -114 -381 -106
rect -330 -106 -322 -97
rect -300 -97 -281 -89
rect -252 -89 -192 -70
rect -252 -97 -233 -89
rect -300 -106 -292 -97
rect -330 -114 -292 -106
rect -241 -106 -233 -97
rect -211 -97 -192 -89
rect -163 -89 -103 -70
rect -163 -97 -144 -89
rect -211 -106 -203 -97
rect -241 -114 -203 -106
rect -152 -106 -144 -97
rect -122 -97 -103 -89
rect -74 -89 -14 -70
rect -74 -97 -55 -89
rect -122 -106 -114 -97
rect -152 -114 -114 -106
rect -63 -106 -55 -97
rect -33 -97 -14 -89
rect 14 -89 74 -70
rect 14 -97 33 -89
rect -33 -106 -25 -97
rect -63 -114 -25 -106
rect 25 -106 33 -97
rect 55 -97 74 -89
rect 103 -89 163 -70
rect 103 -97 122 -89
rect 55 -106 63 -97
rect 25 -114 63 -106
rect 114 -106 122 -97
rect 144 -97 163 -89
rect 192 -89 252 -70
rect 192 -97 211 -89
rect 144 -106 152 -97
rect 114 -114 152 -106
rect 203 -106 211 -97
rect 233 -97 252 -89
rect 281 -89 341 -70
rect 281 -97 300 -89
rect 233 -106 241 -97
rect 203 -114 241 -106
rect 292 -106 300 -97
rect 322 -97 341 -89
rect 370 -89 430 -70
rect 370 -97 389 -89
rect 322 -106 330 -97
rect 292 -114 330 -106
rect 381 -106 389 -97
rect 411 -97 430 -89
rect 459 -89 519 -70
rect 459 -97 478 -89
rect 411 -106 419 -97
rect 381 -114 419 -106
rect 470 -106 478 -97
rect 500 -97 519 -89
rect 548 -89 608 -70
rect 548 -97 567 -89
rect 500 -106 508 -97
rect 470 -114 508 -106
rect 559 -106 567 -97
rect 589 -97 608 -89
rect 637 -89 697 -70
rect 637 -97 656 -89
rect 589 -106 597 -97
rect 559 -114 597 -106
rect 648 -106 656 -97
rect 678 -97 697 -89
rect 678 -106 686 -97
rect 648 -114 686 -106
<< polycont >>
rect -678 89 -656 106
rect -589 89 -567 106
rect -500 89 -478 106
rect -411 89 -389 106
rect -322 89 -300 106
rect -233 89 -211 106
rect -144 89 -122 106
rect -55 89 -33 106
rect 33 89 55 106
rect 122 89 144 106
rect 211 89 233 106
rect 300 89 322 106
rect 389 89 411 106
rect 478 89 500 106
rect 567 89 589 106
rect 656 89 678 106
rect -678 -106 -656 -89
rect -589 -106 -567 -89
rect -500 -106 -478 -89
rect -411 -106 -389 -89
rect -322 -106 -300 -89
rect -233 -106 -211 -89
rect -144 -106 -122 -89
rect -55 -106 -33 -89
rect 33 -106 55 -89
rect 122 -106 144 -89
rect 211 -106 233 -89
rect 300 -106 322 -89
rect 389 -106 411 -89
rect 478 -106 500 -89
rect 567 -106 589 -89
rect 656 -106 678 -89
<< locali >>
rect -686 89 -678 106
rect -656 89 -648 106
rect -597 89 -589 106
rect -567 89 -559 106
rect -508 89 -500 106
rect -478 89 -470 106
rect -419 89 -411 106
rect -389 89 -381 106
rect -330 89 -322 106
rect -300 89 -292 106
rect -241 89 -233 106
rect -211 89 -203 106
rect -152 89 -144 106
rect -122 89 -114 106
rect -63 89 -55 106
rect -33 89 -25 106
rect 25 89 33 106
rect 55 89 63 106
rect 114 89 122 106
rect 144 89 152 106
rect 203 89 211 106
rect 233 89 241 106
rect 292 89 300 106
rect 322 89 330 106
rect 381 89 389 106
rect 411 89 419 106
rect 470 89 478 106
rect 500 89 508 106
rect 559 89 567 106
rect 589 89 597 106
rect 648 89 656 106
rect 678 89 686 106
rect -720 64 -703 72
rect -720 -72 -703 -64
rect -631 64 -614 72
rect -631 -72 -614 -64
rect -542 64 -525 72
rect -542 -72 -525 -64
rect -453 64 -436 72
rect -453 -72 -436 -64
rect -364 64 -347 72
rect -364 -72 -347 -64
rect -275 64 -258 72
rect -275 -72 -258 -64
rect -186 64 -169 72
rect -186 -72 -169 -64
rect -97 64 -80 72
rect -97 -72 -80 -64
rect -8 64 8 72
rect -8 -72 8 -64
rect 80 64 97 72
rect 80 -72 97 -64
rect 169 64 186 72
rect 169 -72 186 -64
rect 258 64 275 72
rect 258 -72 275 -64
rect 347 64 364 72
rect 347 -72 364 -64
rect 436 64 453 72
rect 436 -72 453 -64
rect 525 64 542 72
rect 525 -72 542 -64
rect 614 64 631 72
rect 614 -72 631 -64
rect 703 64 720 72
rect 703 -72 720 -64
rect -686 -106 -678 -89
rect -656 -106 -648 -89
rect -597 -106 -589 -89
rect -567 -106 -559 -89
rect -508 -106 -500 -89
rect -478 -106 -470 -89
rect -419 -106 -411 -89
rect -389 -106 -381 -89
rect -330 -106 -322 -89
rect -300 -106 -292 -89
rect -241 -106 -233 -89
rect -211 -106 -203 -89
rect -152 -106 -144 -89
rect -122 -106 -114 -89
rect -63 -106 -55 -89
rect -33 -106 -25 -89
rect 25 -106 33 -89
rect 55 -106 63 -89
rect 114 -106 122 -89
rect 144 -106 152 -89
rect 203 -106 211 -89
rect 233 -106 241 -89
rect 292 -106 300 -89
rect 322 -106 330 -89
rect 381 -106 389 -89
rect 411 -106 419 -89
rect 470 -106 478 -89
rect 500 -106 508 -89
rect 559 -106 567 -89
rect 589 -106 597 -89
rect 648 -106 656 -89
rect 678 -106 686 -89
<< viali >>
rect -678 89 -656 106
rect -589 89 -567 106
rect -500 89 -478 106
rect -411 89 -389 106
rect -322 89 -300 106
rect -233 89 -211 106
rect -144 89 -122 106
rect -55 89 -33 106
rect 33 89 55 106
rect 122 89 144 106
rect 211 89 233 106
rect 300 89 322 106
rect 389 89 411 106
rect 478 89 500 106
rect 567 89 589 106
rect 656 89 678 106
rect -720 -64 -703 64
rect -631 -64 -614 64
rect -542 -64 -525 64
rect -453 -64 -436 64
rect -364 -64 -347 64
rect -275 -64 -258 64
rect -186 -64 -169 64
rect -97 -64 -80 64
rect -8 -64 8 64
rect 80 -64 97 64
rect 169 -64 186 64
rect 258 -64 275 64
rect 347 -64 364 64
rect 436 -64 453 64
rect 525 -64 542 64
rect 614 -64 631 64
rect 703 -64 720 64
rect -678 -106 -656 -89
rect -589 -106 -567 -89
rect -500 -106 -478 -89
rect -411 -106 -389 -89
rect -322 -106 -300 -89
rect -233 -106 -211 -89
rect -144 -106 -122 -89
rect -55 -106 -33 -89
rect 33 -106 55 -89
rect 122 -106 144 -89
rect 211 -106 233 -89
rect 300 -106 322 -89
rect 389 -106 411 -89
rect 478 -106 500 -89
rect 567 -106 589 -89
rect 656 -106 678 -89
<< metal1 >>
rect -686 106 -648 114
rect -686 89 -678 106
rect -656 89 -648 106
rect -686 86 -648 89
rect -597 106 -559 114
rect -597 89 -589 106
rect -567 89 -559 106
rect -597 86 -559 89
rect -508 106 -470 114
rect -508 89 -500 106
rect -478 89 -470 106
rect -508 86 -470 89
rect -419 106 -381 114
rect -419 89 -411 106
rect -389 89 -381 106
rect -419 86 -381 89
rect -330 106 -292 114
rect -330 89 -322 106
rect -300 89 -292 106
rect -330 86 -292 89
rect -241 106 -203 114
rect -241 89 -233 106
rect -211 89 -203 106
rect -241 86 -203 89
rect -152 106 -114 114
rect -152 89 -144 106
rect -122 89 -114 106
rect -152 86 -114 89
rect -63 106 -25 114
rect -63 89 -55 106
rect -33 89 -25 106
rect -63 86 -25 89
rect 25 106 63 114
rect 25 89 33 106
rect 55 89 63 106
rect 25 86 63 89
rect 114 106 152 114
rect 114 89 122 106
rect 144 89 152 106
rect 114 86 152 89
rect 203 106 241 114
rect 203 89 211 106
rect 233 89 241 106
rect 203 86 241 89
rect 292 106 330 114
rect 292 89 300 106
rect 322 89 330 106
rect 292 86 330 89
rect 381 106 419 114
rect 381 89 389 106
rect 411 89 419 106
rect 381 86 419 89
rect 470 106 508 114
rect 470 89 478 106
rect 500 89 508 106
rect 470 86 508 89
rect 559 106 597 114
rect 559 89 567 106
rect 589 89 597 106
rect 559 86 597 89
rect 648 106 686 114
rect 648 89 656 106
rect 678 89 686 106
rect 648 86 686 89
rect -723 64 -700 70
rect -723 -64 -720 64
rect -703 -64 -700 64
rect -723 -70 -700 -64
rect -634 64 -611 70
rect -634 -64 -631 64
rect -614 -64 -611 64
rect -634 -70 -611 -64
rect -545 64 -522 70
rect -545 -64 -542 64
rect -525 -64 -522 64
rect -545 -70 -522 -64
rect -456 64 -433 70
rect -456 -64 -453 64
rect -436 -64 -433 64
rect -456 -70 -433 -64
rect -367 64 -344 70
rect -367 -64 -364 64
rect -347 -64 -344 64
rect -367 -70 -344 -64
rect -278 64 -255 70
rect -278 -64 -275 64
rect -258 -64 -255 64
rect -278 -70 -255 -64
rect -189 64 -166 70
rect -189 -64 -186 64
rect -169 -64 -166 64
rect -189 -70 -166 -64
rect -100 64 -77 70
rect -100 -64 -97 64
rect -80 -64 -77 64
rect -100 -70 -77 -64
rect -11 64 11 70
rect -11 -64 -8 64
rect 8 -64 11 64
rect -11 -70 11 -64
rect 77 64 100 70
rect 77 -64 80 64
rect 97 -64 100 64
rect 77 -70 100 -64
rect 166 64 189 70
rect 166 -64 169 64
rect 186 -64 189 64
rect 166 -70 189 -64
rect 255 64 278 70
rect 255 -64 258 64
rect 275 -64 278 64
rect 255 -70 278 -64
rect 344 64 367 70
rect 344 -64 347 64
rect 364 -64 367 64
rect 344 -70 367 -64
rect 433 64 456 70
rect 433 -64 436 64
rect 453 -64 456 64
rect 433 -70 456 -64
rect 522 64 545 70
rect 522 -64 525 64
rect 542 -64 545 64
rect 522 -70 545 -64
rect 611 64 634 70
rect 611 -64 614 64
rect 631 -64 634 64
rect 611 -70 634 -64
rect 700 64 723 70
rect 700 -64 703 64
rect 720 -64 723 64
rect 700 -70 723 -64
rect -686 -89 -648 -86
rect -686 -106 -678 -89
rect -656 -106 -648 -89
rect -686 -114 -648 -106
rect -597 -89 -559 -86
rect -597 -106 -589 -89
rect -567 -106 -559 -89
rect -597 -114 -559 -106
rect -508 -89 -470 -86
rect -508 -106 -500 -89
rect -478 -106 -470 -89
rect -508 -114 -470 -106
rect -419 -89 -381 -86
rect -419 -106 -411 -89
rect -389 -106 -381 -89
rect -419 -114 -381 -106
rect -330 -89 -292 -86
rect -330 -106 -322 -89
rect -300 -106 -292 -89
rect -330 -114 -292 -106
rect -241 -89 -203 -86
rect -241 -106 -233 -89
rect -211 -106 -203 -89
rect -241 -114 -203 -106
rect -152 -89 -114 -86
rect -152 -106 -144 -89
rect -122 -106 -114 -89
rect -152 -114 -114 -106
rect -63 -89 -25 -86
rect -63 -106 -55 -89
rect -33 -106 -25 -89
rect -63 -114 -25 -106
rect 25 -89 63 -86
rect 25 -106 33 -89
rect 55 -106 63 -89
rect 25 -114 63 -106
rect 114 -89 152 -86
rect 114 -106 122 -89
rect 144 -106 152 -89
rect 114 -114 152 -106
rect 203 -89 241 -86
rect 203 -106 211 -89
rect 233 -106 241 -89
rect 203 -114 241 -106
rect 292 -89 330 -86
rect 292 -106 300 -89
rect 322 -106 330 -89
rect 292 -114 330 -106
rect 381 -89 419 -86
rect 381 -106 389 -89
rect 411 -106 419 -89
rect 381 -114 419 -106
rect 470 -89 508 -86
rect 470 -106 478 -89
rect 500 -106 508 -89
rect 470 -114 508 -106
rect 559 -89 597 -86
rect 559 -106 567 -89
rect 589 -106 597 -89
rect 559 -114 597 -106
rect 648 -89 686 -86
rect 648 -106 656 -89
rect 678 -106 686 -89
rect 648 -114 686 -106
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 16 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
