* NGSPICE file created from a_mux4_en_flat.ext - technology: sky130A

.subckt a_mux4_en_flat en s1 s0 in0 in1 in2 in3 out VDD VSS
X0 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=1.05536e+13p pd=8.08e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X1 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X2 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X3 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X4 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X5 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X6 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X7 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X8 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X9 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=4.0352e+12p ps=4.048e+07u w=520000u l=150000u
X10 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X11 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X12 a_n499_n2830# sky130_fd_sc_hd__nand2_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=2.439e+12p ps=2.634e+07u w=650000u l=150000u
X13 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X14 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X15 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X16 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X17 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X18 a_n499_n1742# sky130_fd_sc_hd__nand2_1_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X20 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X21 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X22 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X23 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X24 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X25 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X26 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X27 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X28 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X29 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X30 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X31 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X32 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X33 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X34 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X35 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X36 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X37 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X38 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X39 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X40 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X41 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X42 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X43 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X44 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X45 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X46 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X47 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X48 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X49 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X50 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X51 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X52 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X53 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X54 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X55 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X56 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nand2_1_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.9e+12p ps=3.78e+07u w=1e+06u l=150000u
X57 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X58 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X59 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X60 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X61 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X62 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X63 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/en_b VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X64 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X65 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X66 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X67 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X68 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X69 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X70 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X71 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X72 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X73 switch_5t_3/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X74 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X75 VDD s0 switch_5t_2/transmission_gate_0/en_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X76 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X77 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X78 switch_5t_3/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X79 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X80 VDD sky130_fd_sc_hd__nand2_1_3/A switch_5t_1/transmission_gate_0/en_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X81 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X82 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X83 sky130_fd_sc_hd__nand2_1_0/Y s0 a_n499_n3694# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X84 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X85 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X86 VDD s0 sky130_fd_sc_hd__nand2_1_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X87 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X88 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X89 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X90 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X91 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X92 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X93 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X94 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X95 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X96 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X97 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X98 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X99 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X100 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X101 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X102 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X103 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X104 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X105 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X106 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X107 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X108 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X109 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X110 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X111 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X112 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X113 switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X114 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X115 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X116 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X117 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X118 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X119 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X120 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X121 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X122 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X123 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X124 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X125 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X127 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X129 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X130 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X131 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X132 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X133 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X134 a_n499_n3694# s1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X135 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X136 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X137 sky130_fd_sc_hd__nand2_1_3/B s0 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X138 sky130_fd_sc_hd__nand2_1_0/Y s1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X140 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X141 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X142 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X143 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X144 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X145 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X146 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X147 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X148 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X149 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X150 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X151 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X152 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X153 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X154 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X155 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X156 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X157 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X158 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X159 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X160 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X161 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X162 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X163 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X164 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X165 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X166 transmission_gate_0/en_b en VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X167 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X168 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X169 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X170 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X171 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X172 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X173 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X174 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X175 sky130_fd_sc_hd__nand2_1_3/A s1 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X176 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X177 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X178 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X179 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X180 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X181 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X182 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X183 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X184 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X185 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X186 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X187 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X188 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X189 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X190 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X191 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X192 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X193 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X194 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X195 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X196 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X197 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X198 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X199 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X200 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X201 switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/en_b VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X202 sky130_fd_sc_hd__nand2_1_3/B s0 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X203 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X204 sky130_fd_sc_hd__inv_1_3/A s1 a_n499_n2606# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X205 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X206 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X207 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X208 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X209 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X210 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X211 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X212 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X213 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X214 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X215 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X216 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X217 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X218 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X219 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X220 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X221 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X222 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X223 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X224 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X225 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X226 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X227 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X228 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X229 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X230 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X231 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X232 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X233 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X234 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X235 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X236 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X237 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X238 switch_5t_2/transmission_gate_0/en_b s0 a_n499_n2830# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X239 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X240 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X241 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A a_n499_n1742# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X242 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X243 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X244 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X245 transmission_gate_0/en_b en VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X246 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X247 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X248 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X249 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X250 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X251 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X252 a_n499_n2606# sky130_fd_sc_hd__nand2_1_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X253 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X254 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X255 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X256 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X257 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X258 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X259 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X260 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X261 sky130_fd_sc_hd__nand2_1_3/A s1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X262 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X263 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X264 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X265 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X266 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X267 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X268 VDD s1 sky130_fd_sc_hd__inv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X269 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X270 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X271 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X272 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X273 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/en 0.54fF
C1 in2 VDD 1.28fF
C2 sky130_fd_sc_hd__nand2_1_0/Y transmission_gate_0/en_b 0.04fF
C3 switch_5t_2/transmission_gate_0/en_b transmission_gate_0/en_b 0.04fF
C4 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/B 0.07fF
C5 switch_5t_2/transmission_gate_0/in in1 0.06fF
C6 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nand2_1_3/B 0.00fF
C7 en s1 0.66fF
C8 switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in 1.57fF
C9 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/out 7.39fF
C10 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nand2_1_3/A 0.19fF
C11 en switch_5t_1/transmission_gate_0/en 0.07fF
C12 switch_5t_2/transmission_gate_0/out switch_5t_3/transmission_gate_0/in 0.06fF
C13 sky130_fd_sc_hd__inv_1_3/A VDD 3.71fF
C14 transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B 0.04fF
C15 s0 in2 0.00fF
C16 switch_5t_0/transmission_gate_0/out switch_5t_1/transmission_gate_0/out 0.33fF
C17 in1 switch_5t_0/transmission_gate_0/in 6.76fF
C18 switch_5t_0/transmission_gate_0/out switch_5t_1/transmission_gate_0/in 0.07fF
C19 sky130_fd_sc_hd__nand2_1_0/Y s1 0.08fF
C20 switch_5t_2/transmission_gate_0/en_b s1 0.07fF
C21 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/in 7.32fF
C22 switch_5t_2/transmission_gate_0/en switch_5t_3/transmission_gate_0/in 0.04fF
C23 switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out 1.88fF
C24 switch_5t_2/transmission_gate_0/out switch_5t_3/transmission_gate_0/en 0.09fF
C25 switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in 1.39fF
C26 switch_5t_2/transmission_gate_0/in in2 6.62fF
C27 switch_5t_0/transmission_gate_0/in in0 0.06fF
C28 switch_5t_2/transmission_gate_0/out switch_5t_0/transmission_gate_0/out 0.30fF
C29 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en 1.97fF
C30 switch_5t_2/transmission_gate_0/en switch_5t_3/transmission_gate_0/en 0.25fF
C31 VDD sky130_fd_sc_hd__nand2_1_3/A 1.38fF
C32 s0 sky130_fd_sc_hd__inv_1_3/A 0.10fF
C33 en switch_5t_3/transmission_gate_0/in 0.63fF
C34 in3 VDD 1.13fF
C35 switch_5t_1/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/out 0.12fF
C36 in1 transmission_gate_0/en_b 1.29fF
C37 out switch_5t_1/transmission_gate_0/en 0.58fF
C38 switch_5t_2/transmission_gate_0/en switch_5t_0/transmission_gate_0/out 0.09fF
C39 a_n499_n2830# switch_5t_2/transmission_gate_0/en_b 0.01fF
C40 switch_5t_2/transmission_gate_0/out switch_5t_3/transmission_gate_0/out 0.30fF
C41 en switch_5t_1/transmission_gate_0/out 0.00fF
C42 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out 1.96fF
C43 s1 sky130_fd_sc_hd__nand2_1_3/B 0.36fF
C44 en switch_5t_1/transmission_gate_0/in 0.70fF
C45 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A 0.06fF
C46 in0 transmission_gate_0/en_b 1.33fF
C47 switch_5t_2/transmission_gate_0/en switch_5t_3/transmission_gate_0/out 0.02fF
C48 in2 switch_5t_0/transmission_gate_0/in 0.07fF
C49 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in 1.40fF
C50 switch_5t_2/transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in 0.09fF
C51 switch_5t_1/transmission_gate_0/en_b a_n499_n1742# 0.01fF
C52 s0 sky130_fd_sc_hd__nand2_1_3/A 1.04fF
C53 en switch_5t_1/transmission_gate_0/en_b 0.07fF
C54 s0 VDD 1.24fF
C55 switch_5t_2/transmission_gate_0/en en 0.03fF
C56 out switch_5t_3/transmission_gate_0/in 0.43fF
C57 switch_5t_2/transmission_gate_0/en_b switch_5t_3/transmission_gate_0/en 0.46fF
C58 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/en 0.55fF
C59 sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in 1.59fF
C60 in2 transmission_gate_0/en_b 1.30fF
C61 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/A 0.08fF
C62 out switch_5t_1/transmission_gate_0/out 7.54fF
C63 switch_5t_2/transmission_gate_0/in in3 0.07fF
C64 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y 0.62fF
C65 switch_5t_2/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/out 0.02fF
C66 out switch_5t_1/transmission_gate_0/in 0.43fF
C67 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b 1.89fF
C68 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/out 0.06fF
C69 switch_5t_2/transmission_gate_0/in VDD 3.32fF
C70 out switch_5t_3/transmission_gate_0/en 0.63fF
C71 switch_5t_1/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/en_b 0.01fF
C72 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_1/transmission_gate_0/en_b 0.00fF
C73 switch_5t_1/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/B 0.02fF
C74 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out 1.85fF
C75 switch_5t_2/transmission_gate_0/en_b switch_5t_3/transmission_gate_0/out 0.09fF
C76 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/en_b 1.01fF
C77 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/en 0.19fF
C78 out switch_5t_0/transmission_gate_0/out 7.67fF
C79 out switch_5t_2/transmission_gate_0/out 7.67fF
C80 sky130_fd_sc_hd__inv_1_3/A transmission_gate_0/en_b 0.04fF
C81 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/A 0.08fF
C82 out switch_5t_1/transmission_gate_0/en_b 0.50fF
C83 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_3/B 0.02fF
C84 out switch_5t_3/transmission_gate_0/out 7.47fF
C85 switch_5t_2/transmission_gate_0/en out 0.64fF
C86 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C87 en switch_5t_2/transmission_gate_0/en_b 0.03fF
C88 in2 s1 0.00fF
C89 sky130_fd_sc_hd__nand2_1_0/Y en 0.06fF
C90 switch_5t_0/transmission_gate_0/in VDD 2.86fF
C91 switch_5t_2/transmission_gate_0/in s0 0.46fF
C92 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B 0.06fF
C93 sky130_fd_sc_hd__inv_1_3/Y VDD 0.57fF
C94 in1 switch_5t_1/transmission_gate_0/in 0.07fF
C95 transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A 0.10fF
C96 in3 transmission_gate_0/en_b 1.23fF
C97 sky130_fd_sc_hd__inv_1_3/A s1 0.39fF
C98 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/en_b 0.39fF
C99 en sky130_fd_sc_hd__nand2_1_3/B 0.03fF
C100 VDD transmission_gate_0/en_b 5.66fF
C101 switch_5t_1/transmission_gate_0/in in0 6.63fF
C102 s0 switch_5t_0/transmission_gate_0/in 0.07fF
C103 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/en 0.02fF
C104 s0 sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C105 out switch_5t_2/transmission_gate_0/en_b 0.51fF
C106 sky130_fd_sc_hd__nand2_1_0/Y out 0.45fF
C107 in2 switch_5t_3/transmission_gate_0/in 0.06fF
C108 switch_5t_2/transmission_gate_0/in switch_5t_0/transmission_gate_0/in 0.30fF
C109 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B 0.00fF
C110 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C111 s1 sky130_fd_sc_hd__nand2_1_3/A 0.51fF
C112 s0 transmission_gate_0/en_b 0.47fF
C113 en in1 1.35fF
C114 s1 VDD 1.02fF
C115 switch_5t_1/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C116 VDD switch_5t_1/transmission_gate_0/en 0.44fF
C117 en in0 1.35fF
C118 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b 0.58fF
C119 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/out 0.03fF
C120 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/in 0.05fF
C121 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y 1.57fF
C122 sky130_fd_sc_hd__inv_1_3/A a_n499_n2606# 0.02fF
C123 s0 s1 2.22fF
C124 sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out 1.89fF
C125 sky130_fd_sc_hd__inv_1_3/A switch_5t_2/transmission_gate_0/out 0.09fF
C126 s0 switch_5t_1/transmission_gate_0/en 0.03fF
C127 in2 en 1.37fF
C128 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b 0.82fF
C129 in3 switch_5t_3/transmission_gate_0/in 6.62fF
C130 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/en_b 0.47fF
C131 sky130_fd_sc_hd__inv_1_3/Y transmission_gate_0/en_b 0.01fF
C132 switch_5t_2/transmission_gate_0/en sky130_fd_sc_hd__inv_1_3/A 0.42fF
C133 VDD switch_5t_3/transmission_gate_0/in 2.44fF
C134 switch_5t_1/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C135 switch_5t_2/transmission_gate_0/in s1 0.30fF
C136 in1 sky130_fd_sc_hd__nand2_1_3/B 0.01fF
C137 VDD switch_5t_1/transmission_gate_0/out 2.93fF
C138 a_n499_n2830# s0 0.00fF
C139 VDD switch_5t_1/transmission_gate_0/in 3.13fF
C140 switch_5t_3/transmission_gate_0/en VDD 0.58fF
C141 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C142 switch_5t_2/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C143 sky130_fd_sc_hd__inv_1_3/A en 0.03fF
C144 switch_5t_0/transmission_gate_0/out VDD 3.04fF
C145 switch_5t_2/transmission_gate_0/out VDD 3.01fF
C146 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A 0.21fF
C147 s1 switch_5t_0/transmission_gate_0/in 0.08fF
C148 switch_5t_2/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C149 s0 switch_5t_3/transmission_gate_0/in 0.01fF
C150 switch_5t_1/transmission_gate_0/en_b VDD 3.71fF
C151 s1 sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C152 switch_5t_3/transmission_gate_0/out VDD 2.72fF
C153 switch_5t_0/transmission_gate_0/in switch_5t_1/transmission_gate_0/en 0.01fF
C154 switch_5t_2/transmission_gate_0/en VDD 0.57fF
C155 s0 switch_5t_1/transmission_gate_0/in 0.04fF
C156 sky130_fd_sc_hd__inv_1_3/Y switch_5t_1/transmission_gate_0/en 0.20fF
C157 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_3/A 0.01fF
C158 sky130_fd_sc_hd__inv_1_3/A switch_5t_2/transmission_gate_0/en_b 0.23fF
C159 s0 switch_5t_3/transmission_gate_0/en 0.01fF
C160 en sky130_fd_sc_hd__nand2_1_3/A 0.07fF
C161 switch_5t_2/transmission_gate_0/in switch_5t_3/transmission_gate_0/in 0.35fF
C162 in1 in0 0.25fF
C163 en in3 1.34fF
C164 s0 switch_5t_2/transmission_gate_0/out 0.02fF
C165 en VDD 0.48fF
C166 s1 transmission_gate_0/en_b 1.15fF
C167 sky130_fd_sc_hd__inv_1_3/A out 0.51fF
C168 switch_5t_2/transmission_gate_0/in switch_5t_3/transmission_gate_0/en 0.07fF
C169 s0 switch_5t_1/transmission_gate_0/en_b 0.08fF
C170 switch_5t_1/transmission_gate_0/en transmission_gate_0/en_b 0.07fF
C171 switch_5t_2/transmission_gate_0/en s0 0.09fF
C172 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nand2_1_3/B 0.20fF
C173 switch_5t_2/transmission_gate_0/in switch_5t_0/transmission_gate_0/out 0.06fF
C174 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/out 7.32fF
C175 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A 0.09fF
C176 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C177 in2 in1 0.23fF
C178 switch_5t_2/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b 0.00fF
C179 switch_5t_0/transmission_gate_0/in switch_5t_1/transmission_gate_0/out 0.06fF
C180 sky130_fd_sc_hd__nand2_1_0/Y VDD 3.70fF
C181 switch_5t_2/transmission_gate_0/en_b VDD 3.75fF
C182 switch_5t_2/transmission_gate_0/in switch_5t_3/transmission_gate_0/out 0.07fF
C183 switch_5t_0/transmission_gate_0/in switch_5t_1/transmission_gate_0/in 0.45fF
C184 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en 1.51fF
C185 s0 en 0.55fF
C186 sky130_fd_sc_hd__inv_1_3/Y switch_5t_1/transmission_gate_0/out 0.09fF
C187 sky130_fd_sc_hd__inv_1_3/Y switch_5t_1/transmission_gate_0/in 0.12fF
C188 out VDD 6.03fF
C189 switch_5t_0/transmission_gate_0/out switch_5t_0/transmission_gate_0/in 7.36fF
C190 s1 switch_5t_1/transmission_gate_0/en 0.03fF
C191 switch_5t_2/transmission_gate_0/out switch_5t_0/transmission_gate_0/in 0.07fF
C192 sky130_fd_sc_hd__nand2_1_3/B sky130_fd_sc_hd__nand2_1_3/A 0.49fF
C193 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in 0.49fF
C194 switch_5t_2/transmission_gate_0/in en 0.66fF
C195 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y 1.95fF
C196 switch_5t_2/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C197 switch_5t_1/transmission_gate_0/out transmission_gate_0/en_b 0.02fF
C198 VDD sky130_fd_sc_hd__nand2_1_3/B 1.22fF
C199 switch_5t_1/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in 0.13fF
C200 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b 0.73fF
C201 sky130_fd_sc_hd__nand2_1_0/Y s0 0.21fF
C202 s0 switch_5t_2/transmission_gate_0/en_b 0.45fF
C203 switch_5t_2/transmission_gate_0/en switch_5t_0/transmission_gate_0/in 0.05fF
C204 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__inv_1_3/Y 0.67fF
C205 switch_5t_3/transmission_gate_0/en transmission_gate_0/en_b 0.00fF
C206 switch_5t_2/transmission_gate_0/en sky130_fd_sc_hd__inv_1_3/Y 0.16fF
C207 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b 1.46fF
C208 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/in 0.09fF
C209 en switch_5t_0/transmission_gate_0/in 0.68fF
C210 sky130_fd_sc_hd__nand2_1_0/Y a_n499_n3694# 0.02fF
C211 switch_5t_1/transmission_gate_0/en_b transmission_gate_0/en_b 0.06fF
C212 s1 switch_5t_3/transmission_gate_0/in 0.02fF
C213 s0 sky130_fd_sc_hd__nand2_1_3/B 0.34fF
C214 switch_5t_2/transmission_gate_0/en transmission_gate_0/en_b 0.04fF
C215 in1 VDD 1.23fF
C216 switch_5t_2/transmission_gate_0/in out 0.43fF
C217 s1 switch_5t_1/transmission_gate_0/in 0.06fF
C218 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en 2.01fF
C219 VDD in0 1.35fF
C220 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en 1.53fF
C221 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/B 0.02fF
C222 a_n499_n2606# s1 0.00fF
C223 en transmission_gate_0/en_b 3.34fF
C224 switch_5t_2/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in 0.02fF
C225 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C226 switch_5t_2/transmission_gate_0/out s1 0.01fF
C227 switch_5t_0/transmission_gate_0/out switch_5t_1/transmission_gate_0/en 0.03fF
C228 s0 in1 0.00fF
C229 switch_5t_1/transmission_gate_0/en_b s1 0.07fF
C230 out switch_5t_0/transmission_gate_0/in 0.43fF
C231 in2 sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C232 switch_5t_2/transmission_gate_0/en s1 0.03fF
C233 in2 in3 0.23fF
C234 out sky130_fd_sc_hd__inv_1_3/Y 0.64fF
C235 switch_5t_3/transmission_gate_0/out VSS 2.21fF
C236 switch_5t_3/transmission_gate_0/en VSS 3.37fF
C237 in3 VSS 1.22fF
C238 switch_5t_3/transmission_gate_0/in VSS 2.54fF
C239 a_n499_n3694# VSS 0.00fF
C240 sky130_fd_sc_hd__nand2_1_0/Y VSS 1.45fF
C241 switch_5t_2/transmission_gate_0/out VSS 2.35fF
C242 switch_5t_2/transmission_gate_0/en VSS 3.94fF
C243 in2 VSS 1.28fF
C244 switch_5t_2/transmission_gate_0/in VSS 2.87fF
C245 switch_5t_2/transmission_gate_0/en_b VSS 1.41fF
C246 a_n499_n2830# VSS 0.01fF
C247 a_n499_n2606# VSS 0.00fF
C248 s1 VSS 2.28fF
C249 s0 VSS 1.60fF
C250 switch_5t_0/transmission_gate_0/out VSS 2.34fF
C251 a_n499_n1742# VSS 0.01fF
C252 sky130_fd_sc_hd__nand2_1_3/A VSS 0.97fF
C253 sky130_fd_sc_hd__nand2_1_3/B VSS 0.70fF
C254 in1 VSS 1.30fF
C255 switch_5t_0/transmission_gate_0/in VSS 3.43fF
C256 sky130_fd_sc_hd__inv_1_3/Y VSS 3.75fF
C257 sky130_fd_sc_hd__inv_1_3/A VSS 1.52fF
C258 en VSS 9.89fF
C259 out VSS 5.26fF
C260 switch_5t_1/transmission_gate_0/en_b VSS 1.23fF
C261 switch_5t_1/transmission_gate_0/out VSS 2.45fF
C262 switch_5t_1/transmission_gate_0/en VSS 4.40fF
C263 in0 VSS 1.28fF
C264 switch_5t_1/transmission_gate_0/in VSS 3.06fF
C265 transmission_gate_0/en_b VSS 3.07fF
C266 VDD VSS 47.88fF
.ends

