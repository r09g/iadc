* NGSPICE file created from onebit_dac.ext - technology: sky130A

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_n320_n136# a_448_n136# 0.02fF
C1 a_n32_n136# w_n646_n356# 0.05fF
C2 a_n224_n136# a_n320_n136# 0.33fF
C3 a_n128_n136# a_n320_n136# 0.12fF
C4 a_n512_n234# a_n508_n136# 0.03fF
C5 a_160_n136# a_n512_n234# 0.03fF
C6 a_352_n136# a_n512_n234# 0.03fF
C7 a_256_n136# a_n508_n136# 0.02fF
C8 a_256_n136# a_160_n136# 0.33fF
C9 a_352_n136# a_256_n136# 0.33fF
C10 a_n416_n136# a_n512_n234# 0.03fF
C11 a_64_n136# a_n508_n136# 0.03fF
C12 a_160_n136# a_64_n136# 0.33fF
C13 a_352_n136# a_64_n136# 0.07fF
C14 a_n512_n234# w_n646_n356# 1.47fF
C15 a_n512_n234# a_n32_n136# 0.03fF
C16 a_256_n136# a_n416_n136# 0.03fF
C17 a_n416_n136# a_64_n136# 0.04fF
C18 a_256_n136# w_n646_n356# 0.06fF
C19 a_256_n136# a_n32_n136# 0.07fF
C20 a_64_n136# w_n646_n356# 0.05fF
C21 a_n32_n136# a_64_n136# 0.33fF
C22 a_n508_n136# a_448_n136# 0.02fF
C23 a_160_n136# a_448_n136# 0.07fF
C24 a_352_n136# a_448_n136# 0.33fF
C25 a_n224_n136# a_n508_n136# 0.07fF
C26 a_n224_n136# a_160_n136# 0.05fF
C27 a_352_n136# a_n224_n136# 0.03fF
C28 a_n416_n136# a_448_n136# 0.02fF
C29 a_n128_n136# a_n508_n136# 0.05fF
C30 a_160_n136# a_n128_n136# 0.07fF
C31 a_352_n136# a_n128_n136# 0.04fF
C32 a_n224_n136# a_n416_n136# 0.12fF
C33 w_n646_n356# a_448_n136# 0.13fF
C34 a_n32_n136# a_448_n136# 0.04fF
C35 a_n224_n136# w_n646_n356# 0.06fF
C36 a_n224_n136# a_n32_n136# 0.12fF
C37 a_256_n136# a_n512_n234# 0.03fF
C38 a_n512_n234# a_64_n136# 0.03fF
C39 a_n416_n136# a_n128_n136# 0.07fF
C40 w_n646_n356# a_n128_n136# 0.05fF
C41 a_n32_n136# a_n128_n136# 0.33fF
C42 a_256_n136# a_64_n136# 0.12fF
C43 a_n508_n136# a_n320_n136# 0.12fF
C44 a_160_n136# a_n320_n136# 0.04fF
C45 a_352_n136# a_n320_n136# 0.03fF
C46 a_n416_n136# a_n320_n136# 0.33fF
C47 a_n512_n234# a_448_n136# 0.03fF
C48 a_n224_n136# a_n512_n234# 0.03fF
C49 w_n646_n356# a_n320_n136# 0.06fF
C50 a_n32_n136# a_n320_n136# 0.07fF
C51 a_256_n136# a_448_n136# 0.12fF
C52 a_64_n136# a_448_n136# 0.05fF
C53 a_n224_n136# a_256_n136# 0.04fF
C54 a_n512_n234# a_n128_n136# 0.03fF
C55 a_n224_n136# a_64_n136# 0.07fF
C56 a_256_n136# a_n128_n136# 0.05fF
C57 a_64_n136# a_n128_n136# 0.12fF
C58 a_n512_n234# a_n320_n136# 0.03fF
C59 a_n224_n136# a_448_n136# 0.03fF
C60 a_160_n136# a_n508_n136# 0.03fF
C61 a_256_n136# a_n320_n136# 0.03fF
C62 a_352_n136# a_n508_n136# 0.02fF
C63 a_352_n136# a_160_n136# 0.12fF
C64 a_64_n136# a_n320_n136# 0.05fF
C65 a_n128_n136# a_448_n136# 0.03fF
C66 a_n224_n136# a_n128_n136# 0.33fF
C67 a_n416_n136# a_n508_n136# 0.33fF
C68 a_n416_n136# a_160_n136# 0.03fF
C69 a_352_n136# a_n416_n136# 0.02fF
C70 w_n646_n356# a_n508_n136# 0.13fF
C71 a_n32_n136# a_n508_n136# 0.04fF
C72 a_160_n136# w_n646_n356# 0.06fF
C73 a_352_n136# w_n646_n356# 0.08fF
C74 a_160_n136# a_n32_n136# 0.12fF
C75 a_352_n136# a_n32_n136# 0.05fF
C76 a_n416_n136# w_n646_n356# 0.08fF
C77 a_n416_n136# a_n32_n136# 0.05fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# a_448_n52# a_n416_n52# a_160_n52#
+ a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149# a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_448_n52# a_352_n52# 0.13fF
C1 a_n320_n52# a_n32_n52# 0.03fF
C2 a_64_n52# a_160_n52# 0.13fF
C3 a_n416_n52# a_160_n52# 0.01fF
C4 a_256_n52# a_n320_n52# 0.01fF
C5 a_n508_n52# a_n128_n52# 0.02fF
C6 a_352_n52# a_n320_n52# 0.01fF
C7 a_n508_n52# a_n512_n149# 0.03fF
C8 a_448_n52# a_n320_n52# 0.01fF
C9 a_n224_n52# a_n32_n52# 0.05fF
C10 a_64_n52# a_n508_n52# 0.01fF
C11 a_n508_n52# a_n416_n52# 0.13fF
C12 a_n224_n52# a_256_n52# 0.02fF
C13 a_n224_n52# a_352_n52# 0.01fF
C14 a_n224_n52# a_448_n52# 0.01fF
C15 a_n508_n52# a_160_n52# 0.01fF
C16 a_n32_n52# a_n128_n52# 0.13fF
C17 a_n32_n52# a_n512_n149# 0.03fF
C18 a_n224_n52# a_n320_n52# 0.13fF
C19 a_64_n52# a_n32_n52# 0.13fF
C20 a_n416_n52# a_n32_n52# 0.02fF
C21 a_256_n52# a_n128_n52# 0.02fF
C22 a_256_n52# a_n512_n149# 0.03fF
C23 a_352_n52# a_n128_n52# 0.02fF
C24 a_448_n52# a_n128_n52# 0.01fF
C25 a_352_n52# a_n512_n149# 0.03fF
C26 a_448_n52# a_n512_n149# 0.03fF
C27 a_n32_n52# a_160_n52# 0.05fF
C28 a_256_n52# a_64_n52# 0.05fF
C29 a_64_n52# a_352_n52# 0.03fF
C30 a_448_n52# a_64_n52# 0.02fF
C31 a_256_n52# a_n416_n52# 0.01fF
C32 a_352_n52# a_n416_n52# 0.01fF
C33 a_448_n52# a_n416_n52# 0.01fF
C34 a_n320_n52# a_n128_n52# 0.05fF
C35 a_n320_n52# a_n512_n149# 0.03fF
C36 a_256_n52# a_160_n52# 0.13fF
C37 a_352_n52# a_160_n52# 0.05fF
C38 a_448_n52# a_160_n52# 0.03fF
C39 a_n508_n52# a_n32_n52# 0.02fF
C40 a_64_n52# a_n320_n52# 0.02fF
C41 a_n320_n52# a_n416_n52# 0.13fF
C42 a_n224_n52# a_n128_n52# 0.13fF
C43 a_n224_n52# a_n512_n149# 0.03fF
C44 a_256_n52# a_n508_n52# 0.01fF
C45 a_n320_n52# a_160_n52# 0.02fF
C46 a_n508_n52# a_352_n52# 0.01fF
C47 a_448_n52# a_n508_n52# 0.01fF
C48 a_n224_n52# a_64_n52# 0.03fF
C49 a_n224_n52# a_n416_n52# 0.05fF
C50 a_n224_n52# a_160_n52# 0.02fF
C51 a_n508_n52# a_n320_n52# 0.05fF
C52 a_n512_n149# a_n128_n52# 0.03fF
C53 a_256_n52# a_n32_n52# 0.03fF
C54 a_352_n52# a_n32_n52# 0.02fF
C55 a_448_n52# a_n32_n52# 0.02fF
C56 a_64_n52# a_n128_n52# 0.05fF
C57 a_64_n52# a_n512_n149# 0.03fF
C58 a_n416_n52# a_n128_n52# 0.03fF
C59 a_n224_n52# a_n508_n52# 0.03fF
C60 a_n416_n52# a_n512_n149# 0.03fF
C61 a_64_n52# a_n416_n52# 0.02fF
C62 a_160_n52# a_n128_n52# 0.03fF
C63 a_256_n52# a_352_n52# 0.13fF
C64 a_256_n52# a_448_n52# 0.05fF
C65 a_n512_n149# a_160_n52# 0.03fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate in out en en_b VDD VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in out in in VSS out in out out en out nmos_tgate
C0 in en_b 0.15fF
C1 en VDD 0.12fF
C2 VDD out 0.29fF
C3 VDD in 0.70fF
C4 VDD en_b -0.11fF
C5 en out 0.01fF
C6 en in 0.13fF
C7 en en_b 0.07fF
C8 out in 0.77fF
C9 out en_b 0.01fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

.subckt onebit_dac v_hi v_lo v v_b out VDD VSS
Xtransmission_gate_0 v_hi out v v_b VDD VSS transmission_gate
Xtransmission_gate_1 v_lo out v_b v VDD VSS transmission_gate
C0 out v_hi 0.20fF
C1 v_b v_lo 0.40fF
C2 VDD v_lo -0.13fF
C3 out v_lo 0.30fF
C4 v_lo v_hi 0.47fF
C5 v_b v 0.53fF
C6 VDD v 0.33fF
C7 out v 0.29fF
C8 v v_hi 0.49fF
C9 v v_lo 0.46fF
C10 VDD v_b 0.62fF
C11 out v_b 1.55fF
C12 v_b v_hi 0.45fF
C13 VDD out -0.09fF
C14 VDD v_hi 0.20fF
C15 v_b VSS 0.47fF
C16 out VSS 1.99fF
C17 v_lo VSS 1.40fF
C18 v VSS 1.66fF
C19 VDD VSS 7.83fF
C20 v_hi VSS 1.57fF
.ends

