magic
tech sky130A
magscale 1 2
timestamp 1654734873
<< nwell >>
rect 1443 906 1802 1118
rect 1427 468 1802 906
<< pwell >>
rect 1430 323 1686 468
rect 1380 239 1686 323
rect 1430 4 1686 239
<< locali >>
rect 1386 1048 1767 1082
rect 1386 1014 1759 1048
rect 1386 74 1753 108
rect 1368 40 1766 74
<< viali >>
rect 312 946 346 980
rect 1272 946 1306 980
rect 1833 946 1867 980
rect 2793 946 2827 980
rect 1386 223 1420 323
rect 312 135 346 169
rect 1272 135 1306 169
rect 1833 135 1867 169
rect 2793 135 2827 169
<< metal1 >>
rect 293 937 303 989
rect 355 937 365 989
rect 1252 938 1262 990
rect 1314 938 1324 990
rect 1813 938 1823 990
rect 1875 938 1885 990
rect 2773 938 2783 990
rect 2835 938 2845 990
rect 92 441 187 493
rect 1153 451 1717 485
rect 2759 451 2942 485
rect 1517 361 1527 413
rect 1579 361 1589 413
rect 1380 323 1426 335
rect 1380 223 1386 323
rect 1420 223 1526 323
rect 1580 246 1683 323
rect 1580 239 1695 246
rect 1603 223 1695 239
rect 1380 211 1426 223
rect 292 124 302 176
rect 354 124 364 176
rect 1254 126 1264 178
rect 1316 126 1326 178
rect 1815 126 1825 178
rect 1877 126 1887 178
rect 2775 126 2785 178
rect 2837 126 2847 178
<< via1 >>
rect 303 980 355 989
rect 303 946 312 980
rect 312 946 346 980
rect 346 946 355 980
rect 303 937 355 946
rect 1262 980 1314 990
rect 1262 946 1272 980
rect 1272 946 1306 980
rect 1306 946 1314 980
rect 1262 938 1314 946
rect 1823 980 1875 990
rect 1823 946 1833 980
rect 1833 946 1867 980
rect 1867 946 1875 980
rect 1823 938 1875 946
rect 2783 980 2835 990
rect 2783 946 2793 980
rect 2793 946 2827 980
rect 2827 946 2835 980
rect 2783 938 2835 946
rect 1527 361 1579 413
rect 302 169 354 176
rect 302 135 312 169
rect 312 135 346 169
rect 346 135 354 169
rect 302 124 354 135
rect 1264 169 1316 178
rect 1264 135 1272 169
rect 1272 135 1306 169
rect 1306 135 1316 169
rect 1264 126 1316 135
rect 1825 169 1877 178
rect 1825 135 1833 169
rect 1833 135 1867 169
rect 1867 135 1877 169
rect 1825 126 1877 135
rect 2785 169 2837 178
rect 2785 135 2793 169
rect 2793 135 2827 169
rect 2827 135 2837 169
rect 2785 126 2837 135
<< metal2 >>
rect 303 990 355 999
rect 1262 990 1314 1000
rect 1823 990 1875 1000
rect 2783 990 2835 1000
rect 101 989 1262 990
rect 101 938 303 989
rect 355 938 1262 989
rect 1314 938 1823 990
rect 1875 938 2783 990
rect 2835 938 2849 990
rect 303 927 355 937
rect 1262 928 1314 938
rect 1527 413 1579 938
rect 1823 928 1875 938
rect 2783 928 2835 938
rect 1527 351 1579 361
rect 302 183 354 186
rect 394 183 460 185
rect 1264 183 1316 188
rect 1825 183 1877 188
rect 2785 183 2837 188
rect 92 178 2837 183
rect 92 176 1264 178
rect 92 131 302 176
rect 354 131 1264 176
rect 302 114 354 124
rect 394 119 460 131
rect 1316 131 1825 178
rect 1264 116 1316 126
rect 1877 131 2785 178
rect 1825 116 1877 126
rect 2785 116 2837 126
use nmos_PDN_mux2  nmos_PDN_mux2_0
timestamp 1654734873
transform 1 0 1553 0 1 312
box -73 -116 73 98
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1654734873
transform 1 0 215 0 1 55
box -53 -49 1241 1063
use transmission_gate  transmission_gate_1
timestamp 1654734873
transform 1 0 1736 0 1 55
box -53 -49 1241 1063
<< labels >>
flabel locali 1553 1056 1553 1056 1 FreeSans 400 0 0 0 VDD
port 5 n power bidirectional
flabel locali 1553 66 1553 66 1 FreeSans 400 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 114 469 114 469 1 FreeSans 400 0 0 0 in
port 1 n
flabel metal2 120 965 120 965 1 FreeSans 400 0 0 0 en_b
port 4 n
flabel metal2 114 158 114 158 1 FreeSans 400 0 0 0 en
port 3 n
flabel metal1 2927 465 2927 465 1 FreeSans 400 0 0 0 out
port 2 n
<< end >>
