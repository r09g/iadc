magic
tech sky130A
magscale 1 2
timestamp 1654894986
<< error_p >>
rect -6389 18950 -6329 25150
rect -6309 18950 -6249 25150
rect -70 18950 -10 25150
rect 10 18950 70 25150
rect 6249 18950 6309 25150
rect 6329 18950 6389 25150
rect -6389 12650 -6329 18850
rect -6309 12650 -6249 18850
rect -70 12650 -10 18850
rect 10 12650 70 18850
rect 6249 12650 6309 18850
rect 6329 12650 6389 18850
rect -6389 6350 -6329 12550
rect -6309 6350 -6249 12550
rect -70 6350 -10 12550
rect 10 6350 70 12550
rect 6249 6350 6309 12550
rect 6329 6350 6389 12550
rect -6389 50 -6329 6250
rect -6309 50 -6249 6250
rect -70 50 -10 6250
rect 10 50 70 6250
rect 6249 50 6309 6250
rect 6329 50 6389 6250
rect -6389 -6250 -6329 -50
rect -6309 -6250 -6249 -50
rect -70 -6250 -10 -50
rect 10 -6250 70 -50
rect 6249 -6250 6309 -50
rect 6329 -6250 6389 -50
rect -6389 -12550 -6329 -6350
rect -6309 -12550 -6249 -6350
rect -70 -12550 -10 -6350
rect 10 -12550 70 -6350
rect 6249 -12550 6309 -6350
rect 6329 -12550 6389 -6350
rect -6389 -18850 -6329 -12650
rect -6309 -18850 -6249 -12650
rect -70 -18850 -10 -12650
rect 10 -18850 70 -12650
rect 6249 -18850 6309 -12650
rect 6329 -18850 6389 -12650
rect -6389 -25150 -6329 -18950
rect -6309 -25150 -6249 -18950
rect -70 -25150 -10 -18950
rect 10 -25150 70 -18950
rect 6249 -25150 6309 -18950
rect 6329 -25150 6389 -18950
<< metal3 >>
rect -12628 25122 -6329 25150
rect -12628 18978 -6413 25122
rect -6349 18978 -6329 25122
rect -12628 18950 -6329 18978
rect -6309 25122 -10 25150
rect -6309 18978 -94 25122
rect -30 18978 -10 25122
rect -6309 18950 -10 18978
rect 10 25122 6309 25150
rect 10 18978 6225 25122
rect 6289 18978 6309 25122
rect 10 18950 6309 18978
rect 6329 25122 12628 25150
rect 6329 18978 12544 25122
rect 12608 18978 12628 25122
rect 6329 18950 12628 18978
rect -12628 18822 -6329 18850
rect -12628 12678 -6413 18822
rect -6349 12678 -6329 18822
rect -12628 12650 -6329 12678
rect -6309 18822 -10 18850
rect -6309 12678 -94 18822
rect -30 12678 -10 18822
rect -6309 12650 -10 12678
rect 10 18822 6309 18850
rect 10 12678 6225 18822
rect 6289 12678 6309 18822
rect 10 12650 6309 12678
rect 6329 18822 12628 18850
rect 6329 12678 12544 18822
rect 12608 12678 12628 18822
rect 6329 12650 12628 12678
rect -12628 12522 -6329 12550
rect -12628 6378 -6413 12522
rect -6349 6378 -6329 12522
rect -12628 6350 -6329 6378
rect -6309 12522 -10 12550
rect -6309 6378 -94 12522
rect -30 6378 -10 12522
rect -6309 6350 -10 6378
rect 10 12522 6309 12550
rect 10 6378 6225 12522
rect 6289 6378 6309 12522
rect 10 6350 6309 6378
rect 6329 12522 12628 12550
rect 6329 6378 12544 12522
rect 12608 6378 12628 12522
rect 6329 6350 12628 6378
rect -12628 6222 -6329 6250
rect -12628 78 -6413 6222
rect -6349 78 -6329 6222
rect -12628 50 -6329 78
rect -6309 6222 -10 6250
rect -6309 78 -94 6222
rect -30 78 -10 6222
rect -6309 50 -10 78
rect 10 6222 6309 6250
rect 10 78 6225 6222
rect 6289 78 6309 6222
rect 10 50 6309 78
rect 6329 6222 12628 6250
rect 6329 78 12544 6222
rect 12608 78 12628 6222
rect 6329 50 12628 78
rect -12628 -78 -6329 -50
rect -12628 -6222 -6413 -78
rect -6349 -6222 -6329 -78
rect -12628 -6250 -6329 -6222
rect -6309 -78 -10 -50
rect -6309 -6222 -94 -78
rect -30 -6222 -10 -78
rect -6309 -6250 -10 -6222
rect 10 -78 6309 -50
rect 10 -6222 6225 -78
rect 6289 -6222 6309 -78
rect 10 -6250 6309 -6222
rect 6329 -78 12628 -50
rect 6329 -6222 12544 -78
rect 12608 -6222 12628 -78
rect 6329 -6250 12628 -6222
rect -12628 -6378 -6329 -6350
rect -12628 -12522 -6413 -6378
rect -6349 -12522 -6329 -6378
rect -12628 -12550 -6329 -12522
rect -6309 -6378 -10 -6350
rect -6309 -12522 -94 -6378
rect -30 -12522 -10 -6378
rect -6309 -12550 -10 -12522
rect 10 -6378 6309 -6350
rect 10 -12522 6225 -6378
rect 6289 -12522 6309 -6378
rect 10 -12550 6309 -12522
rect 6329 -6378 12628 -6350
rect 6329 -12522 12544 -6378
rect 12608 -12522 12628 -6378
rect 6329 -12550 12628 -12522
rect -12628 -12678 -6329 -12650
rect -12628 -18822 -6413 -12678
rect -6349 -18822 -6329 -12678
rect -12628 -18850 -6329 -18822
rect -6309 -12678 -10 -12650
rect -6309 -18822 -94 -12678
rect -30 -18822 -10 -12678
rect -6309 -18850 -10 -18822
rect 10 -12678 6309 -12650
rect 10 -18822 6225 -12678
rect 6289 -18822 6309 -12678
rect 10 -18850 6309 -18822
rect 6329 -12678 12628 -12650
rect 6329 -18822 12544 -12678
rect 12608 -18822 12628 -12678
rect 6329 -18850 12628 -18822
rect -12628 -18978 -6329 -18950
rect -12628 -25122 -6413 -18978
rect -6349 -25122 -6329 -18978
rect -12628 -25150 -6329 -25122
rect -6309 -18978 -10 -18950
rect -6309 -25122 -94 -18978
rect -30 -25122 -10 -18978
rect -6309 -25150 -10 -25122
rect 10 -18978 6309 -18950
rect 10 -25122 6225 -18978
rect 6289 -25122 6309 -18978
rect 10 -25150 6309 -25122
rect 6329 -18978 12628 -18950
rect 6329 -25122 12544 -18978
rect 12608 -25122 12628 -18978
rect 6329 -25150 12628 -25122
<< via3 >>
rect -6413 18978 -6349 25122
rect -94 18978 -30 25122
rect 6225 18978 6289 25122
rect 12544 18978 12608 25122
rect -6413 12678 -6349 18822
rect -94 12678 -30 18822
rect 6225 12678 6289 18822
rect 12544 12678 12608 18822
rect -6413 6378 -6349 12522
rect -94 6378 -30 12522
rect 6225 6378 6289 12522
rect 12544 6378 12608 12522
rect -6413 78 -6349 6222
rect -94 78 -30 6222
rect 6225 78 6289 6222
rect 12544 78 12608 6222
rect -6413 -6222 -6349 -78
rect -94 -6222 -30 -78
rect 6225 -6222 6289 -78
rect 12544 -6222 12608 -78
rect -6413 -12522 -6349 -6378
rect -94 -12522 -30 -6378
rect 6225 -12522 6289 -6378
rect 12544 -12522 12608 -6378
rect -6413 -18822 -6349 -12678
rect -94 -18822 -30 -12678
rect 6225 -18822 6289 -12678
rect 12544 -18822 12608 -12678
rect -6413 -25122 -6349 -18978
rect -94 -25122 -30 -18978
rect 6225 -25122 6289 -18978
rect 12544 -25122 12608 -18978
<< mimcap >>
rect -12528 25010 -6528 25050
rect -12528 19090 -12488 25010
rect -6568 19090 -6528 25010
rect -12528 19050 -6528 19090
rect -6209 25010 -209 25050
rect -6209 19090 -6169 25010
rect -249 19090 -209 25010
rect -6209 19050 -209 19090
rect 110 25010 6110 25050
rect 110 19090 150 25010
rect 6070 19090 6110 25010
rect 110 19050 6110 19090
rect 6429 25010 12429 25050
rect 6429 19090 6469 25010
rect 12389 19090 12429 25010
rect 6429 19050 12429 19090
rect -12528 18710 -6528 18750
rect -12528 12790 -12488 18710
rect -6568 12790 -6528 18710
rect -12528 12750 -6528 12790
rect -6209 18710 -209 18750
rect -6209 12790 -6169 18710
rect -249 12790 -209 18710
rect -6209 12750 -209 12790
rect 110 18710 6110 18750
rect 110 12790 150 18710
rect 6070 12790 6110 18710
rect 110 12750 6110 12790
rect 6429 18710 12429 18750
rect 6429 12790 6469 18710
rect 12389 12790 12429 18710
rect 6429 12750 12429 12790
rect -12528 12410 -6528 12450
rect -12528 6490 -12488 12410
rect -6568 6490 -6528 12410
rect -12528 6450 -6528 6490
rect -6209 12410 -209 12450
rect -6209 6490 -6169 12410
rect -249 6490 -209 12410
rect -6209 6450 -209 6490
rect 110 12410 6110 12450
rect 110 6490 150 12410
rect 6070 6490 6110 12410
rect 110 6450 6110 6490
rect 6429 12410 12429 12450
rect 6429 6490 6469 12410
rect 12389 6490 12429 12410
rect 6429 6450 12429 6490
rect -12528 6110 -6528 6150
rect -12528 190 -12488 6110
rect -6568 190 -6528 6110
rect -12528 150 -6528 190
rect -6209 6110 -209 6150
rect -6209 190 -6169 6110
rect -249 190 -209 6110
rect -6209 150 -209 190
rect 110 6110 6110 6150
rect 110 190 150 6110
rect 6070 190 6110 6110
rect 110 150 6110 190
rect 6429 6110 12429 6150
rect 6429 190 6469 6110
rect 12389 190 12429 6110
rect 6429 150 12429 190
rect -12528 -190 -6528 -150
rect -12528 -6110 -12488 -190
rect -6568 -6110 -6528 -190
rect -12528 -6150 -6528 -6110
rect -6209 -190 -209 -150
rect -6209 -6110 -6169 -190
rect -249 -6110 -209 -190
rect -6209 -6150 -209 -6110
rect 110 -190 6110 -150
rect 110 -6110 150 -190
rect 6070 -6110 6110 -190
rect 110 -6150 6110 -6110
rect 6429 -190 12429 -150
rect 6429 -6110 6469 -190
rect 12389 -6110 12429 -190
rect 6429 -6150 12429 -6110
rect -12528 -6490 -6528 -6450
rect -12528 -12410 -12488 -6490
rect -6568 -12410 -6528 -6490
rect -12528 -12450 -6528 -12410
rect -6209 -6490 -209 -6450
rect -6209 -12410 -6169 -6490
rect -249 -12410 -209 -6490
rect -6209 -12450 -209 -12410
rect 110 -6490 6110 -6450
rect 110 -12410 150 -6490
rect 6070 -12410 6110 -6490
rect 110 -12450 6110 -12410
rect 6429 -6490 12429 -6450
rect 6429 -12410 6469 -6490
rect 12389 -12410 12429 -6490
rect 6429 -12450 12429 -12410
rect -12528 -12790 -6528 -12750
rect -12528 -18710 -12488 -12790
rect -6568 -18710 -6528 -12790
rect -12528 -18750 -6528 -18710
rect -6209 -12790 -209 -12750
rect -6209 -18710 -6169 -12790
rect -249 -18710 -209 -12790
rect -6209 -18750 -209 -18710
rect 110 -12790 6110 -12750
rect 110 -18710 150 -12790
rect 6070 -18710 6110 -12790
rect 110 -18750 6110 -18710
rect 6429 -12790 12429 -12750
rect 6429 -18710 6469 -12790
rect 12389 -18710 12429 -12790
rect 6429 -18750 12429 -18710
rect -12528 -19090 -6528 -19050
rect -12528 -25010 -12488 -19090
rect -6568 -25010 -6528 -19090
rect -12528 -25050 -6528 -25010
rect -6209 -19090 -209 -19050
rect -6209 -25010 -6169 -19090
rect -249 -25010 -209 -19090
rect -6209 -25050 -209 -25010
rect 110 -19090 6110 -19050
rect 110 -25010 150 -19090
rect 6070 -25010 6110 -19090
rect 110 -25050 6110 -25010
rect 6429 -19090 12429 -19050
rect 6429 -25010 6469 -19090
rect 12389 -25010 12429 -19090
rect 6429 -25050 12429 -25010
<< mimcapcontact >>
rect -12488 19090 -6568 25010
rect -6169 19090 -249 25010
rect 150 19090 6070 25010
rect 6469 19090 12389 25010
rect -12488 12790 -6568 18710
rect -6169 12790 -249 18710
rect 150 12790 6070 18710
rect 6469 12790 12389 18710
rect -12488 6490 -6568 12410
rect -6169 6490 -249 12410
rect 150 6490 6070 12410
rect 6469 6490 12389 12410
rect -12488 190 -6568 6110
rect -6169 190 -249 6110
rect 150 190 6070 6110
rect 6469 190 12389 6110
rect -12488 -6110 -6568 -190
rect -6169 -6110 -249 -190
rect 150 -6110 6070 -190
rect 6469 -6110 12389 -190
rect -12488 -12410 -6568 -6490
rect -6169 -12410 -249 -6490
rect 150 -12410 6070 -6490
rect 6469 -12410 12389 -6490
rect -12488 -18710 -6568 -12790
rect -6169 -18710 -249 -12790
rect 150 -18710 6070 -12790
rect 6469 -18710 12389 -12790
rect -12488 -25010 -6568 -19090
rect -6169 -25010 -249 -19090
rect 150 -25010 6070 -19090
rect 6469 -25010 12389 -19090
<< metal4 >>
rect -9580 25011 -9476 25200
rect -6460 25138 -6356 25200
rect -6460 25122 -6333 25138
rect -12489 25010 -6567 25011
rect -12489 19090 -12488 25010
rect -6568 19090 -6567 25010
rect -12489 19089 -6567 19090
rect -9580 18711 -9476 19089
rect -6460 18978 -6413 25122
rect -6349 18978 -6333 25122
rect -3261 25011 -3157 25200
rect -141 25138 -37 25200
rect -141 25122 -14 25138
rect -6170 25010 -248 25011
rect -6170 19090 -6169 25010
rect -249 19090 -248 25010
rect -6170 19089 -248 19090
rect -6460 18962 -6333 18978
rect -6460 18838 -6356 18962
rect -6460 18822 -6333 18838
rect -12489 18710 -6567 18711
rect -12489 12790 -12488 18710
rect -6568 12790 -6567 18710
rect -12489 12789 -6567 12790
rect -9580 12411 -9476 12789
rect -6460 12678 -6413 18822
rect -6349 12678 -6333 18822
rect -3261 18711 -3157 19089
rect -141 18978 -94 25122
rect -30 18978 -14 25122
rect 3058 25011 3162 25200
rect 6178 25138 6282 25200
rect 6178 25122 6305 25138
rect 149 25010 6071 25011
rect 149 19090 150 25010
rect 6070 19090 6071 25010
rect 149 19089 6071 19090
rect -141 18962 -14 18978
rect -141 18838 -37 18962
rect -141 18822 -14 18838
rect -6170 18710 -248 18711
rect -6170 12790 -6169 18710
rect -249 12790 -248 18710
rect -6170 12789 -248 12790
rect -6460 12662 -6333 12678
rect -6460 12538 -6356 12662
rect -6460 12522 -6333 12538
rect -12489 12410 -6567 12411
rect -12489 6490 -12488 12410
rect -6568 6490 -6567 12410
rect -12489 6489 -6567 6490
rect -9580 6111 -9476 6489
rect -6460 6378 -6413 12522
rect -6349 6378 -6333 12522
rect -3261 12411 -3157 12789
rect -141 12678 -94 18822
rect -30 12678 -14 18822
rect 3058 18711 3162 19089
rect 6178 18978 6225 25122
rect 6289 18978 6305 25122
rect 9377 25011 9481 25200
rect 12497 25138 12601 25200
rect 12497 25122 12624 25138
rect 6468 25010 12390 25011
rect 6468 19090 6469 25010
rect 12389 19090 12390 25010
rect 6468 19089 12390 19090
rect 6178 18962 6305 18978
rect 6178 18838 6282 18962
rect 6178 18822 6305 18838
rect 149 18710 6071 18711
rect 149 12790 150 18710
rect 6070 12790 6071 18710
rect 149 12789 6071 12790
rect -141 12662 -14 12678
rect -141 12538 -37 12662
rect -141 12522 -14 12538
rect -6170 12410 -248 12411
rect -6170 6490 -6169 12410
rect -249 6490 -248 12410
rect -6170 6489 -248 6490
rect -6460 6362 -6333 6378
rect -6460 6238 -6356 6362
rect -6460 6222 -6333 6238
rect -12489 6110 -6567 6111
rect -12489 190 -12488 6110
rect -6568 190 -6567 6110
rect -12489 189 -6567 190
rect -9580 -189 -9476 189
rect -6460 78 -6413 6222
rect -6349 78 -6333 6222
rect -3261 6111 -3157 6489
rect -141 6378 -94 12522
rect -30 6378 -14 12522
rect 3058 12411 3162 12789
rect 6178 12678 6225 18822
rect 6289 12678 6305 18822
rect 9377 18711 9481 19089
rect 12497 18978 12544 25122
rect 12608 18978 12624 25122
rect 12497 18962 12624 18978
rect 12497 18838 12601 18962
rect 12497 18822 12624 18838
rect 6468 18710 12390 18711
rect 6468 12790 6469 18710
rect 12389 12790 12390 18710
rect 6468 12789 12390 12790
rect 6178 12662 6305 12678
rect 6178 12538 6282 12662
rect 6178 12522 6305 12538
rect 149 12410 6071 12411
rect 149 6490 150 12410
rect 6070 6490 6071 12410
rect 149 6489 6071 6490
rect -141 6362 -14 6378
rect -141 6238 -37 6362
rect -141 6222 -14 6238
rect -6170 6110 -248 6111
rect -6170 190 -6169 6110
rect -249 190 -248 6110
rect -6170 189 -248 190
rect -6460 62 -6333 78
rect -6460 -62 -6356 62
rect -6460 -78 -6333 -62
rect -12489 -190 -6567 -189
rect -12489 -6110 -12488 -190
rect -6568 -6110 -6567 -190
rect -12489 -6111 -6567 -6110
rect -9580 -6489 -9476 -6111
rect -6460 -6222 -6413 -78
rect -6349 -6222 -6333 -78
rect -3261 -189 -3157 189
rect -141 78 -94 6222
rect -30 78 -14 6222
rect 3058 6111 3162 6489
rect 6178 6378 6225 12522
rect 6289 6378 6305 12522
rect 9377 12411 9481 12789
rect 12497 12678 12544 18822
rect 12608 12678 12624 18822
rect 12497 12662 12624 12678
rect 12497 12538 12601 12662
rect 12497 12522 12624 12538
rect 6468 12410 12390 12411
rect 6468 6490 6469 12410
rect 12389 6490 12390 12410
rect 6468 6489 12390 6490
rect 6178 6362 6305 6378
rect 6178 6238 6282 6362
rect 6178 6222 6305 6238
rect 149 6110 6071 6111
rect 149 190 150 6110
rect 6070 190 6071 6110
rect 149 189 6071 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -6170 -190 -248 -189
rect -6170 -6110 -6169 -190
rect -249 -6110 -248 -190
rect -6170 -6111 -248 -6110
rect -6460 -6238 -6333 -6222
rect -6460 -6362 -6356 -6238
rect -6460 -6378 -6333 -6362
rect -12489 -6490 -6567 -6489
rect -12489 -12410 -12488 -6490
rect -6568 -12410 -6567 -6490
rect -12489 -12411 -6567 -12410
rect -9580 -12789 -9476 -12411
rect -6460 -12522 -6413 -6378
rect -6349 -12522 -6333 -6378
rect -3261 -6489 -3157 -6111
rect -141 -6222 -94 -78
rect -30 -6222 -14 -78
rect 3058 -189 3162 189
rect 6178 78 6225 6222
rect 6289 78 6305 6222
rect 9377 6111 9481 6489
rect 12497 6378 12544 12522
rect 12608 6378 12624 12522
rect 12497 6362 12624 6378
rect 12497 6238 12601 6362
rect 12497 6222 12624 6238
rect 6468 6110 12390 6111
rect 6468 190 6469 6110
rect 12389 190 12390 6110
rect 6468 189 12390 190
rect 6178 62 6305 78
rect 6178 -62 6282 62
rect 6178 -78 6305 -62
rect 149 -190 6071 -189
rect 149 -6110 150 -190
rect 6070 -6110 6071 -190
rect 149 -6111 6071 -6110
rect -141 -6238 -14 -6222
rect -141 -6362 -37 -6238
rect -141 -6378 -14 -6362
rect -6170 -6490 -248 -6489
rect -6170 -12410 -6169 -6490
rect -249 -12410 -248 -6490
rect -6170 -12411 -248 -12410
rect -6460 -12538 -6333 -12522
rect -6460 -12662 -6356 -12538
rect -6460 -12678 -6333 -12662
rect -12489 -12790 -6567 -12789
rect -12489 -18710 -12488 -12790
rect -6568 -18710 -6567 -12790
rect -12489 -18711 -6567 -18710
rect -9580 -19089 -9476 -18711
rect -6460 -18822 -6413 -12678
rect -6349 -18822 -6333 -12678
rect -3261 -12789 -3157 -12411
rect -141 -12522 -94 -6378
rect -30 -12522 -14 -6378
rect 3058 -6489 3162 -6111
rect 6178 -6222 6225 -78
rect 6289 -6222 6305 -78
rect 9377 -189 9481 189
rect 12497 78 12544 6222
rect 12608 78 12624 6222
rect 12497 62 12624 78
rect 12497 -62 12601 62
rect 12497 -78 12624 -62
rect 6468 -190 12390 -189
rect 6468 -6110 6469 -190
rect 12389 -6110 12390 -190
rect 6468 -6111 12390 -6110
rect 6178 -6238 6305 -6222
rect 6178 -6362 6282 -6238
rect 6178 -6378 6305 -6362
rect 149 -6490 6071 -6489
rect 149 -12410 150 -6490
rect 6070 -12410 6071 -6490
rect 149 -12411 6071 -12410
rect -141 -12538 -14 -12522
rect -141 -12662 -37 -12538
rect -141 -12678 -14 -12662
rect -6170 -12790 -248 -12789
rect -6170 -18710 -6169 -12790
rect -249 -18710 -248 -12790
rect -6170 -18711 -248 -18710
rect -6460 -18838 -6333 -18822
rect -6460 -18962 -6356 -18838
rect -6460 -18978 -6333 -18962
rect -12489 -19090 -6567 -19089
rect -12489 -25010 -12488 -19090
rect -6568 -25010 -6567 -19090
rect -12489 -25011 -6567 -25010
rect -9580 -25200 -9476 -25011
rect -6460 -25122 -6413 -18978
rect -6349 -25122 -6333 -18978
rect -3261 -19089 -3157 -18711
rect -141 -18822 -94 -12678
rect -30 -18822 -14 -12678
rect 3058 -12789 3162 -12411
rect 6178 -12522 6225 -6378
rect 6289 -12522 6305 -6378
rect 9377 -6489 9481 -6111
rect 12497 -6222 12544 -78
rect 12608 -6222 12624 -78
rect 12497 -6238 12624 -6222
rect 12497 -6362 12601 -6238
rect 12497 -6378 12624 -6362
rect 6468 -6490 12390 -6489
rect 6468 -12410 6469 -6490
rect 12389 -12410 12390 -6490
rect 6468 -12411 12390 -12410
rect 6178 -12538 6305 -12522
rect 6178 -12662 6282 -12538
rect 6178 -12678 6305 -12662
rect 149 -12790 6071 -12789
rect 149 -18710 150 -12790
rect 6070 -18710 6071 -12790
rect 149 -18711 6071 -18710
rect -141 -18838 -14 -18822
rect -141 -18962 -37 -18838
rect -141 -18978 -14 -18962
rect -6170 -19090 -248 -19089
rect -6170 -25010 -6169 -19090
rect -249 -25010 -248 -19090
rect -6170 -25011 -248 -25010
rect -6460 -25138 -6333 -25122
rect -6460 -25200 -6356 -25138
rect -3261 -25200 -3157 -25011
rect -141 -25122 -94 -18978
rect -30 -25122 -14 -18978
rect 3058 -19089 3162 -18711
rect 6178 -18822 6225 -12678
rect 6289 -18822 6305 -12678
rect 9377 -12789 9481 -12411
rect 12497 -12522 12544 -6378
rect 12608 -12522 12624 -6378
rect 12497 -12538 12624 -12522
rect 12497 -12662 12601 -12538
rect 12497 -12678 12624 -12662
rect 6468 -12790 12390 -12789
rect 6468 -18710 6469 -12790
rect 12389 -18710 12390 -12790
rect 6468 -18711 12390 -18710
rect 6178 -18838 6305 -18822
rect 6178 -18962 6282 -18838
rect 6178 -18978 6305 -18962
rect 149 -19090 6071 -19089
rect 149 -25010 150 -19090
rect 6070 -25010 6071 -19090
rect 149 -25011 6071 -25010
rect -141 -25138 -14 -25122
rect -141 -25200 -37 -25138
rect 3058 -25200 3162 -25011
rect 6178 -25122 6225 -18978
rect 6289 -25122 6305 -18978
rect 9377 -19089 9481 -18711
rect 12497 -18822 12544 -12678
rect 12608 -18822 12624 -12678
rect 12497 -18838 12624 -18822
rect 12497 -18962 12601 -18838
rect 12497 -18978 12624 -18962
rect 6468 -19090 12390 -19089
rect 6468 -25010 6469 -19090
rect 12389 -25010 12390 -19090
rect 6468 -25011 12390 -25010
rect 6178 -25138 6305 -25122
rect 6178 -25200 6282 -25138
rect 9377 -25200 9481 -25011
rect 12497 -25122 12544 -18978
rect 12608 -25122 12624 -18978
rect 12497 -25138 12624 -25122
rect 12497 -25200 12601 -25138
<< properties >>
string FIXED_BBOX 6329 18950 12529 25150
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
