magic
tech sky130A
timestamp 1654894248
<< metal1 >>
rect -155 13 155 24
rect -155 -13 -141 13
rect -115 -13 -109 13
rect -83 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 83 13
rect 109 -13 115 13
rect 141 -13 155 13
rect -155 -24 155 -13
<< via1 >>
rect -141 -13 -115 13
rect -109 -13 -83 13
rect -77 -13 -51 13
rect -45 -13 -19 13
rect -13 -13 13 13
rect 19 -13 45 13
rect 51 -13 77 13
rect 83 -13 109 13
rect 115 -13 141 13
<< metal2 >>
rect -155 13 155 24
rect -155 -13 -141 13
rect -115 -13 -109 13
rect -83 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 83 13
rect 109 -13 115 13
rect 141 -13 155 13
rect -155 -24 155 -13
<< properties >>
string GDS_END 507862
string GDS_FILE digital_filter_3a.gds
string GDS_START 507154
<< end >>
