magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< metal1 >>
rect -2068 8268 -2022 8360
rect 6932 8182 6978 8360
rect -1032 7689 -948 7695
rect -3494 7647 -2106 7681
rect -3494 -1319 -3419 7647
rect -1032 7637 -1016 7689
rect -964 7637 -948 7689
rect -485 7681 2411 7697
rect -723 7647 2411 7681
rect -1032 7631 -948 7637
rect -485 7633 2411 7647
rect 6681 7691 6765 7697
rect 6681 7639 6697 7691
rect 6749 7681 6765 7691
rect 6749 7647 6899 7681
rect 8265 7647 9310 7681
rect 6749 7639 6765 7647
rect 6681 7633 6765 7639
rect -2068 7160 -2022 7246
rect -2068 6382 -2022 6560
rect 1618 6470 1702 6476
rect 1618 6418 1634 6470
rect 1686 6418 1702 6470
rect 1618 6412 1702 6418
rect -1038 5889 -954 5895
rect -2886 5847 -2090 5881
rect -2886 481 -2811 5847
rect -1038 5837 -1022 5889
rect -970 5837 -954 5889
rect -487 5887 -403 5893
rect -487 5881 -471 5887
rect -739 5847 -471 5881
rect -1038 5831 -954 5837
rect -487 5835 -471 5847
rect -419 5835 -403 5887
rect -487 5829 -403 5835
rect -2068 5360 -2022 5532
rect -2068 4582 -2022 4760
rect -1034 4089 -950 4095
rect -2428 4047 -2100 4081
rect -2428 2281 -2353 4047
rect -1034 4037 -1018 4089
rect -966 4037 -950 4089
rect -444 4088 -360 4094
rect -444 4081 -428 4088
rect -719 4047 -428 4081
rect -1034 4031 -950 4037
rect -444 4036 -428 4047
rect -376 4036 -360 4088
rect -444 4030 -360 4036
rect 1628 3846 1692 6412
rect 2347 4563 2411 7633
rect 6932 7160 6978 7332
rect 6932 6382 6978 6560
rect 6694 5889 6778 5895
rect 6694 5837 6710 5889
rect 6762 5881 6778 5889
rect 6762 5847 6894 5881
rect 8281 5847 8799 5881
rect 6762 5837 6778 5847
rect 6694 5831 6778 5837
rect 3147 5552 3231 5558
rect 3147 5500 3163 5552
rect 3215 5500 3231 5552
rect 3147 5494 3231 5500
rect 3157 5084 3221 5494
rect 6932 5360 6978 5532
rect 3147 5078 3231 5084
rect 3147 5026 3163 5078
rect 3215 5026 3231 5078
rect 3147 5020 3231 5026
rect 3831 4928 6240 4932
rect 3758 4926 6240 4928
rect 3758 4922 6172 4926
rect 3758 4870 3774 4922
rect 3826 4874 6172 4922
rect 6224 4874 6240 4926
rect 3826 4870 6240 4874
rect 3758 4868 6240 4870
rect 3758 4864 3842 4868
rect 6932 4582 6978 4760
rect 2347 4557 3180 4563
rect 2347 4505 3112 4557
rect 3164 4505 3180 4557
rect 2347 4499 3180 4505
rect 4874 4384 5281 4390
rect 4874 4332 5213 4384
rect 5265 4332 5281 4384
rect 4874 4326 5281 4332
rect 3298 4206 3382 4212
rect 3298 4154 3314 4206
rect 3366 4154 3382 4206
rect 3298 4148 3382 4154
rect 3308 4085 3372 4148
rect 1628 3782 1866 3846
rect -2068 3560 -2022 3732
rect 323 3477 1705 3483
rect 323 3425 339 3477
rect 391 3425 1637 3477
rect 1689 3425 1705 3477
rect 323 3419 1705 3425
rect 1802 3154 1866 3782
rect 323 3148 1866 3154
rect 323 3096 339 3148
rect 391 3096 1866 3148
rect 323 3090 1866 3096
rect -2068 2782 -2022 2960
rect -1037 2289 -953 2295
rect -2428 2247 -2106 2281
rect -1037 2237 -1021 2289
rect -969 2237 -953 2289
rect -444 2285 -360 2291
rect -444 2281 -428 2285
rect -719 2247 -428 2281
rect -1037 2231 -953 2237
rect -444 2233 -428 2247
rect -376 2233 -360 2285
rect -444 2227 -360 2233
rect 3308 2223 3371 4085
rect 4874 3642 4938 4326
rect 6749 4089 6833 4095
rect 6749 4037 6765 4089
rect 6817 4081 6833 4089
rect 8724 4081 8799 5847
rect 6817 4047 6894 4081
rect 8271 4047 8799 4081
rect 6817 4037 6833 4047
rect 6749 4031 6833 4037
rect 4864 3636 4948 3642
rect 4864 3584 4880 3636
rect 4932 3584 4948 3636
rect 4864 3578 4948 3584
rect 6932 3560 6978 3732
rect 6932 2782 6978 2960
rect 6754 2291 6838 2297
rect 6754 2239 6770 2291
rect 6822 2281 6838 2291
rect 8724 2281 8799 4047
rect 6822 2247 6894 2281
rect 8275 2247 8799 2281
rect 6822 2239 6838 2247
rect 6754 2233 6838 2239
rect 3298 2217 3382 2223
rect 3298 2165 3314 2217
rect 3366 2165 3382 2217
rect 3298 2159 3382 2165
rect -2068 1760 -2022 1932
rect 6932 1760 6978 1932
rect -364 1634 2404 1640
rect -364 1582 2336 1634
rect 2388 1582 2404 1634
rect -364 1576 2404 1582
rect -2068 982 -2022 1160
rect -1030 491 -946 497
rect -2886 447 -2106 481
rect -1030 439 -1014 491
rect -962 439 -946 491
rect -364 481 -300 1576
rect 3592 1520 6226 1526
rect 3592 1468 3608 1520
rect 3660 1468 6158 1520
rect 6210 1468 6226 1520
rect 3592 1462 6226 1468
rect 160 1335 4400 1341
rect 160 1283 176 1335
rect 228 1283 4332 1335
rect 4384 1283 4400 1335
rect 160 1277 4400 1283
rect 6932 982 6978 1160
rect -729 447 -300 481
rect -364 446 -300 447
rect 6690 487 6774 493
rect -1030 433 -946 439
rect 6690 435 6706 487
rect 6758 481 6774 487
rect 8724 481 8799 2247
rect 6758 447 6895 481
rect 8277 447 8799 481
rect 6758 435 6774 447
rect 6690 429 6774 435
rect -2068 -40 -2022 132
rect 6932 -40 6978 132
rect -2068 -818 -2022 -640
rect 6932 -818 6978 -640
rect -1029 -1310 -945 -1304
rect -3494 -1353 -2106 -1319
rect -1029 -1362 -1013 -1310
rect -961 -1362 -945 -1310
rect -512 -1307 -428 -1301
rect -512 -1319 -496 -1307
rect -720 -1353 -496 -1319
rect -1029 -1368 -945 -1362
rect -512 -1359 -496 -1353
rect -444 -1359 -428 -1307
rect -512 -1365 -428 -1359
rect 6708 -1305 6792 -1299
rect 6708 -1357 6724 -1305
rect 6776 -1319 6792 -1305
rect 9235 -1319 9310 7647
rect 6776 -1353 6894 -1319
rect 8271 -1353 9310 -1319
rect 6776 -1357 6792 -1353
rect 6708 -1363 6792 -1357
rect -2068 -1840 -2022 -1668
rect 6932 -1840 6978 -1668
<< via1 >>
rect -1016 7637 -964 7689
rect 6697 7639 6749 7691
rect 1634 6418 1686 6470
rect -1022 5837 -970 5889
rect -471 5835 -419 5887
rect -1018 4037 -966 4089
rect -428 4036 -376 4088
rect 6710 5837 6762 5889
rect 3163 5500 3215 5552
rect 3163 5026 3215 5078
rect 3774 4870 3826 4922
rect 6172 4874 6224 4926
rect 3112 4505 3164 4557
rect 5213 4332 5265 4384
rect 3314 4154 3366 4206
rect 339 3425 391 3477
rect 1637 3425 1689 3477
rect 339 3096 391 3148
rect -1021 2237 -969 2289
rect -428 2233 -376 2285
rect 6765 4037 6817 4089
rect 4880 3584 4932 3636
rect 6770 2239 6822 2291
rect 3314 2165 3366 2217
rect 2336 1582 2388 1634
rect -1014 439 -962 491
rect 3608 1468 3660 1520
rect 6158 1468 6210 1520
rect 176 1283 228 1335
rect 4332 1283 4384 1335
rect 6706 435 6758 487
rect -1013 -1362 -961 -1310
rect -496 -1359 -444 -1307
rect 6724 -1357 6776 -1305
<< metal2 >>
rect -2651 8194 -2587 8208
rect -2651 8138 -2647 8194
rect -2591 8186 -2587 8194
rect 8848 8194 8912 8208
rect 8848 8186 8852 8194
rect -2591 8138 -1907 8186
rect -2651 8134 -1907 8138
rect 8303 8138 8852 8186
rect 8908 8138 8912 8194
rect 8303 8134 8912 8138
rect -2651 8124 -2587 8134
rect 8848 8124 8912 8134
rect -1022 7855 2060 7919
rect -1022 7689 -958 7855
rect -1022 7637 -1016 7689
rect -964 7637 -958 7689
rect -1022 7621 -958 7637
rect -2398 7386 -2334 7400
rect -2398 7330 -2394 7386
rect -2338 7378 -2334 7386
rect -2338 7330 -1922 7378
rect -2398 7326 -1922 7330
rect -2398 7316 -2334 7326
rect 1996 6752 2060 7855
rect 6691 7693 6755 7707
rect 6691 7637 6695 7693
rect 6751 7637 6755 7693
rect 6691 7623 6755 7637
rect 8595 7387 8659 7401
rect 8595 7379 8599 7387
rect 8279 7331 8599 7379
rect 8655 7331 8659 7387
rect 8279 7327 8659 7331
rect 8595 7317 8659 7327
rect 1996 6696 2000 6752
rect 2056 6696 2060 6752
rect 1996 6682 2060 6696
rect 1628 6472 1692 6486
rect 1628 6416 1632 6472
rect 1688 6416 1692 6472
rect -2651 6394 -2587 6408
rect 1628 6402 1692 6416
rect -2651 6338 -2647 6394
rect -2591 6386 -2587 6394
rect 8848 6394 8912 6408
rect 8848 6386 8852 6394
rect -2591 6338 -1907 6386
rect -2651 6334 -1907 6338
rect 8280 6338 8852 6386
rect 8908 6338 8912 6394
rect 8280 6334 8912 6338
rect -2651 6324 -2587 6334
rect 8848 6324 8912 6334
rect -1028 5889 -964 5905
rect -1028 5837 -1022 5889
rect -970 5837 -964 5889
rect -1028 5726 -964 5837
rect -477 5889 -413 5903
rect -477 5833 -473 5889
rect -417 5833 -413 5889
rect -477 5819 -413 5833
rect 6704 5891 6768 5905
rect 6704 5835 6708 5891
rect 6764 5835 6768 5891
rect 6704 5821 6768 5835
rect 3410 5777 3474 5791
rect -1028 5662 -133 5726
rect -2398 5586 -2334 5600
rect -2398 5530 -2394 5586
rect -2338 5578 -2334 5586
rect -2338 5530 -1906 5578
rect -2398 5526 -1906 5530
rect -2398 5516 -2334 5526
rect -197 5166 -133 5662
rect 3410 5721 3414 5777
rect 3470 5721 3474 5777
rect -197 5110 -193 5166
rect -137 5110 -133 5166
rect -197 5096 -133 5110
rect 1282 5608 1346 5622
rect 1282 5552 1286 5608
rect 1342 5552 1346 5608
rect -2651 4594 -2587 4608
rect -2651 4538 -2647 4594
rect -2591 4586 -2587 4594
rect -2591 4538 -1915 4586
rect -2651 4534 -1915 4538
rect -2651 4524 -2587 4534
rect 1282 4219 1346 5552
rect 1630 5609 1694 5623
rect 1630 5553 1634 5609
rect 1690 5553 1694 5609
rect 1428 4219 1492 4229
rect -434 4215 1492 4219
rect -434 4159 1432 4215
rect 1488 4159 1492 4215
rect -434 4155 1492 4159
rect -1024 4089 -960 4105
rect -1024 4037 -1018 4089
rect -966 4037 -960 4089
rect -1024 3923 -960 4037
rect -434 4088 -370 4155
rect 1428 4145 1492 4155
rect -434 4036 -428 4088
rect -376 4036 -370 4088
rect -434 4020 -370 4036
rect -1024 3859 -369 3923
rect -2398 3786 -2334 3800
rect -2398 3730 -2394 3786
rect -2338 3778 -2334 3786
rect -2338 3730 -1918 3778
rect -2398 3726 -1918 3730
rect -2398 3716 -2334 3726
rect -433 3327 -369 3859
rect 1630 3843 1694 5553
rect 3157 5554 3221 5568
rect 3157 5498 3161 5554
rect 3217 5498 3221 5554
rect 3157 5484 3221 5498
rect 3410 5165 3474 5721
rect 8595 5587 8659 5601
rect 8595 5579 8599 5587
rect 8280 5531 8599 5579
rect 8655 5531 8659 5587
rect 8280 5527 8659 5531
rect 8595 5517 8659 5527
rect 3410 5109 3414 5165
rect 3470 5109 3474 5165
rect 3410 5095 3474 5109
rect 4658 5106 4722 5116
rect 5418 5106 5482 5116
rect 4658 5102 5482 5106
rect 3157 5080 3221 5094
rect 3157 5024 3161 5080
rect 3217 5024 3221 5080
rect 4658 5046 4662 5102
rect 4718 5046 5422 5102
rect 5478 5046 5482 5102
rect 4658 5042 5482 5046
rect 4658 5032 4722 5042
rect 5418 5032 5482 5042
rect 3157 5010 3221 5024
rect 3768 4924 3832 4938
rect 3768 4868 3772 4924
rect 3828 4868 3832 4924
rect 3768 4854 3832 4868
rect 4084 4928 4148 4938
rect 5706 4928 5770 4938
rect 4084 4924 5770 4928
rect 4084 4868 4088 4924
rect 4144 4868 5710 4924
rect 5766 4868 5770 4924
rect 4084 4864 5770 4868
rect 4084 4854 4148 4864
rect 5706 4854 5770 4864
rect 6166 4928 6230 4942
rect 6166 4872 6170 4928
rect 6226 4872 6230 4928
rect 6166 4858 6230 4872
rect 8848 4594 8912 4608
rect 8848 4586 8852 4594
rect 3106 4559 3170 4573
rect 3106 4503 3110 4559
rect 3166 4503 3170 4559
rect 8279 4538 8852 4586
rect 8908 4538 8912 4594
rect 8279 4534 8912 4538
rect 8848 4524 8912 4534
rect 3106 4489 3170 4503
rect 5207 4386 5271 4400
rect 5207 4330 5211 4386
rect 5267 4330 5271 4386
rect 5207 4316 5271 4330
rect 3308 4208 3372 4222
rect 3308 4152 3312 4208
rect 3368 4152 3372 4208
rect 3308 4138 3372 4152
rect 6759 4095 6823 4105
rect 5952 4089 6823 4095
rect 5952 4037 6765 4089
rect 6817 4037 6823 4089
rect 5952 4031 6823 4037
rect 4876 3980 4940 3990
rect 5206 3980 5270 3990
rect 4876 3976 5270 3980
rect 4876 3920 4880 3976
rect 4936 3920 5210 3976
rect 5266 3920 5270 3976
rect 4876 3916 5270 3920
rect 4876 3906 4940 3916
rect 5206 3906 5270 3916
rect 3306 3858 3370 3872
rect 1630 3779 1866 3843
rect 333 3479 397 3493
rect 333 3423 337 3479
rect 393 3423 397 3479
rect 333 3409 397 3423
rect 765 3483 829 3493
rect 1408 3483 1472 3493
rect 765 3479 1472 3483
rect 765 3423 769 3479
rect 825 3423 1412 3479
rect 1468 3423 1472 3479
rect 765 3419 1472 3423
rect 765 3409 829 3419
rect 1408 3409 1472 3419
rect 1631 3479 1695 3493
rect 1631 3423 1635 3479
rect 1691 3423 1695 3479
rect 1631 3409 1695 3423
rect 333 3327 397 3337
rect -433 3323 402 3327
rect -433 3307 337 3323
rect -434 3267 337 3307
rect 393 3267 402 3323
rect -434 3263 402 3267
rect -2651 2794 -2587 2808
rect -2651 2738 -2647 2794
rect -2591 2786 -2587 2794
rect -2591 2738 -1936 2786
rect -2651 2734 -1936 2738
rect -2651 2724 -2587 2734
rect -434 2536 -370 3263
rect 333 3253 397 3263
rect 333 3150 397 3164
rect 333 3094 337 3150
rect 393 3094 397 3150
rect 333 3080 397 3094
rect 764 3153 828 3163
rect 1802 3153 1866 3779
rect 764 3149 1866 3153
rect 764 3093 768 3149
rect 824 3093 1866 3149
rect 764 3089 1866 3093
rect 3306 3802 3310 3858
rect 3366 3802 3370 3858
rect 764 3079 828 3089
rect 3306 2619 3370 3802
rect 4874 3638 4938 3652
rect 4874 3582 4878 3638
rect 4934 3582 4938 3638
rect 4874 3568 4938 3582
rect 4510 3462 4574 3472
rect 5952 3462 6016 4031
rect 6759 4021 6823 4031
rect 8595 3787 8659 3801
rect 8595 3779 8599 3787
rect 8291 3731 8599 3779
rect 8655 3731 8659 3787
rect 8291 3727 8659 3731
rect 8595 3717 8659 3727
rect 4510 3458 6016 3462
rect 4510 3402 4514 3458
rect 4570 3402 6016 3458
rect 4510 3398 6016 3402
rect 4510 3388 4574 3398
rect 4508 3151 4572 3161
rect 4508 3147 6011 3151
rect 4508 3091 4512 3147
rect 4568 3091 6011 3147
rect 4508 3087 6011 3091
rect 4508 3077 4572 3087
rect 3306 2563 3310 2619
rect 3366 2563 3370 2619
rect 3306 2549 3370 2563
rect -1027 2472 -370 2536
rect -1027 2289 -963 2472
rect -1027 2237 -1021 2289
rect -969 2237 -963 2289
rect -1027 2221 -963 2237
rect -434 2285 -370 2301
rect -434 2233 -428 2285
rect -376 2233 -370 2285
rect 5947 2297 6011 3087
rect 8848 2794 8912 2808
rect 8848 2786 8852 2794
rect 8277 2738 8852 2786
rect 8908 2738 8912 2794
rect 8277 2734 8912 2738
rect 8848 2724 8912 2734
rect 6764 2297 6828 2307
rect 5947 2291 6828 2297
rect 5947 2239 6770 2291
rect 6822 2239 6828 2291
rect 5947 2233 6828 2239
rect -2398 1986 -2334 2000
rect -2398 1930 -2394 1986
rect -2338 1978 -2334 1986
rect -2338 1930 -1921 1978
rect -2398 1926 -1921 1930
rect -2398 1916 -2334 1926
rect -434 1674 -370 2233
rect 3308 2219 3372 2233
rect 6764 2223 6828 2233
rect 3308 2163 3312 2219
rect 3368 2163 3372 2219
rect 3308 2149 3372 2163
rect 8595 1987 8659 2001
rect 8595 1979 8599 1987
rect 8292 1931 8599 1979
rect 8655 1931 8659 1987
rect 8292 1927 8659 1931
rect 8595 1917 8659 1927
rect 4437 1704 4501 1714
rect 5426 1704 5490 1714
rect 4437 1700 5490 1704
rect 540 1674 604 1684
rect 1830 1674 1894 1684
rect -434 1670 1894 1674
rect -434 1614 544 1670
rect 600 1614 1834 1670
rect 1890 1614 1894 1670
rect -434 1610 1894 1614
rect 540 1600 604 1610
rect 1830 1600 1894 1610
rect 2330 1636 2394 1650
rect 2330 1580 2334 1636
rect 2390 1580 2394 1636
rect 4437 1644 4441 1700
rect 4497 1644 5430 1700
rect 5486 1644 5490 1700
rect 4437 1640 5490 1644
rect 4437 1630 4501 1640
rect 5426 1630 5490 1640
rect 2330 1566 2394 1580
rect 3602 1522 3666 1536
rect 3602 1466 3606 1522
rect 3662 1466 3666 1522
rect 3602 1452 3666 1466
rect 3894 1522 3958 1532
rect 5736 1522 5800 1532
rect 3894 1518 5800 1522
rect 3894 1462 3898 1518
rect 3954 1462 5740 1518
rect 5796 1462 5800 1518
rect 3894 1458 5800 1462
rect 3894 1448 3958 1458
rect 5736 1448 5800 1458
rect 6152 1522 6216 1536
rect 6152 1466 6156 1522
rect 6212 1466 6216 1522
rect 6152 1452 6216 1466
rect 170 1337 234 1351
rect 170 1281 174 1337
rect 230 1281 234 1337
rect 170 1267 234 1281
rect 930 1341 994 1351
rect 3943 1341 4007 1351
rect 930 1337 4007 1341
rect 930 1281 934 1337
rect 990 1281 3947 1337
rect 4003 1281 4007 1337
rect 930 1277 4007 1281
rect 930 1267 994 1277
rect 3943 1267 4007 1277
rect 4326 1337 4390 1351
rect 4326 1281 4330 1337
rect 4386 1281 4390 1337
rect 4326 1267 4390 1281
rect -2651 994 -2587 1008
rect -2651 938 -2647 994
rect -2591 986 -2587 994
rect 8848 994 8912 1008
rect 8848 986 8852 994
rect -2591 938 -1916 986
rect -2651 934 -1916 938
rect 8292 938 8852 986
rect 8908 938 8912 994
rect 8292 934 8912 938
rect -2651 924 -2587 934
rect 8848 924 8912 934
rect -1020 491 -956 507
rect -1020 439 -1014 491
rect -962 439 -956 491
rect -1020 348 -956 439
rect 6700 489 6764 503
rect 6700 433 6704 489
rect 6760 433 6764 489
rect 6700 419 6764 433
rect 1423 348 1487 359
rect -1020 345 1487 348
rect -1020 289 1427 345
rect 1483 289 1487 345
rect -1020 284 1487 289
rect 1423 275 1487 284
rect -2398 186 -2334 200
rect -2398 130 -2394 186
rect -2338 178 -2334 186
rect 8595 187 8659 201
rect 8595 179 8599 187
rect -2338 130 -1925 178
rect -2398 126 -1925 130
rect 8279 131 8599 179
rect 8655 131 8659 187
rect 8279 127 8659 131
rect -2398 116 -2334 126
rect 8595 117 8659 127
rect 160 -222 224 -208
rect 160 -278 164 -222
rect 220 -278 224 -222
rect -2651 -806 -2587 -792
rect -2651 -862 -2647 -806
rect -2591 -814 -2587 -806
rect -2591 -862 -1906 -814
rect -2651 -866 -1906 -862
rect -2651 -876 -2587 -866
rect -364 -1074 -300 -1064
rect -1019 -1078 -300 -1074
rect -1019 -1134 -360 -1078
rect -304 -1134 -300 -1078
rect -1019 -1138 -300 -1134
rect -1019 -1310 -955 -1138
rect -364 -1148 -300 -1138
rect -1019 -1362 -1013 -1310
rect -961 -1362 -955 -1310
rect -1019 -1378 -955 -1362
rect -502 -1301 -438 -1291
rect 160 -1301 224 -278
rect 8848 -806 8912 -792
rect 8848 -814 8852 -806
rect 8279 -862 8852 -814
rect 8908 -862 8912 -806
rect 8279 -866 8912 -862
rect 8848 -876 8912 -866
rect -502 -1307 224 -1301
rect -502 -1359 -496 -1307
rect -444 -1359 224 -1307
rect -502 -1365 224 -1359
rect 6718 -1303 6782 -1289
rect 6718 -1359 6722 -1303
rect 6778 -1359 6782 -1303
rect -502 -1375 -438 -1365
rect 6718 -1373 6782 -1359
rect -2398 -1614 -2334 -1600
rect -2398 -1670 -2394 -1614
rect -2338 -1622 -2334 -1614
rect 8595 -1613 8659 -1599
rect 8595 -1621 8599 -1613
rect -2338 -1670 -1913 -1622
rect -2398 -1674 -1913 -1670
rect 8300 -1669 8599 -1621
rect 8655 -1669 8659 -1613
rect 8300 -1673 8659 -1669
rect -2398 -1684 -2334 -1674
rect 8595 -1683 8659 -1673
<< via2 >>
rect -2647 8138 -2591 8194
rect 8852 8138 8908 8194
rect -2394 7330 -2338 7386
rect 6695 7691 6751 7693
rect 6695 7639 6697 7691
rect 6697 7639 6749 7691
rect 6749 7639 6751 7691
rect 6695 7637 6751 7639
rect 8599 7331 8655 7387
rect 2000 6696 2056 6752
rect 1632 6470 1688 6472
rect 1632 6418 1634 6470
rect 1634 6418 1686 6470
rect 1686 6418 1688 6470
rect 1632 6416 1688 6418
rect -2647 6338 -2591 6394
rect 8852 6338 8908 6394
rect -473 5887 -417 5889
rect -473 5835 -471 5887
rect -471 5835 -419 5887
rect -419 5835 -417 5887
rect -473 5833 -417 5835
rect 6708 5889 6764 5891
rect 6708 5837 6710 5889
rect 6710 5837 6762 5889
rect 6762 5837 6764 5889
rect 6708 5835 6764 5837
rect -2394 5530 -2338 5586
rect 3414 5721 3470 5777
rect -193 5110 -137 5166
rect 1286 5552 1342 5608
rect -2647 4538 -2591 4594
rect 1634 5553 1690 5609
rect 1432 4159 1488 4215
rect -2394 3730 -2338 3786
rect 3161 5552 3217 5554
rect 3161 5500 3163 5552
rect 3163 5500 3215 5552
rect 3215 5500 3217 5552
rect 3161 5498 3217 5500
rect 8599 5531 8655 5587
rect 3414 5109 3470 5165
rect 3161 5078 3217 5080
rect 3161 5026 3163 5078
rect 3163 5026 3215 5078
rect 3215 5026 3217 5078
rect 3161 5024 3217 5026
rect 4662 5046 4718 5102
rect 5422 5046 5478 5102
rect 3772 4922 3828 4924
rect 3772 4870 3774 4922
rect 3774 4870 3826 4922
rect 3826 4870 3828 4922
rect 3772 4868 3828 4870
rect 4088 4868 4144 4924
rect 5710 4868 5766 4924
rect 6170 4926 6226 4928
rect 6170 4874 6172 4926
rect 6172 4874 6224 4926
rect 6224 4874 6226 4926
rect 6170 4872 6226 4874
rect 3110 4557 3166 4559
rect 3110 4505 3112 4557
rect 3112 4505 3164 4557
rect 3164 4505 3166 4557
rect 3110 4503 3166 4505
rect 8852 4538 8908 4594
rect 5211 4384 5267 4386
rect 5211 4332 5213 4384
rect 5213 4332 5265 4384
rect 5265 4332 5267 4384
rect 5211 4330 5267 4332
rect 3312 4206 3368 4208
rect 3312 4154 3314 4206
rect 3314 4154 3366 4206
rect 3366 4154 3368 4206
rect 3312 4152 3368 4154
rect 4880 3920 4936 3976
rect 5210 3920 5266 3976
rect 337 3477 393 3479
rect 337 3425 339 3477
rect 339 3425 391 3477
rect 391 3425 393 3477
rect 337 3423 393 3425
rect 769 3423 825 3479
rect 1412 3423 1468 3479
rect 1635 3477 1691 3479
rect 1635 3425 1637 3477
rect 1637 3425 1689 3477
rect 1689 3425 1691 3477
rect 1635 3423 1691 3425
rect 337 3267 393 3323
rect -2647 2738 -2591 2794
rect 337 3148 393 3150
rect 337 3096 339 3148
rect 339 3096 391 3148
rect 391 3096 393 3148
rect 337 3094 393 3096
rect 768 3093 824 3149
rect 3310 3802 3366 3858
rect 4878 3636 4934 3638
rect 4878 3584 4880 3636
rect 4880 3584 4932 3636
rect 4932 3584 4934 3636
rect 4878 3582 4934 3584
rect 8599 3731 8655 3787
rect 4514 3402 4570 3458
rect 4512 3091 4568 3147
rect 3310 2563 3366 2619
rect 8852 2738 8908 2794
rect -2394 1930 -2338 1986
rect 3312 2217 3368 2219
rect 3312 2165 3314 2217
rect 3314 2165 3366 2217
rect 3366 2165 3368 2217
rect 3312 2163 3368 2165
rect 8599 1931 8655 1987
rect 544 1614 600 1670
rect 1834 1614 1890 1670
rect 2334 1634 2390 1636
rect 2334 1582 2336 1634
rect 2336 1582 2388 1634
rect 2388 1582 2390 1634
rect 2334 1580 2390 1582
rect 4441 1644 4497 1700
rect 5430 1644 5486 1700
rect 3606 1520 3662 1522
rect 3606 1468 3608 1520
rect 3608 1468 3660 1520
rect 3660 1468 3662 1520
rect 3606 1466 3662 1468
rect 3898 1462 3954 1518
rect 5740 1462 5796 1518
rect 6156 1520 6212 1522
rect 6156 1468 6158 1520
rect 6158 1468 6210 1520
rect 6210 1468 6212 1520
rect 6156 1466 6212 1468
rect 174 1335 230 1337
rect 174 1283 176 1335
rect 176 1283 228 1335
rect 228 1283 230 1335
rect 174 1281 230 1283
rect 934 1281 990 1337
rect 3947 1281 4003 1337
rect 4330 1335 4386 1337
rect 4330 1283 4332 1335
rect 4332 1283 4384 1335
rect 4384 1283 4386 1335
rect 4330 1281 4386 1283
rect -2647 938 -2591 994
rect 8852 938 8908 994
rect 6704 487 6760 489
rect 6704 435 6706 487
rect 6706 435 6758 487
rect 6758 435 6760 487
rect 6704 433 6760 435
rect 1427 289 1483 345
rect -2394 130 -2338 186
rect 8599 131 8655 187
rect 164 -278 220 -222
rect -2647 -862 -2591 -806
rect -360 -1134 -304 -1078
rect 8852 -862 8908 -806
rect 6722 -1305 6778 -1303
rect 6722 -1357 6724 -1305
rect 6724 -1357 6776 -1305
rect 6776 -1357 6778 -1305
rect 6722 -1359 6778 -1357
rect -2394 -1670 -2338 -1614
rect 8599 -1669 8655 -1613
<< metal3 >>
rect -2651 8203 -2587 8208
rect 8848 8203 8912 8208
rect -2661 8194 -2577 8203
rect -2661 8138 -2647 8194
rect -2591 8138 -2577 8194
rect -2661 8129 -2577 8138
rect 8838 8194 8922 8203
rect 8838 8138 8852 8194
rect 8908 8138 8922 8194
rect 8838 8129 8922 8138
rect -2651 6403 -2587 8129
rect 6681 7693 6765 7702
rect 6681 7637 6695 7693
rect 6751 7637 6765 7693
rect 6681 7628 6765 7637
rect -2398 7395 -2334 7400
rect -2408 7386 -2324 7395
rect -2408 7330 -2394 7386
rect -2338 7330 -2324 7386
rect -2408 7321 -2324 7330
rect -2661 6394 -2577 6403
rect -2661 6338 -2647 6394
rect -2591 6338 -2577 6394
rect -2661 6329 -2577 6338
rect -2651 4603 -2587 6329
rect -2398 5595 -2334 7321
rect 1975 6756 2080 6780
rect 6691 6779 6755 7628
rect 8595 7396 8659 7401
rect 8585 7387 8669 7396
rect 8585 7331 8599 7387
rect 8655 7331 8669 7387
rect 8585 7322 8669 7331
rect 1975 6692 1996 6756
rect 2060 6692 2080 6756
rect 1975 6669 2080 6692
rect 6191 6715 6755 6779
rect 6191 6515 6255 6715
rect 1618 6476 1702 6481
rect 1618 6472 1896 6476
rect 1618 6416 1632 6472
rect 1688 6416 1896 6472
rect 1618 6412 1896 6416
rect 1618 6407 1702 6412
rect 3157 6133 3698 6197
rect -497 5893 -391 5915
rect -497 5829 -477 5893
rect -413 5829 -391 5893
rect -497 5808 -391 5829
rect 1272 5612 1356 5617
rect 1110 5608 1356 5612
rect -2408 5586 -2324 5595
rect -2408 5530 -2394 5586
rect -2338 5530 -2324 5586
rect 1110 5552 1286 5608
rect 1342 5552 1356 5608
rect -2408 5521 -2324 5530
rect -2661 4594 -2577 4603
rect -2661 4538 -2647 4594
rect -2591 4538 -2577 4594
rect -2661 4529 -2577 4538
rect -2651 4524 -2587 4529
rect -2398 3795 -2334 5521
rect 544 5311 608 5551
rect 1110 5548 1356 5552
rect 1272 5543 1356 5548
rect 1616 5613 1708 5646
rect 1616 5549 1630 5613
rect 1694 5549 1708 5613
rect 3157 5563 3221 6133
rect 6686 5895 6784 5914
rect 6686 5831 6704 5895
rect 6768 5831 6784 5895
rect 6686 5814 6784 5831
rect 3400 5781 3484 5810
rect 3400 5717 3410 5781
rect 3474 5717 3484 5781
rect 3400 5693 3484 5717
rect 8595 5596 8659 7322
rect 8848 6403 8912 8129
rect 8838 6394 8922 6403
rect 8838 6338 8852 6394
rect 8908 6338 8922 6394
rect 8838 6329 8922 6338
rect 8585 5587 8669 5596
rect 1616 5524 1708 5549
rect 3147 5554 3231 5563
rect 3147 5498 3161 5554
rect 3217 5498 3231 5554
rect 8585 5531 8599 5587
rect 8655 5531 8669 5587
rect 8585 5522 8669 5531
rect 3147 5489 3231 5498
rect 544 5247 5105 5311
rect -238 5170 -98 5201
rect -238 5106 -197 5170
rect -133 5106 -98 5170
rect -238 5072 -98 5106
rect 3379 5169 3508 5177
rect 3379 5105 3410 5169
rect 3474 5105 3508 5169
rect 3379 5097 3508 5105
rect 4648 5102 4732 5111
rect 3147 5084 3231 5089
rect 754 5080 3231 5084
rect 754 5024 3161 5080
rect 3217 5024 3231 5080
rect 4648 5046 4662 5102
rect 4718 5046 4732 5102
rect 4648 5037 4732 5046
rect 754 5020 3231 5024
rect 754 4663 818 5020
rect 3147 5015 3231 5020
rect 3758 4928 3842 4933
rect 1241 4924 3842 4928
rect 1241 4868 3772 4924
rect 3828 4868 3842 4924
rect 1241 4864 3842 4868
rect -2408 3786 -2324 3795
rect -2408 3730 -2394 3786
rect -2338 3730 -2324 3786
rect -2408 3721 -2324 3730
rect 333 3488 397 3761
rect 323 3479 407 3488
rect 323 3423 337 3479
rect 393 3423 407 3479
rect 323 3414 407 3423
rect 743 3483 849 3501
rect 743 3419 765 3483
rect 829 3419 849 3483
rect 333 3332 397 3414
rect 743 3404 849 3419
rect 323 3323 407 3332
rect 323 3267 337 3323
rect 393 3267 407 3323
rect 323 3258 407 3267
rect 333 3159 397 3258
rect 323 3150 407 3159
rect 323 3094 337 3150
rect 393 3094 407 3150
rect 323 3085 407 3094
rect 745 3158 837 3183
rect 745 3153 838 3158
rect 745 3089 764 3153
rect 828 3089 838 3153
rect 333 2812 397 3085
rect 745 3084 838 3089
rect 745 3061 837 3084
rect -2651 2803 -2587 2808
rect -2661 2794 -2577 2803
rect -2661 2738 -2647 2794
rect -2591 2738 -2577 2794
rect -2661 2729 -2577 2738
rect -2651 1003 -2587 2729
rect -2398 1995 -2334 2000
rect -2408 1986 -2324 1995
rect -2408 1930 -2394 1986
rect -2338 1930 -2324 1986
rect -2408 1921 -2324 1930
rect -2661 994 -2577 1003
rect -2661 938 -2647 994
rect -2591 938 -2577 994
rect -2661 929 -2577 938
rect -2651 -797 -2587 929
rect -2398 195 -2334 1921
rect 170 1346 234 1946
rect 530 1670 614 1679
rect 530 1614 544 1670
rect 600 1614 614 1670
rect 530 1605 614 1614
rect 160 1337 244 1346
rect 160 1281 174 1337
rect 230 1281 244 1337
rect 160 1272 244 1281
rect 540 1112 604 1605
rect 910 1341 1011 1357
rect 910 1277 930 1341
rect 994 1277 1011 1341
rect 910 1259 1011 1277
rect 1241 354 1305 4864
rect 3758 4859 3842 4864
rect 4061 4928 4171 4944
rect 4061 4864 4084 4928
rect 4148 4864 4171 4928
rect 4061 4850 4171 4864
rect 4658 4712 4722 5037
rect 3081 4563 3190 4586
rect 3081 4499 3106 4563
rect 3170 4499 3190 4563
rect 3081 4479 3190 4499
rect 1418 4219 1502 4224
rect 1418 4215 1842 4219
rect 1418 4159 1432 4215
rect 1488 4159 1842 4215
rect 1418 4155 1842 4159
rect 3298 4212 3382 4217
rect 3298 4208 3698 4212
rect 1418 4150 1502 4155
rect 3298 4152 3312 4208
rect 3368 4152 3698 4208
rect 3298 4148 3698 4152
rect 3298 4143 3382 4148
rect 4862 3980 4953 4019
rect 4862 3916 4876 3980
rect 4940 3916 4953 3980
rect 3283 3862 3389 3885
rect 4862 3879 4953 3916
rect 3283 3798 3306 3862
rect 3370 3798 3389 3862
rect 3283 3778 3389 3798
rect 1397 3483 1484 3517
rect 1397 3419 1408 3483
rect 1472 3419 1484 3483
rect 1397 3388 1484 3419
rect 1621 3479 1705 3488
rect 1621 3423 1635 3479
rect 1691 3423 1705 3479
rect 1621 3414 1705 3423
rect 2348 3432 2412 3740
rect 4864 3638 4948 3647
rect 4864 3582 4878 3638
rect 4934 3582 4948 3638
rect 4864 3573 4948 3582
rect 4479 3462 4604 3492
rect 999 290 1305 354
rect 1405 349 1503 380
rect 1405 285 1423 349
rect 1487 285 1503 349
rect 1631 365 1695 3414
rect 2348 3368 3912 3432
rect 4479 3398 4510 3462
rect 4574 3398 4604 3462
rect 4479 3371 4604 3398
rect 3848 2819 3912 3368
rect 4486 3151 4590 3171
rect 4486 3087 4508 3151
rect 4572 3087 4590 3151
rect 4486 3071 4590 3087
rect 3284 2623 3390 2645
rect 3284 2559 3306 2623
rect 3370 2559 3390 2623
rect 3284 2538 3390 2559
rect 3298 2223 3382 2228
rect 2887 2219 3382 2223
rect 2887 2163 3312 2219
rect 3368 2163 3382 2219
rect 2887 2159 3382 2163
rect 3298 2154 3382 2159
rect 1830 1679 1894 1868
rect 4437 1709 4501 1893
rect 4427 1700 4511 1709
rect 1820 1670 1904 1679
rect 1820 1614 1834 1670
rect 1890 1614 1904 1670
rect 1820 1605 1904 1614
rect 2307 1640 2415 1666
rect 2307 1576 2330 1640
rect 2394 1576 2415 1640
rect 4427 1644 4441 1700
rect 4497 1644 4511 1700
rect 4427 1635 4511 1644
rect 2307 1553 2415 1576
rect 3592 1526 3676 1531
rect 3083 1522 3676 1526
rect 3083 1466 3606 1522
rect 3662 1466 3676 1522
rect 3083 1462 3676 1466
rect 1631 301 1897 365
rect 3083 363 3147 1462
rect 3592 1457 3676 1462
rect 3873 1522 3978 1546
rect 3873 1458 3894 1522
rect 3958 1458 3978 1522
rect 3873 1437 3978 1458
rect 3923 1341 4024 1360
rect 3923 1277 3943 1341
rect 4007 1277 4024 1341
rect 3923 1262 4024 1277
rect 4316 1337 4400 1346
rect 4316 1281 4330 1337
rect 4386 1281 4400 1337
rect 4316 1272 4400 1281
rect 4326 1060 4390 1272
rect 4874 448 4938 3573
rect 5041 616 5105 5247
rect 5418 5111 5482 5460
rect 5408 5102 5492 5111
rect 5408 5046 5422 5102
rect 5478 5046 5492 5102
rect 5408 5037 5492 5046
rect 5683 4928 5793 4943
rect 6166 4937 6230 5491
rect 5683 4864 5706 4928
rect 5770 4864 5793 4928
rect 5683 4849 5793 4864
rect 6156 4928 6240 4937
rect 6156 4872 6170 4928
rect 6226 4872 6240 4928
rect 6156 4863 6240 4872
rect 5197 4390 5281 4395
rect 5197 4386 5495 4390
rect 5197 4330 5211 4386
rect 5267 4330 5495 4386
rect 5197 4326 5495 4330
rect 5197 4321 5281 4326
rect 5193 3980 5284 4018
rect 5193 3916 5206 3980
rect 5270 3916 5284 3980
rect 5193 3878 5284 3916
rect 8595 3796 8659 5522
rect 8848 4603 8912 6329
rect 8838 4594 8922 4603
rect 8838 4538 8852 4594
rect 8908 4538 8922 4594
rect 8838 4529 8922 4538
rect 8585 3787 8669 3796
rect 8585 3731 8599 3787
rect 8655 3731 8669 3787
rect 8585 3722 8669 3731
rect 8595 3717 8659 3722
rect 8848 2803 8912 2808
rect 8838 2794 8922 2803
rect 8838 2738 8852 2794
rect 8908 2738 8922 2794
rect 8838 2729 8922 2738
rect 8595 1996 8659 2001
rect 8585 1987 8669 1996
rect 8585 1931 8599 1987
rect 8655 1931 8669 1987
rect 8585 1922 8669 1931
rect 5416 1700 5500 1709
rect 5416 1644 5430 1700
rect 5486 1644 5500 1700
rect 5416 1635 5500 1644
rect 5426 1079 5490 1635
rect 5715 1522 5820 1544
rect 6152 1531 6216 1903
rect 5715 1458 5736 1522
rect 5800 1458 5820 1522
rect 5715 1435 5820 1458
rect 6142 1522 6226 1531
rect 6142 1466 6156 1522
rect 6212 1466 6226 1522
rect 6142 1457 6226 1466
rect 5041 552 5566 616
rect 6683 493 6785 514
rect 4610 384 4941 448
rect 6683 429 6700 493
rect 6764 429 6785 493
rect 6683 411 6785 429
rect 2812 299 3147 363
rect 1405 260 1503 285
rect 8595 196 8659 1922
rect 8848 1003 8912 2729
rect 8838 994 8922 1003
rect 8838 938 8852 994
rect 8908 938 8922 994
rect 8838 929 8922 938
rect -2408 186 -2324 195
rect -2408 130 -2394 186
rect -2338 130 -2324 186
rect -2408 121 -2324 130
rect 8585 187 8669 196
rect 8585 131 8599 187
rect 8655 131 8669 187
rect 8585 122 8669 131
rect -2661 -806 -2577 -797
rect -2661 -862 -2647 -806
rect -2591 -862 -2577 -806
rect -2661 -871 -2577 -862
rect -2651 -876 -2587 -871
rect -2398 -1605 -2334 121
rect 139 -218 245 -195
rect 139 -282 160 -218
rect 224 -282 245 -218
rect 139 -299 245 -282
rect 6179 -442 6243 116
rect 6179 -506 6782 -442
rect -378 -1074 -280 -1056
rect -378 -1138 -364 -1074
rect -300 -1138 -280 -1074
rect -378 -1159 -280 -1138
rect 6718 -1294 6782 -506
rect 6708 -1303 6792 -1294
rect 6708 -1359 6722 -1303
rect 6778 -1359 6792 -1303
rect 6708 -1368 6792 -1359
rect 6718 -1372 6782 -1368
rect 8595 -1604 8659 122
rect 8848 -797 8912 929
rect 8838 -806 8922 -797
rect 8838 -862 8852 -806
rect 8908 -862 8922 -806
rect 8838 -871 8922 -862
rect -2408 -1614 -2324 -1605
rect -2408 -1670 -2394 -1614
rect -2338 -1670 -2324 -1614
rect -2408 -1679 -2324 -1670
rect 8585 -1613 8669 -1604
rect 8585 -1669 8599 -1613
rect 8655 -1669 8669 -1613
rect 8585 -1678 8669 -1669
rect -2398 -1684 -2334 -1679
rect 8595 -1683 8659 -1678
<< via3 >>
rect 1996 6752 2060 6756
rect 1996 6696 2000 6752
rect 2000 6696 2056 6752
rect 2056 6696 2060 6752
rect 1996 6692 2060 6696
rect -477 5889 -413 5893
rect -477 5833 -473 5889
rect -473 5833 -417 5889
rect -417 5833 -413 5889
rect -477 5829 -413 5833
rect 1630 5609 1694 5613
rect 1630 5553 1634 5609
rect 1634 5553 1690 5609
rect 1690 5553 1694 5609
rect 1630 5549 1694 5553
rect 6704 5891 6768 5895
rect 6704 5835 6708 5891
rect 6708 5835 6764 5891
rect 6764 5835 6768 5891
rect 6704 5831 6768 5835
rect 3410 5777 3474 5781
rect 3410 5721 3414 5777
rect 3414 5721 3470 5777
rect 3470 5721 3474 5777
rect 3410 5717 3474 5721
rect -197 5166 -133 5170
rect -197 5110 -193 5166
rect -193 5110 -137 5166
rect -137 5110 -133 5166
rect -197 5106 -133 5110
rect 3410 5165 3474 5169
rect 3410 5109 3414 5165
rect 3414 5109 3470 5165
rect 3470 5109 3474 5165
rect 3410 5105 3474 5109
rect 765 3479 829 3483
rect 765 3423 769 3479
rect 769 3423 825 3479
rect 825 3423 829 3479
rect 765 3419 829 3423
rect 764 3149 828 3153
rect 764 3093 768 3149
rect 768 3093 824 3149
rect 824 3093 828 3149
rect 764 3089 828 3093
rect 930 1337 994 1341
rect 930 1281 934 1337
rect 934 1281 990 1337
rect 990 1281 994 1337
rect 930 1277 994 1281
rect 4084 4924 4148 4928
rect 4084 4868 4088 4924
rect 4088 4868 4144 4924
rect 4144 4868 4148 4924
rect 4084 4864 4148 4868
rect 3106 4559 3170 4563
rect 3106 4503 3110 4559
rect 3110 4503 3166 4559
rect 3166 4503 3170 4559
rect 3106 4499 3170 4503
rect 4876 3976 4940 3980
rect 4876 3920 4880 3976
rect 4880 3920 4936 3976
rect 4936 3920 4940 3976
rect 4876 3916 4940 3920
rect 3306 3858 3370 3862
rect 3306 3802 3310 3858
rect 3310 3802 3366 3858
rect 3366 3802 3370 3858
rect 3306 3798 3370 3802
rect 1408 3479 1472 3483
rect 1408 3423 1412 3479
rect 1412 3423 1468 3479
rect 1468 3423 1472 3479
rect 1408 3419 1472 3423
rect 1423 345 1487 349
rect 1423 289 1427 345
rect 1427 289 1483 345
rect 1483 289 1487 345
rect 1423 285 1487 289
rect 4510 3458 4574 3462
rect 4510 3402 4514 3458
rect 4514 3402 4570 3458
rect 4570 3402 4574 3458
rect 4510 3398 4574 3402
rect 4508 3147 4572 3151
rect 4508 3091 4512 3147
rect 4512 3091 4568 3147
rect 4568 3091 4572 3147
rect 4508 3087 4572 3091
rect 3306 2619 3370 2623
rect 3306 2563 3310 2619
rect 3310 2563 3366 2619
rect 3366 2563 3370 2619
rect 3306 2559 3370 2563
rect 2330 1636 2394 1640
rect 2330 1580 2334 1636
rect 2334 1580 2390 1636
rect 2390 1580 2394 1636
rect 2330 1576 2394 1580
rect 3894 1518 3958 1522
rect 3894 1462 3898 1518
rect 3898 1462 3954 1518
rect 3954 1462 3958 1518
rect 3894 1458 3958 1462
rect 3943 1337 4007 1341
rect 3943 1281 3947 1337
rect 3947 1281 4003 1337
rect 4003 1281 4007 1337
rect 3943 1277 4007 1281
rect 5706 4924 5770 4928
rect 5706 4868 5710 4924
rect 5710 4868 5766 4924
rect 5766 4868 5770 4924
rect 5706 4864 5770 4868
rect 5206 3976 5270 3980
rect 5206 3920 5210 3976
rect 5210 3920 5266 3976
rect 5266 3920 5270 3976
rect 5206 3916 5270 3920
rect 5736 1518 5800 1522
rect 5736 1462 5740 1518
rect 5740 1462 5796 1518
rect 5796 1462 5800 1518
rect 5736 1458 5800 1462
rect 6700 489 6764 493
rect 6700 433 6704 489
rect 6704 433 6760 489
rect 6760 433 6764 489
rect 6700 429 6764 433
rect 160 -222 224 -218
rect 160 -278 164 -222
rect 164 -278 220 -222
rect 220 -278 224 -222
rect 160 -282 224 -278
rect -364 -1078 -300 -1074
rect -364 -1134 -360 -1078
rect -360 -1134 -304 -1078
rect -304 -1134 -300 -1078
rect -364 -1138 -300 -1134
<< metal4 >>
rect 1995 6756 2061 6757
rect 1995 6692 1996 6756
rect 2060 6692 2061 6756
rect 1995 6691 2061 6692
rect 1996 6377 2060 6691
rect 6703 5895 6769 5896
rect -478 5893 -412 5894
rect -478 5829 -477 5893
rect -413 5829 155 5893
rect 6322 5831 6704 5895
rect 6768 5831 6769 5895
rect 6703 5830 6769 5831
rect -478 5828 -412 5829
rect 3409 5781 3475 5782
rect 3409 5717 3410 5781
rect 3474 5717 3744 5781
rect 3409 5716 3475 5717
rect 1629 5613 1695 5614
rect 544 5311 608 5551
rect 1629 5549 1630 5613
rect 1694 5549 1949 5613
rect 1629 5548 1695 5549
rect 544 5247 5105 5311
rect -198 5170 -132 5171
rect -198 5106 -197 5170
rect -133 5169 -132 5170
rect 3409 5169 3475 5170
rect -133 5106 3410 5169
rect -198 5105 3410 5106
rect 3474 5105 3475 5169
rect 320 4612 384 5105
rect 3409 5104 3475 5105
rect 4083 4928 4149 4929
rect 1242 4864 4084 4928
rect 4148 4864 4150 4928
rect 765 3484 829 3761
rect 764 3483 830 3484
rect 764 3419 765 3483
rect 829 3419 830 3483
rect 764 3418 830 3419
rect 763 3153 829 3154
rect 763 3089 764 3153
rect 828 3089 829 3153
rect 763 3088 829 3089
rect 764 2811 828 3088
rect -364 1985 213 2049
rect -364 -1073 -300 1985
rect 930 1342 994 1946
rect 929 1341 995 1342
rect 929 1277 930 1341
rect 994 1277 995 1341
rect 929 1276 995 1277
rect 1242 859 1306 4864
rect 4083 4863 4149 4864
rect 3105 4563 3171 4564
rect 2808 4499 3106 4563
rect 3170 4499 3171 4563
rect 3105 4498 3171 4499
rect 4875 3980 4941 3981
rect 4875 3916 4876 3980
rect 4940 3916 4941 3980
rect 4875 3915 4941 3916
rect 3305 3862 3371 3863
rect 3305 3798 3306 3862
rect 3370 3798 3746 3862
rect 3305 3797 3371 3798
rect 1407 3483 1473 3484
rect 1407 3419 1408 3483
rect 1472 3419 1473 3483
rect 1407 3418 1473 3419
rect 2348 3432 2412 3740
rect 4510 3463 4574 3790
rect 4509 3462 4575 3463
rect 998 795 1306 859
rect 1408 813 1472 3418
rect 2348 3368 3912 3432
rect 4509 3398 4510 3462
rect 4574 3398 4575 3462
rect 4509 3397 4575 3398
rect 3848 2820 3912 3368
rect 4507 3151 4573 3152
rect 4507 3087 4508 3151
rect 4572 3087 4573 3151
rect 4507 3086 4573 3087
rect 4508 2788 4572 3086
rect 3305 2623 3371 2624
rect 2816 2559 3306 2623
rect 3370 2559 3371 2623
rect 3305 2558 3371 2559
rect 2330 1641 2394 1961
rect 2329 1640 2395 1641
rect 2329 1576 2330 1640
rect 2394 1576 2395 1640
rect 2329 1575 2395 1576
rect 3893 1522 3959 1523
rect 3083 1458 3894 1522
rect 3958 1458 3959 1522
rect 1408 749 1954 813
rect 3083 812 3147 1458
rect 3893 1457 3959 1458
rect 3943 1342 4007 1345
rect 3942 1341 4008 1342
rect 3942 1277 3943 1341
rect 4007 1277 4008 1341
rect 3942 1276 4008 1277
rect 3943 1007 4007 1276
rect 4876 844 4940 3915
rect 2812 748 3147 812
rect 4609 780 4940 844
rect 5041 616 5105 5247
rect 5706 4929 5770 5552
rect 5705 4928 5771 4929
rect 5705 4864 5706 4928
rect 5770 4864 5771 4928
rect 5705 4863 5771 4864
rect 5205 3980 5271 3981
rect 5205 3916 5206 3980
rect 5270 3916 5546 3980
rect 5205 3915 5271 3916
rect 5736 1523 5800 1953
rect 5735 1522 5801 1523
rect 5735 1458 5736 1522
rect 5800 1458 5801 1522
rect 5735 1457 5801 1458
rect 5041 552 5566 616
rect 6699 493 6765 494
rect 6384 429 6700 493
rect 6764 429 6766 493
rect 6699 428 6765 429
rect 1422 349 1488 350
rect 1420 285 1423 349
rect 1487 285 1953 349
rect 1422 284 1488 285
rect 160 -217 224 179
rect 159 -218 225 -217
rect 159 -282 160 -218
rect 224 -282 225 -218
rect 159 -283 225 -282
rect -365 -1074 -299 -1073
rect -365 -1138 -364 -1074
rect -300 -1138 -299 -1074
rect -365 -1139 -299 -1138
use transmission_gate  transmission_gate_0
timestamp 1654583101
transform -1 0 8143 0 1 7251
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1654583101
transform -1 0 -857 0 1 7251
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1654583101
transform -1 0 8143 0 1 5451
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1654583101
transform -1 0 -857 0 1 5451
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1654583101
transform -1 0 8143 0 1 3651
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1654583101
transform -1 0 -857 0 1 3651
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1654583101
transform -1 0 8143 0 1 1851
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1654583101
transform -1 0 -857 0 1 1851
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1654583101
transform -1 0 8143 0 1 51
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1654583101
transform -1 0 -857 0 1 51
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1654583101
transform -1 0 8143 0 1 -1749
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1654583101
transform -1 0 -857 0 1 -1749
box -216 -51 1283 1063
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_0
timestamp 1654583101
transform 1 0 7830 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_1
timestamp 1654583101
transform 1 0 6030 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_2
timestamp 1654583101
transform 1 0 4230 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_3
timestamp 1654583101
transform 1 0 2430 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_4
timestamp 1654583101
transform 1 0 630 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_5
timestamp 1654583101
transform 1 0 -1170 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_6
timestamp 1654583101
transform 1 0 7830 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_7
timestamp 1654583101
transform 1 0 6030 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_8
timestamp 1654583101
transform 1 0 4230 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_9
timestamp 1654583101
transform 1 0 2430 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_10
timestamp 1654583101
transform 1 0 630 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_11
timestamp 1654583101
transform 1 0 -1170 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_12
timestamp 1654583101
transform 1 0 7830 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_13
timestamp 1654583101
transform 1 0 6030 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_14
timestamp 1654583101
transform 1 0 4230 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_15
timestamp 1654583101
transform 1 0 2430 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_16
timestamp 1654583101
transform 1 0 630 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_17
timestamp 1654583101
transform 1 0 -1170 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_18
timestamp 1654583101
transform 1 0 7830 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_19
timestamp 1654583101
transform 1 0 6030 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_20
timestamp 1654583101
transform 1 0 4230 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_21
timestamp 1654583101
transform 1 0 2430 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_22
timestamp 1654583101
transform 1 0 630 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_23
timestamp 1654583101
transform 1 0 -1170 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_24
timestamp 1654583101
transform 1 0 7830 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_25
timestamp 1654583101
transform 1 0 6030 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_26
timestamp 1654583101
transform 1 0 4230 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_27
timestamp 1654583101
transform 1 0 2430 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_28
timestamp 1654583101
transform 1 0 630 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_29
timestamp 1654583101
transform 1 0 -1170 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_30
timestamp 1654583101
transform 1 0 7830 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_31
timestamp 1654583101
transform 1 0 6030 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_32
timestamp 1654583101
transform 1 0 4230 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_33
timestamp 1654583101
transform 1 0 2430 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_34
timestamp 1654583101
transform 1 0 630 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_35
timestamp 1654583101
transform 1 0 -1170 0 1 -1220
box -630 -580 528 580
<< labels >>
flabel metal3 s -2642 8019 -2642 8019 1 FreeSans 500 0 0 0 p2_b
port 1 nsew
flabel metal3 s -2389 7236 -2389 7236 1 FreeSans 500 0 0 0 p2
port 2 nsew
flabel metal3 s -2639 2626 -2639 2626 1 FreeSans 500 0 0 0 p1_b
port 3 nsew
flabel metal3 s -2389 1840 -2389 1840 1 FreeSans 500 0 0 0 p1
port 4 nsew
flabel metal3 s 8645 -1537 8645 -1537 1 FreeSans 500 0 0 0 p1
port 4 nsew
flabel metal3 s 8898 -670 8898 -670 1 FreeSans 500 0 0 0 p1_b
port 3 nsew
flabel metal3 s 8648 7246 8648 7246 1 FreeSans 500 0 0 0 p2
port 2 nsew
flabel metal3 s 8904 8016 8904 8016 1 FreeSans 500 0 0 0 p2_b
port 1 nsew
flabel metal1 s -3484 3369 -3484 3369 1 FreeSans 500 0 0 0 op
port 5 nsew
flabel metal1 s -2872 3368 -2872 3368 1 FreeSans 500 0 0 0 on
port 6 nsew
flabel metal1 s -2412 3371 -2412 3371 1 FreeSans 500 0 0 0 cmc
port 7 nsew
flabel metal1 s 8790 3295 8790 3295 1 FreeSans 500 0 0 0 cm
port 8 nsew
flabel metal1 s 9292 3298 9292 3298 1 FreeSans 500 0 0 0 bias_a
port 9 nsew
flabel metal1 s -2046 8350 -2046 8350 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s -2045 7178 -2045 7178 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s -2043 6543 -2043 6543 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s -2045 5370 -2045 5370 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s -2043 4743 -2043 4743 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s -2047 3574 -2047 3574 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s -2047 2942 -2047 2942 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s -2045 1776 -2045 1776 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s -2043 1146 -2043 1146 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s -2047 -27 -2047 -27 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s -2045 -659 -2045 -659 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s -2045 -1822 -2045 -1822 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6957 -1822 6957 -1822 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6954 -659 6954 -659 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s 6957 -26 6957 -26 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6952 1141 6952 1141 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s 6952 1776 6952 1776 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6954 2944 6954 2944 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s 6954 3579 6954 3579 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6957 4740 6957 4740 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s 6954 5375 6954 5375 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6952 6547 6952 6547 1 FreeSans 500 0 0 0 VDD
port 10 nsew
flabel metal1 s 6954 7180 6954 7180 1 FreeSans 500 0 0 0 VSS
port 11 nsew
flabel metal1 s 6954 8345 6954 8345 1 FreeSans 500 0 0 0 VDD
port 10 nsew
<< end >>
