magic
tech sky130A
timestamp 1654720150
<< error_p >>
rect -2062 90 -2033 93
rect -1852 90 -1823 93
rect -1642 90 -1613 93
rect -1432 90 -1403 93
rect -1222 90 -1193 93
rect -1012 90 -983 93
rect -802 90 -773 93
rect -592 90 -563 93
rect -382 90 -353 93
rect -172 90 -143 93
rect 38 90 67 93
rect 248 90 277 93
rect 458 90 487 93
rect 668 90 697 93
rect 878 90 907 93
rect 1088 90 1117 93
rect 1298 90 1327 93
rect 1508 90 1537 93
rect 1718 90 1747 93
rect 1928 90 1957 93
rect -2062 73 -2056 90
rect -1852 73 -1846 90
rect -1642 73 -1636 90
rect -1432 73 -1426 90
rect -1222 73 -1216 90
rect -1012 73 -1006 90
rect -802 73 -796 90
rect -592 73 -586 90
rect -382 73 -376 90
rect -172 73 -166 90
rect 38 73 44 90
rect 248 73 254 90
rect 458 73 464 90
rect 668 73 674 90
rect 878 73 884 90
rect 1088 73 1094 90
rect 1298 73 1304 90
rect 1508 73 1514 90
rect 1718 73 1724 90
rect 1928 73 1934 90
rect -2062 70 -2033 73
rect -1852 70 -1823 73
rect -1642 70 -1613 73
rect -1432 70 -1403 73
rect -1222 70 -1193 73
rect -1012 70 -983 73
rect -802 70 -773 73
rect -592 70 -563 73
rect -382 70 -353 73
rect -172 70 -143 73
rect 38 70 67 73
rect 248 70 277 73
rect 458 70 487 73
rect 668 70 697 73
rect 878 70 907 73
rect 1088 70 1117 73
rect 1298 70 1327 73
rect 1508 70 1537 73
rect 1718 70 1747 73
rect 1928 70 1957 73
rect -1957 -73 -1928 -70
rect -1747 -73 -1718 -70
rect -1537 -73 -1508 -70
rect -1327 -73 -1298 -70
rect -1117 -73 -1088 -70
rect -907 -73 -878 -70
rect -697 -73 -668 -70
rect -487 -73 -458 -70
rect -277 -73 -248 -70
rect -67 -73 -38 -70
rect 143 -73 172 -70
rect 353 -73 382 -70
rect 563 -73 592 -70
rect 773 -73 802 -70
rect 983 -73 1012 -70
rect 1193 -73 1222 -70
rect 1403 -73 1432 -70
rect 1613 -73 1642 -70
rect 1823 -73 1852 -70
rect 2033 -73 2062 -70
rect -1957 -90 -1951 -73
rect -1747 -90 -1741 -73
rect -1537 -90 -1531 -73
rect -1327 -90 -1321 -73
rect -1117 -90 -1111 -73
rect -907 -90 -901 -73
rect -697 -90 -691 -73
rect -487 -90 -481 -73
rect -277 -90 -271 -73
rect -67 -90 -61 -73
rect 143 -90 149 -73
rect 353 -90 359 -73
rect 563 -90 569 -73
rect 773 -90 779 -73
rect 983 -90 989 -73
rect 1193 -90 1199 -73
rect 1403 -90 1409 -73
rect 1613 -90 1619 -73
rect 1823 -90 1829 -73
rect 2033 -90 2039 -73
rect -1957 -93 -1928 -90
rect -1747 -93 -1718 -90
rect -1537 -93 -1508 -90
rect -1327 -93 -1298 -90
rect -1117 -93 -1088 -90
rect -907 -93 -878 -90
rect -697 -93 -668 -90
rect -487 -93 -458 -90
rect -277 -93 -248 -90
rect -67 -93 -38 -90
rect 143 -93 172 -90
rect 353 -93 382 -90
rect 563 -93 592 -90
rect 773 -93 802 -90
rect 983 -93 1012 -90
rect 1193 -93 1222 -90
rect 1403 -93 1432 -90
rect 1613 -93 1642 -90
rect 1823 -93 1852 -90
rect 2033 -93 2062 -90
rect -2061 -175 -2032 -172
rect -1851 -175 -1822 -172
rect -1641 -175 -1612 -172
rect -1431 -175 -1402 -172
rect -1221 -175 -1192 -172
rect -1011 -175 -982 -172
rect -801 -175 -772 -172
rect -591 -175 -562 -172
rect -381 -175 -352 -172
rect -171 -175 -142 -172
rect 39 -175 68 -172
rect 249 -175 278 -172
rect 459 -175 488 -172
rect 669 -175 698 -172
rect 879 -175 908 -172
rect 1089 -175 1118 -172
rect 1299 -175 1328 -172
rect 1509 -175 1538 -172
rect 1719 -175 1748 -172
rect 1929 -175 1958 -172
rect -2061 -192 -2055 -175
rect -1851 -192 -1845 -175
rect -1641 -192 -1635 -175
rect -1431 -192 -1425 -175
rect -1221 -192 -1215 -175
rect -1011 -192 -1005 -175
rect -801 -192 -795 -175
rect -591 -192 -585 -175
rect -381 -192 -375 -175
rect -171 -192 -165 -175
rect 39 -192 45 -175
rect 249 -192 255 -175
rect 459 -192 465 -175
rect 669 -192 675 -175
rect 879 -192 885 -175
rect 1089 -192 1095 -175
rect 1299 -192 1305 -175
rect 1509 -192 1515 -175
rect 1719 -192 1725 -175
rect 1929 -192 1935 -175
rect -2061 -195 -2032 -192
rect -1851 -195 -1822 -192
rect -1641 -195 -1612 -192
rect -1431 -195 -1402 -192
rect -1221 -195 -1192 -192
rect -1011 -195 -982 -192
rect -801 -195 -772 -192
rect -591 -195 -562 -192
rect -381 -195 -352 -192
rect -171 -195 -142 -192
rect 39 -195 68 -192
rect 249 -195 278 -192
rect 459 -195 488 -192
rect 669 -195 698 -192
rect 879 -195 908 -192
rect 1089 -195 1118 -192
rect 1299 -195 1328 -192
rect 1509 -195 1538 -192
rect 1719 -195 1748 -192
rect 1929 -195 1958 -192
rect -1956 -339 -1927 -336
rect -1746 -339 -1717 -336
rect -1536 -339 -1507 -336
rect -1326 -339 -1297 -336
rect -1116 -339 -1087 -336
rect -906 -339 -877 -336
rect -696 -339 -667 -336
rect -486 -339 -457 -336
rect -276 -339 -247 -336
rect -66 -339 -37 -336
rect 144 -339 173 -336
rect 354 -339 383 -336
rect 564 -339 593 -336
rect 774 -339 803 -336
rect 984 -339 1013 -336
rect 1194 -339 1223 -336
rect 1404 -339 1433 -336
rect 1614 -339 1643 -336
rect 1824 -339 1853 -336
rect 2034 -339 2063 -336
rect -1956 -356 -1950 -339
rect -1746 -356 -1740 -339
rect -1536 -356 -1530 -339
rect -1326 -356 -1320 -339
rect -1116 -356 -1110 -339
rect -906 -356 -900 -339
rect -696 -356 -690 -339
rect -486 -356 -480 -339
rect -276 -356 -270 -339
rect -66 -356 -60 -339
rect 144 -356 150 -339
rect 354 -356 360 -339
rect 564 -356 570 -339
rect 774 -356 780 -339
rect 984 -356 990 -339
rect 1194 -356 1200 -339
rect 1404 -356 1410 -339
rect 1614 -356 1620 -339
rect 1824 -356 1830 -339
rect 2034 -356 2040 -339
rect -1956 -359 -1927 -356
rect -1746 -359 -1717 -356
rect -1536 -359 -1507 -356
rect -1326 -359 -1297 -356
rect -1116 -359 -1087 -356
rect -906 -359 -877 -356
rect -696 -359 -667 -356
rect -486 -359 -457 -356
rect -276 -359 -247 -356
rect -66 -359 -37 -356
rect 144 -359 173 -356
rect 354 -359 383 -356
rect 564 -359 593 -356
rect 774 -359 803 -356
rect 984 -359 1013 -356
rect 1194 -359 1223 -356
rect 1404 -359 1433 -356
rect 1614 -359 1643 -356
rect 1824 -359 1853 -356
rect 2034 -359 2063 -356
<< nwell >>
rect -2260 -425 2260 159
<< pmos >>
rect -2160 -50 -2145 50
rect -2055 -50 -2040 50
rect -1950 -50 -1935 50
rect -1845 -50 -1830 50
rect -1740 -50 -1725 50
rect -1635 -50 -1620 50
rect -1530 -50 -1515 50
rect -1425 -50 -1410 50
rect -1320 -50 -1305 50
rect -1215 -50 -1200 50
rect -1110 -50 -1095 50
rect -1005 -50 -990 50
rect -900 -50 -885 50
rect -795 -50 -780 50
rect -690 -50 -675 50
rect -585 -50 -570 50
rect -480 -50 -465 50
rect -375 -50 -360 50
rect -270 -50 -255 50
rect -165 -50 -150 50
rect -60 -50 -45 50
rect 45 -50 60 50
rect 150 -50 165 50
rect 255 -50 270 50
rect 360 -50 375 50
rect 465 -50 480 50
rect 570 -50 585 50
rect 675 -50 690 50
rect 780 -50 795 50
rect 885 -50 900 50
rect 990 -50 1005 50
rect 1095 -50 1110 50
rect 1200 -50 1215 50
rect 1305 -50 1320 50
rect 1410 -50 1425 50
rect 1515 -50 1530 50
rect 1620 -50 1635 50
rect 1725 -50 1740 50
rect 1830 -50 1845 50
rect 1935 -50 1950 50
rect 2040 -50 2055 50
rect 2145 -50 2160 50
rect -2159 -316 -2144 -216
rect -2054 -316 -2039 -216
rect -1949 -316 -1934 -216
rect -1844 -316 -1829 -216
rect -1739 -316 -1724 -216
rect -1634 -316 -1619 -216
rect -1529 -316 -1514 -216
rect -1424 -316 -1409 -216
rect -1319 -316 -1304 -216
rect -1214 -316 -1199 -216
rect -1109 -316 -1094 -216
rect -1004 -316 -989 -216
rect -899 -316 -884 -216
rect -794 -316 -779 -216
rect -689 -316 -674 -216
rect -584 -316 -569 -216
rect -479 -316 -464 -216
rect -374 -316 -359 -216
rect -269 -316 -254 -216
rect -164 -316 -149 -216
rect -59 -316 -44 -216
rect 46 -316 61 -216
rect 151 -316 166 -216
rect 256 -316 271 -216
rect 361 -316 376 -216
rect 466 -316 481 -216
rect 571 -316 586 -216
rect 676 -316 691 -216
rect 781 -316 796 -216
rect 886 -316 901 -216
rect 991 -316 1006 -216
rect 1096 -316 1111 -216
rect 1201 -316 1216 -216
rect 1306 -316 1321 -216
rect 1411 -316 1426 -216
rect 1516 -316 1531 -216
rect 1621 -316 1636 -216
rect 1726 -316 1741 -216
rect 1831 -316 1846 -216
rect 1936 -316 1951 -216
rect 2041 -316 2056 -216
rect 2146 -316 2161 -216
<< pdiff >>
rect -2191 44 -2160 50
rect -2191 -44 -2185 44
rect -2168 -44 -2160 44
rect -2191 -50 -2160 -44
rect -2145 44 -2114 50
rect -2145 -44 -2137 44
rect -2120 -44 -2114 44
rect -2145 -50 -2114 -44
rect -2086 44 -2055 50
rect -2086 -44 -2080 44
rect -2063 -44 -2055 44
rect -2086 -50 -2055 -44
rect -2040 44 -2009 50
rect -2040 -44 -2032 44
rect -2015 -44 -2009 44
rect -2040 -50 -2009 -44
rect -1981 44 -1950 50
rect -1981 -44 -1975 44
rect -1958 -44 -1950 44
rect -1981 -50 -1950 -44
rect -1935 44 -1904 50
rect -1935 -44 -1927 44
rect -1910 -44 -1904 44
rect -1935 -50 -1904 -44
rect -1876 44 -1845 50
rect -1876 -44 -1870 44
rect -1853 -44 -1845 44
rect -1876 -50 -1845 -44
rect -1830 44 -1799 50
rect -1830 -44 -1822 44
rect -1805 -44 -1799 44
rect -1830 -50 -1799 -44
rect -1771 44 -1740 50
rect -1771 -44 -1765 44
rect -1748 -44 -1740 44
rect -1771 -50 -1740 -44
rect -1725 44 -1694 50
rect -1725 -44 -1717 44
rect -1700 -44 -1694 44
rect -1725 -50 -1694 -44
rect -1666 44 -1635 50
rect -1666 -44 -1660 44
rect -1643 -44 -1635 44
rect -1666 -50 -1635 -44
rect -1620 44 -1589 50
rect -1620 -44 -1612 44
rect -1595 -44 -1589 44
rect -1620 -50 -1589 -44
rect -1561 44 -1530 50
rect -1561 -44 -1555 44
rect -1538 -44 -1530 44
rect -1561 -50 -1530 -44
rect -1515 44 -1484 50
rect -1515 -44 -1507 44
rect -1490 -44 -1484 44
rect -1515 -50 -1484 -44
rect -1456 44 -1425 50
rect -1456 -44 -1450 44
rect -1433 -44 -1425 44
rect -1456 -50 -1425 -44
rect -1410 44 -1379 50
rect -1410 -44 -1402 44
rect -1385 -44 -1379 44
rect -1410 -50 -1379 -44
rect -1351 44 -1320 50
rect -1351 -44 -1345 44
rect -1328 -44 -1320 44
rect -1351 -50 -1320 -44
rect -1305 44 -1274 50
rect -1305 -44 -1297 44
rect -1280 -44 -1274 44
rect -1305 -50 -1274 -44
rect -1246 44 -1215 50
rect -1246 -44 -1240 44
rect -1223 -44 -1215 44
rect -1246 -50 -1215 -44
rect -1200 44 -1169 50
rect -1200 -44 -1192 44
rect -1175 -44 -1169 44
rect -1200 -50 -1169 -44
rect -1141 44 -1110 50
rect -1141 -44 -1135 44
rect -1118 -44 -1110 44
rect -1141 -50 -1110 -44
rect -1095 44 -1064 50
rect -1095 -44 -1087 44
rect -1070 -44 -1064 44
rect -1095 -50 -1064 -44
rect -1036 44 -1005 50
rect -1036 -44 -1030 44
rect -1013 -44 -1005 44
rect -1036 -50 -1005 -44
rect -990 44 -959 50
rect -990 -44 -982 44
rect -965 -44 -959 44
rect -990 -50 -959 -44
rect -931 44 -900 50
rect -931 -44 -925 44
rect -908 -44 -900 44
rect -931 -50 -900 -44
rect -885 44 -854 50
rect -885 -44 -877 44
rect -860 -44 -854 44
rect -885 -50 -854 -44
rect -826 44 -795 50
rect -826 -44 -820 44
rect -803 -44 -795 44
rect -826 -50 -795 -44
rect -780 44 -749 50
rect -780 -44 -772 44
rect -755 -44 -749 44
rect -780 -50 -749 -44
rect -721 44 -690 50
rect -721 -44 -715 44
rect -698 -44 -690 44
rect -721 -50 -690 -44
rect -675 44 -644 50
rect -675 -44 -667 44
rect -650 -44 -644 44
rect -675 -50 -644 -44
rect -616 44 -585 50
rect -616 -44 -610 44
rect -593 -44 -585 44
rect -616 -50 -585 -44
rect -570 44 -539 50
rect -570 -44 -562 44
rect -545 -44 -539 44
rect -570 -50 -539 -44
rect -511 44 -480 50
rect -511 -44 -505 44
rect -488 -44 -480 44
rect -511 -50 -480 -44
rect -465 44 -434 50
rect -465 -44 -457 44
rect -440 -44 -434 44
rect -465 -50 -434 -44
rect -406 44 -375 50
rect -406 -44 -400 44
rect -383 -44 -375 44
rect -406 -50 -375 -44
rect -360 44 -329 50
rect -360 -44 -352 44
rect -335 -44 -329 44
rect -360 -50 -329 -44
rect -301 44 -270 50
rect -301 -44 -295 44
rect -278 -44 -270 44
rect -301 -50 -270 -44
rect -255 44 -224 50
rect -255 -44 -247 44
rect -230 -44 -224 44
rect -255 -50 -224 -44
rect -196 44 -165 50
rect -196 -44 -190 44
rect -173 -44 -165 44
rect -196 -50 -165 -44
rect -150 44 -119 50
rect -150 -44 -142 44
rect -125 -44 -119 44
rect -150 -50 -119 -44
rect -91 44 -60 50
rect -91 -44 -85 44
rect -68 -44 -60 44
rect -91 -50 -60 -44
rect -45 44 -14 50
rect -45 -44 -37 44
rect -20 -44 -14 44
rect -45 -50 -14 -44
rect 14 44 45 50
rect 14 -44 20 44
rect 37 -44 45 44
rect 14 -50 45 -44
rect 60 44 91 50
rect 60 -44 68 44
rect 85 -44 91 44
rect 60 -50 91 -44
rect 119 44 150 50
rect 119 -44 125 44
rect 142 -44 150 44
rect 119 -50 150 -44
rect 165 44 196 50
rect 165 -44 173 44
rect 190 -44 196 44
rect 165 -50 196 -44
rect 224 44 255 50
rect 224 -44 230 44
rect 247 -44 255 44
rect 224 -50 255 -44
rect 270 44 301 50
rect 270 -44 278 44
rect 295 -44 301 44
rect 270 -50 301 -44
rect 329 44 360 50
rect 329 -44 335 44
rect 352 -44 360 44
rect 329 -50 360 -44
rect 375 44 406 50
rect 375 -44 383 44
rect 400 -44 406 44
rect 375 -50 406 -44
rect 434 44 465 50
rect 434 -44 440 44
rect 457 -44 465 44
rect 434 -50 465 -44
rect 480 44 511 50
rect 480 -44 488 44
rect 505 -44 511 44
rect 480 -50 511 -44
rect 539 44 570 50
rect 539 -44 545 44
rect 562 -44 570 44
rect 539 -50 570 -44
rect 585 44 616 50
rect 585 -44 593 44
rect 610 -44 616 44
rect 585 -50 616 -44
rect 644 44 675 50
rect 644 -44 650 44
rect 667 -44 675 44
rect 644 -50 675 -44
rect 690 44 721 50
rect 690 -44 698 44
rect 715 -44 721 44
rect 690 -50 721 -44
rect 749 44 780 50
rect 749 -44 755 44
rect 772 -44 780 44
rect 749 -50 780 -44
rect 795 44 826 50
rect 795 -44 803 44
rect 820 -44 826 44
rect 795 -50 826 -44
rect 854 44 885 50
rect 854 -44 860 44
rect 877 -44 885 44
rect 854 -50 885 -44
rect 900 44 931 50
rect 900 -44 908 44
rect 925 -44 931 44
rect 900 -50 931 -44
rect 959 44 990 50
rect 959 -44 965 44
rect 982 -44 990 44
rect 959 -50 990 -44
rect 1005 44 1036 50
rect 1005 -44 1013 44
rect 1030 -44 1036 44
rect 1005 -50 1036 -44
rect 1064 44 1095 50
rect 1064 -44 1070 44
rect 1087 -44 1095 44
rect 1064 -50 1095 -44
rect 1110 44 1141 50
rect 1110 -44 1118 44
rect 1135 -44 1141 44
rect 1110 -50 1141 -44
rect 1169 44 1200 50
rect 1169 -44 1175 44
rect 1192 -44 1200 44
rect 1169 -50 1200 -44
rect 1215 44 1246 50
rect 1215 -44 1223 44
rect 1240 -44 1246 44
rect 1215 -50 1246 -44
rect 1274 44 1305 50
rect 1274 -44 1280 44
rect 1297 -44 1305 44
rect 1274 -50 1305 -44
rect 1320 44 1351 50
rect 1320 -44 1328 44
rect 1345 -44 1351 44
rect 1320 -50 1351 -44
rect 1379 44 1410 50
rect 1379 -44 1385 44
rect 1402 -44 1410 44
rect 1379 -50 1410 -44
rect 1425 44 1456 50
rect 1425 -44 1433 44
rect 1450 -44 1456 44
rect 1425 -50 1456 -44
rect 1484 44 1515 50
rect 1484 -44 1490 44
rect 1507 -44 1515 44
rect 1484 -50 1515 -44
rect 1530 44 1561 50
rect 1530 -44 1538 44
rect 1555 -44 1561 44
rect 1530 -50 1561 -44
rect 1589 44 1620 50
rect 1589 -44 1595 44
rect 1612 -44 1620 44
rect 1589 -50 1620 -44
rect 1635 44 1666 50
rect 1635 -44 1643 44
rect 1660 -44 1666 44
rect 1635 -50 1666 -44
rect 1694 44 1725 50
rect 1694 -44 1700 44
rect 1717 -44 1725 44
rect 1694 -50 1725 -44
rect 1740 44 1771 50
rect 1740 -44 1748 44
rect 1765 -44 1771 44
rect 1740 -50 1771 -44
rect 1799 44 1830 50
rect 1799 -44 1805 44
rect 1822 -44 1830 44
rect 1799 -50 1830 -44
rect 1845 44 1876 50
rect 1845 -44 1853 44
rect 1870 -44 1876 44
rect 1845 -50 1876 -44
rect 1904 44 1935 50
rect 1904 -44 1910 44
rect 1927 -44 1935 44
rect 1904 -50 1935 -44
rect 1950 44 1981 50
rect 1950 -44 1958 44
rect 1975 -44 1981 44
rect 1950 -50 1981 -44
rect 2009 44 2040 50
rect 2009 -44 2015 44
rect 2032 -44 2040 44
rect 2009 -50 2040 -44
rect 2055 44 2086 50
rect 2055 -44 2063 44
rect 2080 -44 2086 44
rect 2055 -50 2086 -44
rect 2114 44 2145 50
rect 2114 -44 2120 44
rect 2137 -44 2145 44
rect 2114 -50 2145 -44
rect 2160 44 2191 50
rect 2160 -44 2168 44
rect 2185 -44 2191 44
rect 2160 -50 2191 -44
rect -2190 -222 -2159 -216
rect -2190 -310 -2184 -222
rect -2167 -310 -2159 -222
rect -2190 -316 -2159 -310
rect -2144 -222 -2113 -216
rect -2144 -310 -2136 -222
rect -2119 -310 -2113 -222
rect -2144 -316 -2113 -310
rect -2085 -222 -2054 -216
rect -2085 -310 -2079 -222
rect -2062 -310 -2054 -222
rect -2085 -316 -2054 -310
rect -2039 -222 -2008 -216
rect -2039 -310 -2031 -222
rect -2014 -310 -2008 -222
rect -2039 -316 -2008 -310
rect -1980 -222 -1949 -216
rect -1980 -310 -1974 -222
rect -1957 -310 -1949 -222
rect -1980 -316 -1949 -310
rect -1934 -222 -1903 -216
rect -1934 -310 -1926 -222
rect -1909 -310 -1903 -222
rect -1934 -316 -1903 -310
rect -1875 -222 -1844 -216
rect -1875 -310 -1869 -222
rect -1852 -310 -1844 -222
rect -1875 -316 -1844 -310
rect -1829 -222 -1798 -216
rect -1829 -310 -1821 -222
rect -1804 -310 -1798 -222
rect -1829 -316 -1798 -310
rect -1770 -222 -1739 -216
rect -1770 -310 -1764 -222
rect -1747 -310 -1739 -222
rect -1770 -316 -1739 -310
rect -1724 -222 -1693 -216
rect -1724 -310 -1716 -222
rect -1699 -310 -1693 -222
rect -1724 -316 -1693 -310
rect -1665 -222 -1634 -216
rect -1665 -310 -1659 -222
rect -1642 -310 -1634 -222
rect -1665 -316 -1634 -310
rect -1619 -222 -1588 -216
rect -1619 -310 -1611 -222
rect -1594 -310 -1588 -222
rect -1619 -316 -1588 -310
rect -1560 -222 -1529 -216
rect -1560 -310 -1554 -222
rect -1537 -310 -1529 -222
rect -1560 -316 -1529 -310
rect -1514 -222 -1483 -216
rect -1514 -310 -1506 -222
rect -1489 -310 -1483 -222
rect -1514 -316 -1483 -310
rect -1455 -222 -1424 -216
rect -1455 -310 -1449 -222
rect -1432 -310 -1424 -222
rect -1455 -316 -1424 -310
rect -1409 -222 -1378 -216
rect -1409 -310 -1401 -222
rect -1384 -310 -1378 -222
rect -1409 -316 -1378 -310
rect -1350 -222 -1319 -216
rect -1350 -310 -1344 -222
rect -1327 -310 -1319 -222
rect -1350 -316 -1319 -310
rect -1304 -222 -1273 -216
rect -1304 -310 -1296 -222
rect -1279 -310 -1273 -222
rect -1304 -316 -1273 -310
rect -1245 -222 -1214 -216
rect -1245 -310 -1239 -222
rect -1222 -310 -1214 -222
rect -1245 -316 -1214 -310
rect -1199 -222 -1168 -216
rect -1199 -310 -1191 -222
rect -1174 -310 -1168 -222
rect -1199 -316 -1168 -310
rect -1140 -222 -1109 -216
rect -1140 -310 -1134 -222
rect -1117 -310 -1109 -222
rect -1140 -316 -1109 -310
rect -1094 -222 -1063 -216
rect -1094 -310 -1086 -222
rect -1069 -310 -1063 -222
rect -1094 -316 -1063 -310
rect -1035 -222 -1004 -216
rect -1035 -310 -1029 -222
rect -1012 -310 -1004 -222
rect -1035 -316 -1004 -310
rect -989 -222 -958 -216
rect -989 -310 -981 -222
rect -964 -310 -958 -222
rect -989 -316 -958 -310
rect -930 -222 -899 -216
rect -930 -310 -924 -222
rect -907 -310 -899 -222
rect -930 -316 -899 -310
rect -884 -222 -853 -216
rect -884 -310 -876 -222
rect -859 -310 -853 -222
rect -884 -316 -853 -310
rect -825 -222 -794 -216
rect -825 -310 -819 -222
rect -802 -310 -794 -222
rect -825 -316 -794 -310
rect -779 -222 -748 -216
rect -779 -310 -771 -222
rect -754 -310 -748 -222
rect -779 -316 -748 -310
rect -720 -222 -689 -216
rect -720 -310 -714 -222
rect -697 -310 -689 -222
rect -720 -316 -689 -310
rect -674 -222 -643 -216
rect -674 -310 -666 -222
rect -649 -310 -643 -222
rect -674 -316 -643 -310
rect -615 -222 -584 -216
rect -615 -310 -609 -222
rect -592 -310 -584 -222
rect -615 -316 -584 -310
rect -569 -222 -538 -216
rect -569 -310 -561 -222
rect -544 -310 -538 -222
rect -569 -316 -538 -310
rect -510 -222 -479 -216
rect -510 -310 -504 -222
rect -487 -310 -479 -222
rect -510 -316 -479 -310
rect -464 -222 -433 -216
rect -464 -310 -456 -222
rect -439 -310 -433 -222
rect -464 -316 -433 -310
rect -405 -222 -374 -216
rect -405 -310 -399 -222
rect -382 -310 -374 -222
rect -405 -316 -374 -310
rect -359 -222 -328 -216
rect -359 -310 -351 -222
rect -334 -310 -328 -222
rect -359 -316 -328 -310
rect -300 -222 -269 -216
rect -300 -310 -294 -222
rect -277 -310 -269 -222
rect -300 -316 -269 -310
rect -254 -222 -223 -216
rect -254 -310 -246 -222
rect -229 -310 -223 -222
rect -254 -316 -223 -310
rect -195 -222 -164 -216
rect -195 -310 -189 -222
rect -172 -310 -164 -222
rect -195 -316 -164 -310
rect -149 -222 -118 -216
rect -149 -310 -141 -222
rect -124 -310 -118 -222
rect -149 -316 -118 -310
rect -90 -222 -59 -216
rect -90 -310 -84 -222
rect -67 -310 -59 -222
rect -90 -316 -59 -310
rect -44 -222 -13 -216
rect -44 -310 -36 -222
rect -19 -310 -13 -222
rect -44 -316 -13 -310
rect 15 -222 46 -216
rect 15 -310 21 -222
rect 38 -310 46 -222
rect 15 -316 46 -310
rect 61 -222 92 -216
rect 61 -310 69 -222
rect 86 -310 92 -222
rect 61 -316 92 -310
rect 120 -222 151 -216
rect 120 -310 126 -222
rect 143 -310 151 -222
rect 120 -316 151 -310
rect 166 -222 197 -216
rect 166 -310 174 -222
rect 191 -310 197 -222
rect 166 -316 197 -310
rect 225 -222 256 -216
rect 225 -310 231 -222
rect 248 -310 256 -222
rect 225 -316 256 -310
rect 271 -222 302 -216
rect 271 -310 279 -222
rect 296 -310 302 -222
rect 271 -316 302 -310
rect 330 -222 361 -216
rect 330 -310 336 -222
rect 353 -310 361 -222
rect 330 -316 361 -310
rect 376 -222 407 -216
rect 376 -310 384 -222
rect 401 -310 407 -222
rect 376 -316 407 -310
rect 435 -222 466 -216
rect 435 -310 441 -222
rect 458 -310 466 -222
rect 435 -316 466 -310
rect 481 -222 512 -216
rect 481 -310 489 -222
rect 506 -310 512 -222
rect 481 -316 512 -310
rect 540 -222 571 -216
rect 540 -310 546 -222
rect 563 -310 571 -222
rect 540 -316 571 -310
rect 586 -222 617 -216
rect 586 -310 594 -222
rect 611 -310 617 -222
rect 586 -316 617 -310
rect 645 -222 676 -216
rect 645 -310 651 -222
rect 668 -310 676 -222
rect 645 -316 676 -310
rect 691 -222 722 -216
rect 691 -310 699 -222
rect 716 -310 722 -222
rect 691 -316 722 -310
rect 750 -222 781 -216
rect 750 -310 756 -222
rect 773 -310 781 -222
rect 750 -316 781 -310
rect 796 -222 827 -216
rect 796 -310 804 -222
rect 821 -310 827 -222
rect 796 -316 827 -310
rect 855 -222 886 -216
rect 855 -310 861 -222
rect 878 -310 886 -222
rect 855 -316 886 -310
rect 901 -222 932 -216
rect 901 -310 909 -222
rect 926 -310 932 -222
rect 901 -316 932 -310
rect 960 -222 991 -216
rect 960 -310 966 -222
rect 983 -310 991 -222
rect 960 -316 991 -310
rect 1006 -222 1037 -216
rect 1006 -310 1014 -222
rect 1031 -310 1037 -222
rect 1006 -316 1037 -310
rect 1065 -222 1096 -216
rect 1065 -310 1071 -222
rect 1088 -310 1096 -222
rect 1065 -316 1096 -310
rect 1111 -222 1142 -216
rect 1111 -310 1119 -222
rect 1136 -310 1142 -222
rect 1111 -316 1142 -310
rect 1170 -222 1201 -216
rect 1170 -310 1176 -222
rect 1193 -310 1201 -222
rect 1170 -316 1201 -310
rect 1216 -222 1247 -216
rect 1216 -310 1224 -222
rect 1241 -310 1247 -222
rect 1216 -316 1247 -310
rect 1275 -222 1306 -216
rect 1275 -310 1281 -222
rect 1298 -310 1306 -222
rect 1275 -316 1306 -310
rect 1321 -222 1352 -216
rect 1321 -310 1329 -222
rect 1346 -310 1352 -222
rect 1321 -316 1352 -310
rect 1380 -222 1411 -216
rect 1380 -310 1386 -222
rect 1403 -310 1411 -222
rect 1380 -316 1411 -310
rect 1426 -222 1457 -216
rect 1426 -310 1434 -222
rect 1451 -310 1457 -222
rect 1426 -316 1457 -310
rect 1485 -222 1516 -216
rect 1485 -310 1491 -222
rect 1508 -310 1516 -222
rect 1485 -316 1516 -310
rect 1531 -222 1562 -216
rect 1531 -310 1539 -222
rect 1556 -310 1562 -222
rect 1531 -316 1562 -310
rect 1590 -222 1621 -216
rect 1590 -310 1596 -222
rect 1613 -310 1621 -222
rect 1590 -316 1621 -310
rect 1636 -222 1667 -216
rect 1636 -310 1644 -222
rect 1661 -310 1667 -222
rect 1636 -316 1667 -310
rect 1695 -222 1726 -216
rect 1695 -310 1701 -222
rect 1718 -310 1726 -222
rect 1695 -316 1726 -310
rect 1741 -222 1772 -216
rect 1741 -310 1749 -222
rect 1766 -310 1772 -222
rect 1741 -316 1772 -310
rect 1800 -222 1831 -216
rect 1800 -310 1806 -222
rect 1823 -310 1831 -222
rect 1800 -316 1831 -310
rect 1846 -222 1877 -216
rect 1846 -310 1854 -222
rect 1871 -310 1877 -222
rect 1846 -316 1877 -310
rect 1905 -222 1936 -216
rect 1905 -310 1911 -222
rect 1928 -310 1936 -222
rect 1905 -316 1936 -310
rect 1951 -222 1982 -216
rect 1951 -310 1959 -222
rect 1976 -310 1982 -222
rect 1951 -316 1982 -310
rect 2010 -222 2041 -216
rect 2010 -310 2016 -222
rect 2033 -310 2041 -222
rect 2010 -316 2041 -310
rect 2056 -222 2087 -216
rect 2056 -310 2064 -222
rect 2081 -310 2087 -222
rect 2056 -316 2087 -310
rect 2115 -222 2146 -216
rect 2115 -310 2121 -222
rect 2138 -310 2146 -222
rect 2115 -316 2146 -310
rect 2161 -222 2192 -216
rect 2161 -310 2169 -222
rect 2186 -310 2192 -222
rect 2161 -316 2192 -310
<< pdiffc >>
rect -2185 -44 -2168 44
rect -2137 -44 -2120 44
rect -2080 -44 -2063 44
rect -2032 -44 -2015 44
rect -1975 -44 -1958 44
rect -1927 -44 -1910 44
rect -1870 -44 -1853 44
rect -1822 -44 -1805 44
rect -1765 -44 -1748 44
rect -1717 -44 -1700 44
rect -1660 -44 -1643 44
rect -1612 -44 -1595 44
rect -1555 -44 -1538 44
rect -1507 -44 -1490 44
rect -1450 -44 -1433 44
rect -1402 -44 -1385 44
rect -1345 -44 -1328 44
rect -1297 -44 -1280 44
rect -1240 -44 -1223 44
rect -1192 -44 -1175 44
rect -1135 -44 -1118 44
rect -1087 -44 -1070 44
rect -1030 -44 -1013 44
rect -982 -44 -965 44
rect -925 -44 -908 44
rect -877 -44 -860 44
rect -820 -44 -803 44
rect -772 -44 -755 44
rect -715 -44 -698 44
rect -667 -44 -650 44
rect -610 -44 -593 44
rect -562 -44 -545 44
rect -505 -44 -488 44
rect -457 -44 -440 44
rect -400 -44 -383 44
rect -352 -44 -335 44
rect -295 -44 -278 44
rect -247 -44 -230 44
rect -190 -44 -173 44
rect -142 -44 -125 44
rect -85 -44 -68 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 68 -44 85 44
rect 125 -44 142 44
rect 173 -44 190 44
rect 230 -44 247 44
rect 278 -44 295 44
rect 335 -44 352 44
rect 383 -44 400 44
rect 440 -44 457 44
rect 488 -44 505 44
rect 545 -44 562 44
rect 593 -44 610 44
rect 650 -44 667 44
rect 698 -44 715 44
rect 755 -44 772 44
rect 803 -44 820 44
rect 860 -44 877 44
rect 908 -44 925 44
rect 965 -44 982 44
rect 1013 -44 1030 44
rect 1070 -44 1087 44
rect 1118 -44 1135 44
rect 1175 -44 1192 44
rect 1223 -44 1240 44
rect 1280 -44 1297 44
rect 1328 -44 1345 44
rect 1385 -44 1402 44
rect 1433 -44 1450 44
rect 1490 -44 1507 44
rect 1538 -44 1555 44
rect 1595 -44 1612 44
rect 1643 -44 1660 44
rect 1700 -44 1717 44
rect 1748 -44 1765 44
rect 1805 -44 1822 44
rect 1853 -44 1870 44
rect 1910 -44 1927 44
rect 1958 -44 1975 44
rect 2015 -44 2032 44
rect 2063 -44 2080 44
rect 2120 -44 2137 44
rect 2168 -44 2185 44
rect -2184 -310 -2167 -222
rect -2136 -310 -2119 -222
rect -2079 -310 -2062 -222
rect -2031 -310 -2014 -222
rect -1974 -310 -1957 -222
rect -1926 -310 -1909 -222
rect -1869 -310 -1852 -222
rect -1821 -310 -1804 -222
rect -1764 -310 -1747 -222
rect -1716 -310 -1699 -222
rect -1659 -310 -1642 -222
rect -1611 -310 -1594 -222
rect -1554 -310 -1537 -222
rect -1506 -310 -1489 -222
rect -1449 -310 -1432 -222
rect -1401 -310 -1384 -222
rect -1344 -310 -1327 -222
rect -1296 -310 -1279 -222
rect -1239 -310 -1222 -222
rect -1191 -310 -1174 -222
rect -1134 -310 -1117 -222
rect -1086 -310 -1069 -222
rect -1029 -310 -1012 -222
rect -981 -310 -964 -222
rect -924 -310 -907 -222
rect -876 -310 -859 -222
rect -819 -310 -802 -222
rect -771 -310 -754 -222
rect -714 -310 -697 -222
rect -666 -310 -649 -222
rect -609 -310 -592 -222
rect -561 -310 -544 -222
rect -504 -310 -487 -222
rect -456 -310 -439 -222
rect -399 -310 -382 -222
rect -351 -310 -334 -222
rect -294 -310 -277 -222
rect -246 -310 -229 -222
rect -189 -310 -172 -222
rect -141 -310 -124 -222
rect -84 -310 -67 -222
rect -36 -310 -19 -222
rect 21 -310 38 -222
rect 69 -310 86 -222
rect 126 -310 143 -222
rect 174 -310 191 -222
rect 231 -310 248 -222
rect 279 -310 296 -222
rect 336 -310 353 -222
rect 384 -310 401 -222
rect 441 -310 458 -222
rect 489 -310 506 -222
rect 546 -310 563 -222
rect 594 -310 611 -222
rect 651 -310 668 -222
rect 699 -310 716 -222
rect 756 -310 773 -222
rect 804 -310 821 -222
rect 861 -310 878 -222
rect 909 -310 926 -222
rect 966 -310 983 -222
rect 1014 -310 1031 -222
rect 1071 -310 1088 -222
rect 1119 -310 1136 -222
rect 1176 -310 1193 -222
rect 1224 -310 1241 -222
rect 1281 -310 1298 -222
rect 1329 -310 1346 -222
rect 1386 -310 1403 -222
rect 1434 -310 1451 -222
rect 1491 -310 1508 -222
rect 1539 -310 1556 -222
rect 1596 -310 1613 -222
rect 1644 -310 1661 -222
rect 1701 -310 1718 -222
rect 1749 -310 1766 -222
rect 1806 -310 1823 -222
rect 1854 -310 1871 -222
rect 1911 -310 1928 -222
rect 1959 -310 1976 -222
rect 2016 -310 2033 -222
rect 2064 -310 2081 -222
rect 2121 -310 2138 -222
rect 2169 -310 2186 -222
<< nsubdiff >>
rect -2242 124 -2194 141
rect 2194 124 2242 141
rect -2242 93 -2225 124
rect 2225 93 2242 124
rect -2242 -172 -2225 -93
rect 2225 -172 2242 -93
rect -2242 -390 -2225 -359
rect 2225 -390 2242 -359
rect -2242 -407 -2194 -390
rect 2194 -407 2242 -390
<< nsubdiffcont >>
rect -2194 124 2194 141
rect -2242 -93 -2225 93
rect 2225 -93 2242 93
rect -2242 -359 -2225 -172
rect 2225 -359 2242 -172
rect -2194 -407 2194 -390
<< poly >>
rect -2064 90 -2031 98
rect -2064 73 -2056 90
rect -2039 73 -2031 90
rect -2064 65 -2031 73
rect -1854 90 -1821 98
rect -1854 73 -1846 90
rect -1829 73 -1821 90
rect -1854 65 -1821 73
rect -1644 90 -1611 98
rect -1644 73 -1636 90
rect -1619 73 -1611 90
rect -1644 65 -1611 73
rect -1434 90 -1401 98
rect -1434 73 -1426 90
rect -1409 73 -1401 90
rect -1434 65 -1401 73
rect -1224 90 -1191 98
rect -1224 73 -1216 90
rect -1199 73 -1191 90
rect -1224 65 -1191 73
rect -1014 90 -981 98
rect -1014 73 -1006 90
rect -989 73 -981 90
rect -1014 65 -981 73
rect -804 90 -771 98
rect -804 73 -796 90
rect -779 73 -771 90
rect -804 65 -771 73
rect -594 90 -561 98
rect -594 73 -586 90
rect -569 73 -561 90
rect -594 65 -561 73
rect -384 90 -351 98
rect -384 73 -376 90
rect -359 73 -351 90
rect -384 65 -351 73
rect -174 90 -141 98
rect -174 73 -166 90
rect -149 73 -141 90
rect -174 65 -141 73
rect 36 90 69 98
rect 36 73 44 90
rect 61 73 69 90
rect 36 65 69 73
rect 246 90 279 98
rect 246 73 254 90
rect 271 73 279 90
rect 246 65 279 73
rect 456 90 489 98
rect 456 73 464 90
rect 481 73 489 90
rect 456 65 489 73
rect 666 90 699 98
rect 666 73 674 90
rect 691 73 699 90
rect 666 65 699 73
rect 876 90 909 98
rect 876 73 884 90
rect 901 73 909 90
rect 876 65 909 73
rect 1086 90 1119 98
rect 1086 73 1094 90
rect 1111 73 1119 90
rect 1086 65 1119 73
rect 1296 90 1329 98
rect 1296 73 1304 90
rect 1321 73 1329 90
rect 1296 65 1329 73
rect 1506 90 1539 98
rect 1506 73 1514 90
rect 1531 73 1539 90
rect 1506 65 1539 73
rect 1716 90 1749 98
rect 1716 73 1724 90
rect 1741 73 1749 90
rect 1716 65 1749 73
rect 1926 90 1959 98
rect 1926 73 1934 90
rect 1951 73 1959 90
rect 1926 65 1959 73
rect 2136 90 2169 98
rect 2136 73 2144 90
rect 2161 73 2169 90
rect 2136 65 2169 73
rect -2160 50 -2145 63
rect -2055 50 -2040 65
rect -1950 50 -1935 63
rect -1845 50 -1830 65
rect -1740 50 -1725 63
rect -1635 50 -1620 65
rect -1530 50 -1515 63
rect -1425 50 -1410 65
rect -1320 50 -1305 63
rect -1215 50 -1200 65
rect -1110 50 -1095 63
rect -1005 50 -990 65
rect -900 50 -885 63
rect -795 50 -780 65
rect -690 50 -675 63
rect -585 50 -570 65
rect -480 50 -465 63
rect -375 50 -360 65
rect -270 50 -255 63
rect -165 50 -150 65
rect -60 50 -45 63
rect 45 50 60 65
rect 150 50 165 63
rect 255 50 270 65
rect 360 50 375 63
rect 465 50 480 65
rect 570 50 585 63
rect 675 50 690 65
rect 780 50 795 63
rect 885 50 900 65
rect 990 50 1005 63
rect 1095 50 1110 65
rect 1200 50 1215 63
rect 1305 50 1320 65
rect 1410 50 1425 63
rect 1515 50 1530 65
rect 1620 50 1635 63
rect 1725 50 1740 65
rect 1830 50 1845 63
rect 1935 50 1950 65
rect 2040 50 2055 63
rect 2145 50 2160 65
rect -2160 -65 -2145 -50
rect -2055 -63 -2040 -50
rect -1950 -65 -1935 -50
rect -1845 -63 -1830 -50
rect -1740 -65 -1725 -50
rect -1635 -63 -1620 -50
rect -1530 -65 -1515 -50
rect -1425 -63 -1410 -50
rect -1320 -65 -1305 -50
rect -1215 -63 -1200 -50
rect -1110 -65 -1095 -50
rect -1005 -63 -990 -50
rect -900 -65 -885 -50
rect -795 -63 -780 -50
rect -690 -65 -675 -50
rect -585 -63 -570 -50
rect -480 -65 -465 -50
rect -375 -63 -360 -50
rect -270 -65 -255 -50
rect -165 -63 -150 -50
rect -60 -65 -45 -50
rect 45 -63 60 -50
rect 150 -65 165 -50
rect 255 -63 270 -50
rect 360 -65 375 -50
rect 465 -63 480 -50
rect 570 -65 585 -50
rect 675 -63 690 -50
rect 780 -65 795 -50
rect 885 -63 900 -50
rect 990 -65 1005 -50
rect 1095 -63 1110 -50
rect 1200 -65 1215 -50
rect 1305 -63 1320 -50
rect 1410 -65 1425 -50
rect 1515 -63 1530 -50
rect 1620 -65 1635 -50
rect 1725 -63 1740 -50
rect 1830 -65 1845 -50
rect 1935 -63 1950 -50
rect 2040 -65 2055 -50
rect 2145 -63 2160 -50
rect -2169 -73 -2136 -65
rect -2169 -90 -2161 -73
rect -2144 -90 -2136 -73
rect -2169 -98 -2136 -90
rect -1959 -73 -1926 -65
rect -1959 -90 -1951 -73
rect -1934 -90 -1926 -73
rect -1959 -98 -1926 -90
rect -1749 -73 -1716 -65
rect -1749 -90 -1741 -73
rect -1724 -90 -1716 -73
rect -1749 -98 -1716 -90
rect -1539 -73 -1506 -65
rect -1539 -90 -1531 -73
rect -1514 -90 -1506 -73
rect -1539 -98 -1506 -90
rect -1329 -73 -1296 -65
rect -1329 -90 -1321 -73
rect -1304 -90 -1296 -73
rect -1329 -98 -1296 -90
rect -1119 -73 -1086 -65
rect -1119 -90 -1111 -73
rect -1094 -90 -1086 -73
rect -1119 -98 -1086 -90
rect -909 -73 -876 -65
rect -909 -90 -901 -73
rect -884 -90 -876 -73
rect -909 -98 -876 -90
rect -699 -73 -666 -65
rect -699 -90 -691 -73
rect -674 -90 -666 -73
rect -699 -98 -666 -90
rect -489 -73 -456 -65
rect -489 -90 -481 -73
rect -464 -90 -456 -73
rect -489 -98 -456 -90
rect -279 -73 -246 -65
rect -279 -90 -271 -73
rect -254 -90 -246 -73
rect -279 -98 -246 -90
rect -69 -73 -36 -65
rect -69 -90 -61 -73
rect -44 -90 -36 -73
rect -69 -98 -36 -90
rect 141 -73 174 -65
rect 141 -90 149 -73
rect 166 -90 174 -73
rect 141 -98 174 -90
rect 351 -73 384 -65
rect 351 -90 359 -73
rect 376 -90 384 -73
rect 351 -98 384 -90
rect 561 -73 594 -65
rect 561 -90 569 -73
rect 586 -90 594 -73
rect 561 -98 594 -90
rect 771 -73 804 -65
rect 771 -90 779 -73
rect 796 -90 804 -73
rect 771 -98 804 -90
rect 981 -73 1014 -65
rect 981 -90 989 -73
rect 1006 -90 1014 -73
rect 981 -98 1014 -90
rect 1191 -73 1224 -65
rect 1191 -90 1199 -73
rect 1216 -90 1224 -73
rect 1191 -98 1224 -90
rect 1401 -73 1434 -65
rect 1401 -90 1409 -73
rect 1426 -90 1434 -73
rect 1401 -98 1434 -90
rect 1611 -73 1644 -65
rect 1611 -90 1619 -73
rect 1636 -90 1644 -73
rect 1611 -98 1644 -90
rect 1821 -73 1854 -65
rect 1821 -90 1829 -73
rect 1846 -90 1854 -73
rect 1821 -98 1854 -90
rect 2031 -73 2064 -65
rect 2031 -90 2039 -73
rect 2056 -90 2064 -73
rect 2031 -98 2064 -90
rect -2063 -175 -2030 -167
rect -2063 -192 -2055 -175
rect -2038 -192 -2030 -175
rect -2063 -200 -2030 -192
rect -1853 -175 -1820 -167
rect -1853 -192 -1845 -175
rect -1828 -192 -1820 -175
rect -1853 -200 -1820 -192
rect -1643 -175 -1610 -167
rect -1643 -192 -1635 -175
rect -1618 -192 -1610 -175
rect -1643 -200 -1610 -192
rect -1433 -175 -1400 -167
rect -1433 -192 -1425 -175
rect -1408 -192 -1400 -175
rect -1433 -200 -1400 -192
rect -1223 -175 -1190 -167
rect -1223 -192 -1215 -175
rect -1198 -192 -1190 -175
rect -1223 -200 -1190 -192
rect -1013 -175 -980 -167
rect -1013 -192 -1005 -175
rect -988 -192 -980 -175
rect -1013 -200 -980 -192
rect -803 -175 -770 -167
rect -803 -192 -795 -175
rect -778 -192 -770 -175
rect -803 -200 -770 -192
rect -593 -175 -560 -167
rect -593 -192 -585 -175
rect -568 -192 -560 -175
rect -593 -200 -560 -192
rect -383 -175 -350 -167
rect -383 -192 -375 -175
rect -358 -192 -350 -175
rect -383 -200 -350 -192
rect -173 -175 -140 -167
rect -173 -192 -165 -175
rect -148 -192 -140 -175
rect -173 -200 -140 -192
rect 37 -175 70 -167
rect 37 -192 45 -175
rect 62 -192 70 -175
rect 37 -200 70 -192
rect 247 -175 280 -167
rect 247 -192 255 -175
rect 272 -192 280 -175
rect 247 -200 280 -192
rect 457 -175 490 -167
rect 457 -192 465 -175
rect 482 -192 490 -175
rect 457 -200 490 -192
rect 667 -175 700 -167
rect 667 -192 675 -175
rect 692 -192 700 -175
rect 667 -200 700 -192
rect 877 -175 910 -167
rect 877 -192 885 -175
rect 902 -192 910 -175
rect 877 -200 910 -192
rect 1087 -175 1120 -167
rect 1087 -192 1095 -175
rect 1112 -192 1120 -175
rect 1087 -200 1120 -192
rect 1297 -175 1330 -167
rect 1297 -192 1305 -175
rect 1322 -192 1330 -175
rect 1297 -200 1330 -192
rect 1507 -175 1540 -167
rect 1507 -192 1515 -175
rect 1532 -192 1540 -175
rect 1507 -200 1540 -192
rect 1717 -175 1750 -167
rect 1717 -192 1725 -175
rect 1742 -192 1750 -175
rect 1717 -200 1750 -192
rect 1927 -175 1960 -167
rect 1927 -192 1935 -175
rect 1952 -192 1960 -175
rect 1927 -200 1960 -192
rect 2137 -175 2170 -167
rect 2137 -192 2145 -175
rect 2162 -192 2170 -175
rect 2137 -200 2170 -192
rect -2159 -216 -2144 -203
rect -2054 -216 -2039 -200
rect -1949 -216 -1934 -203
rect -1844 -216 -1829 -200
rect -1739 -216 -1724 -203
rect -1634 -216 -1619 -200
rect -1529 -216 -1514 -203
rect -1424 -216 -1409 -200
rect -1319 -216 -1304 -203
rect -1214 -216 -1199 -200
rect -1109 -216 -1094 -203
rect -1004 -216 -989 -200
rect -899 -216 -884 -203
rect -794 -216 -779 -200
rect -689 -216 -674 -203
rect -584 -216 -569 -200
rect -479 -216 -464 -203
rect -374 -216 -359 -200
rect -269 -216 -254 -203
rect -164 -216 -149 -200
rect -59 -216 -44 -203
rect 46 -216 61 -200
rect 151 -216 166 -203
rect 256 -216 271 -200
rect 361 -216 376 -203
rect 466 -216 481 -200
rect 571 -216 586 -203
rect 676 -216 691 -200
rect 781 -216 796 -203
rect 886 -216 901 -200
rect 991 -216 1006 -203
rect 1096 -216 1111 -200
rect 1201 -216 1216 -203
rect 1306 -216 1321 -200
rect 1411 -216 1426 -203
rect 1516 -216 1531 -200
rect 1621 -216 1636 -203
rect 1726 -216 1741 -200
rect 1831 -216 1846 -203
rect 1936 -216 1951 -200
rect 2041 -216 2056 -203
rect 2146 -216 2161 -200
rect -2159 -331 -2144 -316
rect -2054 -329 -2039 -316
rect -1949 -331 -1934 -316
rect -1844 -329 -1829 -316
rect -1739 -331 -1724 -316
rect -1634 -329 -1619 -316
rect -1529 -331 -1514 -316
rect -1424 -329 -1409 -316
rect -1319 -331 -1304 -316
rect -1214 -329 -1199 -316
rect -1109 -331 -1094 -316
rect -1004 -329 -989 -316
rect -899 -331 -884 -316
rect -794 -329 -779 -316
rect -689 -331 -674 -316
rect -584 -329 -569 -316
rect -479 -331 -464 -316
rect -374 -329 -359 -316
rect -269 -331 -254 -316
rect -164 -329 -149 -316
rect -59 -331 -44 -316
rect 46 -329 61 -316
rect 151 -331 166 -316
rect 256 -329 271 -316
rect 361 -331 376 -316
rect 466 -329 481 -316
rect 571 -331 586 -316
rect 676 -329 691 -316
rect 781 -331 796 -316
rect 886 -329 901 -316
rect 991 -331 1006 -316
rect 1096 -329 1111 -316
rect 1201 -331 1216 -316
rect 1306 -329 1321 -316
rect 1411 -331 1426 -316
rect 1516 -329 1531 -316
rect 1621 -331 1636 -316
rect 1726 -329 1741 -316
rect 1831 -331 1846 -316
rect 1936 -329 1951 -316
rect 2041 -331 2056 -316
rect 2146 -329 2161 -316
rect -2168 -339 -2135 -331
rect -2168 -356 -2160 -339
rect -2143 -356 -2135 -339
rect -2168 -364 -2135 -356
rect -1958 -339 -1925 -331
rect -1958 -356 -1950 -339
rect -1933 -356 -1925 -339
rect -1958 -364 -1925 -356
rect -1748 -339 -1715 -331
rect -1748 -356 -1740 -339
rect -1723 -356 -1715 -339
rect -1748 -364 -1715 -356
rect -1538 -339 -1505 -331
rect -1538 -356 -1530 -339
rect -1513 -356 -1505 -339
rect -1538 -364 -1505 -356
rect -1328 -339 -1295 -331
rect -1328 -356 -1320 -339
rect -1303 -356 -1295 -339
rect -1328 -364 -1295 -356
rect -1118 -339 -1085 -331
rect -1118 -356 -1110 -339
rect -1093 -356 -1085 -339
rect -1118 -364 -1085 -356
rect -908 -339 -875 -331
rect -908 -356 -900 -339
rect -883 -356 -875 -339
rect -908 -364 -875 -356
rect -698 -339 -665 -331
rect -698 -356 -690 -339
rect -673 -356 -665 -339
rect -698 -364 -665 -356
rect -488 -339 -455 -331
rect -488 -356 -480 -339
rect -463 -356 -455 -339
rect -488 -364 -455 -356
rect -278 -339 -245 -331
rect -278 -356 -270 -339
rect -253 -356 -245 -339
rect -278 -364 -245 -356
rect -68 -339 -35 -331
rect -68 -356 -60 -339
rect -43 -356 -35 -339
rect -68 -364 -35 -356
rect 142 -339 175 -331
rect 142 -356 150 -339
rect 167 -356 175 -339
rect 142 -364 175 -356
rect 352 -339 385 -331
rect 352 -356 360 -339
rect 377 -356 385 -339
rect 352 -364 385 -356
rect 562 -339 595 -331
rect 562 -356 570 -339
rect 587 -356 595 -339
rect 562 -364 595 -356
rect 772 -339 805 -331
rect 772 -356 780 -339
rect 797 -356 805 -339
rect 772 -364 805 -356
rect 982 -339 1015 -331
rect 982 -356 990 -339
rect 1007 -356 1015 -339
rect 982 -364 1015 -356
rect 1192 -339 1225 -331
rect 1192 -356 1200 -339
rect 1217 -356 1225 -339
rect 1192 -364 1225 -356
rect 1402 -339 1435 -331
rect 1402 -356 1410 -339
rect 1427 -356 1435 -339
rect 1402 -364 1435 -356
rect 1612 -339 1645 -331
rect 1612 -356 1620 -339
rect 1637 -356 1645 -339
rect 1612 -364 1645 -356
rect 1822 -339 1855 -331
rect 1822 -356 1830 -339
rect 1847 -356 1855 -339
rect 1822 -364 1855 -356
rect 2032 -339 2065 -331
rect 2032 -356 2040 -339
rect 2057 -356 2065 -339
rect 2032 -364 2065 -356
<< polycont >>
rect -2056 73 -2039 90
rect -1846 73 -1829 90
rect -1636 73 -1619 90
rect -1426 73 -1409 90
rect -1216 73 -1199 90
rect -1006 73 -989 90
rect -796 73 -779 90
rect -586 73 -569 90
rect -376 73 -359 90
rect -166 73 -149 90
rect 44 73 61 90
rect 254 73 271 90
rect 464 73 481 90
rect 674 73 691 90
rect 884 73 901 90
rect 1094 73 1111 90
rect 1304 73 1321 90
rect 1514 73 1531 90
rect 1724 73 1741 90
rect 1934 73 1951 90
rect 2144 73 2161 90
rect -2161 -90 -2144 -73
rect -1951 -90 -1934 -73
rect -1741 -90 -1724 -73
rect -1531 -90 -1514 -73
rect -1321 -90 -1304 -73
rect -1111 -90 -1094 -73
rect -901 -90 -884 -73
rect -691 -90 -674 -73
rect -481 -90 -464 -73
rect -271 -90 -254 -73
rect -61 -90 -44 -73
rect 149 -90 166 -73
rect 359 -90 376 -73
rect 569 -90 586 -73
rect 779 -90 796 -73
rect 989 -90 1006 -73
rect 1199 -90 1216 -73
rect 1409 -90 1426 -73
rect 1619 -90 1636 -73
rect 1829 -90 1846 -73
rect 2039 -90 2056 -73
rect -2055 -192 -2038 -175
rect -1845 -192 -1828 -175
rect -1635 -192 -1618 -175
rect -1425 -192 -1408 -175
rect -1215 -192 -1198 -175
rect -1005 -192 -988 -175
rect -795 -192 -778 -175
rect -585 -192 -568 -175
rect -375 -192 -358 -175
rect -165 -192 -148 -175
rect 45 -192 62 -175
rect 255 -192 272 -175
rect 465 -192 482 -175
rect 675 -192 692 -175
rect 885 -192 902 -175
rect 1095 -192 1112 -175
rect 1305 -192 1322 -175
rect 1515 -192 1532 -175
rect 1725 -192 1742 -175
rect 1935 -192 1952 -175
rect 2145 -192 2162 -175
rect -2160 -356 -2143 -339
rect -1950 -356 -1933 -339
rect -1740 -356 -1723 -339
rect -1530 -356 -1513 -339
rect -1320 -356 -1303 -339
rect -1110 -356 -1093 -339
rect -900 -356 -883 -339
rect -690 -356 -673 -339
rect -480 -356 -463 -339
rect -270 -356 -253 -339
rect -60 -356 -43 -339
rect 150 -356 167 -339
rect 360 -356 377 -339
rect 570 -356 587 -339
rect 780 -356 797 -339
rect 990 -356 1007 -339
rect 1200 -356 1217 -339
rect 1410 -356 1427 -339
rect 1620 -356 1637 -339
rect 1830 -356 1847 -339
rect 2040 -356 2057 -339
<< locali >>
rect -2242 124 -2194 141
rect 2194 124 2242 141
rect -2242 93 -2225 124
rect 2225 93 2242 124
rect -2064 73 -2056 90
rect -2039 73 -2031 90
rect -1854 73 -1846 90
rect -1829 73 -1821 90
rect -1644 73 -1636 90
rect -1619 73 -1611 90
rect -1434 73 -1426 90
rect -1409 73 -1401 90
rect -1224 73 -1216 90
rect -1199 73 -1191 90
rect -1014 73 -1006 90
rect -989 73 -981 90
rect -804 73 -796 90
rect -779 73 -771 90
rect -594 73 -586 90
rect -569 73 -561 90
rect -384 73 -376 90
rect -359 73 -351 90
rect -174 73 -166 90
rect -149 73 -141 90
rect 36 73 44 90
rect 61 73 69 90
rect 246 73 254 90
rect 271 73 279 90
rect 456 73 464 90
rect 481 73 489 90
rect 666 73 674 90
rect 691 73 699 90
rect 876 73 884 90
rect 901 73 909 90
rect 1086 73 1094 90
rect 1111 73 1119 90
rect 1296 73 1304 90
rect 1321 73 1329 90
rect 1506 73 1514 90
rect 1531 73 1539 90
rect 1716 73 1724 90
rect 1741 73 1749 90
rect 1926 73 1934 90
rect 1951 73 1959 90
rect 2120 73 2144 90
rect 2161 73 2225 90
rect -2185 44 -2168 52
rect -2185 -73 -2168 -44
rect -2137 44 -2120 52
rect -2137 -73 -2120 -44
rect -2080 44 -2063 52
rect -2080 -52 -2063 -44
rect -2032 44 -2015 52
rect -2032 -52 -2015 -44
rect -1975 44 -1958 52
rect -1975 -52 -1958 -44
rect -1927 44 -1910 52
rect -1927 -52 -1910 -44
rect -1870 44 -1853 52
rect -1870 -52 -1853 -44
rect -1822 44 -1805 52
rect -1822 -52 -1805 -44
rect -1765 44 -1748 52
rect -1765 -52 -1748 -44
rect -1717 44 -1700 52
rect -1717 -52 -1700 -44
rect -1660 44 -1643 52
rect -1660 -52 -1643 -44
rect -1612 44 -1595 52
rect -1612 -52 -1595 -44
rect -1555 44 -1538 52
rect -1555 -52 -1538 -44
rect -1507 44 -1490 52
rect -1507 -52 -1490 -44
rect -1450 44 -1433 52
rect -1450 -52 -1433 -44
rect -1402 44 -1385 52
rect -1402 -52 -1385 -44
rect -1345 44 -1328 52
rect -1345 -52 -1328 -44
rect -1297 44 -1280 52
rect -1297 -52 -1280 -44
rect -1240 44 -1223 52
rect -1240 -52 -1223 -44
rect -1192 44 -1175 52
rect -1192 -52 -1175 -44
rect -1135 44 -1118 52
rect -1135 -52 -1118 -44
rect -1087 44 -1070 52
rect -1087 -52 -1070 -44
rect -1030 44 -1013 52
rect -1030 -52 -1013 -44
rect -982 44 -965 52
rect -982 -52 -965 -44
rect -925 44 -908 52
rect -925 -52 -908 -44
rect -877 44 -860 52
rect -877 -52 -860 -44
rect -820 44 -803 52
rect -820 -52 -803 -44
rect -772 44 -755 52
rect -772 -52 -755 -44
rect -715 44 -698 52
rect -715 -52 -698 -44
rect -667 44 -650 52
rect -667 -52 -650 -44
rect -610 44 -593 52
rect -610 -52 -593 -44
rect -562 44 -545 52
rect -562 -52 -545 -44
rect -505 44 -488 52
rect -505 -52 -488 -44
rect -457 44 -440 52
rect -457 -52 -440 -44
rect -400 44 -383 52
rect -400 -52 -383 -44
rect -352 44 -335 52
rect -352 -52 -335 -44
rect -295 44 -278 52
rect -295 -52 -278 -44
rect -247 44 -230 52
rect -247 -52 -230 -44
rect -190 44 -173 52
rect -190 -52 -173 -44
rect -142 44 -125 52
rect -142 -52 -125 -44
rect -85 44 -68 52
rect -85 -52 -68 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 68 44 85 52
rect 68 -52 85 -44
rect 125 44 142 52
rect 125 -52 142 -44
rect 173 44 190 52
rect 173 -52 190 -44
rect 230 44 247 52
rect 230 -52 247 -44
rect 278 44 295 52
rect 278 -52 295 -44
rect 335 44 352 52
rect 335 -52 352 -44
rect 383 44 400 52
rect 383 -52 400 -44
rect 440 44 457 52
rect 440 -52 457 -44
rect 488 44 505 52
rect 488 -52 505 -44
rect 545 44 562 52
rect 545 -52 562 -44
rect 593 44 610 52
rect 593 -52 610 -44
rect 650 44 667 52
rect 650 -52 667 -44
rect 698 44 715 52
rect 698 -52 715 -44
rect 755 44 772 52
rect 755 -52 772 -44
rect 803 44 820 52
rect 803 -52 820 -44
rect 860 44 877 52
rect 860 -52 877 -44
rect 908 44 925 52
rect 908 -52 925 -44
rect 965 44 982 52
rect 965 -52 982 -44
rect 1013 44 1030 52
rect 1013 -52 1030 -44
rect 1070 44 1087 52
rect 1070 -52 1087 -44
rect 1118 44 1135 52
rect 1118 -52 1135 -44
rect 1175 44 1192 52
rect 1175 -52 1192 -44
rect 1223 44 1240 52
rect 1223 -52 1240 -44
rect 1280 44 1297 52
rect 1280 -52 1297 -44
rect 1328 44 1345 52
rect 1328 -52 1345 -44
rect 1385 44 1402 52
rect 1385 -52 1402 -44
rect 1433 44 1450 52
rect 1433 -52 1450 -44
rect 1490 44 1507 52
rect 1490 -52 1507 -44
rect 1538 44 1555 52
rect 1538 -52 1555 -44
rect 1595 44 1612 52
rect 1595 -52 1612 -44
rect 1643 44 1660 52
rect 1643 -52 1660 -44
rect 1700 44 1717 52
rect 1700 -52 1717 -44
rect 1748 44 1765 52
rect 1748 -52 1765 -44
rect 1805 44 1822 52
rect 1805 -52 1822 -44
rect 1853 44 1870 52
rect 1853 -52 1870 -44
rect 1910 44 1927 52
rect 1910 -52 1927 -44
rect 1958 44 1975 52
rect 1958 -52 1975 -44
rect 2015 44 2032 52
rect 2015 -52 2032 -44
rect 2063 44 2080 52
rect 2063 -52 2080 -44
rect 2120 44 2137 73
rect 2120 -52 2137 -44
rect 2168 44 2185 73
rect 2168 -52 2185 -44
rect -2225 -90 -2161 -73
rect -2144 -90 -2120 -73
rect -1959 -90 -1951 -73
rect -1934 -90 -1926 -73
rect -1749 -90 -1741 -73
rect -1724 -90 -1716 -73
rect -1539 -90 -1531 -73
rect -1514 -90 -1506 -73
rect -1329 -90 -1321 -73
rect -1304 -90 -1296 -73
rect -1119 -90 -1111 -73
rect -1094 -90 -1086 -73
rect -909 -90 -901 -73
rect -884 -90 -876 -73
rect -699 -90 -691 -73
rect -674 -90 -666 -73
rect -489 -90 -481 -73
rect -464 -90 -456 -73
rect -279 -90 -271 -73
rect -254 -90 -246 -73
rect -69 -90 -61 -73
rect -44 -90 -36 -73
rect 141 -90 149 -73
rect 166 -90 174 -73
rect 351 -90 359 -73
rect 376 -90 384 -73
rect 561 -90 569 -73
rect 586 -90 594 -73
rect 771 -90 779 -73
rect 796 -90 804 -73
rect 981 -90 989 -73
rect 1006 -90 1014 -73
rect 1191 -90 1199 -73
rect 1216 -90 1224 -73
rect 1401 -90 1409 -73
rect 1426 -90 1434 -73
rect 1611 -90 1619 -73
rect 1636 -90 1644 -73
rect 1821 -90 1829 -73
rect 1846 -90 1854 -73
rect 2031 -90 2039 -73
rect 2056 -90 2064 -73
rect -2242 -172 -2225 -93
rect 2225 -172 2242 -93
rect -2063 -192 -2055 -175
rect -2038 -192 -2030 -175
rect -1853 -192 -1845 -175
rect -1828 -192 -1820 -175
rect -1643 -192 -1635 -175
rect -1618 -192 -1610 -175
rect -1433 -192 -1425 -175
rect -1408 -192 -1400 -175
rect -1223 -192 -1215 -175
rect -1198 -192 -1190 -175
rect -1013 -192 -1005 -175
rect -988 -192 -980 -175
rect -803 -192 -795 -175
rect -778 -192 -770 -175
rect -593 -192 -585 -175
rect -568 -192 -560 -175
rect -383 -192 -375 -175
rect -358 -192 -350 -175
rect -173 -192 -165 -175
rect -148 -192 -140 -175
rect 37 -192 45 -175
rect 62 -192 70 -175
rect 247 -192 255 -175
rect 272 -192 280 -175
rect 457 -192 465 -175
rect 482 -192 490 -175
rect 667 -192 675 -175
rect 692 -192 700 -175
rect 877 -192 885 -175
rect 902 -192 910 -175
rect 1087 -192 1095 -175
rect 1112 -192 1120 -175
rect 1297 -192 1305 -175
rect 1322 -192 1330 -175
rect 1507 -192 1515 -175
rect 1532 -192 1540 -175
rect 1717 -192 1725 -175
rect 1742 -192 1750 -175
rect 1927 -192 1935 -175
rect 1952 -192 1960 -175
rect 2121 -192 2145 -175
rect 2162 -192 2225 -175
rect -2184 -222 -2167 -214
rect -2184 -339 -2167 -310
rect -2136 -222 -2119 -214
rect -2136 -339 -2119 -310
rect -2079 -222 -2062 -214
rect -2079 -318 -2062 -310
rect -2031 -222 -2014 -214
rect -2031 -318 -2014 -310
rect -1974 -222 -1957 -214
rect -1974 -318 -1957 -310
rect -1926 -222 -1909 -214
rect -1926 -318 -1909 -310
rect -1869 -222 -1852 -214
rect -1869 -318 -1852 -310
rect -1821 -222 -1804 -214
rect -1821 -318 -1804 -310
rect -1764 -222 -1747 -214
rect -1764 -318 -1747 -310
rect -1716 -222 -1699 -214
rect -1716 -318 -1699 -310
rect -1659 -222 -1642 -214
rect -1659 -318 -1642 -310
rect -1611 -222 -1594 -214
rect -1611 -318 -1594 -310
rect -1554 -222 -1537 -214
rect -1554 -318 -1537 -310
rect -1506 -222 -1489 -214
rect -1506 -318 -1489 -310
rect -1449 -222 -1432 -214
rect -1449 -318 -1432 -310
rect -1401 -222 -1384 -214
rect -1401 -318 -1384 -310
rect -1344 -222 -1327 -214
rect -1344 -318 -1327 -310
rect -1296 -222 -1279 -214
rect -1296 -318 -1279 -310
rect -1239 -222 -1222 -214
rect -1239 -318 -1222 -310
rect -1191 -222 -1174 -214
rect -1191 -318 -1174 -310
rect -1134 -222 -1117 -214
rect -1134 -318 -1117 -310
rect -1086 -222 -1069 -214
rect -1086 -318 -1069 -310
rect -1029 -222 -1012 -214
rect -1029 -318 -1012 -310
rect -981 -222 -964 -214
rect -981 -318 -964 -310
rect -924 -222 -907 -214
rect -924 -318 -907 -310
rect -876 -222 -859 -214
rect -876 -318 -859 -310
rect -819 -222 -802 -214
rect -819 -318 -802 -310
rect -771 -222 -754 -214
rect -771 -318 -754 -310
rect -714 -222 -697 -214
rect -714 -318 -697 -310
rect -666 -222 -649 -214
rect -666 -318 -649 -310
rect -609 -222 -592 -214
rect -609 -318 -592 -310
rect -561 -222 -544 -214
rect -561 -318 -544 -310
rect -504 -222 -487 -214
rect -504 -318 -487 -310
rect -456 -222 -439 -214
rect -456 -318 -439 -310
rect -399 -222 -382 -214
rect -399 -318 -382 -310
rect -351 -222 -334 -214
rect -351 -318 -334 -310
rect -294 -222 -277 -214
rect -294 -318 -277 -310
rect -246 -222 -229 -214
rect -246 -318 -229 -310
rect -189 -222 -172 -214
rect -189 -318 -172 -310
rect -141 -222 -124 -214
rect -141 -318 -124 -310
rect -84 -222 -67 -214
rect -84 -318 -67 -310
rect -36 -222 -19 -214
rect -36 -318 -19 -310
rect 21 -222 38 -214
rect 21 -318 38 -310
rect 69 -222 86 -214
rect 69 -318 86 -310
rect 126 -222 143 -214
rect 126 -318 143 -310
rect 174 -222 191 -214
rect 174 -318 191 -310
rect 231 -222 248 -214
rect 231 -318 248 -310
rect 279 -222 296 -214
rect 279 -318 296 -310
rect 336 -222 353 -214
rect 336 -318 353 -310
rect 384 -222 401 -214
rect 384 -318 401 -310
rect 441 -222 458 -214
rect 441 -318 458 -310
rect 489 -222 506 -214
rect 489 -318 506 -310
rect 546 -222 563 -214
rect 546 -318 563 -310
rect 594 -222 611 -214
rect 594 -318 611 -310
rect 651 -222 668 -214
rect 651 -318 668 -310
rect 699 -222 716 -214
rect 699 -318 716 -310
rect 756 -222 773 -214
rect 756 -318 773 -310
rect 804 -222 821 -214
rect 804 -318 821 -310
rect 861 -222 878 -214
rect 861 -318 878 -310
rect 909 -222 926 -214
rect 909 -318 926 -310
rect 966 -222 983 -214
rect 966 -318 983 -310
rect 1014 -222 1031 -214
rect 1014 -318 1031 -310
rect 1071 -222 1088 -214
rect 1071 -318 1088 -310
rect 1119 -222 1136 -214
rect 1119 -318 1136 -310
rect 1176 -222 1193 -214
rect 1176 -318 1193 -310
rect 1224 -222 1241 -214
rect 1224 -318 1241 -310
rect 1281 -222 1298 -214
rect 1281 -318 1298 -310
rect 1329 -222 1346 -214
rect 1329 -318 1346 -310
rect 1386 -222 1403 -214
rect 1386 -318 1403 -310
rect 1434 -222 1451 -214
rect 1434 -318 1451 -310
rect 1491 -222 1508 -214
rect 1491 -318 1508 -310
rect 1539 -222 1556 -214
rect 1539 -318 1556 -310
rect 1596 -222 1613 -214
rect 1596 -318 1613 -310
rect 1644 -222 1661 -214
rect 1644 -318 1661 -310
rect 1701 -222 1718 -214
rect 1701 -318 1718 -310
rect 1749 -222 1766 -214
rect 1749 -318 1766 -310
rect 1806 -222 1823 -214
rect 1806 -318 1823 -310
rect 1854 -222 1871 -214
rect 1854 -318 1871 -310
rect 1911 -222 1928 -214
rect 1911 -318 1928 -310
rect 1959 -222 1976 -214
rect 1959 -318 1976 -310
rect 2016 -222 2033 -214
rect 2016 -318 2033 -310
rect 2064 -222 2081 -214
rect 2064 -318 2081 -310
rect 2121 -222 2138 -192
rect 2121 -318 2138 -310
rect 2169 -222 2186 -192
rect 2169 -318 2186 -310
rect -2225 -356 -2160 -339
rect -2143 -356 -2119 -339
rect -1958 -356 -1950 -339
rect -1933 -356 -1925 -339
rect -1748 -356 -1740 -339
rect -1723 -356 -1715 -339
rect -1538 -356 -1530 -339
rect -1513 -356 -1505 -339
rect -1328 -356 -1320 -339
rect -1303 -356 -1295 -339
rect -1118 -356 -1110 -339
rect -1093 -356 -1085 -339
rect -908 -356 -900 -339
rect -883 -356 -875 -339
rect -698 -356 -690 -339
rect -673 -356 -665 -339
rect -488 -356 -480 -339
rect -463 -356 -455 -339
rect -278 -356 -270 -339
rect -253 -356 -245 -339
rect -68 -356 -60 -339
rect -43 -356 -35 -339
rect 142 -356 150 -339
rect 167 -356 175 -339
rect 352 -356 360 -339
rect 377 -356 385 -339
rect 562 -356 570 -339
rect 587 -356 595 -339
rect 772 -356 780 -339
rect 797 -356 805 -339
rect 982 -356 990 -339
rect 1007 -356 1015 -339
rect 1192 -356 1200 -339
rect 1217 -356 1225 -339
rect 1402 -356 1410 -339
rect 1427 -356 1435 -339
rect 1612 -356 1620 -339
rect 1637 -356 1645 -339
rect 1822 -356 1830 -339
rect 1847 -356 1855 -339
rect 2032 -356 2040 -339
rect 2057 -356 2065 -339
rect -2242 -390 -2225 -359
rect 2225 -390 2242 -359
rect -2242 -407 -2194 -390
rect 2194 -407 2242 -390
<< viali >>
rect -2056 73 -2039 90
rect -1846 73 -1829 90
rect -1636 73 -1619 90
rect -1426 73 -1409 90
rect -1216 73 -1199 90
rect -1006 73 -989 90
rect -796 73 -779 90
rect -586 73 -569 90
rect -376 73 -359 90
rect -166 73 -149 90
rect 44 73 61 90
rect 254 73 271 90
rect 464 73 481 90
rect 674 73 691 90
rect 884 73 901 90
rect 1094 73 1111 90
rect 1304 73 1321 90
rect 1514 73 1531 90
rect 1724 73 1741 90
rect 1934 73 1951 90
rect -1951 -90 -1934 -73
rect -1741 -90 -1724 -73
rect -1531 -90 -1514 -73
rect -1321 -90 -1304 -73
rect -1111 -90 -1094 -73
rect -901 -90 -884 -73
rect -691 -90 -674 -73
rect -481 -90 -464 -73
rect -271 -90 -254 -73
rect -61 -90 -44 -73
rect 149 -90 166 -73
rect 359 -90 376 -73
rect 569 -90 586 -73
rect 779 -90 796 -73
rect 989 -90 1006 -73
rect 1199 -90 1216 -73
rect 1409 -90 1426 -73
rect 1619 -90 1636 -73
rect 1829 -90 1846 -73
rect 2039 -90 2056 -73
rect -2055 -192 -2038 -175
rect -1845 -192 -1828 -175
rect -1635 -192 -1618 -175
rect -1425 -192 -1408 -175
rect -1215 -192 -1198 -175
rect -1005 -192 -988 -175
rect -795 -192 -778 -175
rect -585 -192 -568 -175
rect -375 -192 -358 -175
rect -165 -192 -148 -175
rect 45 -192 62 -175
rect 255 -192 272 -175
rect 465 -192 482 -175
rect 675 -192 692 -175
rect 885 -192 902 -175
rect 1095 -192 1112 -175
rect 1305 -192 1322 -175
rect 1515 -192 1532 -175
rect 1725 -192 1742 -175
rect 1935 -192 1952 -175
rect -1950 -356 -1933 -339
rect -1740 -356 -1723 -339
rect -1530 -356 -1513 -339
rect -1320 -356 -1303 -339
rect -1110 -356 -1093 -339
rect -900 -356 -883 -339
rect -690 -356 -673 -339
rect -480 -356 -463 -339
rect -270 -356 -253 -339
rect -60 -356 -43 -339
rect 150 -356 167 -339
rect 360 -356 377 -339
rect 570 -356 587 -339
rect 780 -356 797 -339
rect 990 -356 1007 -339
rect 1200 -356 1217 -339
rect 1410 -356 1427 -339
rect 1620 -356 1637 -339
rect 1830 -356 1847 -339
rect 2040 -356 2057 -339
<< metal1 >>
rect -2062 90 -2033 93
rect -2062 73 -2056 90
rect -2039 73 -2033 90
rect -2062 70 -2033 73
rect -1852 90 -1823 93
rect -1852 73 -1846 90
rect -1829 73 -1823 90
rect -1852 70 -1823 73
rect -1642 90 -1613 93
rect -1642 73 -1636 90
rect -1619 73 -1613 90
rect -1642 70 -1613 73
rect -1432 90 -1403 93
rect -1432 73 -1426 90
rect -1409 73 -1403 90
rect -1432 70 -1403 73
rect -1222 90 -1193 93
rect -1222 73 -1216 90
rect -1199 73 -1193 90
rect -1222 70 -1193 73
rect -1012 90 -983 93
rect -1012 73 -1006 90
rect -989 73 -983 90
rect -1012 70 -983 73
rect -802 90 -773 93
rect -802 73 -796 90
rect -779 73 -773 90
rect -802 70 -773 73
rect -592 90 -563 93
rect -592 73 -586 90
rect -569 73 -563 90
rect -592 70 -563 73
rect -382 90 -353 93
rect -382 73 -376 90
rect -359 73 -353 90
rect -382 70 -353 73
rect -172 90 -143 93
rect -172 73 -166 90
rect -149 73 -143 90
rect -172 70 -143 73
rect 38 90 67 93
rect 38 73 44 90
rect 61 73 67 90
rect 38 70 67 73
rect 248 90 277 93
rect 248 73 254 90
rect 271 73 277 90
rect 248 70 277 73
rect 458 90 487 93
rect 458 73 464 90
rect 481 73 487 90
rect 458 70 487 73
rect 668 90 697 93
rect 668 73 674 90
rect 691 73 697 90
rect 668 70 697 73
rect 878 90 907 93
rect 878 73 884 90
rect 901 73 907 90
rect 878 70 907 73
rect 1088 90 1117 93
rect 1088 73 1094 90
rect 1111 73 1117 90
rect 1088 70 1117 73
rect 1298 90 1327 93
rect 1298 73 1304 90
rect 1321 73 1327 90
rect 1298 70 1327 73
rect 1508 90 1537 93
rect 1508 73 1514 90
rect 1531 73 1537 90
rect 1508 70 1537 73
rect 1718 90 1747 93
rect 1718 73 1724 90
rect 1741 73 1747 90
rect 1718 70 1747 73
rect 1928 90 1957 93
rect 1928 73 1934 90
rect 1951 73 1957 90
rect 1928 70 1957 73
rect -1957 -73 -1928 -70
rect -1957 -90 -1951 -73
rect -1934 -90 -1928 -73
rect -1957 -93 -1928 -90
rect -1747 -73 -1718 -70
rect -1747 -90 -1741 -73
rect -1724 -90 -1718 -73
rect -1747 -93 -1718 -90
rect -1537 -73 -1508 -70
rect -1537 -90 -1531 -73
rect -1514 -90 -1508 -73
rect -1537 -93 -1508 -90
rect -1327 -73 -1298 -70
rect -1327 -90 -1321 -73
rect -1304 -90 -1298 -73
rect -1327 -93 -1298 -90
rect -1117 -73 -1088 -70
rect -1117 -90 -1111 -73
rect -1094 -90 -1088 -73
rect -1117 -93 -1088 -90
rect -907 -73 -878 -70
rect -907 -90 -901 -73
rect -884 -90 -878 -73
rect -907 -93 -878 -90
rect -697 -73 -668 -70
rect -697 -90 -691 -73
rect -674 -90 -668 -73
rect -697 -93 -668 -90
rect -487 -73 -458 -70
rect -487 -90 -481 -73
rect -464 -90 -458 -73
rect -487 -93 -458 -90
rect -277 -73 -248 -70
rect -277 -90 -271 -73
rect -254 -90 -248 -73
rect -277 -93 -248 -90
rect -67 -73 -38 -70
rect -67 -90 -61 -73
rect -44 -90 -38 -73
rect -67 -93 -38 -90
rect 143 -73 172 -70
rect 143 -90 149 -73
rect 166 -90 172 -73
rect 143 -93 172 -90
rect 353 -73 382 -70
rect 353 -90 359 -73
rect 376 -90 382 -73
rect 353 -93 382 -90
rect 563 -73 592 -70
rect 563 -90 569 -73
rect 586 -90 592 -73
rect 563 -93 592 -90
rect 773 -73 802 -70
rect 773 -90 779 -73
rect 796 -90 802 -73
rect 773 -93 802 -90
rect 983 -73 1012 -70
rect 983 -90 989 -73
rect 1006 -90 1012 -73
rect 983 -93 1012 -90
rect 1193 -73 1222 -70
rect 1193 -90 1199 -73
rect 1216 -90 1222 -73
rect 1193 -93 1222 -90
rect 1403 -73 1432 -70
rect 1403 -90 1409 -73
rect 1426 -90 1432 -73
rect 1403 -93 1432 -90
rect 1613 -73 1642 -70
rect 1613 -90 1619 -73
rect 1636 -90 1642 -73
rect 1613 -93 1642 -90
rect 1823 -73 1852 -70
rect 1823 -90 1829 -73
rect 1846 -90 1852 -73
rect 1823 -93 1852 -90
rect 2033 -73 2062 -70
rect 2033 -90 2039 -73
rect 2056 -90 2062 -73
rect 2033 -93 2062 -90
rect -2061 -175 -2032 -172
rect -2061 -192 -2055 -175
rect -2038 -192 -2032 -175
rect -2061 -195 -2032 -192
rect -1851 -175 -1822 -172
rect -1851 -192 -1845 -175
rect -1828 -192 -1822 -175
rect -1851 -195 -1822 -192
rect -1641 -175 -1612 -172
rect -1641 -192 -1635 -175
rect -1618 -192 -1612 -175
rect -1641 -195 -1612 -192
rect -1431 -175 -1402 -172
rect -1431 -192 -1425 -175
rect -1408 -192 -1402 -175
rect -1431 -195 -1402 -192
rect -1221 -175 -1192 -172
rect -1221 -192 -1215 -175
rect -1198 -192 -1192 -175
rect -1221 -195 -1192 -192
rect -1011 -175 -982 -172
rect -1011 -192 -1005 -175
rect -988 -192 -982 -175
rect -1011 -195 -982 -192
rect -801 -175 -772 -172
rect -801 -192 -795 -175
rect -778 -192 -772 -175
rect -801 -195 -772 -192
rect -591 -175 -562 -172
rect -591 -192 -585 -175
rect -568 -192 -562 -175
rect -591 -195 -562 -192
rect -381 -175 -352 -172
rect -381 -192 -375 -175
rect -358 -192 -352 -175
rect -381 -195 -352 -192
rect -171 -175 -142 -172
rect -171 -192 -165 -175
rect -148 -192 -142 -175
rect -171 -195 -142 -192
rect 39 -175 68 -172
rect 39 -192 45 -175
rect 62 -192 68 -175
rect 39 -195 68 -192
rect 249 -175 278 -172
rect 249 -192 255 -175
rect 272 -192 278 -175
rect 249 -195 278 -192
rect 459 -175 488 -172
rect 459 -192 465 -175
rect 482 -192 488 -175
rect 459 -195 488 -192
rect 669 -175 698 -172
rect 669 -192 675 -175
rect 692 -192 698 -175
rect 669 -195 698 -192
rect 879 -175 908 -172
rect 879 -192 885 -175
rect 902 -192 908 -175
rect 879 -195 908 -192
rect 1089 -175 1118 -172
rect 1089 -192 1095 -175
rect 1112 -192 1118 -175
rect 1089 -195 1118 -192
rect 1299 -175 1328 -172
rect 1299 -192 1305 -175
rect 1322 -192 1328 -175
rect 1299 -195 1328 -192
rect 1509 -175 1538 -172
rect 1509 -192 1515 -175
rect 1532 -192 1538 -175
rect 1509 -195 1538 -192
rect 1719 -175 1748 -172
rect 1719 -192 1725 -175
rect 1742 -192 1748 -175
rect 1719 -195 1748 -192
rect 1929 -175 1958 -172
rect 1929 -192 1935 -175
rect 1952 -192 1958 -175
rect 1929 -195 1958 -192
rect -1956 -339 -1927 -336
rect -1956 -356 -1950 -339
rect -1933 -356 -1927 -339
rect -1956 -359 -1927 -356
rect -1746 -339 -1717 -336
rect -1746 -356 -1740 -339
rect -1723 -356 -1717 -339
rect -1746 -359 -1717 -356
rect -1536 -339 -1507 -336
rect -1536 -356 -1530 -339
rect -1513 -356 -1507 -339
rect -1536 -359 -1507 -356
rect -1326 -339 -1297 -336
rect -1326 -356 -1320 -339
rect -1303 -356 -1297 -339
rect -1326 -359 -1297 -356
rect -1116 -339 -1087 -336
rect -1116 -356 -1110 -339
rect -1093 -356 -1087 -339
rect -1116 -359 -1087 -356
rect -906 -339 -877 -336
rect -906 -356 -900 -339
rect -883 -356 -877 -339
rect -906 -359 -877 -356
rect -696 -339 -667 -336
rect -696 -356 -690 -339
rect -673 -356 -667 -339
rect -696 -359 -667 -356
rect -486 -339 -457 -336
rect -486 -356 -480 -339
rect -463 -356 -457 -339
rect -486 -359 -457 -356
rect -276 -339 -247 -336
rect -276 -356 -270 -339
rect -253 -356 -247 -339
rect -276 -359 -247 -356
rect -66 -339 -37 -336
rect -66 -356 -60 -339
rect -43 -356 -37 -339
rect -66 -359 -37 -356
rect 144 -339 173 -336
rect 144 -356 150 -339
rect 167 -356 173 -339
rect 144 -359 173 -356
rect 354 -339 383 -336
rect 354 -356 360 -339
rect 377 -356 383 -339
rect 354 -359 383 -356
rect 564 -339 593 -336
rect 564 -356 570 -339
rect 587 -356 593 -339
rect 564 -359 593 -356
rect 774 -339 803 -336
rect 774 -356 780 -339
rect 797 -356 803 -339
rect 774 -359 803 -356
rect 984 -339 1013 -336
rect 984 -356 990 -339
rect 1007 -356 1013 -339
rect 984 -359 1013 -356
rect 1194 -339 1223 -336
rect 1194 -356 1200 -339
rect 1217 -356 1223 -339
rect 1194 -359 1223 -356
rect 1404 -339 1433 -336
rect 1404 -356 1410 -339
rect 1427 -356 1433 -339
rect 1404 -359 1433 -356
rect 1614 -339 1643 -336
rect 1614 -356 1620 -339
rect 1637 -356 1643 -339
rect 1614 -359 1643 -356
rect 1824 -339 1853 -336
rect 1824 -356 1830 -339
rect 1847 -356 1853 -339
rect 1824 -359 1853 -356
rect 2034 -339 2063 -336
rect 2034 -356 2040 -339
rect 2057 -356 2063 -339
rect 2034 -359 2063 -356
<< properties >>
string FIXED_BBOX -2233 -133 2233 133
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 42 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
