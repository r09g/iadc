magic
tech sky130A
magscale 1 2
timestamp 1654637878
<< nwell >>
rect 10352 6149 11405 6374
rect 8209 5669 13518 6149
rect 10352 5317 11342 5669
rect 13038 5316 13518 5669
rect 10047 4608 12103 4916
rect 8566 4128 13162 4608
rect 8566 3866 9046 4128
rect 10047 3866 12103 4128
<< viali >>
rect 8436 6228 8470 6262
rect 8792 6228 8826 6262
rect 9148 6228 9182 6262
rect 9504 6228 9538 6262
rect 9860 6228 9894 6262
rect 10216 6228 10250 6262
rect 10572 6228 10606 6262
rect 11122 6228 11156 6262
rect 11478 6228 11512 6262
rect 11834 6228 11868 6262
rect 12190 6228 12224 6262
rect 12546 6228 12580 6262
rect 12902 6228 12936 6262
rect 13258 6228 13292 6262
rect 8614 6006 8648 6040
rect 8970 6006 9004 6040
rect 9326 6006 9360 6040
rect 9682 6006 9716 6040
rect 10038 6006 10072 6040
rect 10394 6006 10428 6040
rect 11300 6006 11334 6040
rect 11656 6006 11690 6040
rect 12012 6006 12046 6040
rect 12368 6006 12402 6040
rect 12724 6006 12758 6040
rect 13080 6006 13114 6040
rect 8436 5651 8470 5685
rect 8792 5651 8826 5685
rect 9148 5651 9182 5685
rect 9504 5651 9538 5685
rect 9860 5651 9894 5685
rect 10216 5651 10250 5685
rect 10572 5651 10606 5685
rect 11122 5650 11156 5684
rect 11478 5650 11512 5684
rect 11834 5650 11868 5684
rect 12190 5650 12224 5684
rect 12546 5650 12580 5684
rect 12902 5650 12936 5684
rect 13258 5650 13292 5684
rect 8614 5429 8648 5463
rect 8970 5429 9004 5463
rect 9326 5429 9360 5463
rect 9682 5429 9716 5463
rect 10038 5429 10072 5463
rect 10394 5429 10428 5463
rect 11300 5428 11334 5462
rect 11656 5428 11690 5462
rect 12012 5428 12046 5462
rect 12368 5428 12402 5462
rect 12724 5428 12758 5462
rect 13080 5428 13114 5462
rect 8792 4770 8826 4804
rect 9148 4770 9182 4804
rect 9504 4770 9538 4804
rect 9860 4770 9894 4804
rect 10216 4770 10250 4804
rect 10572 4770 10606 4804
rect 11122 4770 11156 4804
rect 11478 4770 11512 4804
rect 11834 4770 11868 4804
rect 12190 4770 12224 4804
rect 12546 4770 12580 4804
rect 12902 4770 12936 4804
rect 8970 4548 9004 4582
rect 9326 4548 9360 4582
rect 9682 4548 9716 4582
rect 10038 4548 10072 4582
rect 10394 4548 10428 4582
rect 11300 4548 11334 4582
rect 11656 4548 11690 4582
rect 12012 4548 12046 4582
rect 12368 4548 12402 4582
rect 12724 4548 12758 4582
rect 8792 4200 8826 4234
rect 9148 4200 9182 4234
rect 9504 4200 9538 4234
rect 9860 4200 9894 4234
rect 10216 4200 10250 4234
rect 10572 4200 10606 4234
rect 11122 4200 11156 4234
rect 11478 4200 11512 4234
rect 11834 4200 11868 4234
rect 12190 4200 12224 4234
rect 12546 4200 12580 4234
rect 12902 4200 12936 4234
rect 8970 3978 9004 4012
rect 9326 3978 9360 4012
rect 9682 3978 9716 4012
rect 10038 3978 10072 4012
rect 10394 3978 10428 4012
rect 11300 3978 11334 4012
rect 11656 3978 11690 4012
rect 12012 3978 12046 4012
rect 12368 3978 12402 4012
rect 12724 3978 12758 4012
rect 15792 3850 15826 3884
rect 16004 3850 16038 3884
rect 16216 3850 16250 3884
rect 16428 3850 16462 3884
rect 16640 3850 16674 3884
rect 16852 3850 16886 3884
rect 17572 3850 17606 3884
rect 17784 3850 17818 3884
rect 17996 3850 18030 3884
rect 18208 3850 18242 3884
rect 18420 3850 18454 3884
rect 18632 3850 18666 3884
rect 15890 3668 15924 3702
rect 16102 3668 16136 3702
rect 16314 3668 16348 3702
rect 16526 3668 16560 3702
rect 16738 3668 16772 3702
rect 16950 3668 16984 3702
rect 17670 3668 17704 3702
rect 17882 3668 17916 3702
rect 18094 3668 18128 3702
rect 18306 3668 18340 3702
rect 18518 3668 18552 3702
rect 18730 3668 18764 3702
rect 8434 3370 8468 3404
rect 8790 3370 8824 3404
rect 9146 3370 9180 3404
rect 9502 3370 9536 3404
rect 9858 3370 9892 3404
rect 10214 3370 10248 3404
rect 10570 3370 10604 3404
rect 11121 3370 11155 3404
rect 11477 3370 11511 3404
rect 11833 3370 11867 3404
rect 12189 3370 12223 3404
rect 12545 3370 12579 3404
rect 12901 3370 12935 3404
rect 13257 3370 13291 3404
rect 8612 3148 8646 3182
rect 8968 3148 9002 3182
rect 9324 3148 9358 3182
rect 9680 3148 9714 3182
rect 10036 3148 10070 3182
rect 10392 3148 10426 3182
rect 11299 3148 11333 3182
rect 11655 3148 11689 3182
rect 12011 3148 12045 3182
rect 12367 3148 12401 3182
rect 12723 3148 12757 3182
rect 13079 3148 13113 3182
rect 14138 3170 14172 3204
rect 14494 3170 14528 3204
rect 14850 3170 14884 3204
rect 15206 3170 15240 3204
rect 15562 3170 15596 3204
rect 15918 3170 15952 3204
rect 16274 3170 16308 3204
rect 16630 3170 16664 3204
rect 16986 3170 17020 3204
rect 17538 3170 17572 3204
rect 17894 3170 17928 3204
rect 18250 3170 18284 3204
rect 18606 3170 18640 3204
rect 18962 3170 18996 3204
rect 19318 3170 19352 3204
rect 19674 3170 19708 3204
rect 20030 3170 20064 3204
rect 20386 3170 20420 3204
rect 14316 2948 14350 2982
rect 14672 2948 14706 2982
rect 15028 2948 15062 2982
rect 15384 2948 15418 2982
rect 15740 2948 15774 2982
rect 16096 2948 16130 2982
rect 16452 2948 16486 2982
rect 16808 2948 16842 2982
rect 17716 2948 17750 2982
rect 18072 2948 18106 2982
rect 18428 2948 18462 2982
rect 18784 2948 18818 2982
rect 19140 2948 19174 2982
rect 19496 2948 19530 2982
rect 19852 2948 19886 2982
rect 20208 2948 20242 2982
rect 8434 2870 8468 2904
rect 8790 2870 8824 2904
rect 9146 2870 9180 2904
rect 9502 2870 9536 2904
rect 9858 2870 9892 2904
rect 10214 2870 10248 2904
rect 10570 2870 10604 2904
rect 11121 2870 11155 2904
rect 11477 2870 11511 2904
rect 11833 2870 11867 2904
rect 12189 2870 12223 2904
rect 12545 2870 12579 2904
rect 12901 2870 12935 2904
rect 13257 2870 13291 2904
rect 8612 2648 8646 2682
rect 8968 2648 9002 2682
rect 9324 2648 9358 2682
rect 9680 2648 9714 2682
rect 10036 2648 10070 2682
rect 10392 2648 10426 2682
rect 11299 2648 11333 2682
rect 11655 2648 11689 2682
rect 12011 2648 12045 2682
rect 12367 2648 12401 2682
rect 12723 2648 12757 2682
rect 13079 2648 13113 2682
rect 14138 2670 14172 2704
rect 14494 2670 14528 2704
rect 14850 2670 14884 2704
rect 15206 2670 15240 2704
rect 15562 2670 15596 2704
rect 15918 2670 15952 2704
rect 16274 2670 16308 2704
rect 16630 2670 16664 2704
rect 16986 2670 17020 2704
rect 17538 2670 17572 2704
rect 17894 2670 17928 2704
rect 18250 2670 18284 2704
rect 18606 2670 18640 2704
rect 18962 2670 18996 2704
rect 19318 2670 19352 2704
rect 19674 2670 19708 2704
rect 20030 2670 20064 2704
rect 20386 2670 20420 2704
rect 14316 2448 14350 2482
rect 14672 2448 14706 2482
rect 15028 2448 15062 2482
rect 15384 2448 15418 2482
rect 15740 2448 15774 2482
rect 16096 2448 16130 2482
rect 16452 2448 16486 2482
rect 16808 2448 16842 2482
rect 17716 2448 17750 2482
rect 18072 2448 18106 2482
rect 18428 2448 18462 2482
rect 18784 2448 18818 2482
rect 19140 2448 19174 2482
rect 19496 2448 19530 2482
rect 19852 2448 19886 2482
rect 20208 2448 20242 2482
rect 8434 2370 8468 2404
rect 8790 2370 8824 2404
rect 9146 2370 9180 2404
rect 9502 2370 9536 2404
rect 9858 2370 9892 2404
rect 10214 2370 10248 2404
rect 10570 2370 10604 2404
rect 11121 2370 11155 2404
rect 11477 2370 11511 2404
rect 11833 2370 11867 2404
rect 12189 2370 12223 2404
rect 12545 2370 12579 2404
rect 12901 2370 12935 2404
rect 13257 2370 13291 2404
rect 8612 2148 8646 2182
rect 8968 2148 9002 2182
rect 9324 2148 9358 2182
rect 9680 2148 9714 2182
rect 10036 2148 10070 2182
rect 10392 2148 10426 2182
rect 11299 2148 11333 2182
rect 11655 2148 11689 2182
rect 12011 2148 12045 2182
rect 12367 2148 12401 2182
rect 12723 2148 12757 2182
rect 13079 2148 13113 2182
rect 14138 2170 14172 2204
rect 14494 2170 14528 2204
rect 14850 2170 14884 2204
rect 15206 2170 15240 2204
rect 15562 2170 15596 2204
rect 15918 2170 15952 2204
rect 16274 2170 16308 2204
rect 16630 2170 16664 2204
rect 16986 2170 17020 2204
rect 17538 2170 17572 2204
rect 17894 2170 17928 2204
rect 18250 2170 18284 2204
rect 18606 2170 18640 2204
rect 18962 2170 18996 2204
rect 19318 2170 19352 2204
rect 19674 2170 19708 2204
rect 20030 2170 20064 2204
rect 20386 2170 20420 2204
rect 14316 1948 14350 1982
rect 14672 1948 14706 1982
rect 15028 1948 15062 1982
rect 15384 1948 15418 1982
rect 15740 1948 15774 1982
rect 16096 1948 16130 1982
rect 16452 1948 16486 1982
rect 16808 1948 16842 1982
rect 17716 1948 17750 1982
rect 18072 1948 18106 1982
rect 18428 1948 18462 1982
rect 18784 1948 18818 1982
rect 19140 1948 19174 1982
rect 19496 1948 19530 1982
rect 19852 1948 19886 1982
rect 20208 1948 20242 1982
rect 8434 1670 8468 1704
rect 8790 1670 8824 1704
rect 9146 1670 9180 1704
rect 9502 1670 9536 1704
rect 9858 1670 9892 1704
rect 10214 1670 10248 1704
rect 10570 1670 10604 1704
rect 11121 1670 11155 1704
rect 11477 1670 11511 1704
rect 11833 1670 11867 1704
rect 12189 1670 12223 1704
rect 12545 1670 12579 1704
rect 12901 1670 12935 1704
rect 13257 1670 13291 1704
rect 14138 1670 14172 1704
rect 14494 1670 14528 1704
rect 14850 1670 14884 1704
rect 15206 1670 15240 1704
rect 15562 1670 15596 1704
rect 15918 1670 15952 1704
rect 16274 1670 16308 1704
rect 16630 1670 16664 1704
rect 16986 1670 17020 1704
rect 17538 1670 17572 1704
rect 17894 1670 17928 1704
rect 18250 1670 18284 1704
rect 18606 1670 18640 1704
rect 18962 1670 18996 1704
rect 19318 1670 19352 1704
rect 19674 1670 19708 1704
rect 20030 1670 20064 1704
rect 20386 1670 20420 1704
rect 8612 1448 8646 1482
rect 8968 1448 9002 1482
rect 9324 1448 9358 1482
rect 9680 1448 9714 1482
rect 10036 1448 10070 1482
rect 10392 1448 10426 1482
rect 11299 1448 11333 1482
rect 11655 1448 11689 1482
rect 12011 1448 12045 1482
rect 12367 1448 12401 1482
rect 12723 1448 12757 1482
rect 13079 1448 13113 1482
rect 14316 1448 14350 1482
rect 14672 1448 14706 1482
rect 15028 1448 15062 1482
rect 15384 1448 15418 1482
rect 15740 1448 15774 1482
rect 16096 1448 16130 1482
rect 16452 1448 16486 1482
rect 16808 1448 16842 1482
rect 17716 1448 17750 1482
rect 18072 1448 18106 1482
rect 18428 1448 18462 1482
rect 18784 1448 18818 1482
rect 19140 1448 19174 1482
rect 19496 1448 19530 1482
rect 19852 1448 19886 1482
rect 20208 1448 20242 1482
rect 8434 1170 8468 1204
rect 8790 1170 8824 1204
rect 9146 1170 9180 1204
rect 9502 1170 9536 1204
rect 9858 1170 9892 1204
rect 10214 1170 10248 1204
rect 10570 1170 10604 1204
rect 11121 1170 11155 1204
rect 11477 1170 11511 1204
rect 11833 1170 11867 1204
rect 12189 1170 12223 1204
rect 12545 1170 12579 1204
rect 12901 1170 12935 1204
rect 13257 1170 13291 1204
rect 14138 1170 14172 1204
rect 14494 1170 14528 1204
rect 14850 1170 14884 1204
rect 15206 1170 15240 1204
rect 15562 1170 15596 1204
rect 15918 1170 15952 1204
rect 16274 1170 16308 1204
rect 16630 1170 16664 1204
rect 16986 1170 17020 1204
rect 17538 1170 17572 1204
rect 17894 1170 17928 1204
rect 18250 1170 18284 1204
rect 18606 1170 18640 1204
rect 18962 1170 18996 1204
rect 19318 1170 19352 1204
rect 19674 1170 19708 1204
rect 20030 1170 20064 1204
rect 20386 1170 20420 1204
rect 8612 948 8646 982
rect 8968 948 9002 982
rect 9324 948 9358 982
rect 9680 948 9714 982
rect 10036 948 10070 982
rect 10392 948 10426 982
rect 11299 948 11333 982
rect 11655 948 11689 982
rect 12011 948 12045 982
rect 12367 948 12401 982
rect 12723 948 12757 982
rect 13079 948 13113 982
rect 14316 948 14350 982
rect 14672 948 14706 982
rect 15028 948 15062 982
rect 15384 948 15418 982
rect 15740 948 15774 982
rect 16096 948 16130 982
rect 16452 948 16486 982
rect 16808 948 16842 982
rect 17716 948 17750 982
rect 18072 948 18106 982
rect 18428 948 18462 982
rect 18784 948 18818 982
rect 19140 948 19174 982
rect 19496 948 19530 982
rect 19852 948 19886 982
rect 20208 948 20242 982
rect 8434 670 8468 704
rect 8790 670 8824 704
rect 9146 670 9180 704
rect 9502 670 9536 704
rect 9858 670 9892 704
rect 10214 670 10248 704
rect 10570 670 10604 704
rect 11121 670 11155 704
rect 11477 670 11511 704
rect 11833 670 11867 704
rect 12189 670 12223 704
rect 12545 670 12579 704
rect 12901 670 12935 704
rect 13257 670 13291 704
rect 14138 670 14172 704
rect 14494 670 14528 704
rect 14850 670 14884 704
rect 15206 670 15240 704
rect 15562 670 15596 704
rect 15918 670 15952 704
rect 16274 670 16308 704
rect 16630 670 16664 704
rect 16986 670 17020 704
rect 17538 670 17572 704
rect 17894 670 17928 704
rect 18250 670 18284 704
rect 18606 670 18640 704
rect 18962 670 18996 704
rect 19318 670 19352 704
rect 19674 670 19708 704
rect 20030 670 20064 704
rect 20386 670 20420 704
rect 8612 448 8646 482
rect 8968 448 9002 482
rect 9324 448 9358 482
rect 9680 448 9714 482
rect 10036 448 10070 482
rect 10392 448 10426 482
rect 11299 448 11333 482
rect 11655 448 11689 482
rect 12011 448 12045 482
rect 12367 448 12401 482
rect 12723 448 12757 482
rect 13079 448 13113 482
rect 14316 448 14350 482
rect 14672 448 14706 482
rect 15028 448 15062 482
rect 15384 448 15418 482
rect 15740 448 15774 482
rect 16096 448 16130 482
rect 16452 448 16486 482
rect 16808 448 16842 482
rect 17716 448 17750 482
rect 18072 448 18106 482
rect 18428 448 18462 482
rect 18784 448 18818 482
rect 19140 448 19174 482
rect 19496 448 19530 482
rect 19852 448 19886 482
rect 20208 448 20242 482
<< metal1 >>
rect 8770 6268 8780 6269
rect 8424 6262 8780 6268
rect 8838 6268 8848 6269
rect 8838 6262 10618 6268
rect 8424 6228 8436 6262
rect 8470 6228 8780 6262
rect 8838 6228 9148 6262
rect 9182 6228 9504 6262
rect 9538 6228 9860 6262
rect 9894 6228 10204 6262
rect 10262 6228 10572 6262
rect 10606 6228 10618 6262
rect 8424 6222 8780 6228
rect 8770 6211 8780 6222
rect 8838 6222 10204 6228
rect 8838 6211 8848 6222
rect 10194 6204 10204 6222
rect 10262 6222 10618 6228
rect 11110 6262 11466 6268
rect 11524 6263 13304 6268
rect 11524 6262 12890 6263
rect 12948 6262 13304 6263
rect 11110 6228 11122 6262
rect 11156 6228 11466 6262
rect 11524 6228 11834 6262
rect 11868 6228 12190 6262
rect 12224 6228 12546 6262
rect 12580 6228 12890 6262
rect 12948 6228 13258 6262
rect 13292 6228 13304 6262
rect 11110 6222 11466 6228
rect 10262 6204 10272 6222
rect 11456 6210 11466 6222
rect 11524 6222 12890 6228
rect 11524 6210 11534 6222
rect 12880 6205 12890 6222
rect 12948 6222 13304 6228
rect 12948 6205 12958 6222
rect 8948 6046 8958 6058
rect 8602 6040 8958 6046
rect 9016 6046 9026 6058
rect 10016 6046 10026 6058
rect 9016 6040 10026 6046
rect 10084 6046 10094 6058
rect 11634 6046 11644 6058
rect 10084 6040 10440 6046
rect 8602 6006 8614 6040
rect 8648 6006 8958 6040
rect 9016 6006 9326 6040
rect 9360 6006 9682 6040
rect 9716 6006 10026 6040
rect 10084 6006 10394 6040
rect 10428 6006 10440 6040
rect 8602 6000 8958 6006
rect 9016 6000 10026 6006
rect 10084 6000 10440 6006
rect 11288 6040 11644 6046
rect 11702 6046 11712 6058
rect 12702 6046 12712 6058
rect 11702 6040 12712 6046
rect 12770 6046 12780 6058
rect 12770 6040 13126 6046
rect 11288 6006 11300 6040
rect 11334 6006 11644 6040
rect 11702 6006 12012 6040
rect 12046 6006 12368 6040
rect 12402 6006 12712 6040
rect 12770 6006 13080 6040
rect 13114 6006 13126 6040
rect 11288 6000 11644 6006
rect 11702 6000 12712 6006
rect 12770 6000 13126 6006
rect 8568 5944 10511 5947
rect 8568 5937 10538 5944
rect 11229 5937 13172 5947
rect 8504 5913 10538 5937
rect 8504 5877 8580 5913
rect 8074 5819 8084 5877
rect 8142 5819 8152 5877
rect 8504 5819 8514 5877
rect 8572 5819 8582 5877
rect 10462 5874 10538 5913
rect 11190 5936 13172 5937
rect 11190 5913 13224 5936
rect 11190 5874 11266 5913
rect 8504 5778 8580 5819
rect 10461 5816 10471 5874
rect 10529 5816 10539 5874
rect 11190 5816 11200 5874
rect 11258 5816 11268 5874
rect 10462 5778 10538 5816
rect 8504 5759 10538 5778
rect 11190 5777 11266 5816
rect 13148 5777 13224 5913
rect 8504 5752 10512 5759
rect 11190 5752 13224 5777
rect 8560 5744 10512 5752
rect 11234 5751 13224 5752
rect 11234 5743 13177 5751
rect 8424 5685 8780 5691
rect 8838 5685 9492 5691
rect 9550 5685 10204 5691
rect 10262 5685 10618 5691
rect 8424 5651 8436 5685
rect 8470 5651 8780 5685
rect 8838 5651 9148 5685
rect 9182 5651 9492 5685
rect 9550 5651 9860 5685
rect 9894 5651 10204 5685
rect 10262 5651 10572 5685
rect 10606 5651 10618 5685
rect 8424 5645 8780 5651
rect 8770 5633 8780 5645
rect 8838 5645 9492 5651
rect 8838 5633 8848 5645
rect 9482 5633 9492 5645
rect 9550 5645 10204 5651
rect 9550 5633 9560 5645
rect 10194 5633 10204 5645
rect 10262 5645 10618 5651
rect 11110 5684 11466 5690
rect 11524 5684 12178 5690
rect 12236 5684 12890 5690
rect 12948 5684 13304 5690
rect 11110 5650 11122 5684
rect 11156 5650 11466 5684
rect 11524 5650 11834 5684
rect 11868 5650 12178 5684
rect 12236 5650 12546 5684
rect 12580 5650 12890 5684
rect 12948 5650 13258 5684
rect 13292 5650 13304 5684
rect 10262 5633 10272 5645
rect 11110 5644 11466 5650
rect 11456 5632 11466 5644
rect 11524 5644 12178 5650
rect 11524 5632 11534 5644
rect 12168 5632 12178 5644
rect 12236 5644 12890 5650
rect 12236 5632 12246 5644
rect 12880 5632 12890 5644
rect 12948 5644 13304 5650
rect 12948 5632 12958 5644
rect 8948 5469 8958 5481
rect 8602 5463 8958 5469
rect 9016 5469 9026 5481
rect 10016 5469 10026 5481
rect 9016 5463 10026 5469
rect 10084 5469 10094 5481
rect 10084 5463 10440 5469
rect 11634 5468 11644 5480
rect 8602 5429 8614 5463
rect 8648 5429 8958 5463
rect 9016 5429 9326 5463
rect 9360 5429 9682 5463
rect 9716 5429 10026 5463
rect 10084 5429 10394 5463
rect 10428 5429 10440 5463
rect 8602 5423 8958 5429
rect 9016 5423 10026 5429
rect 10084 5423 10440 5429
rect 11288 5462 11644 5468
rect 11702 5468 11712 5480
rect 12702 5468 12712 5480
rect 11702 5462 12712 5468
rect 12770 5468 12780 5480
rect 12770 5462 13126 5468
rect 11288 5428 11300 5462
rect 11334 5428 11644 5462
rect 11702 5428 12012 5462
rect 12046 5428 12368 5462
rect 12402 5428 12712 5462
rect 12770 5428 13080 5462
rect 13114 5428 13126 5462
rect 11288 5422 11644 5428
rect 11702 5422 12712 5428
rect 12770 5422 13126 5428
rect 7980 5010 11266 5127
rect 10462 4903 10538 5010
rect 11190 4897 11266 5010
rect 8924 4863 9645 4897
rect 9762 4863 10512 4897
rect 11190 4864 11969 4897
rect 11229 4863 11969 4864
rect 12086 4863 12817 4897
rect 8770 4752 8780 4810
rect 8838 4804 10560 4810
rect 8838 4770 9148 4804
rect 9182 4770 9504 4804
rect 9538 4770 9860 4804
rect 9894 4770 10216 4804
rect 10250 4770 10560 4804
rect 8838 4764 10560 4770
rect 8838 4752 8848 4764
rect 10550 4752 10560 4764
rect 10618 4752 10628 4810
rect 11100 4752 11110 4810
rect 11168 4804 12890 4810
rect 11168 4770 11478 4804
rect 11512 4770 11834 4804
rect 11868 4770 12190 4804
rect 12224 4770 12546 4804
rect 12580 4770 12890 4804
rect 11168 4764 12890 4770
rect 11168 4752 11178 4764
rect 12880 4752 12890 4764
rect 12948 4752 12958 4810
rect 8948 4542 8958 4600
rect 9016 4588 9026 4600
rect 9482 4588 9492 4600
rect 9016 4582 9492 4588
rect 9016 4548 9326 4582
rect 9360 4548 9492 4582
rect 9016 4542 9492 4548
rect 9550 4588 9560 4600
rect 10372 4588 10382 4600
rect 9550 4582 10382 4588
rect 9550 4548 9682 4582
rect 9716 4548 10038 4582
rect 10072 4548 10382 4582
rect 9550 4542 10382 4548
rect 10440 4542 10450 4600
rect 11278 4542 11288 4600
rect 11346 4588 11356 4600
rect 12168 4588 12178 4600
rect 11346 4582 12178 4588
rect 11346 4548 11656 4582
rect 11690 4548 12012 4582
rect 12046 4548 12178 4582
rect 11346 4542 12178 4548
rect 12236 4588 12246 4600
rect 12702 4588 12712 4600
rect 12236 4582 12712 4588
rect 12236 4548 12368 4582
rect 12402 4548 12712 4582
rect 12236 4542 12712 4548
rect 12770 4542 12780 4600
rect 8860 4327 8936 4484
rect 10462 4327 10538 4483
rect 8860 4299 10538 4327
rect 8913 4298 10538 4299
rect 11190 4327 11266 4479
rect 12792 4327 12868 4485
rect 11190 4300 12868 4327
rect 8913 4293 10501 4298
rect 11190 4294 12832 4300
rect 11244 4293 12832 4294
rect 8770 4182 8780 4240
rect 8838 4234 9490 4240
rect 9548 4234 10560 4240
rect 8838 4200 9148 4234
rect 9182 4200 9490 4234
rect 9548 4200 9860 4234
rect 9894 4200 10216 4234
rect 10250 4200 10560 4234
rect 8838 4194 9490 4200
rect 8838 4182 8848 4194
rect 9480 4182 9490 4194
rect 9548 4194 10560 4200
rect 9548 4182 9558 4194
rect 10550 4182 10560 4194
rect 10618 4182 10628 4240
rect 11100 4182 11110 4240
rect 11168 4234 12178 4240
rect 12236 4234 12890 4240
rect 11168 4200 11478 4234
rect 11512 4200 11834 4234
rect 11868 4200 12178 4234
rect 12236 4200 12546 4234
rect 12580 4200 12890 4234
rect 11168 4194 12178 4200
rect 11168 4182 11178 4194
rect 12168 4182 12178 4194
rect 12236 4194 12890 4200
rect 12236 4182 12246 4194
rect 12880 4182 12890 4194
rect 12948 4182 12958 4240
rect 8948 3972 8958 4030
rect 9016 4018 9026 4030
rect 10372 4018 10382 4030
rect 9016 4012 10382 4018
rect 9016 3978 9326 4012
rect 9360 3978 9682 4012
rect 9716 3978 10038 4012
rect 10072 3978 10382 4012
rect 9016 3972 10382 3978
rect 10440 3972 10450 4030
rect 11278 3972 11288 4030
rect 11346 4018 11356 4030
rect 12702 4018 12712 4030
rect 11346 4012 12712 4018
rect 11346 3978 11656 4012
rect 11690 3978 12012 4012
rect 12046 3978 12368 4012
rect 12402 3978 12712 4012
rect 11346 3972 12712 3978
rect 12770 3972 12780 4030
rect 16249 3984 16315 4631
rect 16349 3984 16359 3986
rect 15825 3928 16359 3984
rect 16417 3984 16427 3986
rect 18029 3984 18095 4631
rect 18129 3984 18139 3986
rect 16417 3928 16739 3984
rect 17097 3928 17163 3984
rect 17605 3928 18139 3984
rect 18197 3984 18207 3986
rect 18197 3928 18519 3984
rect 18877 3928 18943 3984
rect 15780 3884 16898 3890
rect 15780 3850 15792 3884
rect 15826 3850 16004 3884
rect 16038 3850 16216 3884
rect 16250 3850 16428 3884
rect 16462 3850 16640 3884
rect 16674 3850 16783 3884
rect 15780 3844 16783 3850
rect 16773 3826 16783 3844
rect 16841 3850 16852 3884
rect 16886 3850 16898 3884
rect 16841 3844 16898 3850
rect 17446 3884 18678 3890
rect 17446 3844 17503 3884
rect 16841 3826 16851 3844
rect 17493 3826 17503 3844
rect 17561 3850 17572 3884
rect 17606 3850 17784 3884
rect 17818 3850 17996 3884
rect 18030 3850 18208 3884
rect 18242 3850 18420 3884
rect 18454 3850 18632 3884
rect 18666 3850 18678 3884
rect 17561 3844 18678 3850
rect 17561 3826 17571 3844
rect 8071 3673 11265 3790
rect 10460 3488 10536 3673
rect 8566 3458 10536 3488
rect 11189 3488 11265 3673
rect 15868 3668 15878 3726
rect 15936 3708 15946 3726
rect 18708 3708 18718 3720
rect 15936 3702 16996 3708
rect 15936 3668 16102 3702
rect 16136 3668 16314 3702
rect 16348 3668 16526 3702
rect 16560 3668 16738 3702
rect 16772 3668 16950 3702
rect 16984 3668 16996 3702
rect 15878 3662 16996 3668
rect 17658 3702 18718 3708
rect 17658 3668 17670 3702
rect 17704 3668 17882 3702
rect 17916 3668 18094 3702
rect 18128 3668 18306 3702
rect 18340 3668 18518 3702
rect 18552 3668 18718 3702
rect 17658 3662 18718 3668
rect 18776 3662 18786 3720
rect 16349 3624 16359 3626
rect 15613 3568 15679 3624
rect 16037 3568 16359 3624
rect 16417 3624 16427 3626
rect 18129 3624 18139 3626
rect 16417 3568 16951 3624
rect 17393 3568 17459 3624
rect 17817 3568 18139 3624
rect 18197 3624 18207 3626
rect 18197 3568 18731 3624
rect 11189 3469 13211 3488
rect 8566 3454 10524 3458
rect 11253 3454 13211 3469
rect 8412 3352 8422 3410
rect 8480 3404 9490 3410
rect 9548 3404 10558 3410
rect 8480 3370 8790 3404
rect 8824 3370 9146 3404
rect 9180 3370 9490 3404
rect 9548 3370 9858 3404
rect 9892 3370 10214 3404
rect 10248 3370 10558 3404
rect 8480 3364 9490 3370
rect 8480 3352 8490 3364
rect 9480 3352 9490 3364
rect 9548 3364 10558 3370
rect 9548 3352 9558 3364
rect 10548 3352 10558 3364
rect 10616 3352 10626 3410
rect 11099 3352 11109 3410
rect 11167 3404 12177 3410
rect 12235 3404 13245 3410
rect 11167 3370 11477 3404
rect 11511 3370 11833 3404
rect 11867 3370 12177 3404
rect 12235 3370 12545 3404
rect 12579 3370 12901 3404
rect 12935 3370 13245 3404
rect 11167 3364 12177 3370
rect 11167 3352 11177 3364
rect 12167 3352 12177 3364
rect 12235 3364 13245 3370
rect 12235 3352 12245 3364
rect 13235 3352 13245 3364
rect 13303 3352 13313 3410
rect 20276 3288 20352 3519
rect 14218 3254 16940 3288
rect 17664 3254 19030 3288
rect 19106 3255 20352 3288
rect 19106 3254 20346 3255
rect 8946 3188 8956 3200
rect 8600 3182 8956 3188
rect 9014 3188 9024 3200
rect 10014 3188 10024 3200
rect 9014 3182 10024 3188
rect 10082 3188 10092 3200
rect 11633 3188 11643 3200
rect 10082 3182 10438 3188
rect 8600 3148 8612 3182
rect 8646 3148 8956 3182
rect 9014 3148 9324 3182
rect 9358 3148 9680 3182
rect 9714 3148 10024 3182
rect 10082 3148 10392 3182
rect 10426 3148 10438 3182
rect 8600 3142 8956 3148
rect 9014 3142 10024 3148
rect 10082 3142 10438 3148
rect 11287 3182 11643 3188
rect 11701 3188 11711 3200
rect 12701 3188 12711 3200
rect 11701 3182 12711 3188
rect 12769 3188 12779 3200
rect 12769 3182 13125 3188
rect 11287 3148 11299 3182
rect 11333 3148 11643 3182
rect 11701 3148 12011 3182
rect 12045 3148 12367 3182
rect 12401 3148 12711 3182
rect 12769 3148 13079 3182
rect 13113 3148 13125 3182
rect 14116 3152 14126 3210
rect 14184 3204 15550 3210
rect 14184 3170 14494 3204
rect 14528 3170 14850 3204
rect 14884 3170 15206 3204
rect 15240 3170 15550 3204
rect 14184 3164 15550 3170
rect 14184 3152 14194 3164
rect 15540 3152 15550 3164
rect 15608 3164 15878 3210
rect 15936 3204 16974 3210
rect 15952 3170 16274 3204
rect 16308 3170 16630 3204
rect 16664 3170 16974 3204
rect 15608 3152 15618 3164
rect 15868 3152 15878 3164
rect 15936 3164 16974 3170
rect 15936 3152 15946 3164
rect 16964 3152 16974 3164
rect 17032 3164 17526 3210
rect 17584 3204 18718 3210
rect 17584 3170 17894 3204
rect 17928 3170 18250 3204
rect 18284 3170 18606 3204
rect 18640 3170 18718 3204
rect 17032 3152 17042 3164
rect 17516 3152 17526 3164
rect 17584 3164 18718 3170
rect 17584 3152 17594 3164
rect 18708 3152 18718 3164
rect 18776 3164 18950 3210
rect 19008 3204 20374 3210
rect 19008 3170 19318 3204
rect 19352 3170 19674 3204
rect 19708 3170 20030 3204
rect 20064 3170 20374 3204
rect 18776 3152 18786 3164
rect 18940 3152 18950 3164
rect 19008 3164 20374 3170
rect 19008 3152 19018 3164
rect 20364 3152 20374 3164
rect 20432 3152 20442 3210
rect 11287 3142 11643 3148
rect 11701 3142 12711 3148
rect 12769 3142 13125 3148
rect 8502 2988 8578 3086
rect 10460 2988 10536 3085
rect 8502 2963 10536 2988
rect 11189 2988 11265 3086
rect 13147 2988 13223 3085
rect 15006 2988 15016 3000
rect 11189 2963 13223 2988
rect 8566 2962 10536 2963
rect 11253 2962 13223 2963
rect 14304 2982 15016 2988
rect 15074 2988 15084 3000
rect 16074 2988 16084 3000
rect 15074 2982 16084 2988
rect 16142 2988 16152 3000
rect 18406 2988 18416 3000
rect 16142 2982 16854 2988
rect 8566 2954 10519 2962
rect 11253 2954 13206 2962
rect 14304 2948 14316 2982
rect 14350 2948 14672 2982
rect 14706 2948 15016 2982
rect 15074 2948 15384 2982
rect 15418 2948 15740 2982
rect 15774 2948 16084 2982
rect 16142 2948 16452 2982
rect 16486 2948 16808 2982
rect 16842 2948 16854 2982
rect 14304 2942 15016 2948
rect 15074 2942 16084 2948
rect 16142 2942 16854 2948
rect 17704 2982 18416 2988
rect 18474 2988 18484 3000
rect 19474 2988 19484 3000
rect 18474 2982 19484 2988
rect 19542 2988 19552 3000
rect 19542 2982 20254 2988
rect 17704 2948 17716 2982
rect 17750 2948 18072 2982
rect 18106 2948 18416 2982
rect 18474 2948 18784 2982
rect 18818 2948 19140 2982
rect 19174 2948 19484 2982
rect 19542 2948 19852 2982
rect 19886 2948 20208 2982
rect 20242 2948 20254 2982
rect 17704 2942 18416 2948
rect 18474 2942 19484 2948
rect 19542 2942 20254 2948
rect 8412 2852 8422 2910
rect 8480 2904 9490 2910
rect 9548 2904 10558 2910
rect 8480 2870 8790 2904
rect 8824 2870 9146 2904
rect 9180 2870 9490 2904
rect 9548 2870 9858 2904
rect 9892 2870 10214 2904
rect 10248 2870 10558 2904
rect 8480 2864 9490 2870
rect 8480 2852 8490 2864
rect 9480 2852 9490 2864
rect 9548 2864 10558 2870
rect 9548 2852 9558 2864
rect 10548 2852 10558 2864
rect 10616 2852 10626 2910
rect 11099 2852 11109 2910
rect 11167 2904 12177 2910
rect 12235 2904 13245 2910
rect 11167 2870 11477 2904
rect 11511 2870 11833 2904
rect 11867 2870 12177 2904
rect 12235 2870 12545 2904
rect 12579 2870 12901 2904
rect 12935 2870 13245 2904
rect 11167 2864 12177 2870
rect 11167 2852 11177 2864
rect 12167 2852 12177 2864
rect 12235 2864 13245 2870
rect 12235 2852 12245 2864
rect 13235 2852 13245 2864
rect 13303 2852 13313 2910
rect 14206 2791 14282 2865
rect 16876 2790 16952 2867
rect 17606 2790 17682 2870
rect 20276 2789 20352 2871
rect 14270 2754 16940 2788
rect 17660 2754 20342 2788
rect 8946 2688 8956 2700
rect 8600 2682 8956 2688
rect 9014 2688 9024 2700
rect 10014 2688 10024 2700
rect 9014 2682 10024 2688
rect 10082 2688 10092 2700
rect 11633 2688 11643 2700
rect 10082 2682 10438 2688
rect 8600 2648 8612 2682
rect 8646 2648 8956 2682
rect 9014 2648 9324 2682
rect 9358 2648 9680 2682
rect 9714 2648 10024 2682
rect 10082 2648 10392 2682
rect 10426 2648 10438 2682
rect 8600 2642 8956 2648
rect 9014 2642 10024 2648
rect 10082 2642 10438 2648
rect 11287 2682 11643 2688
rect 11701 2688 11711 2700
rect 12701 2688 12711 2700
rect 11701 2682 12711 2688
rect 12769 2688 12779 2700
rect 12769 2682 13125 2688
rect 11287 2648 11299 2682
rect 11333 2648 11643 2682
rect 11701 2648 12011 2682
rect 12045 2648 12367 2682
rect 12401 2648 12711 2682
rect 12769 2648 13079 2682
rect 13113 2648 13125 2682
rect 14116 2652 14126 2710
rect 14184 2704 15550 2710
rect 15608 2704 16974 2710
rect 14184 2670 14494 2704
rect 14528 2670 14850 2704
rect 14884 2670 15206 2704
rect 15240 2670 15550 2704
rect 15608 2670 15918 2704
rect 15952 2670 16274 2704
rect 16308 2670 16630 2704
rect 16664 2670 16974 2704
rect 14184 2664 15550 2670
rect 14184 2652 14194 2664
rect 15540 2652 15550 2664
rect 15608 2664 16974 2670
rect 15608 2652 15618 2664
rect 16964 2652 16974 2664
rect 17032 2652 17042 2710
rect 17516 2652 17526 2710
rect 17584 2704 18950 2710
rect 19008 2704 20374 2710
rect 17584 2670 17894 2704
rect 17928 2670 18250 2704
rect 18284 2670 18606 2704
rect 18640 2670 18950 2704
rect 19008 2670 19318 2704
rect 19352 2670 19674 2704
rect 19708 2670 20030 2704
rect 20064 2670 20374 2704
rect 17584 2664 18950 2670
rect 17584 2652 17594 2664
rect 18940 2652 18950 2664
rect 19008 2664 20374 2670
rect 19008 2652 19018 2664
rect 20364 2652 20374 2664
rect 20432 2652 20442 2710
rect 11287 2642 11643 2648
rect 11701 2642 12711 2648
rect 12769 2642 13125 2648
rect 8502 2488 8578 2581
rect 10460 2488 10536 2590
rect 8502 2467 10536 2488
rect 11189 2488 11265 2581
rect 13147 2488 13223 2590
rect 15006 2488 15016 2501
rect 11189 2467 13223 2488
rect 14304 2482 15016 2488
rect 15074 2488 15084 2501
rect 16074 2488 16084 2500
rect 15074 2482 16084 2488
rect 16142 2488 16152 2500
rect 18406 2488 18416 2500
rect 16142 2482 16854 2488
rect 8502 2458 10497 2467
rect 11189 2458 13184 2467
rect 8544 2454 10497 2458
rect 11231 2454 13184 2458
rect 14304 2448 14316 2482
rect 14350 2448 14672 2482
rect 14706 2448 15016 2482
rect 15074 2448 15384 2482
rect 15418 2448 15740 2482
rect 15774 2448 16084 2482
rect 16142 2448 16452 2482
rect 16486 2448 16808 2482
rect 16842 2448 16854 2482
rect 14304 2443 15016 2448
rect 15074 2443 16084 2448
rect 14304 2442 16084 2443
rect 16142 2442 16854 2448
rect 17704 2482 18416 2488
rect 18474 2488 18484 2500
rect 19474 2488 19484 2500
rect 18474 2482 19484 2488
rect 19542 2488 19552 2500
rect 19542 2482 20254 2488
rect 17704 2448 17716 2482
rect 17750 2448 18072 2482
rect 18106 2448 18416 2482
rect 18474 2448 18784 2482
rect 18818 2448 19140 2482
rect 19174 2448 19484 2482
rect 19542 2448 19852 2482
rect 19886 2448 20208 2482
rect 20242 2448 20254 2482
rect 17704 2442 18416 2448
rect 18474 2442 19484 2448
rect 19542 2442 20254 2448
rect 8412 2352 8422 2410
rect 8480 2404 9490 2410
rect 9548 2404 10558 2410
rect 8480 2370 8790 2404
rect 8824 2370 9146 2404
rect 9180 2370 9490 2404
rect 9548 2370 9858 2404
rect 9892 2370 10214 2404
rect 10248 2370 10558 2404
rect 8480 2364 9490 2370
rect 8480 2352 8490 2364
rect 9480 2352 9490 2364
rect 9548 2364 10558 2370
rect 9548 2352 9558 2364
rect 10548 2352 10558 2364
rect 10616 2352 10626 2410
rect 11099 2352 11109 2410
rect 11167 2404 12177 2410
rect 12235 2404 13245 2410
rect 11167 2370 11477 2404
rect 11511 2370 11833 2404
rect 11867 2370 12177 2404
rect 12235 2370 12545 2404
rect 12579 2370 12901 2404
rect 12935 2370 13245 2404
rect 11167 2364 12177 2370
rect 11167 2352 11177 2364
rect 12167 2352 12177 2364
rect 12235 2364 13245 2370
rect 12235 2352 12245 2364
rect 13235 2352 13245 2364
rect 13303 2352 13313 2410
rect 14206 2288 14282 2365
rect 16876 2291 16952 2368
rect 17606 2291 17682 2371
rect 20276 2288 20352 2370
rect 14257 2254 16939 2288
rect 17660 2254 20342 2288
rect 8946 2188 8956 2200
rect 8600 2182 8956 2188
rect 9014 2188 9024 2200
rect 9302 2188 9312 2200
rect 8600 2148 8612 2182
rect 8646 2148 8956 2182
rect 8600 2142 8956 2148
rect 9014 2142 9312 2188
rect 9370 2188 9380 2200
rect 10014 2188 10024 2200
rect 9370 2182 10024 2188
rect 10082 2188 10092 2200
rect 11633 2188 11643 2200
rect 10082 2182 10438 2188
rect 9370 2148 9680 2182
rect 9714 2148 10024 2182
rect 10082 2148 10392 2182
rect 10426 2148 10438 2182
rect 9370 2142 10024 2148
rect 10082 2142 10438 2148
rect 11287 2182 11643 2188
rect 11701 2188 11711 2200
rect 12345 2188 12355 2200
rect 11701 2182 12355 2188
rect 12413 2188 12423 2200
rect 12701 2188 12711 2200
rect 11287 2148 11299 2182
rect 11333 2148 11643 2182
rect 11701 2148 12011 2182
rect 12045 2148 12355 2182
rect 11287 2142 11643 2148
rect 11701 2142 12355 2148
rect 12413 2142 12711 2188
rect 12769 2188 12779 2200
rect 12769 2182 13125 2188
rect 12769 2148 13079 2182
rect 13113 2148 13125 2182
rect 14116 2152 14126 2210
rect 14184 2204 15550 2210
rect 15608 2204 16974 2210
rect 14184 2170 14494 2204
rect 14528 2170 14850 2204
rect 14884 2170 15206 2204
rect 15240 2170 15550 2204
rect 15608 2170 15918 2204
rect 15952 2170 16274 2204
rect 16308 2170 16630 2204
rect 16664 2170 16974 2204
rect 14184 2164 15550 2170
rect 14184 2152 14194 2164
rect 15540 2152 15550 2164
rect 15608 2164 16974 2170
rect 15608 2152 15618 2164
rect 16964 2152 16974 2164
rect 17032 2152 17042 2210
rect 17516 2152 17526 2210
rect 17584 2204 18950 2210
rect 19008 2204 20374 2210
rect 17584 2170 17894 2204
rect 17928 2170 18250 2204
rect 18284 2170 18606 2204
rect 18640 2170 18950 2204
rect 19008 2170 19318 2204
rect 19352 2170 19674 2204
rect 19708 2170 20030 2204
rect 20064 2170 20374 2204
rect 17584 2164 18950 2170
rect 17584 2152 17594 2164
rect 18940 2152 18950 2164
rect 19008 2164 20374 2170
rect 19008 2152 19018 2164
rect 20364 2152 20374 2164
rect 20432 2152 20442 2210
rect 12769 2142 13125 2148
rect 15006 1988 15016 2000
rect 14304 1982 15016 1988
rect 15074 1988 15084 2000
rect 16074 1988 16084 2000
rect 15074 1982 16084 1988
rect 16142 1988 16152 2000
rect 18406 1988 18416 2000
rect 16142 1982 16854 1988
rect 14304 1948 14316 1982
rect 14350 1948 14672 1982
rect 14706 1948 15016 1982
rect 15074 1948 15384 1982
rect 15418 1948 15740 1982
rect 15774 1948 16084 1982
rect 16142 1948 16452 1982
rect 16486 1948 16808 1982
rect 16842 1948 16854 1982
rect 14304 1942 15016 1948
rect 15074 1942 16084 1948
rect 16142 1942 16854 1948
rect 17704 1982 18416 1988
rect 18474 1988 18484 2000
rect 19474 1988 19484 2000
rect 18474 1982 19484 1988
rect 19542 1988 19552 2000
rect 19542 1982 20254 1988
rect 17704 1948 17716 1982
rect 17750 1948 18072 1982
rect 18106 1948 18416 1982
rect 18474 1948 18784 1982
rect 18818 1948 19140 1982
rect 19174 1948 19484 1982
rect 19542 1948 19852 1982
rect 19886 1948 20208 1982
rect 20242 1948 20254 1982
rect 17704 1942 18416 1948
rect 18474 1942 19484 1948
rect 19542 1942 20254 1948
rect 14206 1789 14282 1866
rect 16876 1791 16952 1868
rect 17606 1790 17682 1870
rect 20276 1789 20352 1871
rect 8566 1754 10524 1788
rect 11253 1754 13211 1788
rect 14253 1754 16935 1788
rect 17659 1754 20341 1788
rect 8412 1652 8422 1710
rect 8480 1704 9312 1710
rect 8480 1670 8790 1704
rect 8824 1670 9146 1704
rect 9180 1670 9312 1704
rect 8480 1664 9312 1670
rect 8480 1652 8490 1664
rect 9302 1652 9312 1664
rect 9370 1664 9490 1710
rect 9548 1704 10558 1710
rect 9548 1670 9858 1704
rect 9892 1670 10214 1704
rect 10248 1670 10558 1704
rect 9370 1652 9380 1664
rect 9480 1652 9490 1664
rect 9548 1664 10558 1670
rect 9548 1652 9558 1664
rect 10548 1652 10558 1664
rect 10616 1652 10626 1710
rect 11099 1652 11109 1710
rect 11167 1704 12177 1710
rect 11167 1670 11477 1704
rect 11511 1670 11833 1704
rect 11867 1670 12177 1704
rect 11167 1664 12177 1670
rect 11167 1652 11177 1664
rect 12167 1652 12177 1664
rect 12235 1664 12355 1710
rect 12235 1652 12245 1664
rect 12345 1652 12355 1664
rect 12413 1704 13245 1710
rect 12413 1670 12545 1704
rect 12579 1670 12901 1704
rect 12935 1670 13245 1704
rect 12413 1664 13245 1670
rect 12413 1652 12423 1664
rect 13235 1652 13245 1664
rect 13303 1652 13313 1710
rect 14116 1652 14126 1710
rect 14184 1704 15550 1710
rect 15608 1704 16974 1710
rect 14184 1670 14494 1704
rect 14528 1670 14850 1704
rect 14884 1670 15206 1704
rect 15240 1670 15550 1704
rect 15608 1670 15918 1704
rect 15952 1670 16274 1704
rect 16308 1670 16630 1704
rect 16664 1670 16974 1704
rect 14184 1664 15550 1670
rect 14184 1652 14194 1664
rect 15540 1652 15550 1664
rect 15608 1664 16974 1670
rect 15608 1652 15618 1664
rect 16964 1652 16974 1664
rect 17032 1652 17042 1710
rect 17516 1652 17526 1710
rect 17584 1704 18950 1710
rect 19008 1704 20374 1710
rect 17584 1670 17894 1704
rect 17928 1670 18250 1704
rect 18284 1670 18606 1704
rect 18640 1670 18950 1704
rect 19008 1670 19318 1704
rect 19352 1670 19674 1704
rect 19708 1670 20030 1704
rect 20064 1670 20374 1704
rect 17584 1664 18950 1670
rect 17584 1652 17594 1664
rect 18940 1652 18950 1664
rect 19008 1664 20374 1670
rect 19008 1652 19018 1664
rect 20364 1652 20374 1664
rect 20432 1652 20442 1710
rect 8946 1488 8956 1500
rect 8600 1482 8956 1488
rect 9014 1488 9024 1500
rect 10014 1488 10024 1500
rect 9014 1482 10024 1488
rect 10082 1488 10092 1500
rect 11633 1488 11643 1500
rect 10082 1482 10438 1488
rect 8600 1448 8612 1482
rect 8646 1448 8956 1482
rect 9014 1448 9324 1482
rect 9358 1448 9680 1482
rect 9714 1448 10024 1482
rect 10082 1448 10392 1482
rect 10426 1448 10438 1482
rect 8600 1442 8956 1448
rect 9014 1442 10024 1448
rect 10082 1442 10438 1448
rect 11287 1482 11643 1488
rect 11701 1488 11711 1500
rect 12701 1488 12711 1500
rect 11701 1482 12711 1488
rect 12769 1488 12779 1500
rect 15006 1488 15016 1500
rect 12769 1482 13125 1488
rect 11287 1448 11299 1482
rect 11333 1448 11643 1482
rect 11701 1448 12011 1482
rect 12045 1448 12367 1482
rect 12401 1448 12711 1482
rect 12769 1448 13079 1482
rect 13113 1448 13125 1482
rect 11287 1442 11643 1448
rect 11701 1442 12711 1448
rect 12769 1442 13125 1448
rect 14304 1482 15016 1488
rect 15074 1488 15084 1500
rect 16074 1488 16084 1500
rect 15074 1482 16084 1488
rect 16142 1488 16152 1500
rect 18406 1488 18416 1500
rect 16142 1482 16854 1488
rect 14304 1448 14316 1482
rect 14350 1448 14672 1482
rect 14706 1448 15016 1482
rect 15074 1448 15384 1482
rect 15418 1448 15740 1482
rect 15774 1448 16084 1482
rect 16142 1448 16452 1482
rect 16486 1448 16808 1482
rect 16842 1448 16854 1482
rect 14304 1442 15016 1448
rect 15074 1442 16084 1448
rect 16142 1442 16854 1448
rect 17704 1482 18416 1488
rect 18474 1488 18484 1500
rect 19474 1488 19484 1500
rect 18474 1482 19484 1488
rect 19542 1488 19552 1500
rect 19542 1482 20254 1488
rect 17704 1448 17716 1482
rect 17750 1448 18072 1482
rect 18106 1448 18416 1482
rect 18474 1448 18784 1482
rect 18818 1448 19140 1482
rect 19174 1448 19484 1482
rect 19542 1448 19852 1482
rect 19886 1448 20208 1482
rect 20242 1448 20254 1482
rect 17704 1442 18416 1448
rect 18474 1442 19484 1448
rect 19542 1442 20254 1448
rect 8502 1288 8578 1386
rect 10460 1288 10536 1385
rect 8502 1263 10536 1288
rect 11189 1288 11265 1386
rect 13147 1288 13223 1385
rect 14206 1290 14282 1367
rect 16876 1290 16952 1367
rect 17606 1291 17682 1371
rect 20276 1289 20352 1371
rect 11189 1263 13223 1288
rect 8566 1262 10536 1263
rect 11253 1262 13223 1263
rect 8566 1254 10519 1262
rect 11253 1254 13206 1262
rect 14252 1254 16934 1288
rect 17662 1254 20344 1288
rect 8412 1152 8422 1210
rect 8480 1204 9490 1210
rect 9548 1204 10558 1210
rect 8480 1170 8790 1204
rect 8824 1170 9146 1204
rect 9180 1170 9490 1204
rect 9548 1170 9858 1204
rect 9892 1170 10214 1204
rect 10248 1170 10558 1204
rect 8480 1164 9490 1170
rect 8480 1152 8490 1164
rect 9480 1152 9490 1164
rect 9548 1164 10558 1170
rect 9548 1152 9558 1164
rect 10548 1152 10558 1164
rect 10616 1152 10626 1210
rect 11099 1152 11109 1210
rect 11167 1204 12177 1210
rect 12235 1204 13245 1210
rect 11167 1170 11477 1204
rect 11511 1170 11833 1204
rect 11867 1170 12177 1204
rect 12235 1170 12545 1204
rect 12579 1170 12901 1204
rect 12935 1170 13245 1204
rect 11167 1164 12177 1170
rect 11167 1152 11177 1164
rect 12167 1152 12177 1164
rect 12235 1164 13245 1170
rect 12235 1152 12245 1164
rect 13235 1152 13245 1164
rect 13303 1152 13313 1210
rect 14116 1152 14126 1210
rect 14184 1204 15550 1210
rect 15608 1204 16974 1210
rect 14184 1170 14494 1204
rect 14528 1170 14850 1204
rect 14884 1170 15206 1204
rect 15240 1170 15550 1204
rect 15608 1170 15918 1204
rect 15952 1170 16274 1204
rect 16308 1170 16630 1204
rect 16664 1170 16974 1204
rect 14184 1164 15550 1170
rect 14184 1152 14194 1164
rect 15540 1152 15550 1164
rect 15608 1164 16974 1170
rect 15608 1152 15618 1164
rect 16964 1152 16974 1164
rect 17032 1152 17042 1210
rect 17516 1152 17526 1210
rect 17584 1204 18950 1210
rect 19008 1204 20374 1210
rect 17584 1170 17894 1204
rect 17928 1170 18250 1204
rect 18284 1170 18606 1204
rect 18640 1170 18950 1204
rect 19008 1170 19318 1204
rect 19352 1170 19674 1204
rect 19708 1170 20030 1204
rect 20064 1170 20374 1204
rect 17584 1164 18950 1170
rect 17584 1152 17594 1164
rect 18940 1152 18950 1164
rect 19008 1164 20374 1170
rect 19008 1152 19018 1164
rect 20364 1152 20374 1164
rect 20432 1152 20442 1210
rect 8946 988 8956 1000
rect 8600 982 8956 988
rect 9014 988 9024 1000
rect 10014 988 10024 1000
rect 9014 982 10024 988
rect 10082 988 10092 1000
rect 11633 988 11643 1000
rect 10082 982 10438 988
rect 8600 948 8612 982
rect 8646 948 8956 982
rect 9014 948 9324 982
rect 9358 948 9680 982
rect 9714 948 10024 982
rect 10082 948 10392 982
rect 10426 948 10438 982
rect 8600 942 8956 948
rect 9014 942 10024 948
rect 10082 942 10438 948
rect 11287 982 11643 988
rect 11701 988 11711 1000
rect 12701 988 12711 1000
rect 11701 982 12711 988
rect 12769 988 12779 1000
rect 15006 988 15016 1000
rect 12769 982 13125 988
rect 11287 948 11299 982
rect 11333 948 11643 982
rect 11701 948 12011 982
rect 12045 948 12367 982
rect 12401 948 12711 982
rect 12769 948 13079 982
rect 13113 948 13125 982
rect 11287 942 11643 948
rect 11701 942 12711 948
rect 12769 942 13125 948
rect 14304 982 15016 988
rect 15074 988 15084 1000
rect 16074 988 16084 1000
rect 15074 982 16084 988
rect 16142 988 16152 1000
rect 18406 988 18416 1000
rect 16142 982 16854 988
rect 14304 948 14316 982
rect 14350 948 14672 982
rect 14706 948 15016 982
rect 15074 948 15384 982
rect 15418 948 15740 982
rect 15774 948 16084 982
rect 16142 948 16452 982
rect 16486 948 16808 982
rect 16842 948 16854 982
rect 14304 942 15016 948
rect 15074 942 16084 948
rect 16142 942 16854 948
rect 17704 982 18416 988
rect 18474 988 18484 1000
rect 19474 988 19484 1000
rect 18474 982 19484 988
rect 19542 988 19552 1000
rect 19542 982 20254 988
rect 17704 948 17716 982
rect 17750 948 18072 982
rect 18106 948 18416 982
rect 18474 948 18784 982
rect 18818 948 19140 982
rect 19174 948 19484 982
rect 19542 948 19852 982
rect 19886 948 20208 982
rect 20242 948 20254 982
rect 17704 942 18416 948
rect 18474 942 19484 948
rect 19542 942 20254 948
rect 8502 788 8578 881
rect 10460 788 10536 890
rect 8502 767 10536 788
rect 11189 788 11265 881
rect 13147 788 13223 890
rect 14206 790 14282 867
rect 16876 791 16952 868
rect 17606 790 17682 870
rect 20276 788 20352 870
rect 11189 767 13223 788
rect 8502 758 10497 767
rect 11189 758 13184 767
rect 8544 754 10497 758
rect 11231 754 13184 758
rect 14255 754 16937 788
rect 17659 754 20341 788
rect 8412 652 8422 710
rect 8480 704 9490 710
rect 9548 704 10558 710
rect 8480 670 8790 704
rect 8824 670 9146 704
rect 9180 670 9490 704
rect 9548 670 9858 704
rect 9892 670 10214 704
rect 10248 670 10558 704
rect 8480 664 9490 670
rect 8480 652 8490 664
rect 9480 652 9490 664
rect 9548 664 10558 670
rect 9548 652 9558 664
rect 10548 652 10558 664
rect 10616 652 10626 710
rect 11099 652 11109 710
rect 11167 704 12177 710
rect 12235 704 13245 710
rect 11167 670 11477 704
rect 11511 670 11833 704
rect 11867 670 12177 704
rect 12235 670 12545 704
rect 12579 670 12901 704
rect 12935 670 13245 704
rect 11167 664 12177 670
rect 11167 652 11177 664
rect 12167 652 12177 664
rect 12235 664 13245 670
rect 12235 652 12245 664
rect 13235 652 13245 664
rect 13303 652 13313 710
rect 14116 652 14126 710
rect 14184 704 15550 710
rect 15608 704 16974 710
rect 14184 670 14494 704
rect 14528 670 14850 704
rect 14884 670 15206 704
rect 15240 670 15550 704
rect 15608 670 15918 704
rect 15952 670 16274 704
rect 16308 670 16630 704
rect 16664 670 16974 704
rect 14184 664 15550 670
rect 14184 652 14194 664
rect 15540 652 15550 664
rect 15608 664 16974 670
rect 15608 652 15618 664
rect 16964 652 16974 664
rect 17032 664 17526 710
rect 17584 704 18950 710
rect 19008 704 20374 710
rect 17584 670 17894 704
rect 17928 670 18250 704
rect 18284 670 18606 704
rect 18640 670 18950 704
rect 19008 670 19318 704
rect 19352 670 19674 704
rect 19708 670 20030 704
rect 20064 670 20374 704
rect 17032 652 17042 664
rect 17516 652 17526 664
rect 17584 664 18950 670
rect 17584 652 17594 664
rect 18940 652 18950 664
rect 19008 664 20374 670
rect 19008 652 19018 664
rect 20364 652 20374 664
rect 20432 652 20442 710
rect 8946 488 8956 500
rect 8600 482 8956 488
rect 9014 488 9024 500
rect 10014 488 10024 500
rect 9014 482 10024 488
rect 10082 488 10092 500
rect 11633 488 11643 500
rect 10082 482 10438 488
rect 8600 448 8612 482
rect 8646 448 8956 482
rect 9014 448 9324 482
rect 9358 448 9680 482
rect 9714 448 10024 482
rect 10082 448 10392 482
rect 10426 448 10438 482
rect 8600 442 8956 448
rect 9014 442 10024 448
rect 10082 442 10438 448
rect 11287 482 11643 488
rect 11701 488 11711 500
rect 12701 488 12711 500
rect 11701 482 12711 488
rect 12769 488 12779 500
rect 15006 488 15016 500
rect 12769 482 13125 488
rect 11287 448 11299 482
rect 11333 448 11643 482
rect 11701 448 12011 482
rect 12045 448 12367 482
rect 12401 448 12711 482
rect 12769 448 13079 482
rect 13113 448 13125 482
rect 11287 442 11643 448
rect 11701 442 12711 448
rect 12769 442 13125 448
rect 14304 482 15016 488
rect 15074 488 15084 500
rect 16074 488 16084 500
rect 15074 482 16084 488
rect 16142 488 16152 500
rect 18406 488 18416 500
rect 16142 482 16854 488
rect 14304 448 14316 482
rect 14350 448 14672 482
rect 14706 448 15016 482
rect 15074 448 15384 482
rect 15418 448 15740 482
rect 15774 448 16084 482
rect 16142 448 16452 482
rect 16486 448 16808 482
rect 16842 448 16854 482
rect 14304 442 15016 448
rect 15074 442 16084 448
rect 16142 442 16854 448
rect 17704 482 18416 488
rect 18474 488 18484 500
rect 19474 488 19484 500
rect 18474 482 19484 488
rect 19542 488 19552 500
rect 19542 482 20254 488
rect 17704 448 17716 482
rect 17750 448 18072 482
rect 18106 448 18416 482
rect 18474 448 18784 482
rect 18818 448 19140 482
rect 19174 448 19484 482
rect 19542 448 19852 482
rect 19886 448 20208 482
rect 20242 448 20254 482
rect 17704 442 18416 448
rect 18474 442 19484 448
rect 19542 442 20254 448
rect 8560 364 10513 398
rect 11230 374 13183 398
rect 11188 364 13183 374
rect 14254 364 16936 398
rect 10460 75 10536 360
rect 11188 75 11264 364
rect 15630 75 15706 358
rect 8272 -42 15706 75
<< via1 >>
rect 8780 6262 8838 6269
rect 8780 6228 8792 6262
rect 8792 6228 8826 6262
rect 8826 6228 8838 6262
rect 10204 6228 10216 6262
rect 10216 6228 10250 6262
rect 10250 6228 10262 6262
rect 8780 6211 8838 6228
rect 10204 6204 10262 6228
rect 11466 6262 11524 6268
rect 12890 6262 12948 6263
rect 11466 6228 11478 6262
rect 11478 6228 11512 6262
rect 11512 6228 11524 6262
rect 12890 6228 12902 6262
rect 12902 6228 12936 6262
rect 12936 6228 12948 6262
rect 11466 6210 11524 6228
rect 12890 6205 12948 6228
rect 8958 6040 9016 6058
rect 10026 6040 10084 6058
rect 8958 6006 8970 6040
rect 8970 6006 9004 6040
rect 9004 6006 9016 6040
rect 10026 6006 10038 6040
rect 10038 6006 10072 6040
rect 10072 6006 10084 6040
rect 8958 6000 9016 6006
rect 10026 6000 10084 6006
rect 11644 6040 11702 6058
rect 12712 6040 12770 6058
rect 11644 6006 11656 6040
rect 11656 6006 11690 6040
rect 11690 6006 11702 6040
rect 12712 6006 12724 6040
rect 12724 6006 12758 6040
rect 12758 6006 12770 6040
rect 11644 6000 11702 6006
rect 12712 6000 12770 6006
rect 8084 5819 8142 5877
rect 8514 5819 8572 5877
rect 10471 5816 10529 5874
rect 11200 5816 11258 5874
rect 8780 5685 8838 5691
rect 9492 5685 9550 5691
rect 10204 5685 10262 5691
rect 8780 5651 8792 5685
rect 8792 5651 8826 5685
rect 8826 5651 8838 5685
rect 9492 5651 9504 5685
rect 9504 5651 9538 5685
rect 9538 5651 9550 5685
rect 10204 5651 10216 5685
rect 10216 5651 10250 5685
rect 10250 5651 10262 5685
rect 8780 5633 8838 5651
rect 9492 5633 9550 5651
rect 10204 5633 10262 5651
rect 11466 5684 11524 5690
rect 12178 5684 12236 5690
rect 12890 5684 12948 5690
rect 11466 5650 11478 5684
rect 11478 5650 11512 5684
rect 11512 5650 11524 5684
rect 12178 5650 12190 5684
rect 12190 5650 12224 5684
rect 12224 5650 12236 5684
rect 12890 5650 12902 5684
rect 12902 5650 12936 5684
rect 12936 5650 12948 5684
rect 11466 5632 11524 5650
rect 12178 5632 12236 5650
rect 12890 5632 12948 5650
rect 8958 5463 9016 5481
rect 10026 5463 10084 5481
rect 8958 5429 8970 5463
rect 8970 5429 9004 5463
rect 9004 5429 9016 5463
rect 10026 5429 10038 5463
rect 10038 5429 10072 5463
rect 10072 5429 10084 5463
rect 8958 5423 9016 5429
rect 10026 5423 10084 5429
rect 11644 5462 11702 5480
rect 12712 5462 12770 5480
rect 11644 5428 11656 5462
rect 11656 5428 11690 5462
rect 11690 5428 11702 5462
rect 12712 5428 12724 5462
rect 12724 5428 12758 5462
rect 12758 5428 12770 5462
rect 11644 5422 11702 5428
rect 12712 5422 12770 5428
rect 8780 4804 8838 4810
rect 10560 4804 10618 4810
rect 8780 4770 8792 4804
rect 8792 4770 8826 4804
rect 8826 4770 8838 4804
rect 10560 4770 10572 4804
rect 10572 4770 10606 4804
rect 10606 4770 10618 4804
rect 8780 4752 8838 4770
rect 10560 4752 10618 4770
rect 11110 4804 11168 4810
rect 12890 4804 12948 4810
rect 11110 4770 11122 4804
rect 11122 4770 11156 4804
rect 11156 4770 11168 4804
rect 12890 4770 12902 4804
rect 12902 4770 12936 4804
rect 12936 4770 12948 4804
rect 11110 4752 11168 4770
rect 12890 4752 12948 4770
rect 8958 4582 9016 4600
rect 8958 4548 8970 4582
rect 8970 4548 9004 4582
rect 9004 4548 9016 4582
rect 8958 4542 9016 4548
rect 9492 4542 9550 4600
rect 10382 4582 10440 4600
rect 10382 4548 10394 4582
rect 10394 4548 10428 4582
rect 10428 4548 10440 4582
rect 10382 4542 10440 4548
rect 11288 4582 11346 4600
rect 11288 4548 11300 4582
rect 11300 4548 11334 4582
rect 11334 4548 11346 4582
rect 11288 4542 11346 4548
rect 12178 4542 12236 4600
rect 12712 4582 12770 4600
rect 12712 4548 12724 4582
rect 12724 4548 12758 4582
rect 12758 4548 12770 4582
rect 12712 4542 12770 4548
rect 8780 4234 8838 4240
rect 9490 4234 9548 4240
rect 10560 4234 10618 4240
rect 8780 4200 8792 4234
rect 8792 4200 8826 4234
rect 8826 4200 8838 4234
rect 9490 4200 9504 4234
rect 9504 4200 9538 4234
rect 9538 4200 9548 4234
rect 10560 4200 10572 4234
rect 10572 4200 10606 4234
rect 10606 4200 10618 4234
rect 8780 4182 8838 4200
rect 9490 4182 9548 4200
rect 10560 4182 10618 4200
rect 11110 4234 11168 4240
rect 12178 4234 12236 4240
rect 12890 4234 12948 4240
rect 11110 4200 11122 4234
rect 11122 4200 11156 4234
rect 11156 4200 11168 4234
rect 12178 4200 12190 4234
rect 12190 4200 12224 4234
rect 12224 4200 12236 4234
rect 12890 4200 12902 4234
rect 12902 4200 12936 4234
rect 12936 4200 12948 4234
rect 11110 4182 11168 4200
rect 12178 4182 12236 4200
rect 12890 4182 12948 4200
rect 8958 4012 9016 4030
rect 10382 4012 10440 4030
rect 8958 3978 8970 4012
rect 8970 3978 9004 4012
rect 9004 3978 9016 4012
rect 10382 3978 10394 4012
rect 10394 3978 10428 4012
rect 10428 3978 10440 4012
rect 8958 3972 9016 3978
rect 10382 3972 10440 3978
rect 11288 4012 11346 4030
rect 12712 4012 12770 4030
rect 11288 3978 11300 4012
rect 11300 3978 11334 4012
rect 11334 3978 11346 4012
rect 12712 3978 12724 4012
rect 12724 3978 12758 4012
rect 12758 3978 12770 4012
rect 11288 3972 11346 3978
rect 12712 3972 12770 3978
rect 16359 3928 16417 3986
rect 18139 3928 18197 3986
rect 16783 3826 16841 3884
rect 17503 3826 17561 3884
rect 15878 3702 15936 3726
rect 15878 3668 15890 3702
rect 15890 3668 15924 3702
rect 15924 3668 15936 3702
rect 18718 3702 18776 3720
rect 18718 3668 18730 3702
rect 18730 3668 18764 3702
rect 18764 3668 18776 3702
rect 18718 3662 18776 3668
rect 16359 3568 16417 3626
rect 18139 3568 18197 3626
rect 8422 3404 8480 3410
rect 9490 3404 9548 3410
rect 10558 3404 10616 3410
rect 8422 3370 8434 3404
rect 8434 3370 8468 3404
rect 8468 3370 8480 3404
rect 9490 3370 9502 3404
rect 9502 3370 9536 3404
rect 9536 3370 9548 3404
rect 10558 3370 10570 3404
rect 10570 3370 10604 3404
rect 10604 3370 10616 3404
rect 8422 3352 8480 3370
rect 9490 3352 9548 3370
rect 10558 3352 10616 3370
rect 11109 3404 11167 3410
rect 12177 3404 12235 3410
rect 13245 3404 13303 3410
rect 11109 3370 11121 3404
rect 11121 3370 11155 3404
rect 11155 3370 11167 3404
rect 12177 3370 12189 3404
rect 12189 3370 12223 3404
rect 12223 3370 12235 3404
rect 13245 3370 13257 3404
rect 13257 3370 13291 3404
rect 13291 3370 13303 3404
rect 11109 3352 11167 3370
rect 12177 3352 12235 3370
rect 13245 3352 13303 3370
rect 8956 3182 9014 3200
rect 10024 3182 10082 3200
rect 8956 3148 8968 3182
rect 8968 3148 9002 3182
rect 9002 3148 9014 3182
rect 10024 3148 10036 3182
rect 10036 3148 10070 3182
rect 10070 3148 10082 3182
rect 8956 3142 9014 3148
rect 10024 3142 10082 3148
rect 11643 3182 11701 3200
rect 12711 3182 12769 3200
rect 11643 3148 11655 3182
rect 11655 3148 11689 3182
rect 11689 3148 11701 3182
rect 12711 3148 12723 3182
rect 12723 3148 12757 3182
rect 12757 3148 12769 3182
rect 14126 3204 14184 3210
rect 15550 3204 15608 3210
rect 14126 3170 14138 3204
rect 14138 3170 14172 3204
rect 14172 3170 14184 3204
rect 15550 3170 15562 3204
rect 15562 3170 15596 3204
rect 15596 3170 15608 3204
rect 14126 3152 14184 3170
rect 15550 3152 15608 3170
rect 15878 3204 15936 3210
rect 16974 3204 17032 3210
rect 15878 3170 15918 3204
rect 15918 3170 15936 3204
rect 16974 3170 16986 3204
rect 16986 3170 17020 3204
rect 17020 3170 17032 3204
rect 15878 3152 15936 3170
rect 16974 3152 17032 3170
rect 17526 3204 17584 3210
rect 17526 3170 17538 3204
rect 17538 3170 17572 3204
rect 17572 3170 17584 3204
rect 17526 3152 17584 3170
rect 18718 3152 18776 3210
rect 18950 3204 19008 3210
rect 20374 3204 20432 3210
rect 18950 3170 18962 3204
rect 18962 3170 18996 3204
rect 18996 3170 19008 3204
rect 20374 3170 20386 3204
rect 20386 3170 20420 3204
rect 20420 3170 20432 3204
rect 18950 3152 19008 3170
rect 20374 3152 20432 3170
rect 11643 3142 11701 3148
rect 12711 3142 12769 3148
rect 15016 2982 15074 3000
rect 16084 2982 16142 3000
rect 15016 2948 15028 2982
rect 15028 2948 15062 2982
rect 15062 2948 15074 2982
rect 16084 2948 16096 2982
rect 16096 2948 16130 2982
rect 16130 2948 16142 2982
rect 15016 2942 15074 2948
rect 16084 2942 16142 2948
rect 18416 2982 18474 3000
rect 19484 2982 19542 3000
rect 18416 2948 18428 2982
rect 18428 2948 18462 2982
rect 18462 2948 18474 2982
rect 19484 2948 19496 2982
rect 19496 2948 19530 2982
rect 19530 2948 19542 2982
rect 18416 2942 18474 2948
rect 19484 2942 19542 2948
rect 8422 2904 8480 2910
rect 9490 2904 9548 2910
rect 10558 2904 10616 2910
rect 8422 2870 8434 2904
rect 8434 2870 8468 2904
rect 8468 2870 8480 2904
rect 9490 2870 9502 2904
rect 9502 2870 9536 2904
rect 9536 2870 9548 2904
rect 10558 2870 10570 2904
rect 10570 2870 10604 2904
rect 10604 2870 10616 2904
rect 8422 2852 8480 2870
rect 9490 2852 9548 2870
rect 10558 2852 10616 2870
rect 11109 2904 11167 2910
rect 12177 2904 12235 2910
rect 13245 2904 13303 2910
rect 11109 2870 11121 2904
rect 11121 2870 11155 2904
rect 11155 2870 11167 2904
rect 12177 2870 12189 2904
rect 12189 2870 12223 2904
rect 12223 2870 12235 2904
rect 13245 2870 13257 2904
rect 13257 2870 13291 2904
rect 13291 2870 13303 2904
rect 11109 2852 11167 2870
rect 12177 2852 12235 2870
rect 13245 2852 13303 2870
rect 8956 2682 9014 2700
rect 10024 2682 10082 2700
rect 8956 2648 8968 2682
rect 8968 2648 9002 2682
rect 9002 2648 9014 2682
rect 10024 2648 10036 2682
rect 10036 2648 10070 2682
rect 10070 2648 10082 2682
rect 8956 2642 9014 2648
rect 10024 2642 10082 2648
rect 11643 2682 11701 2700
rect 12711 2682 12769 2700
rect 11643 2648 11655 2682
rect 11655 2648 11689 2682
rect 11689 2648 11701 2682
rect 12711 2648 12723 2682
rect 12723 2648 12757 2682
rect 12757 2648 12769 2682
rect 14126 2704 14184 2710
rect 15550 2704 15608 2710
rect 16974 2704 17032 2710
rect 14126 2670 14138 2704
rect 14138 2670 14172 2704
rect 14172 2670 14184 2704
rect 15550 2670 15562 2704
rect 15562 2670 15596 2704
rect 15596 2670 15608 2704
rect 16974 2670 16986 2704
rect 16986 2670 17020 2704
rect 17020 2670 17032 2704
rect 14126 2652 14184 2670
rect 15550 2652 15608 2670
rect 16974 2652 17032 2670
rect 17526 2704 17584 2710
rect 18950 2704 19008 2710
rect 20374 2704 20432 2710
rect 17526 2670 17538 2704
rect 17538 2670 17572 2704
rect 17572 2670 17584 2704
rect 18950 2670 18962 2704
rect 18962 2670 18996 2704
rect 18996 2670 19008 2704
rect 20374 2670 20386 2704
rect 20386 2670 20420 2704
rect 20420 2670 20432 2704
rect 17526 2652 17584 2670
rect 18950 2652 19008 2670
rect 20374 2652 20432 2670
rect 11643 2642 11701 2648
rect 12711 2642 12769 2648
rect 15016 2482 15074 2501
rect 16084 2482 16142 2500
rect 15016 2448 15028 2482
rect 15028 2448 15062 2482
rect 15062 2448 15074 2482
rect 16084 2448 16096 2482
rect 16096 2448 16130 2482
rect 16130 2448 16142 2482
rect 15016 2443 15074 2448
rect 16084 2442 16142 2448
rect 18416 2482 18474 2500
rect 19484 2482 19542 2500
rect 18416 2448 18428 2482
rect 18428 2448 18462 2482
rect 18462 2448 18474 2482
rect 19484 2448 19496 2482
rect 19496 2448 19530 2482
rect 19530 2448 19542 2482
rect 18416 2442 18474 2448
rect 19484 2442 19542 2448
rect 8422 2404 8480 2410
rect 9490 2404 9548 2410
rect 10558 2404 10616 2410
rect 8422 2370 8434 2404
rect 8434 2370 8468 2404
rect 8468 2370 8480 2404
rect 9490 2370 9502 2404
rect 9502 2370 9536 2404
rect 9536 2370 9548 2404
rect 10558 2370 10570 2404
rect 10570 2370 10604 2404
rect 10604 2370 10616 2404
rect 8422 2352 8480 2370
rect 9490 2352 9548 2370
rect 10558 2352 10616 2370
rect 11109 2404 11167 2410
rect 12177 2404 12235 2410
rect 13245 2404 13303 2410
rect 11109 2370 11121 2404
rect 11121 2370 11155 2404
rect 11155 2370 11167 2404
rect 12177 2370 12189 2404
rect 12189 2370 12223 2404
rect 12223 2370 12235 2404
rect 13245 2370 13257 2404
rect 13257 2370 13291 2404
rect 13291 2370 13303 2404
rect 11109 2352 11167 2370
rect 12177 2352 12235 2370
rect 13245 2352 13303 2370
rect 8956 2182 9014 2200
rect 8956 2148 8968 2182
rect 8968 2148 9002 2182
rect 9002 2148 9014 2182
rect 8956 2142 9014 2148
rect 9312 2182 9370 2200
rect 10024 2182 10082 2200
rect 9312 2148 9324 2182
rect 9324 2148 9358 2182
rect 9358 2148 9370 2182
rect 10024 2148 10036 2182
rect 10036 2148 10070 2182
rect 10070 2148 10082 2182
rect 9312 2142 9370 2148
rect 10024 2142 10082 2148
rect 11643 2182 11701 2200
rect 12355 2182 12413 2200
rect 11643 2148 11655 2182
rect 11655 2148 11689 2182
rect 11689 2148 11701 2182
rect 12355 2148 12367 2182
rect 12367 2148 12401 2182
rect 12401 2148 12413 2182
rect 11643 2142 11701 2148
rect 12355 2142 12413 2148
rect 12711 2182 12769 2200
rect 12711 2148 12723 2182
rect 12723 2148 12757 2182
rect 12757 2148 12769 2182
rect 14126 2204 14184 2210
rect 15550 2204 15608 2210
rect 16974 2204 17032 2210
rect 14126 2170 14138 2204
rect 14138 2170 14172 2204
rect 14172 2170 14184 2204
rect 15550 2170 15562 2204
rect 15562 2170 15596 2204
rect 15596 2170 15608 2204
rect 16974 2170 16986 2204
rect 16986 2170 17020 2204
rect 17020 2170 17032 2204
rect 14126 2152 14184 2170
rect 15550 2152 15608 2170
rect 16974 2152 17032 2170
rect 17526 2204 17584 2210
rect 18950 2204 19008 2210
rect 20374 2204 20432 2210
rect 17526 2170 17538 2204
rect 17538 2170 17572 2204
rect 17572 2170 17584 2204
rect 18950 2170 18962 2204
rect 18962 2170 18996 2204
rect 18996 2170 19008 2204
rect 20374 2170 20386 2204
rect 20386 2170 20420 2204
rect 20420 2170 20432 2204
rect 17526 2152 17584 2170
rect 18950 2152 19008 2170
rect 20374 2152 20432 2170
rect 12711 2142 12769 2148
rect 15016 1982 15074 2000
rect 16084 1982 16142 2000
rect 15016 1948 15028 1982
rect 15028 1948 15062 1982
rect 15062 1948 15074 1982
rect 16084 1948 16096 1982
rect 16096 1948 16130 1982
rect 16130 1948 16142 1982
rect 15016 1942 15074 1948
rect 16084 1942 16142 1948
rect 18416 1982 18474 2000
rect 19484 1982 19542 2000
rect 18416 1948 18428 1982
rect 18428 1948 18462 1982
rect 18462 1948 18474 1982
rect 19484 1948 19496 1982
rect 19496 1948 19530 1982
rect 19530 1948 19542 1982
rect 18416 1942 18474 1948
rect 19484 1942 19542 1948
rect 8422 1704 8480 1710
rect 8422 1670 8434 1704
rect 8434 1670 8468 1704
rect 8468 1670 8480 1704
rect 8422 1652 8480 1670
rect 9312 1652 9370 1710
rect 9490 1704 9548 1710
rect 10558 1704 10616 1710
rect 9490 1670 9502 1704
rect 9502 1670 9536 1704
rect 9536 1670 9548 1704
rect 10558 1670 10570 1704
rect 10570 1670 10604 1704
rect 10604 1670 10616 1704
rect 9490 1652 9548 1670
rect 10558 1652 10616 1670
rect 11109 1704 11167 1710
rect 12177 1704 12235 1710
rect 11109 1670 11121 1704
rect 11121 1670 11155 1704
rect 11155 1670 11167 1704
rect 12177 1670 12189 1704
rect 12189 1670 12223 1704
rect 12223 1670 12235 1704
rect 11109 1652 11167 1670
rect 12177 1652 12235 1670
rect 12355 1652 12413 1710
rect 13245 1704 13303 1710
rect 13245 1670 13257 1704
rect 13257 1670 13291 1704
rect 13291 1670 13303 1704
rect 13245 1652 13303 1670
rect 14126 1704 14184 1710
rect 15550 1704 15608 1710
rect 16974 1704 17032 1710
rect 14126 1670 14138 1704
rect 14138 1670 14172 1704
rect 14172 1670 14184 1704
rect 15550 1670 15562 1704
rect 15562 1670 15596 1704
rect 15596 1670 15608 1704
rect 16974 1670 16986 1704
rect 16986 1670 17020 1704
rect 17020 1670 17032 1704
rect 14126 1652 14184 1670
rect 15550 1652 15608 1670
rect 16974 1652 17032 1670
rect 17526 1704 17584 1710
rect 18950 1704 19008 1710
rect 20374 1704 20432 1710
rect 17526 1670 17538 1704
rect 17538 1670 17572 1704
rect 17572 1670 17584 1704
rect 18950 1670 18962 1704
rect 18962 1670 18996 1704
rect 18996 1670 19008 1704
rect 20374 1670 20386 1704
rect 20386 1670 20420 1704
rect 20420 1670 20432 1704
rect 17526 1652 17584 1670
rect 18950 1652 19008 1670
rect 20374 1652 20432 1670
rect 8956 1482 9014 1500
rect 10024 1482 10082 1500
rect 8956 1448 8968 1482
rect 8968 1448 9002 1482
rect 9002 1448 9014 1482
rect 10024 1448 10036 1482
rect 10036 1448 10070 1482
rect 10070 1448 10082 1482
rect 8956 1442 9014 1448
rect 10024 1442 10082 1448
rect 11643 1482 11701 1500
rect 12711 1482 12769 1500
rect 11643 1448 11655 1482
rect 11655 1448 11689 1482
rect 11689 1448 11701 1482
rect 12711 1448 12723 1482
rect 12723 1448 12757 1482
rect 12757 1448 12769 1482
rect 11643 1442 11701 1448
rect 12711 1442 12769 1448
rect 15016 1482 15074 1500
rect 16084 1482 16142 1500
rect 15016 1448 15028 1482
rect 15028 1448 15062 1482
rect 15062 1448 15074 1482
rect 16084 1448 16096 1482
rect 16096 1448 16130 1482
rect 16130 1448 16142 1482
rect 15016 1442 15074 1448
rect 16084 1442 16142 1448
rect 18416 1482 18474 1500
rect 19484 1482 19542 1500
rect 18416 1448 18428 1482
rect 18428 1448 18462 1482
rect 18462 1448 18474 1482
rect 19484 1448 19496 1482
rect 19496 1448 19530 1482
rect 19530 1448 19542 1482
rect 18416 1442 18474 1448
rect 19484 1442 19542 1448
rect 8422 1204 8480 1210
rect 9490 1204 9548 1210
rect 10558 1204 10616 1210
rect 8422 1170 8434 1204
rect 8434 1170 8468 1204
rect 8468 1170 8480 1204
rect 9490 1170 9502 1204
rect 9502 1170 9536 1204
rect 9536 1170 9548 1204
rect 10558 1170 10570 1204
rect 10570 1170 10604 1204
rect 10604 1170 10616 1204
rect 8422 1152 8480 1170
rect 9490 1152 9548 1170
rect 10558 1152 10616 1170
rect 11109 1204 11167 1210
rect 12177 1204 12235 1210
rect 13245 1204 13303 1210
rect 11109 1170 11121 1204
rect 11121 1170 11155 1204
rect 11155 1170 11167 1204
rect 12177 1170 12189 1204
rect 12189 1170 12223 1204
rect 12223 1170 12235 1204
rect 13245 1170 13257 1204
rect 13257 1170 13291 1204
rect 13291 1170 13303 1204
rect 11109 1152 11167 1170
rect 12177 1152 12235 1170
rect 13245 1152 13303 1170
rect 14126 1204 14184 1210
rect 15550 1204 15608 1210
rect 16974 1204 17032 1210
rect 14126 1170 14138 1204
rect 14138 1170 14172 1204
rect 14172 1170 14184 1204
rect 15550 1170 15562 1204
rect 15562 1170 15596 1204
rect 15596 1170 15608 1204
rect 16974 1170 16986 1204
rect 16986 1170 17020 1204
rect 17020 1170 17032 1204
rect 14126 1152 14184 1170
rect 15550 1152 15608 1170
rect 16974 1152 17032 1170
rect 17526 1204 17584 1210
rect 18950 1204 19008 1210
rect 20374 1204 20432 1210
rect 17526 1170 17538 1204
rect 17538 1170 17572 1204
rect 17572 1170 17584 1204
rect 18950 1170 18962 1204
rect 18962 1170 18996 1204
rect 18996 1170 19008 1204
rect 20374 1170 20386 1204
rect 20386 1170 20420 1204
rect 20420 1170 20432 1204
rect 17526 1152 17584 1170
rect 18950 1152 19008 1170
rect 20374 1152 20432 1170
rect 8956 982 9014 1000
rect 10024 982 10082 1000
rect 8956 948 8968 982
rect 8968 948 9002 982
rect 9002 948 9014 982
rect 10024 948 10036 982
rect 10036 948 10070 982
rect 10070 948 10082 982
rect 8956 942 9014 948
rect 10024 942 10082 948
rect 11643 982 11701 1000
rect 12711 982 12769 1000
rect 11643 948 11655 982
rect 11655 948 11689 982
rect 11689 948 11701 982
rect 12711 948 12723 982
rect 12723 948 12757 982
rect 12757 948 12769 982
rect 11643 942 11701 948
rect 12711 942 12769 948
rect 15016 982 15074 1000
rect 16084 982 16142 1000
rect 15016 948 15028 982
rect 15028 948 15062 982
rect 15062 948 15074 982
rect 16084 948 16096 982
rect 16096 948 16130 982
rect 16130 948 16142 982
rect 15016 942 15074 948
rect 16084 942 16142 948
rect 18416 982 18474 1000
rect 19484 982 19542 1000
rect 18416 948 18428 982
rect 18428 948 18462 982
rect 18462 948 18474 982
rect 19484 948 19496 982
rect 19496 948 19530 982
rect 19530 948 19542 982
rect 18416 942 18474 948
rect 19484 942 19542 948
rect 8422 704 8480 710
rect 9490 704 9548 710
rect 10558 704 10616 710
rect 8422 670 8434 704
rect 8434 670 8468 704
rect 8468 670 8480 704
rect 9490 670 9502 704
rect 9502 670 9536 704
rect 9536 670 9548 704
rect 10558 670 10570 704
rect 10570 670 10604 704
rect 10604 670 10616 704
rect 8422 652 8480 670
rect 9490 652 9548 670
rect 10558 652 10616 670
rect 11109 704 11167 710
rect 12177 704 12235 710
rect 13245 704 13303 710
rect 11109 670 11121 704
rect 11121 670 11155 704
rect 11155 670 11167 704
rect 12177 670 12189 704
rect 12189 670 12223 704
rect 12223 670 12235 704
rect 13245 670 13257 704
rect 13257 670 13291 704
rect 13291 670 13303 704
rect 11109 652 11167 670
rect 12177 652 12235 670
rect 13245 652 13303 670
rect 14126 704 14184 710
rect 15550 704 15608 710
rect 16974 704 17032 710
rect 14126 670 14138 704
rect 14138 670 14172 704
rect 14172 670 14184 704
rect 15550 670 15562 704
rect 15562 670 15596 704
rect 15596 670 15608 704
rect 16974 670 16986 704
rect 16986 670 17020 704
rect 17020 670 17032 704
rect 14126 652 14184 670
rect 15550 652 15608 670
rect 16974 652 17032 670
rect 17526 704 17584 710
rect 18950 704 19008 710
rect 20374 704 20432 710
rect 17526 670 17538 704
rect 17538 670 17572 704
rect 17572 670 17584 704
rect 18950 670 18962 704
rect 18962 670 18996 704
rect 18996 670 19008 704
rect 20374 670 20386 704
rect 20386 670 20420 704
rect 20420 670 20432 704
rect 17526 652 17584 670
rect 18950 652 19008 670
rect 20374 652 20432 670
rect 8956 482 9014 500
rect 10024 482 10082 500
rect 8956 448 8968 482
rect 8968 448 9002 482
rect 9002 448 9014 482
rect 10024 448 10036 482
rect 10036 448 10070 482
rect 10070 448 10082 482
rect 8956 442 9014 448
rect 10024 442 10082 448
rect 11643 482 11701 500
rect 12711 482 12769 500
rect 11643 448 11655 482
rect 11655 448 11689 482
rect 11689 448 11701 482
rect 12711 448 12723 482
rect 12723 448 12757 482
rect 12757 448 12769 482
rect 11643 442 11701 448
rect 12711 442 12769 448
rect 15016 482 15074 500
rect 16084 482 16142 500
rect 15016 448 15028 482
rect 15028 448 15062 482
rect 15062 448 15074 482
rect 16084 448 16096 482
rect 16096 448 16130 482
rect 16130 448 16142 482
rect 15016 442 15074 448
rect 16084 442 16142 448
rect 18416 482 18474 500
rect 19484 482 19542 500
rect 18416 448 18428 482
rect 18428 448 18462 482
rect 18462 448 18474 482
rect 19484 448 19496 482
rect 19496 448 19530 482
rect 19530 448 19542 482
rect 18416 442 18474 448
rect 19484 442 19542 448
<< metal2 >>
rect 8780 6269 8838 6279
rect 8084 5877 8572 5893
rect 8142 5819 8514 5877
rect 8084 5776 8572 5819
rect 8780 5691 8838 6211
rect 8780 5623 8838 5633
rect 8958 6058 9016 6546
rect 8958 5481 9016 6000
rect 10026 6058 10084 6544
rect 8958 5413 9016 5423
rect 9492 5691 9550 5701
rect 8780 4810 8838 4820
rect 8780 4240 8838 4752
rect 8780 4172 8838 4182
rect 8958 4600 9016 4610
rect 8958 4030 9016 4542
rect 9492 4600 9550 5633
rect 10026 5481 10084 6000
rect 10204 6262 10262 6272
rect 10204 5691 10262 6204
rect 11466 6268 11524 6278
rect 10471 5874 10529 5884
rect 11200 5874 11258 5884
rect 10529 5816 11200 5874
rect 10471 5806 10529 5816
rect 11200 5806 11258 5816
rect 10204 5623 10262 5633
rect 11466 5690 11524 6210
rect 11466 5622 11524 5632
rect 11644 6058 11702 6578
rect 10026 5413 10084 5423
rect 11644 5480 11702 6000
rect 12712 6058 12770 6573
rect 11644 5412 11702 5422
rect 12178 5690 12236 5700
rect 10560 4810 10618 4820
rect 9492 4532 9550 4542
rect 10382 4600 10440 4610
rect 8958 3962 9016 3972
rect 9490 4240 9548 4250
rect 8422 3410 8480 3420
rect 8422 2910 8480 3352
rect 9490 3410 9548 4182
rect 10382 4123 10440 4542
rect 10560 4240 10618 4752
rect 10560 4172 10618 4182
rect 11110 4810 11168 4820
rect 11110 4240 11168 4752
rect 11288 4600 11346 4610
rect 11288 4333 11346 4542
rect 12178 4600 12236 5632
rect 12712 5480 12770 6000
rect 12890 6263 12948 6273
rect 12890 5690 12948 6205
rect 12890 5622 12948 5632
rect 12712 5412 12770 5422
rect 12890 4810 12948 4820
rect 12178 4532 12236 4542
rect 12712 4600 12770 4610
rect 11281 4323 11354 4333
rect 11281 4240 11354 4250
rect 12178 4240 12236 4250
rect 11110 4172 11168 4182
rect 10382 4030 10440 4065
rect 10382 3962 10440 3972
rect 11288 4030 11346 4240
rect 11288 3962 11346 3972
rect 12178 3420 12236 4182
rect 12712 4030 12770 4542
rect 12890 4240 12948 4752
rect 12890 4172 12948 4182
rect 17503 4313 17561 4323
rect 16783 4120 16841 4130
rect 12712 3962 12770 3972
rect 16359 3986 16417 3996
rect 15878 3726 15936 3736
rect 8422 2410 8480 2852
rect 8422 2342 8480 2352
rect 8956 3200 9014 3210
rect 8956 2700 9014 3142
rect 8956 2200 9014 2642
rect 9490 2910 9548 3352
rect 10558 3410 10616 3420
rect 9490 2410 9548 2852
rect 9490 2342 9548 2352
rect 10024 3200 10082 3210
rect 10024 2700 10082 3142
rect 8956 2132 9014 2142
rect 9312 2200 9370 2210
rect 8422 1710 8480 1720
rect 8422 1210 8480 1652
rect 9312 1710 9370 2142
rect 10024 2200 10082 2642
rect 10558 2910 10616 3352
rect 10558 2410 10616 2852
rect 10558 2342 10616 2352
rect 11109 3410 11167 3420
rect 11109 2910 11167 3352
rect 12177 3410 12236 3420
rect 12235 3352 12236 3410
rect 12177 3301 12236 3352
rect 13245 3410 13303 3420
rect 11109 2410 11167 2852
rect 11109 2342 11167 2352
rect 11643 3200 11701 3210
rect 11643 2700 11701 3142
rect 10024 2132 10082 2142
rect 11643 2200 11701 2642
rect 12177 2910 12235 3301
rect 12177 2410 12235 2852
rect 12177 2342 12235 2352
rect 12711 3200 12769 3210
rect 12711 2700 12769 3142
rect 11643 2132 11701 2142
rect 12355 2200 12413 2210
rect 9312 1642 9370 1652
rect 9490 1710 9548 1720
rect 8422 710 8480 1152
rect 8422 642 8480 652
rect 8956 1500 9014 1510
rect 8956 1000 9014 1442
rect 8956 500 9014 942
rect 9490 1210 9548 1652
rect 10558 1710 10616 1720
rect 9490 710 9548 1152
rect 9490 642 9548 652
rect 10024 1500 10082 1510
rect 10024 1000 10082 1442
rect 8956 155 9014 442
rect 10024 500 10082 942
rect 10558 1210 10616 1652
rect 10558 710 10616 1152
rect 10558 642 10616 652
rect 11109 1710 11167 1720
rect 11109 1210 11167 1652
rect 12177 1710 12235 1720
rect 11109 710 11167 1152
rect 11109 642 11167 652
rect 11643 1500 11701 1510
rect 11643 1000 11701 1442
rect 10024 155 10082 442
rect 11643 500 11701 942
rect 12177 1210 12235 1652
rect 12355 1710 12413 2142
rect 12711 2200 12769 2642
rect 13245 2910 13303 3352
rect 13245 2410 13303 2852
rect 13245 2342 13303 2352
rect 14126 3210 14184 3220
rect 14126 2710 14184 3152
rect 15550 3210 15608 3220
rect 12711 2132 12769 2142
rect 14126 2210 14184 2652
rect 12355 1642 12413 1652
rect 13245 1710 13303 1720
rect 12177 710 12235 1152
rect 12177 642 12235 652
rect 12711 1500 12769 1510
rect 12711 1000 12769 1442
rect 11643 155 11701 442
rect 12711 500 12769 942
rect 13245 1210 13303 1652
rect 13245 710 13303 1152
rect 13245 642 13303 652
rect 14126 1710 14184 2152
rect 14126 1210 14184 1652
rect 14126 710 14184 1152
rect 14126 642 14184 652
rect 15016 3000 15074 3010
rect 15016 2501 15074 2942
rect 15016 2000 15074 2443
rect 15016 1500 15074 1942
rect 15016 1000 15074 1442
rect 12711 173 12769 442
rect 15016 500 15074 942
rect 15550 2710 15608 3152
rect 15878 3210 15936 3668
rect 16359 3626 16417 3928
rect 16783 3884 16841 4062
rect 16783 3816 16841 3826
rect 17503 3884 17561 4255
rect 17503 3816 17561 3826
rect 18139 3986 18197 3996
rect 16359 3558 16417 3568
rect 18139 3626 18197 3928
rect 18139 3558 18197 3568
rect 18718 3720 18776 3730
rect 15878 3142 15936 3152
rect 16974 3210 17032 3220
rect 15550 2210 15608 2652
rect 15550 1710 15608 2152
rect 15550 1210 15608 1652
rect 15550 710 15608 1152
rect 15550 642 15608 652
rect 16084 3000 16142 3010
rect 16084 2500 16142 2942
rect 16084 2000 16142 2442
rect 16084 1500 16142 1942
rect 16084 1000 16142 1442
rect 15016 135 15074 442
rect 16084 500 16142 942
rect 16974 2710 17032 3152
rect 16974 2210 17032 2652
rect 16974 1710 17032 2152
rect 16974 1210 17032 1652
rect 16974 710 17032 1152
rect 16974 642 17032 652
rect 17526 3210 17584 3220
rect 17526 2710 17584 3152
rect 18718 3210 18776 3662
rect 18718 3142 18776 3152
rect 18950 3210 19008 3220
rect 17526 2210 17584 2652
rect 17526 1710 17584 2152
rect 17526 1210 17584 1652
rect 17526 710 17584 1152
rect 17526 642 17584 652
rect 18416 3000 18474 3010
rect 18416 2500 18474 2942
rect 18416 2000 18474 2442
rect 18416 1500 18474 1942
rect 18416 1000 18474 1442
rect 16084 135 16142 442
rect 18416 500 18474 942
rect 18950 2710 19008 3152
rect 20374 3210 20432 3220
rect 18950 2210 19008 2652
rect 18950 1710 19008 2152
rect 18950 1210 19008 1652
rect 18950 710 19008 1152
rect 18950 642 19008 652
rect 19484 3000 19542 3010
rect 19484 2500 19542 2942
rect 19484 2000 19542 2442
rect 19484 1500 19542 1942
rect 19484 1000 19542 1442
rect 18416 135 18474 442
rect 19484 500 19542 942
rect 20374 2710 20432 3152
rect 20374 2210 20432 2652
rect 20374 1710 20432 2152
rect 20374 1210 20432 1652
rect 20374 710 20432 1152
rect 20374 642 20432 652
rect 19484 135 19542 442
<< via2 >>
rect 11281 4250 11354 4323
rect 10382 4065 10440 4123
rect 17503 4255 17561 4313
rect 16783 4062 16841 4120
<< metal3 >>
rect 11271 4323 11364 4328
rect 11271 4250 11281 4323
rect 11354 4313 17571 4323
rect 11354 4255 17503 4313
rect 17561 4255 17571 4313
rect 11354 4250 17571 4255
rect 11271 4245 11364 4250
rect 10367 4123 16851 4130
rect 10367 4065 10382 4123
rect 10440 4120 16851 4123
rect 10440 4065 16783 4120
rect 10367 4062 16783 4065
rect 16841 4062 16851 4120
rect 10367 4057 16851 4062
use bias_circuit  bias_circuit_0
timestamp 1654598202
transform 1 0 -215 0 1 276
box -400 -318 8604 6523
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_0
timestamp 1654558846
transform 1 0 9519 0 1 576
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_1
timestamp 1654558846
transform 1 0 9519 0 1 1076
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_2
timestamp 1654558846
transform 1 0 9519 0 1 1576
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_3
timestamp 1654558846
transform 1 0 12206 0 1 1576
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_4
timestamp 1654558846
transform 1 0 12206 0 1 1076
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_5
timestamp 1654558846
transform 1 0 12206 0 1 576
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_6
timestamp 1654558846
transform 1 0 9519 0 1 2276
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_7
timestamp 1654558846
transform 1 0 9519 0 1 2776
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_8
timestamp 1654558846
transform 1 0 9519 0 1 3276
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_9
timestamp 1654558846
transform 1 0 12206 0 1 3276
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_10
timestamp 1654558846
transform 1 0 12206 0 1 2776
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_11
timestamp 1654558846
transform 1 0 12206 0 1 2276
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_0
timestamp 1654557735
transform 1 0 15579 0 1 2576
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_1
timestamp 1654557735
transform 1 0 18979 0 1 576
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_2
timestamp 1654557735
transform 1 0 18979 0 1 1076
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_3
timestamp 1654557735
transform 1 0 18979 0 1 1576
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_4
timestamp 1654557735
transform 1 0 18979 0 1 2076
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_5
timestamp 1654557735
transform 1 0 18979 0 1 2576
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_6
timestamp 1654557735
transform 1 0 18979 0 1 3076
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_7
timestamp 1654557735
transform 1 0 15579 0 1 3076
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_8
timestamp 1654557735
transform 1 0 15579 0 1 2076
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_9
timestamp 1654557735
transform 1 0 15579 0 1 1576
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_10
timestamp 1654557735
transform 1 0 15579 0 1 1076
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_11
timestamp 1654557735
transform 1 0 15579 0 1 576
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_lvt_K7HVMB  sky130_fd_pr__nfet_01v8_lvt_K7HVMB_0
timestamp 1654599767
transform 1 0 16388 0 1 3776
box -820 -208 820 208
use sky130_fd_pr__nfet_01v8_lvt_K7HVMB  sky130_fd_pr__nfet_01v8_lvt_K7HVMB_1
timestamp 1654599767
transform 1 0 18168 0 1 3776
box -820 -208 820 208
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_0
timestamp 1654568132
transform 1 0 9699 0 1 4106
box -1133 -240 1133 240
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_1
timestamp 1654568132
transform 1 0 9699 0 1 4676
box -1133 -240 1133 240
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_2
timestamp 1654568132
transform 1 0 12029 0 1 4676
box -1133 -240 1133 240
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_3
timestamp 1654568132
transform 1 0 12029 0 1 4106
box -1133 -240 1133 240
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_0
timestamp 1654590681
transform 1 0 9521 0 1 5557
box -1311 -240 1311 240
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_1
timestamp 1654590681
transform 1 0 12207 0 1 5556
box -1311 -240 1311 240
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_2
timestamp 1654590681
transform 1 0 9521 0 1 6134
box -1311 -240 1311 240
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_3
timestamp 1654590681
transform 1 0 12207 0 1 6134
box -1311 -240 1311 240
<< labels >>
flabel metal1 20312 3483 20312 3483 1 FreeSans 800 0 0 0 cmc
flabel metal1 16281 4596 16281 4596 1 FreeSans 800 0 0 0 ip
flabel metal1 18061 4602 18061 4602 1 FreeSans 800 0 0 0 in
<< end >>
