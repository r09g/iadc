magic
tech sky130A
magscale 1 2
timestamp 1654583406
<< locali >>
rect 11189 76664 11223 76698
rect 11189 76592 11223 76630
rect 11189 76520 11223 76558
rect 11189 76448 11223 76486
rect 11189 76376 11223 76414
rect 11189 76304 11223 76342
rect 11189 76232 11223 76270
rect 11189 76160 11223 76198
rect 11189 76088 11223 76126
rect 11189 76016 11223 76054
rect 11189 75944 11223 75982
rect 11189 75872 11223 75910
rect 11189 75800 11223 75838
rect 11189 75728 11223 75766
rect 11189 75656 11223 75694
rect 11189 75584 11223 75622
rect 11189 75512 11223 75550
rect 11189 75440 11223 75478
rect 11189 75368 11223 75406
rect 11189 75296 11223 75334
rect 11189 75224 11223 75262
rect 11189 75152 11223 75190
rect 11189 75080 11223 75118
rect 11189 75008 11223 75046
rect 11189 74936 11223 74974
rect 11189 74864 11223 74902
rect 11189 74792 11223 74830
rect 11189 74720 11223 74758
rect 11189 74648 11223 74686
rect 11189 74576 11223 74614
rect 11189 74504 11223 74542
rect 11189 74432 11223 74470
rect 11189 74360 11223 74398
rect 11189 74288 11223 74326
rect 11189 74216 11223 74254
rect 11189 74144 11223 74182
rect 11189 74072 11223 74110
rect 11189 74000 11223 74038
rect 11189 73928 11223 73966
rect 11189 73856 11223 73894
rect 11189 73784 11223 73822
rect 11189 73712 11223 73750
rect 11189 73640 11223 73678
rect 11189 73568 11223 73606
rect 11189 73496 11223 73534
rect 11189 73428 11223 73462
rect 377 60746 477 60758
rect 377 60712 410 60746
rect 444 60712 477 60746
rect 377 60674 477 60712
rect 377 60640 410 60674
rect 444 60640 477 60674
rect 377 60602 477 60640
rect 377 60568 410 60602
rect 444 60568 477 60602
rect 377 60530 477 60568
rect 377 60496 410 60530
rect 444 60496 477 60530
rect 377 60458 477 60496
rect 377 60424 410 60458
rect 444 60424 477 60458
rect 377 60386 477 60424
rect 377 60352 410 60386
rect 444 60352 477 60386
rect 377 60314 477 60352
rect 377 60280 410 60314
rect 444 60280 477 60314
rect 377 60242 477 60280
rect 377 60208 410 60242
rect 444 60208 477 60242
rect 377 60170 477 60208
rect 377 60136 410 60170
rect 444 60136 477 60170
rect 377 60098 477 60136
rect 377 60064 410 60098
rect 444 60064 477 60098
rect 377 60026 477 60064
rect 377 59992 410 60026
rect 444 59992 477 60026
rect 377 59954 477 59992
rect 377 59920 410 59954
rect 444 59920 477 59954
rect 377 59882 477 59920
rect 377 59848 410 59882
rect 444 59848 477 59882
rect 377 59810 477 59848
rect 377 59776 410 59810
rect 444 59776 477 59810
rect 377 59738 477 59776
rect 377 59704 410 59738
rect 444 59704 477 59738
rect 377 59666 477 59704
rect 377 59632 410 59666
rect 444 59632 477 59666
rect 377 59594 477 59632
rect 377 59560 410 59594
rect 444 59560 477 59594
rect 377 59522 477 59560
rect 377 59488 410 59522
rect 444 59488 477 59522
rect 377 59450 477 59488
rect 377 59416 410 59450
rect 444 59416 477 59450
rect 377 59378 477 59416
rect 377 59344 410 59378
rect 444 59344 477 59378
rect 377 59306 477 59344
rect 377 59272 410 59306
rect 444 59272 477 59306
rect 377 59234 477 59272
rect 377 59200 410 59234
rect 444 59200 477 59234
rect 377 59162 477 59200
rect 377 59128 410 59162
rect 444 59128 477 59162
rect 377 59090 477 59128
rect 377 59056 410 59090
rect 444 59056 477 59090
rect 377 59018 477 59056
rect 377 58984 410 59018
rect 444 58984 477 59018
rect 377 58946 477 58984
rect 377 58912 410 58946
rect 444 58912 477 58946
rect 377 58874 477 58912
rect 377 58840 410 58874
rect 444 58840 477 58874
rect 377 58802 477 58840
rect 377 58768 410 58802
rect 444 58768 477 58802
rect 377 58730 477 58768
rect 377 58696 410 58730
rect 444 58696 477 58730
rect 377 58658 477 58696
rect 377 58624 410 58658
rect 444 58624 477 58658
rect 377 58586 477 58624
rect 377 58552 410 58586
rect 444 58552 477 58586
rect 377 58514 477 58552
rect 377 58480 410 58514
rect 444 58480 477 58514
rect 377 58442 477 58480
rect 377 58408 410 58442
rect 444 58408 477 58442
rect 377 58370 477 58408
rect 377 58336 410 58370
rect 444 58336 477 58370
rect 377 58298 477 58336
rect 377 58264 410 58298
rect 444 58264 477 58298
rect 377 58226 477 58264
rect 377 58192 410 58226
rect 444 58192 477 58226
rect 377 58154 477 58192
rect 377 58120 410 58154
rect 444 58120 477 58154
rect 377 58082 477 58120
rect 377 58048 410 58082
rect 444 58048 477 58082
rect 377 58010 477 58048
rect 377 57976 410 58010
rect 444 57976 477 58010
rect 377 57938 477 57976
rect 377 57904 410 57938
rect 444 57904 477 57938
rect 377 57866 477 57904
rect 377 57832 410 57866
rect 444 57832 477 57866
rect 377 57794 477 57832
rect 377 57760 410 57794
rect 444 57760 477 57794
rect 377 57722 477 57760
rect 377 57688 410 57722
rect 444 57688 477 57722
rect 377 57650 477 57688
rect 377 57616 410 57650
rect 444 57616 477 57650
rect 377 57578 477 57616
rect 377 57544 410 57578
rect 444 57544 477 57578
rect 377 57506 477 57544
rect 377 57472 410 57506
rect 444 57472 477 57506
rect 377 57434 477 57472
rect 377 57400 410 57434
rect 444 57400 477 57434
rect 377 57362 477 57400
rect 377 57328 410 57362
rect 444 57328 477 57362
rect 377 57290 477 57328
rect 377 57256 410 57290
rect 444 57256 477 57290
rect 377 57218 477 57256
rect 377 57184 410 57218
rect 444 57184 477 57218
rect 377 57146 477 57184
rect 377 57112 410 57146
rect 444 57112 477 57146
rect 377 57074 477 57112
rect 377 57040 410 57074
rect 444 57040 477 57074
rect 377 57002 477 57040
rect 377 56968 410 57002
rect 444 56968 477 57002
rect 377 56930 477 56968
rect 377 56896 410 56930
rect 444 56896 477 56930
rect 377 56858 477 56896
rect 377 56824 410 56858
rect 444 56824 477 56858
rect 377 56786 477 56824
rect 377 56752 410 56786
rect 444 56752 477 56786
rect 377 56714 477 56752
rect 377 56680 410 56714
rect 444 56680 477 56714
rect 377 56642 477 56680
rect 377 56608 410 56642
rect 444 56608 477 56642
rect 377 56570 477 56608
rect 377 56536 410 56570
rect 444 56536 477 56570
rect 377 56498 477 56536
rect 377 56464 410 56498
rect 444 56464 477 56498
rect 377 56426 477 56464
rect 377 56392 410 56426
rect 444 56392 477 56426
rect 377 56354 477 56392
rect 377 56320 410 56354
rect 444 56320 477 56354
rect 377 56282 477 56320
rect 377 56248 410 56282
rect 444 56248 477 56282
rect 377 56210 477 56248
rect 377 56176 410 56210
rect 444 56176 477 56210
rect 377 56138 477 56176
rect 377 56104 410 56138
rect 444 56104 477 56138
rect 377 56066 477 56104
rect 377 56032 410 56066
rect 444 56032 477 56066
rect 377 55994 477 56032
rect 377 55960 410 55994
rect 444 55960 477 55994
rect 377 55922 477 55960
rect 377 55888 410 55922
rect 444 55888 477 55922
rect 377 55850 477 55888
rect 377 55816 410 55850
rect 444 55816 477 55850
rect 377 55778 477 55816
rect 377 55744 410 55778
rect 444 55744 477 55778
rect 377 55706 477 55744
rect 377 55672 410 55706
rect 444 55672 477 55706
rect 377 55634 477 55672
rect 377 55600 410 55634
rect 444 55600 477 55634
rect 377 55562 477 55600
rect 377 55528 410 55562
rect 444 55528 477 55562
rect 377 55490 477 55528
rect 377 55456 410 55490
rect 444 55456 477 55490
rect 377 55418 477 55456
rect 377 55384 410 55418
rect 444 55384 477 55418
rect 377 55346 477 55384
rect 377 55312 410 55346
rect 444 55312 477 55346
rect 377 55274 477 55312
rect 377 55240 410 55274
rect 444 55240 477 55274
rect 377 55202 477 55240
rect 377 55168 410 55202
rect 444 55168 477 55202
rect 377 55130 477 55168
rect 377 55096 410 55130
rect 444 55096 477 55130
rect 377 55058 477 55096
rect 377 55024 410 55058
rect 444 55024 477 55058
rect 377 54986 477 55024
rect 377 54952 410 54986
rect 444 54952 477 54986
rect 377 54914 477 54952
rect 377 54880 410 54914
rect 444 54880 477 54914
rect 377 54842 477 54880
rect 377 54808 410 54842
rect 444 54808 477 54842
rect 377 54770 477 54808
rect 377 54736 410 54770
rect 444 54736 477 54770
rect 377 54698 477 54736
rect 377 54664 410 54698
rect 444 54664 477 54698
rect 377 54626 477 54664
rect 377 54592 410 54626
rect 444 54592 477 54626
rect 377 54554 477 54592
rect 377 54520 410 54554
rect 444 54520 477 54554
rect 377 54482 477 54520
rect 377 54448 410 54482
rect 444 54448 477 54482
rect 377 54410 477 54448
rect 377 54376 410 54410
rect 444 54376 477 54410
rect 377 54338 477 54376
rect 377 54304 410 54338
rect 444 54304 477 54338
rect 377 54266 477 54304
rect 377 54232 410 54266
rect 444 54232 477 54266
rect 377 54194 477 54232
rect 377 54160 410 54194
rect 444 54160 477 54194
rect 377 54122 477 54160
rect 377 54088 410 54122
rect 444 54088 477 54122
rect 377 54050 477 54088
rect 377 54016 410 54050
rect 444 54016 477 54050
rect 377 53978 477 54016
rect 377 53944 410 53978
rect 444 53944 477 53978
rect 377 53906 477 53944
rect 377 53872 410 53906
rect 444 53872 477 53906
rect 377 53834 477 53872
rect 377 53800 410 53834
rect 444 53800 477 53834
rect 377 53762 477 53800
rect 377 53728 410 53762
rect 444 53728 477 53762
rect 377 53690 477 53728
rect 377 53656 410 53690
rect 444 53656 477 53690
rect 377 53618 477 53656
rect 377 53584 410 53618
rect 444 53584 477 53618
rect 377 53546 477 53584
rect 377 53512 410 53546
rect 444 53512 477 53546
rect 377 53474 477 53512
rect 377 53440 410 53474
rect 444 53440 477 53474
rect 377 53402 477 53440
rect 377 53368 410 53402
rect 444 53368 477 53402
rect 377 53330 477 53368
rect 377 53296 410 53330
rect 444 53296 477 53330
rect 377 53258 477 53296
rect 377 53224 410 53258
rect 444 53224 477 53258
rect 377 53186 477 53224
rect 377 53152 410 53186
rect 444 53152 477 53186
rect 377 53140 477 53152
rect -5624 50988 -155 51018
rect -5624 50954 -5607 50988
rect -5573 50954 -5535 50988
rect -5501 50954 -5463 50988
rect -5429 50954 -5391 50988
rect -5357 50954 -5319 50988
rect -5285 50954 -5247 50988
rect -5213 50954 -5175 50988
rect -5141 50954 -5103 50988
rect -5069 50954 -5031 50988
rect -4997 50954 -4959 50988
rect -4925 50954 -4887 50988
rect -4853 50954 -4815 50988
rect -4781 50954 -4743 50988
rect -4709 50954 -4671 50988
rect -4637 50954 -4599 50988
rect -4565 50954 -4527 50988
rect -4493 50954 -4455 50988
rect -4421 50954 -4383 50988
rect -4349 50954 -4311 50988
rect -4277 50954 -4239 50988
rect -4205 50954 -4167 50988
rect -4133 50954 -4095 50988
rect -4061 50954 -4023 50988
rect -3989 50954 -3951 50988
rect -3917 50954 -3879 50988
rect -3845 50954 -3807 50988
rect -3773 50954 -3735 50988
rect -3701 50954 -3663 50988
rect -3629 50954 -3591 50988
rect -3557 50954 -3519 50988
rect -3485 50954 -3447 50988
rect -3413 50954 -3375 50988
rect -3341 50954 -3303 50988
rect -3269 50954 -3231 50988
rect -3197 50954 -3159 50988
rect -3125 50954 -3087 50988
rect -3053 50954 -3015 50988
rect -2981 50954 -2943 50988
rect -2909 50954 -2871 50988
rect -2837 50954 -2799 50988
rect -2765 50954 -2727 50988
rect -2693 50954 -2655 50988
rect -2621 50954 -2583 50988
rect -2549 50954 -2511 50988
rect -2477 50954 -2439 50988
rect -2405 50954 -2367 50988
rect -2333 50954 -2295 50988
rect -2261 50954 -2223 50988
rect -2189 50954 -2151 50988
rect -2117 50954 -2079 50988
rect -2045 50954 -2007 50988
rect -1973 50954 -1935 50988
rect -1901 50954 -1863 50988
rect -1829 50954 -1791 50988
rect -1757 50954 -1719 50988
rect -1685 50954 -1647 50988
rect -1613 50954 -1575 50988
rect -1541 50954 -1503 50988
rect -1469 50954 -1431 50988
rect -1397 50954 -1359 50988
rect -1325 50954 -1287 50988
rect -1253 50954 -1215 50988
rect -1181 50954 -1143 50988
rect -1109 50954 -1071 50988
rect -1037 50954 -999 50988
rect -965 50954 -927 50988
rect -893 50954 -855 50988
rect -821 50954 -783 50988
rect -749 50954 -711 50988
rect -677 50954 -639 50988
rect -605 50954 -567 50988
rect -533 50954 -495 50988
rect -461 50954 -423 50988
rect -389 50954 -351 50988
rect -317 50954 -279 50988
rect -245 50954 -207 50988
rect -173 50954 -155 50988
rect -5624 50925 -155 50954
rect -4 50713 89 50741
rect -4 50679 25 50713
rect 59 50679 89 50713
rect -4 50641 89 50679
rect -4 50607 25 50641
rect 59 50607 89 50641
rect -4 50569 89 50607
rect -4 50535 25 50569
rect 59 50535 89 50569
rect -4 50497 89 50535
rect -4 50463 25 50497
rect 59 50463 89 50497
rect -4 50425 89 50463
rect -4 50391 25 50425
rect 59 50391 89 50425
rect -4 50353 89 50391
rect -4 50319 25 50353
rect 59 50319 89 50353
rect -4 50281 89 50319
rect -4 50247 25 50281
rect 59 50247 89 50281
rect -4 50209 89 50247
rect -4 50175 25 50209
rect 59 50175 89 50209
rect -4 50137 89 50175
rect -4 50103 25 50137
rect 59 50103 89 50137
rect -4 50065 89 50103
rect -4 50031 25 50065
rect 59 50031 89 50065
rect -4 49993 89 50031
rect -4 49959 25 49993
rect 59 49959 89 49993
rect -4 49921 89 49959
rect -4 49887 25 49921
rect 59 49887 89 49921
rect -4 49849 89 49887
rect -4 49815 25 49849
rect 59 49815 89 49849
rect -4 49777 89 49815
rect -4 49743 25 49777
rect 59 49743 89 49777
rect -4 49705 89 49743
rect -4 49671 25 49705
rect 59 49671 89 49705
rect -4 49633 89 49671
rect -4 49599 25 49633
rect 59 49599 89 49633
rect -4 49561 89 49599
rect -4 49527 25 49561
rect 59 49527 89 49561
rect -4 49489 89 49527
rect -4 49455 25 49489
rect 59 49455 89 49489
rect -4 49417 89 49455
rect -26399 49398 -26176 49404
rect -26399 49364 -26377 49398
rect -26343 49364 -26305 49398
rect -26271 49364 -26233 49398
rect -26199 49364 -26176 49398
rect -26399 49359 -26176 49364
rect -4 49383 25 49417
rect 59 49383 89 49417
rect -4 49345 89 49383
rect -4 49311 25 49345
rect 59 49311 89 49345
rect -4 49273 89 49311
rect -4 49239 25 49273
rect 59 49239 89 49273
rect -4 49201 89 49239
rect -4 49167 25 49201
rect 59 49167 89 49201
rect -4 49129 89 49167
rect -4 49095 25 49129
rect 59 49095 89 49129
rect -4 49057 89 49095
rect -4 49023 25 49057
rect 59 49023 89 49057
rect -4 48985 89 49023
rect -4 48951 25 48985
rect 59 48951 89 48985
rect -4 48913 89 48951
rect -4 48879 25 48913
rect 59 48879 89 48913
rect -4 48841 89 48879
rect -4 48807 25 48841
rect 59 48807 89 48841
rect -4 48769 89 48807
rect -4 48735 25 48769
rect 59 48735 89 48769
rect -4 48697 89 48735
rect -4 48663 25 48697
rect 59 48663 89 48697
rect -4 48625 89 48663
rect -4 48591 25 48625
rect 59 48591 89 48625
rect -4 48553 89 48591
rect -4 48519 25 48553
rect 59 48519 89 48553
rect -4 48481 89 48519
rect -4 48447 25 48481
rect 59 48447 89 48481
rect -4 48409 89 48447
rect -4 48375 25 48409
rect 59 48375 89 48409
rect -4 48337 89 48375
rect -4 48303 25 48337
rect 59 48303 89 48337
rect -4 48265 89 48303
rect -4 48231 25 48265
rect 59 48231 89 48265
rect -4 48193 89 48231
rect -4 48159 25 48193
rect 59 48159 89 48193
rect -4 48121 89 48159
rect -4 48087 25 48121
rect 59 48087 89 48121
rect -4 48049 89 48087
rect -4 48015 25 48049
rect 59 48015 89 48049
rect -4 47977 89 48015
rect -4 47943 25 47977
rect 59 47943 89 47977
rect -4 47905 89 47943
rect -4 47871 25 47905
rect 59 47871 89 47905
rect -4 47833 89 47871
rect -4 47799 25 47833
rect 59 47799 89 47833
rect -4 47771 89 47799
rect 377 45785 477 45818
rect 377 45751 410 45785
rect 444 45751 477 45785
rect 377 45713 477 45751
rect 377 45679 410 45713
rect 444 45679 477 45713
rect 377 45641 477 45679
rect 377 45607 410 45641
rect 444 45607 477 45641
rect 377 45569 477 45607
rect 377 45535 410 45569
rect 444 45535 477 45569
rect 377 45497 477 45535
rect 377 45463 410 45497
rect 444 45463 477 45497
rect 377 45425 477 45463
rect 377 45391 410 45425
rect 444 45391 477 45425
rect 377 45353 477 45391
rect 377 45319 410 45353
rect 444 45319 477 45353
rect 377 45281 477 45319
rect 377 45247 410 45281
rect 444 45247 477 45281
rect 377 45209 477 45247
rect 377 45175 410 45209
rect 444 45175 477 45209
rect 377 45137 477 45175
rect 377 45103 410 45137
rect 444 45103 477 45137
rect 377 45065 477 45103
rect 377 45031 410 45065
rect 444 45031 477 45065
rect 377 44993 477 45031
rect 377 44959 410 44993
rect 444 44959 477 44993
rect 377 44921 477 44959
rect 377 44887 410 44921
rect 444 44887 477 44921
rect 377 44849 477 44887
rect 377 44815 410 44849
rect 444 44815 477 44849
rect 41808 44927 41842 44936
rect 41808 44855 41842 44893
rect 377 44777 477 44815
rect 377 44743 410 44777
rect 444 44743 477 44777
rect 41808 44783 41842 44821
rect 377 44705 477 44743
rect 377 44671 410 44705
rect 444 44671 477 44705
rect 41808 44711 41842 44749
rect 43003 44786 43038 44818
rect 43037 44752 43038 44786
rect 42537 44713 42539 44747
rect 42573 44713 42611 44747
rect 42645 44713 42683 44747
rect 42717 44713 42755 44747
rect 42789 44713 42827 44747
rect 42861 44713 42899 44747
rect 42933 44713 42936 44747
rect 43003 44714 43038 44752
rect 43253 44716 43277 44750
rect 43311 44716 43349 44750
rect 43383 44716 43408 44750
rect 377 44633 477 44671
rect 377 44599 410 44633
rect 444 44599 477 44633
rect 377 44561 477 44599
rect 41808 44639 41842 44677
rect 43037 44680 43038 44714
rect 43003 44648 43038 44680
rect 41808 44596 41842 44605
rect 377 44527 410 44561
rect 444 44527 477 44561
rect 377 44489 477 44527
rect 377 44455 410 44489
rect 444 44455 477 44489
rect 377 44417 477 44455
rect 377 44383 410 44417
rect 444 44383 477 44417
rect 377 44350 477 44383
rect 41808 43777 41842 43786
rect 41808 43705 41842 43743
rect 41808 43633 41842 43671
rect 41808 43561 41842 43599
rect 43003 43636 43038 43668
rect 43037 43602 43038 43636
rect 42537 43563 42539 43597
rect 42573 43563 42611 43597
rect 42645 43563 42683 43597
rect 42717 43563 42755 43597
rect 42789 43563 42827 43597
rect 42861 43563 42899 43597
rect 42933 43563 42936 43597
rect 43003 43564 43038 43602
rect 43253 43566 43277 43600
rect 43311 43566 43349 43600
rect 43383 43566 43408 43600
rect 41808 43489 41842 43527
rect 43037 43530 43038 43564
rect 43003 43498 43038 43530
rect 41808 43446 41842 43455
rect 377 41326 477 41343
rect 377 41292 410 41326
rect 444 41292 477 41326
rect 377 41254 477 41292
rect 377 41220 410 41254
rect 444 41220 477 41254
rect 377 41182 477 41220
rect 377 41148 410 41182
rect 444 41148 477 41182
rect 377 41110 477 41148
rect 41808 41237 41842 41246
rect 41808 41165 41842 41203
rect 377 41076 410 41110
rect 444 41076 477 41110
rect 41808 41093 41842 41131
rect 377 41038 477 41076
rect 377 41004 410 41038
rect 444 41004 477 41038
rect 41808 41021 41842 41059
rect 43003 41096 43038 41128
rect 43037 41062 43038 41096
rect 42537 41023 42539 41057
rect 42573 41023 42611 41057
rect 42645 41023 42683 41057
rect 42717 41023 42755 41057
rect 42789 41023 42827 41057
rect 42861 41023 42899 41057
rect 42933 41023 42936 41057
rect 43003 41024 43038 41062
rect 43253 41026 43277 41060
rect 43311 41026 43349 41060
rect 43383 41026 43408 41060
rect 377 40966 477 41004
rect 377 40932 410 40966
rect 444 40932 477 40966
rect 377 40894 477 40932
rect 41808 40949 41842 40987
rect 43037 40990 43038 41024
rect 43003 40958 43038 40990
rect 41808 40906 41842 40915
rect 377 40860 410 40894
rect 444 40860 477 40894
rect 377 40822 477 40860
rect 377 40788 410 40822
rect 444 40788 477 40822
rect 377 40750 477 40788
rect 377 40716 410 40750
rect 444 40716 477 40750
rect 377 40678 477 40716
rect 377 40644 410 40678
rect 444 40644 477 40678
rect 377 40606 477 40644
rect 377 40572 410 40606
rect 444 40572 477 40606
rect 377 40534 477 40572
rect 377 40500 410 40534
rect 444 40500 477 40534
rect 377 40462 477 40500
rect 377 40428 410 40462
rect 444 40428 477 40462
rect 377 40390 477 40428
rect 377 40356 410 40390
rect 444 40356 477 40390
rect 377 40318 477 40356
rect 377 40284 410 40318
rect 444 40284 477 40318
rect 377 40246 477 40284
rect 377 40212 410 40246
rect 444 40212 477 40246
rect 377 40174 477 40212
rect 377 40140 410 40174
rect 444 40140 477 40174
rect 377 40102 477 40140
rect 377 40068 410 40102
rect 444 40068 477 40102
rect 377 40051 477 40068
rect 41808 39967 41842 39976
rect 41808 39895 41842 39933
rect 41808 39823 41842 39861
rect -5637 39773 -168 39803
rect -5637 39739 -5620 39773
rect -5586 39739 -5548 39773
rect -5514 39739 -5476 39773
rect -5442 39739 -5404 39773
rect -5370 39739 -5332 39773
rect -5298 39739 -5260 39773
rect -5226 39739 -5188 39773
rect -5154 39739 -5116 39773
rect -5082 39739 -5044 39773
rect -5010 39739 -4972 39773
rect -4938 39739 -4900 39773
rect -4866 39739 -4828 39773
rect -4794 39739 -4756 39773
rect -4722 39739 -4684 39773
rect -4650 39739 -4612 39773
rect -4578 39739 -4540 39773
rect -4506 39739 -4468 39773
rect -4434 39739 -4396 39773
rect -4362 39739 -4324 39773
rect -4290 39739 -4252 39773
rect -4218 39739 -4180 39773
rect -4146 39739 -4108 39773
rect -4074 39739 -4036 39773
rect -4002 39739 -3964 39773
rect -3930 39739 -3892 39773
rect -3858 39739 -3820 39773
rect -3786 39739 -3748 39773
rect -3714 39739 -3676 39773
rect -3642 39739 -3604 39773
rect -3570 39739 -3532 39773
rect -3498 39739 -3460 39773
rect -3426 39739 -3388 39773
rect -3354 39739 -3316 39773
rect -3282 39739 -3244 39773
rect -3210 39739 -3172 39773
rect -3138 39739 -3100 39773
rect -3066 39739 -3028 39773
rect -2994 39739 -2956 39773
rect -2922 39739 -2884 39773
rect -2850 39739 -2812 39773
rect -2778 39739 -2740 39773
rect -2706 39739 -2668 39773
rect -2634 39739 -2596 39773
rect -2562 39739 -2524 39773
rect -2490 39739 -2452 39773
rect -2418 39739 -2380 39773
rect -2346 39739 -2308 39773
rect -2274 39739 -2236 39773
rect -2202 39739 -2164 39773
rect -2130 39739 -2092 39773
rect -2058 39739 -2020 39773
rect -1986 39739 -1948 39773
rect -1914 39739 -1876 39773
rect -1842 39739 -1804 39773
rect -1770 39739 -1732 39773
rect -1698 39739 -1660 39773
rect -1626 39739 -1588 39773
rect -1554 39739 -1516 39773
rect -1482 39739 -1444 39773
rect -1410 39739 -1372 39773
rect -1338 39739 -1300 39773
rect -1266 39739 -1228 39773
rect -1194 39739 -1156 39773
rect -1122 39739 -1084 39773
rect -1050 39739 -1012 39773
rect -978 39739 -940 39773
rect -906 39739 -868 39773
rect -834 39739 -796 39773
rect -762 39739 -724 39773
rect -690 39739 -652 39773
rect -618 39739 -580 39773
rect -546 39739 -508 39773
rect -474 39739 -436 39773
rect -402 39739 -364 39773
rect -330 39739 -292 39773
rect -258 39739 -220 39773
rect -186 39739 -168 39773
rect 41808 39751 41842 39789
rect 43003 39826 43038 39858
rect 43037 39792 43038 39826
rect 42537 39753 42539 39787
rect 42573 39753 42611 39787
rect 42645 39753 42683 39787
rect 42717 39753 42755 39787
rect 42789 39753 42827 39787
rect 42861 39753 42899 39787
rect 42933 39753 42936 39787
rect 43003 39754 43038 39792
rect 43253 39756 43277 39790
rect 43311 39756 43349 39790
rect 43383 39756 43408 39790
rect -5637 39710 -168 39739
rect 41808 39679 41842 39717
rect 43037 39720 43038 39754
rect 43003 39688 43038 39720
rect 41808 39636 41842 39645
rect -31795 39114 -31761 39132
rect -31795 39042 -31761 39080
rect -31795 38970 -31761 39008
rect -31795 38898 -31761 38936
rect -31795 38846 -31761 38864
rect -31795 38550 -31761 38576
rect -31795 38478 -31761 38516
rect -31795 38406 -31761 38444
rect -31795 38334 -31761 38372
rect -31795 38262 -31761 38300
rect -31795 38202 -31761 38228
rect 59 16117 152 16135
rect 59 16083 88 16117
rect 122 16083 152 16117
rect 59 16045 152 16083
rect 59 16011 88 16045
rect 122 16011 152 16045
rect 59 15973 152 16011
rect 59 15939 88 15973
rect 122 15939 152 15973
rect 59 15901 152 15939
rect 59 15867 88 15901
rect 122 15867 152 15901
rect 59 15829 152 15867
rect 59 15795 88 15829
rect 122 15795 152 15829
rect 59 15757 152 15795
rect 59 15723 88 15757
rect 122 15723 152 15757
rect 59 15685 152 15723
rect 59 15651 88 15685
rect 122 15651 152 15685
rect 59 15613 152 15651
rect 59 15579 88 15613
rect 122 15579 152 15613
rect 59 15541 152 15579
rect 59 15507 88 15541
rect 122 15507 152 15541
rect 59 15469 152 15507
rect 59 15435 88 15469
rect 122 15435 152 15469
rect 59 15397 152 15435
rect 59 15363 88 15397
rect 122 15363 152 15397
rect 59 15325 152 15363
rect 59 15291 88 15325
rect 122 15291 152 15325
rect 59 15253 152 15291
rect 59 15219 88 15253
rect 122 15219 152 15253
rect 59 15181 152 15219
rect 59 15147 88 15181
rect 122 15147 152 15181
rect 59 15109 152 15147
rect 59 15075 88 15109
rect 122 15075 152 15109
rect 59 15037 152 15075
rect 59 15003 88 15037
rect 122 15003 152 15037
rect 59 14965 152 15003
rect 59 14931 88 14965
rect 122 14931 152 14965
rect 59 14893 152 14931
rect 59 14859 88 14893
rect 122 14859 152 14893
rect 59 14821 152 14859
rect 59 14787 88 14821
rect 122 14787 152 14821
rect 59 14749 152 14787
rect 59 14715 88 14749
rect 122 14715 152 14749
rect 59 14677 152 14715
rect 59 14643 88 14677
rect 122 14643 152 14677
rect 59 14605 152 14643
rect 59 14571 88 14605
rect 122 14571 152 14605
rect 59 14533 152 14571
rect 59 14499 88 14533
rect 122 14499 152 14533
rect 59 14461 152 14499
rect 59 14427 88 14461
rect 122 14427 152 14461
rect 11274 16088 11303 16122
rect 11337 16088 11367 16122
rect 11274 16050 11367 16088
rect 11274 16016 11303 16050
rect 11337 16016 11367 16050
rect 11274 15978 11367 16016
rect 11274 15944 11303 15978
rect 11337 15944 11367 15978
rect 11274 15906 11367 15944
rect 11274 15872 11303 15906
rect 11337 15872 11367 15906
rect 11274 15834 11367 15872
rect 11274 15800 11303 15834
rect 11337 15800 11367 15834
rect 11274 15762 11367 15800
rect 11274 15728 11303 15762
rect 11337 15728 11367 15762
rect 11274 15690 11367 15728
rect 11274 15656 11303 15690
rect 11337 15656 11367 15690
rect 11274 15618 11367 15656
rect 11274 15584 11303 15618
rect 11337 15584 11367 15618
rect 11274 15546 11367 15584
rect 11274 15512 11303 15546
rect 11337 15512 11367 15546
rect 11274 15474 11367 15512
rect 11274 15440 11303 15474
rect 11337 15440 11367 15474
rect 11274 15402 11367 15440
rect 11274 15368 11303 15402
rect 11337 15368 11367 15402
rect 11274 15330 11367 15368
rect 11274 15296 11303 15330
rect 11337 15296 11367 15330
rect 11274 15258 11367 15296
rect 11274 15224 11303 15258
rect 11337 15224 11367 15258
rect 11274 15186 11367 15224
rect 11274 15152 11303 15186
rect 11337 15152 11367 15186
rect 11274 15114 11367 15152
rect 11274 15080 11303 15114
rect 11337 15080 11367 15114
rect 11274 15042 11367 15080
rect 11274 15008 11303 15042
rect 11337 15008 11367 15042
rect 11274 14970 11367 15008
rect 11274 14936 11303 14970
rect 11337 14936 11367 14970
rect 11274 14898 11367 14936
rect 11274 14864 11303 14898
rect 11337 14864 11367 14898
rect 11274 14826 11367 14864
rect 11274 14792 11303 14826
rect 11337 14792 11367 14826
rect 11274 14754 11367 14792
rect 11274 14720 11303 14754
rect 11337 14720 11367 14754
rect 11274 14682 11367 14720
rect 11274 14648 11303 14682
rect 11337 14648 11367 14682
rect 11274 14610 11367 14648
rect 11274 14576 11303 14610
rect 11337 14576 11367 14610
rect 11274 14538 11367 14576
rect 11274 14504 11303 14538
rect 11337 14504 11367 14538
rect 11274 14466 11367 14504
rect 11274 14432 11303 14466
rect 11337 14432 11367 14466
rect 59 14389 152 14427
rect 59 14355 88 14389
rect 122 14355 152 14389
rect 59 14317 152 14355
rect 59 14283 88 14317
rect 122 14283 152 14317
rect 59 14245 152 14283
rect 59 14211 88 14245
rect 122 14211 152 14245
rect 59 14173 152 14211
rect 59 14139 88 14173
rect 122 14139 152 14173
rect 59 14101 152 14139
rect 59 14067 88 14101
rect 122 14067 152 14101
rect 59 14029 152 14067
rect 59 13995 88 14029
rect 122 13995 152 14029
rect 59 13957 152 13995
rect 59 13923 88 13957
rect 122 13923 152 13957
rect 59 13885 152 13923
rect 59 13851 88 13885
rect 122 13851 152 13885
rect 59 13813 152 13851
rect 59 13779 88 13813
rect 122 13779 152 13813
rect 59 13741 152 13779
rect 59 13707 88 13741
rect 122 13707 152 13741
rect 59 13669 152 13707
rect 59 13635 88 13669
rect 122 13635 152 13669
rect 59 13597 152 13635
rect 59 13563 88 13597
rect 122 13563 152 13597
rect 59 13525 152 13563
rect 59 13491 88 13525
rect 122 13491 152 13525
rect 59 13453 152 13491
rect 59 13419 88 13453
rect 122 13419 152 13453
rect 59 13381 152 13419
rect 59 13347 88 13381
rect 122 13347 152 13381
rect 59 13309 152 13347
rect 59 13275 88 13309
rect 122 13275 152 13309
rect 59 13237 152 13275
rect 59 13203 88 13237
rect 122 13203 152 13237
rect 59 13165 152 13203
rect 59 13131 88 13165
rect 122 13131 152 13165
rect 59 13093 152 13131
rect 59 13059 88 13093
rect 122 13059 152 13093
rect 59 13021 152 13059
rect 59 12987 88 13021
rect 122 12987 152 13021
rect 11274 13920 11367 13953
rect 11274 13886 11303 13920
rect 11337 13886 11367 13920
rect 11274 13848 11367 13886
rect 11274 13814 11303 13848
rect 11337 13814 11367 13848
rect 11274 13776 11367 13814
rect 11274 13742 11303 13776
rect 11337 13742 11367 13776
rect 11274 13704 11367 13742
rect 11274 13670 11303 13704
rect 11337 13670 11367 13704
rect 11274 13632 11367 13670
rect 11274 13598 11303 13632
rect 11337 13598 11367 13632
rect 11274 13560 11367 13598
rect 11274 13526 11303 13560
rect 11337 13526 11367 13560
rect 11274 13488 11367 13526
rect 11274 13454 11303 13488
rect 11337 13454 11367 13488
rect 11274 13416 11367 13454
rect 11274 13382 11303 13416
rect 11337 13382 11367 13416
rect 11274 13344 11367 13382
rect 11274 13310 11303 13344
rect 11337 13310 11367 13344
rect 11274 13272 11367 13310
rect 11274 13238 11303 13272
rect 11337 13238 11367 13272
rect 11274 13200 11367 13238
rect 11274 13166 11303 13200
rect 11337 13166 11367 13200
rect 11274 13128 11367 13166
rect 11274 13094 11303 13128
rect 11337 13094 11367 13128
rect 11274 13056 11367 13094
rect 11274 13022 11303 13056
rect 11337 13022 11367 13056
rect 11274 12989 11367 13022
rect 59 12949 152 12987
rect 59 12915 88 12949
rect 122 12915 152 12949
rect 59 12877 152 12915
rect 59 12843 88 12877
rect 122 12843 152 12877
rect 59 12805 152 12843
rect 59 12771 88 12805
rect 122 12771 152 12805
rect 59 12733 152 12771
rect 59 12699 88 12733
rect 122 12699 152 12733
rect 59 12661 152 12699
rect 59 12627 88 12661
rect 122 12627 152 12661
rect 59 12589 152 12627
rect 59 12555 88 12589
rect 122 12555 152 12589
rect 59 12517 152 12555
rect 59 12483 88 12517
rect 122 12483 152 12517
rect 59 12445 152 12483
rect 59 12411 88 12445
rect 122 12411 152 12445
rect 59 12373 152 12411
rect 59 12339 88 12373
rect 122 12339 152 12373
rect 59 12301 152 12339
rect 59 12267 88 12301
rect 122 12267 152 12301
rect 59 12229 152 12267
rect 59 12195 88 12229
rect 122 12195 152 12229
rect 59 12157 152 12195
rect 59 12123 88 12157
rect 122 12123 152 12157
rect 59 12085 152 12123
rect 59 12051 88 12085
rect 122 12051 152 12085
rect 59 12013 152 12051
rect 59 11979 88 12013
rect 122 11979 152 12013
rect 59 11941 152 11979
rect 59 11907 88 11941
rect 122 11907 152 11941
rect 59 11869 152 11907
rect 59 11835 88 11869
rect 122 11835 152 11869
rect 59 11797 152 11835
rect 59 11763 88 11797
rect 122 11763 152 11797
rect 59 11725 152 11763
rect 59 11691 88 11725
rect 122 11691 152 11725
rect 59 11653 152 11691
rect 59 11619 88 11653
rect 122 11619 152 11653
rect 59 11581 152 11619
rect 59 11547 88 11581
rect 122 11547 152 11581
rect 59 11509 152 11547
rect 59 11475 88 11509
rect 122 11475 152 11509
rect 59 11437 152 11475
rect 59 11403 88 11437
rect 122 11403 152 11437
rect 59 11365 152 11403
rect 59 11331 88 11365
rect 122 11331 152 11365
rect 59 11293 152 11331
rect 11274 12091 11367 12105
rect 11274 12057 11303 12091
rect 11337 12057 11367 12091
rect 11274 12019 11367 12057
rect 11274 11985 11303 12019
rect 11337 11985 11367 12019
rect 11274 11947 11367 11985
rect 11274 11913 11303 11947
rect 11337 11913 11367 11947
rect 11274 11875 11367 11913
rect 11274 11841 11303 11875
rect 11337 11841 11367 11875
rect 11274 11803 11367 11841
rect 11274 11769 11303 11803
rect 11337 11769 11367 11803
rect 11274 11731 11367 11769
rect 11274 11697 11303 11731
rect 11337 11697 11367 11731
rect 11274 11659 11367 11697
rect 11274 11625 11303 11659
rect 11337 11625 11367 11659
rect 11274 11587 11367 11625
rect 11274 11553 11303 11587
rect 11337 11553 11367 11587
rect 11274 11515 11367 11553
rect 11274 11481 11303 11515
rect 11337 11481 11367 11515
rect 11274 11443 11367 11481
rect 11274 11409 11303 11443
rect 11337 11409 11367 11443
rect 11274 11371 11367 11409
rect 11274 11337 11303 11371
rect 11337 11337 11367 11371
rect 11274 11323 11367 11337
rect 59 11259 88 11293
rect 122 11259 152 11293
rect 59 11221 152 11259
rect 59 11187 88 11221
rect 122 11187 152 11221
rect 59 11149 152 11187
rect 59 11115 88 11149
rect 122 11115 152 11149
rect 59 11077 152 11115
rect 59 11043 88 11077
rect 122 11043 152 11077
rect 59 11005 152 11043
rect 59 10971 88 11005
rect 122 10971 152 11005
rect 59 10933 152 10971
rect 59 10899 88 10933
rect 122 10899 152 10933
rect 59 10861 152 10899
rect 59 10827 88 10861
rect 122 10827 152 10861
rect 59 10789 152 10827
rect 59 10755 88 10789
rect 122 10755 152 10789
rect 59 10717 152 10755
rect 59 10683 88 10717
rect 122 10683 152 10717
rect 59 10666 152 10683
rect 6553 10472 11090 10502
rect 6553 10438 6572 10472
rect 6606 10438 6644 10472
rect 6678 10438 6716 10472
rect 6750 10438 6788 10472
rect 6822 10438 6860 10472
rect 6894 10438 6932 10472
rect 6966 10438 7004 10472
rect 7038 10438 7076 10472
rect 7110 10438 7148 10472
rect 7182 10438 7220 10472
rect 7254 10438 7292 10472
rect 7326 10438 7364 10472
rect 7398 10438 7436 10472
rect 7470 10438 7508 10472
rect 7542 10438 7580 10472
rect 7614 10438 7652 10472
rect 7686 10438 7724 10472
rect 7758 10438 7796 10472
rect 7830 10438 7868 10472
rect 7902 10438 7940 10472
rect 7974 10438 8012 10472
rect 8046 10438 8084 10472
rect 8118 10438 8156 10472
rect 8190 10438 8228 10472
rect 8262 10438 8300 10472
rect 8334 10438 8372 10472
rect 8406 10438 8444 10472
rect 8478 10438 8516 10472
rect 8550 10438 8588 10472
rect 8622 10438 8660 10472
rect 8694 10438 8732 10472
rect 8766 10438 8804 10472
rect 8838 10438 8876 10472
rect 8910 10438 8948 10472
rect 8982 10438 9020 10472
rect 9054 10438 9092 10472
rect 9126 10438 9164 10472
rect 9198 10438 9236 10472
rect 9270 10438 9308 10472
rect 9342 10438 9380 10472
rect 9414 10438 9452 10472
rect 9486 10438 9524 10472
rect 9558 10438 9596 10472
rect 9630 10438 9668 10472
rect 9702 10438 9740 10472
rect 9774 10438 9812 10472
rect 9846 10438 9884 10472
rect 9918 10438 9956 10472
rect 9990 10438 10028 10472
rect 10062 10438 10100 10472
rect 10134 10438 10172 10472
rect 10206 10438 10244 10472
rect 10278 10438 10316 10472
rect 10350 10438 10388 10472
rect 10422 10438 10460 10472
rect 10494 10438 10532 10472
rect 10566 10438 10604 10472
rect 10638 10438 10676 10472
rect 10710 10438 10748 10472
rect 10782 10438 10820 10472
rect 10854 10438 10892 10472
rect 10926 10438 10964 10472
rect 10998 10438 11036 10472
rect 11070 10438 11090 10472
rect 6553 10409 11090 10438
<< viali >>
rect 11189 76630 11223 76664
rect 11189 76558 11223 76592
rect 11189 76486 11223 76520
rect 11189 76414 11223 76448
rect 11189 76342 11223 76376
rect 11189 76270 11223 76304
rect 11189 76198 11223 76232
rect 11189 76126 11223 76160
rect 11189 76054 11223 76088
rect 11189 75982 11223 76016
rect 11189 75910 11223 75944
rect 11189 75838 11223 75872
rect 11189 75766 11223 75800
rect 11189 75694 11223 75728
rect 11189 75622 11223 75656
rect 11189 75550 11223 75584
rect 11189 75478 11223 75512
rect 11189 75406 11223 75440
rect 11189 75334 11223 75368
rect 11189 75262 11223 75296
rect 11189 75190 11223 75224
rect 11189 75118 11223 75152
rect 11189 75046 11223 75080
rect 11189 74974 11223 75008
rect 11189 74902 11223 74936
rect 11189 74830 11223 74864
rect 11189 74758 11223 74792
rect 11189 74686 11223 74720
rect 11189 74614 11223 74648
rect 11189 74542 11223 74576
rect 11189 74470 11223 74504
rect 11189 74398 11223 74432
rect 11189 74326 11223 74360
rect 11189 74254 11223 74288
rect 11189 74182 11223 74216
rect 11189 74110 11223 74144
rect 11189 74038 11223 74072
rect 11189 73966 11223 74000
rect 11189 73894 11223 73928
rect 11189 73822 11223 73856
rect 11189 73750 11223 73784
rect 11189 73678 11223 73712
rect 11189 73606 11223 73640
rect 11189 73534 11223 73568
rect 11189 73462 11223 73496
rect 410 60712 444 60746
rect 410 60640 444 60674
rect 410 60568 444 60602
rect 410 60496 444 60530
rect 410 60424 444 60458
rect 410 60352 444 60386
rect 410 60280 444 60314
rect 410 60208 444 60242
rect 410 60136 444 60170
rect 410 60064 444 60098
rect 410 59992 444 60026
rect 410 59920 444 59954
rect 410 59848 444 59882
rect 410 59776 444 59810
rect 410 59704 444 59738
rect 410 59632 444 59666
rect 410 59560 444 59594
rect 410 59488 444 59522
rect 410 59416 444 59450
rect 410 59344 444 59378
rect 410 59272 444 59306
rect 410 59200 444 59234
rect 410 59128 444 59162
rect 410 59056 444 59090
rect 410 58984 444 59018
rect 410 58912 444 58946
rect 410 58840 444 58874
rect 410 58768 444 58802
rect 410 58696 444 58730
rect 410 58624 444 58658
rect 410 58552 444 58586
rect 410 58480 444 58514
rect 410 58408 444 58442
rect 410 58336 444 58370
rect 410 58264 444 58298
rect 410 58192 444 58226
rect 410 58120 444 58154
rect 410 58048 444 58082
rect 410 57976 444 58010
rect 410 57904 444 57938
rect 410 57832 444 57866
rect 410 57760 444 57794
rect 410 57688 444 57722
rect 410 57616 444 57650
rect 410 57544 444 57578
rect 410 57472 444 57506
rect 410 57400 444 57434
rect 410 57328 444 57362
rect 410 57256 444 57290
rect 410 57184 444 57218
rect 410 57112 444 57146
rect 410 57040 444 57074
rect 410 56968 444 57002
rect 410 56896 444 56930
rect 410 56824 444 56858
rect 410 56752 444 56786
rect 410 56680 444 56714
rect 410 56608 444 56642
rect 410 56536 444 56570
rect 410 56464 444 56498
rect 410 56392 444 56426
rect 410 56320 444 56354
rect 410 56248 444 56282
rect 410 56176 444 56210
rect 410 56104 444 56138
rect 410 56032 444 56066
rect 410 55960 444 55994
rect 410 55888 444 55922
rect 410 55816 444 55850
rect 410 55744 444 55778
rect 410 55672 444 55706
rect 410 55600 444 55634
rect 410 55528 444 55562
rect 410 55456 444 55490
rect 410 55384 444 55418
rect 410 55312 444 55346
rect 410 55240 444 55274
rect 410 55168 444 55202
rect 410 55096 444 55130
rect 410 55024 444 55058
rect 410 54952 444 54986
rect 410 54880 444 54914
rect 410 54808 444 54842
rect 410 54736 444 54770
rect 410 54664 444 54698
rect 410 54592 444 54626
rect 410 54520 444 54554
rect 410 54448 444 54482
rect 410 54376 444 54410
rect 410 54304 444 54338
rect 410 54232 444 54266
rect 410 54160 444 54194
rect 410 54088 444 54122
rect 410 54016 444 54050
rect 410 53944 444 53978
rect 410 53872 444 53906
rect 410 53800 444 53834
rect 410 53728 444 53762
rect 410 53656 444 53690
rect 410 53584 444 53618
rect 410 53512 444 53546
rect 410 53440 444 53474
rect 410 53368 444 53402
rect 410 53296 444 53330
rect 410 53224 444 53258
rect 410 53152 444 53186
rect -5607 50954 -5573 50988
rect -5535 50954 -5501 50988
rect -5463 50954 -5429 50988
rect -5391 50954 -5357 50988
rect -5319 50954 -5285 50988
rect -5247 50954 -5213 50988
rect -5175 50954 -5141 50988
rect -5103 50954 -5069 50988
rect -5031 50954 -4997 50988
rect -4959 50954 -4925 50988
rect -4887 50954 -4853 50988
rect -4815 50954 -4781 50988
rect -4743 50954 -4709 50988
rect -4671 50954 -4637 50988
rect -4599 50954 -4565 50988
rect -4527 50954 -4493 50988
rect -4455 50954 -4421 50988
rect -4383 50954 -4349 50988
rect -4311 50954 -4277 50988
rect -4239 50954 -4205 50988
rect -4167 50954 -4133 50988
rect -4095 50954 -4061 50988
rect -4023 50954 -3989 50988
rect -3951 50954 -3917 50988
rect -3879 50954 -3845 50988
rect -3807 50954 -3773 50988
rect -3735 50954 -3701 50988
rect -3663 50954 -3629 50988
rect -3591 50954 -3557 50988
rect -3519 50954 -3485 50988
rect -3447 50954 -3413 50988
rect -3375 50954 -3341 50988
rect -3303 50954 -3269 50988
rect -3231 50954 -3197 50988
rect -3159 50954 -3125 50988
rect -3087 50954 -3053 50988
rect -3015 50954 -2981 50988
rect -2943 50954 -2909 50988
rect -2871 50954 -2837 50988
rect -2799 50954 -2765 50988
rect -2727 50954 -2693 50988
rect -2655 50954 -2621 50988
rect -2583 50954 -2549 50988
rect -2511 50954 -2477 50988
rect -2439 50954 -2405 50988
rect -2367 50954 -2333 50988
rect -2295 50954 -2261 50988
rect -2223 50954 -2189 50988
rect -2151 50954 -2117 50988
rect -2079 50954 -2045 50988
rect -2007 50954 -1973 50988
rect -1935 50954 -1901 50988
rect -1863 50954 -1829 50988
rect -1791 50954 -1757 50988
rect -1719 50954 -1685 50988
rect -1647 50954 -1613 50988
rect -1575 50954 -1541 50988
rect -1503 50954 -1469 50988
rect -1431 50954 -1397 50988
rect -1359 50954 -1325 50988
rect -1287 50954 -1253 50988
rect -1215 50954 -1181 50988
rect -1143 50954 -1109 50988
rect -1071 50954 -1037 50988
rect -999 50954 -965 50988
rect -927 50954 -893 50988
rect -855 50954 -821 50988
rect -783 50954 -749 50988
rect -711 50954 -677 50988
rect -639 50954 -605 50988
rect -567 50954 -533 50988
rect -495 50954 -461 50988
rect -423 50954 -389 50988
rect -351 50954 -317 50988
rect -279 50954 -245 50988
rect -207 50954 -173 50988
rect 25 50679 59 50713
rect 25 50607 59 50641
rect 25 50535 59 50569
rect 25 50463 59 50497
rect 25 50391 59 50425
rect 25 50319 59 50353
rect 25 50247 59 50281
rect 25 50175 59 50209
rect 25 50103 59 50137
rect 25 50031 59 50065
rect 25 49959 59 49993
rect 25 49887 59 49921
rect 25 49815 59 49849
rect 25 49743 59 49777
rect 25 49671 59 49705
rect 25 49599 59 49633
rect 25 49527 59 49561
rect 25 49455 59 49489
rect -26047 49413 -26013 49447
rect -26377 49364 -26343 49398
rect -26305 49364 -26271 49398
rect -26233 49364 -26199 49398
rect 25 49383 59 49417
rect -26047 49327 -26013 49361
rect 25 49311 59 49345
rect 25 49239 59 49273
rect 25 49167 59 49201
rect 25 49095 59 49129
rect 25 49023 59 49057
rect 25 48951 59 48985
rect 25 48879 59 48913
rect 25 48807 59 48841
rect 25 48735 59 48769
rect 25 48663 59 48697
rect 25 48591 59 48625
rect 25 48519 59 48553
rect 25 48447 59 48481
rect 25 48375 59 48409
rect 25 48303 59 48337
rect 25 48231 59 48265
rect 25 48159 59 48193
rect 25 48087 59 48121
rect 25 48015 59 48049
rect 25 47943 59 47977
rect 25 47871 59 47905
rect 25 47799 59 47833
rect 410 45751 444 45785
rect 410 45679 444 45713
rect 410 45607 444 45641
rect 410 45535 444 45569
rect 410 45463 444 45497
rect 410 45391 444 45425
rect 410 45319 444 45353
rect 410 45247 444 45281
rect 410 45175 444 45209
rect 410 45103 444 45137
rect 410 45031 444 45065
rect 410 44959 444 44993
rect 410 44887 444 44921
rect 410 44815 444 44849
rect 41808 44893 41842 44927
rect 41808 44821 41842 44855
rect 39984 44783 40018 44817
rect 40603 44782 40637 44816
rect 410 44743 444 44777
rect 41005 44776 41039 44810
rect 41161 44782 41195 44816
rect 410 44671 444 44705
rect 40128 44702 40162 44736
rect 40905 44717 40939 44751
rect 41808 44749 41842 44783
rect 43281 44802 43315 44836
rect 43453 44802 43487 44836
rect 43625 44802 43659 44836
rect 43797 44802 43831 44836
rect 43969 44802 44003 44836
rect 44174 44802 44208 44836
rect 44351 44802 44385 44836
rect 44523 44802 44557 44836
rect 44695 44802 44729 44836
rect 44867 44802 44901 44836
rect 45039 44802 45073 44836
rect 45211 44802 45245 44836
rect 43003 44752 43037 44786
rect 42539 44713 42573 44747
rect 42611 44713 42645 44747
rect 42683 44713 42717 44747
rect 42755 44713 42789 44747
rect 42827 44713 42861 44747
rect 42899 44713 42933 44747
rect 43277 44716 43311 44750
rect 43349 44716 43383 44750
rect 410 44599 444 44633
rect 41808 44677 41842 44711
rect 43003 44680 43037 44714
rect 41808 44605 41842 44639
rect 410 44527 444 44561
rect 410 44455 444 44489
rect 410 44383 444 44417
rect 41808 43743 41842 43777
rect 41808 43671 41842 43705
rect 39984 43633 40018 43667
rect 40603 43632 40637 43666
rect 41005 43626 41039 43660
rect 41161 43632 41195 43666
rect 40128 43552 40162 43586
rect 40905 43567 40939 43601
rect 41808 43599 41842 43633
rect 43281 43652 43315 43686
rect 43453 43652 43487 43686
rect 43625 43652 43659 43686
rect 43797 43652 43831 43686
rect 43969 43652 44003 43686
rect 44174 43652 44208 43686
rect 44351 43652 44385 43686
rect 44523 43652 44557 43686
rect 44695 43652 44729 43686
rect 44867 43652 44901 43686
rect 45039 43652 45073 43686
rect 45211 43652 45245 43686
rect 43003 43602 43037 43636
rect 42539 43563 42573 43597
rect 42611 43563 42645 43597
rect 42683 43563 42717 43597
rect 42755 43563 42789 43597
rect 42827 43563 42861 43597
rect 42899 43563 42933 43597
rect 43277 43566 43311 43600
rect 43349 43566 43383 43600
rect 41808 43527 41842 43561
rect 43003 43530 43037 43564
rect 41808 43455 41842 43489
rect 410 41292 444 41326
rect 410 41220 444 41254
rect 410 41148 444 41182
rect 41808 41203 41842 41237
rect 41808 41131 41842 41165
rect 410 41076 444 41110
rect 39984 41093 40018 41127
rect 40603 41092 40637 41126
rect 41005 41086 41039 41120
rect 41161 41092 41195 41126
rect 410 41004 444 41038
rect 40128 41012 40162 41046
rect 40905 41027 40939 41061
rect 41808 41059 41842 41093
rect 43281 41112 43315 41146
rect 43453 41112 43487 41146
rect 43625 41112 43659 41146
rect 43797 41112 43831 41146
rect 43969 41112 44003 41146
rect 44174 41112 44208 41146
rect 44351 41112 44385 41146
rect 44523 41112 44557 41146
rect 44695 41112 44729 41146
rect 44867 41112 44901 41146
rect 45039 41112 45073 41146
rect 45211 41112 45245 41146
rect 43003 41062 43037 41096
rect 42539 41023 42573 41057
rect 42611 41023 42645 41057
rect 42683 41023 42717 41057
rect 42755 41023 42789 41057
rect 42827 41023 42861 41057
rect 42899 41023 42933 41057
rect 43277 41026 43311 41060
rect 43349 41026 43383 41060
rect 410 40932 444 40966
rect 41808 40987 41842 41021
rect 43003 40990 43037 41024
rect 41808 40915 41842 40949
rect 410 40860 444 40894
rect 410 40788 444 40822
rect 410 40716 444 40750
rect 410 40644 444 40678
rect 410 40572 444 40606
rect 410 40500 444 40534
rect 410 40428 444 40462
rect 410 40356 444 40390
rect 410 40284 444 40318
rect 410 40212 444 40246
rect 410 40140 444 40174
rect 410 40068 444 40102
rect 41808 39933 41842 39967
rect 41808 39861 41842 39895
rect 39984 39823 40018 39857
rect 40603 39822 40637 39856
rect 41005 39816 41039 39850
rect 41161 39822 41195 39856
rect -5620 39739 -5586 39773
rect -5548 39739 -5514 39773
rect -5476 39739 -5442 39773
rect -5404 39739 -5370 39773
rect -5332 39739 -5298 39773
rect -5260 39739 -5226 39773
rect -5188 39739 -5154 39773
rect -5116 39739 -5082 39773
rect -5044 39739 -5010 39773
rect -4972 39739 -4938 39773
rect -4900 39739 -4866 39773
rect -4828 39739 -4794 39773
rect -4756 39739 -4722 39773
rect -4684 39739 -4650 39773
rect -4612 39739 -4578 39773
rect -4540 39739 -4506 39773
rect -4468 39739 -4434 39773
rect -4396 39739 -4362 39773
rect -4324 39739 -4290 39773
rect -4252 39739 -4218 39773
rect -4180 39739 -4146 39773
rect -4108 39739 -4074 39773
rect -4036 39739 -4002 39773
rect -3964 39739 -3930 39773
rect -3892 39739 -3858 39773
rect -3820 39739 -3786 39773
rect -3748 39739 -3714 39773
rect -3676 39739 -3642 39773
rect -3604 39739 -3570 39773
rect -3532 39739 -3498 39773
rect -3460 39739 -3426 39773
rect -3388 39739 -3354 39773
rect -3316 39739 -3282 39773
rect -3244 39739 -3210 39773
rect -3172 39739 -3138 39773
rect -3100 39739 -3066 39773
rect -3028 39739 -2994 39773
rect -2956 39739 -2922 39773
rect -2884 39739 -2850 39773
rect -2812 39739 -2778 39773
rect -2740 39739 -2706 39773
rect -2668 39739 -2634 39773
rect -2596 39739 -2562 39773
rect -2524 39739 -2490 39773
rect -2452 39739 -2418 39773
rect -2380 39739 -2346 39773
rect -2308 39739 -2274 39773
rect -2236 39739 -2202 39773
rect -2164 39739 -2130 39773
rect -2092 39739 -2058 39773
rect -2020 39739 -1986 39773
rect -1948 39739 -1914 39773
rect -1876 39739 -1842 39773
rect -1804 39739 -1770 39773
rect -1732 39739 -1698 39773
rect -1660 39739 -1626 39773
rect -1588 39739 -1554 39773
rect -1516 39739 -1482 39773
rect -1444 39739 -1410 39773
rect -1372 39739 -1338 39773
rect -1300 39739 -1266 39773
rect -1228 39739 -1194 39773
rect -1156 39739 -1122 39773
rect -1084 39739 -1050 39773
rect -1012 39739 -978 39773
rect -940 39739 -906 39773
rect -868 39739 -834 39773
rect -796 39739 -762 39773
rect -724 39739 -690 39773
rect -652 39739 -618 39773
rect -580 39739 -546 39773
rect -508 39739 -474 39773
rect -436 39739 -402 39773
rect -364 39739 -330 39773
rect -292 39739 -258 39773
rect -220 39739 -186 39773
rect 40128 39742 40162 39776
rect 40905 39757 40939 39791
rect 41808 39789 41842 39823
rect 43281 39842 43315 39876
rect 43453 39842 43487 39876
rect 43625 39842 43659 39876
rect 43797 39842 43831 39876
rect 43969 39842 44003 39876
rect 44174 39842 44208 39876
rect 44351 39842 44385 39876
rect 44523 39842 44557 39876
rect 44695 39842 44729 39876
rect 44867 39842 44901 39876
rect 45039 39842 45073 39876
rect 45211 39842 45245 39876
rect 43003 39792 43037 39826
rect 42539 39753 42573 39787
rect 42611 39753 42645 39787
rect 42683 39753 42717 39787
rect 42755 39753 42789 39787
rect 42827 39753 42861 39787
rect 42899 39753 42933 39787
rect 43277 39756 43311 39790
rect 43349 39756 43383 39790
rect 41808 39717 41842 39751
rect 43003 39720 43037 39754
rect 41808 39645 41842 39679
rect -31795 39080 -31761 39114
rect -31795 39008 -31761 39042
rect -31795 38936 -31761 38970
rect -31795 38864 -31761 38898
rect -31795 38516 -31761 38550
rect -31795 38444 -31761 38478
rect -31795 38372 -31761 38406
rect -31795 38300 -31761 38334
rect -31795 38228 -31761 38262
rect 88 16083 122 16117
rect 88 16011 122 16045
rect 88 15939 122 15973
rect 88 15867 122 15901
rect 88 15795 122 15829
rect 88 15723 122 15757
rect 88 15651 122 15685
rect 88 15579 122 15613
rect 88 15507 122 15541
rect 88 15435 122 15469
rect 88 15363 122 15397
rect 88 15291 122 15325
rect 88 15219 122 15253
rect 88 15147 122 15181
rect 88 15075 122 15109
rect 88 15003 122 15037
rect 88 14931 122 14965
rect 88 14859 122 14893
rect 88 14787 122 14821
rect 88 14715 122 14749
rect 88 14643 122 14677
rect 88 14571 122 14605
rect 88 14499 122 14533
rect 88 14427 122 14461
rect 11303 16088 11337 16122
rect 11303 16016 11337 16050
rect 11303 15944 11337 15978
rect 11303 15872 11337 15906
rect 11303 15800 11337 15834
rect 11303 15728 11337 15762
rect 11303 15656 11337 15690
rect 11303 15584 11337 15618
rect 11303 15512 11337 15546
rect 11303 15440 11337 15474
rect 11303 15368 11337 15402
rect 11303 15296 11337 15330
rect 11303 15224 11337 15258
rect 11303 15152 11337 15186
rect 11303 15080 11337 15114
rect 11303 15008 11337 15042
rect 11303 14936 11337 14970
rect 11303 14864 11337 14898
rect 11303 14792 11337 14826
rect 11303 14720 11337 14754
rect 11303 14648 11337 14682
rect 11303 14576 11337 14610
rect 11303 14504 11337 14538
rect 11303 14432 11337 14466
rect 88 14355 122 14389
rect 88 14283 122 14317
rect 88 14211 122 14245
rect 88 14139 122 14173
rect 88 14067 122 14101
rect 88 13995 122 14029
rect 88 13923 122 13957
rect 88 13851 122 13885
rect 88 13779 122 13813
rect 88 13707 122 13741
rect 88 13635 122 13669
rect 88 13563 122 13597
rect 88 13491 122 13525
rect 88 13419 122 13453
rect 88 13347 122 13381
rect 88 13275 122 13309
rect 88 13203 122 13237
rect 88 13131 122 13165
rect 88 13059 122 13093
rect 88 12987 122 13021
rect 11303 13886 11337 13920
rect 11303 13814 11337 13848
rect 11303 13742 11337 13776
rect 11303 13670 11337 13704
rect 11303 13598 11337 13632
rect 11303 13526 11337 13560
rect 11303 13454 11337 13488
rect 11303 13382 11337 13416
rect 11303 13310 11337 13344
rect 11303 13238 11337 13272
rect 11303 13166 11337 13200
rect 11303 13094 11337 13128
rect 11303 13022 11337 13056
rect 88 12915 122 12949
rect 88 12843 122 12877
rect 88 12771 122 12805
rect 88 12699 122 12733
rect 88 12627 122 12661
rect 88 12555 122 12589
rect 88 12483 122 12517
rect 88 12411 122 12445
rect 88 12339 122 12373
rect 88 12267 122 12301
rect 88 12195 122 12229
rect 88 12123 122 12157
rect 88 12051 122 12085
rect 88 11979 122 12013
rect 88 11907 122 11941
rect 88 11835 122 11869
rect 88 11763 122 11797
rect 88 11691 122 11725
rect 88 11619 122 11653
rect 88 11547 122 11581
rect 88 11475 122 11509
rect 88 11403 122 11437
rect 88 11331 122 11365
rect 11303 12057 11337 12091
rect 11303 11985 11337 12019
rect 11303 11913 11337 11947
rect 11303 11841 11337 11875
rect 11303 11769 11337 11803
rect 11303 11697 11337 11731
rect 11303 11625 11337 11659
rect 11303 11553 11337 11587
rect 11303 11481 11337 11515
rect 11303 11409 11337 11443
rect 11303 11337 11337 11371
rect 88 11259 122 11293
rect 88 11187 122 11221
rect 88 11115 122 11149
rect 88 11043 122 11077
rect 88 10971 122 11005
rect 88 10899 122 10933
rect 88 10827 122 10861
rect 88 10755 122 10789
rect 88 10683 122 10717
rect 6572 10438 6606 10472
rect 6644 10438 6678 10472
rect 6716 10438 6750 10472
rect 6788 10438 6822 10472
rect 6860 10438 6894 10472
rect 6932 10438 6966 10472
rect 7004 10438 7038 10472
rect 7076 10438 7110 10472
rect 7148 10438 7182 10472
rect 7220 10438 7254 10472
rect 7292 10438 7326 10472
rect 7364 10438 7398 10472
rect 7436 10438 7470 10472
rect 7508 10438 7542 10472
rect 7580 10438 7614 10472
rect 7652 10438 7686 10472
rect 7724 10438 7758 10472
rect 7796 10438 7830 10472
rect 7868 10438 7902 10472
rect 7940 10438 7974 10472
rect 8012 10438 8046 10472
rect 8084 10438 8118 10472
rect 8156 10438 8190 10472
rect 8228 10438 8262 10472
rect 8300 10438 8334 10472
rect 8372 10438 8406 10472
rect 8444 10438 8478 10472
rect 8516 10438 8550 10472
rect 8588 10438 8622 10472
rect 8660 10438 8694 10472
rect 8732 10438 8766 10472
rect 8804 10438 8838 10472
rect 8876 10438 8910 10472
rect 8948 10438 8982 10472
rect 9020 10438 9054 10472
rect 9092 10438 9126 10472
rect 9164 10438 9198 10472
rect 9236 10438 9270 10472
rect 9308 10438 9342 10472
rect 9380 10438 9414 10472
rect 9452 10438 9486 10472
rect 9524 10438 9558 10472
rect 9596 10438 9630 10472
rect 9668 10438 9702 10472
rect 9740 10438 9774 10472
rect 9812 10438 9846 10472
rect 9884 10438 9918 10472
rect 9956 10438 9990 10472
rect 10028 10438 10062 10472
rect 10100 10438 10134 10472
rect 10172 10438 10206 10472
rect 10244 10438 10278 10472
rect 10316 10438 10350 10472
rect 10388 10438 10422 10472
rect 10460 10438 10494 10472
rect 10532 10438 10566 10472
rect 10604 10438 10638 10472
rect 10676 10438 10710 10472
rect 10748 10438 10782 10472
rect 10820 10438 10854 10472
rect 10892 10438 10926 10472
rect 10964 10438 10998 10472
rect 11036 10438 11070 10472
<< metal1 >>
rect -15420 78112 -15164 78140
rect -15420 77932 -15382 78112
rect -15202 77932 -15164 78112
rect -15420 77904 -15164 77932
rect 12596 78083 12852 78111
rect -16859 76718 -16738 76723
rect -16859 76666 -16825 76718
rect -16773 76666 -16738 76718
rect -16859 76654 -16738 76666
rect -16859 76602 -16825 76654
rect -16773 76602 -16738 76654
rect -16859 76590 -16738 76602
rect -16859 76538 -16825 76590
rect -16773 76538 -16738 76590
rect -16859 76526 -16738 76538
rect -16859 76474 -16825 76526
rect -16773 76474 -16738 76526
rect -16859 76462 -16738 76474
rect -16859 76410 -16825 76462
rect -16773 76410 -16738 76462
rect -16859 76398 -16738 76410
rect -16859 76346 -16825 76398
rect -16773 76346 -16738 76398
rect -16859 76334 -16738 76346
rect -16859 76282 -16825 76334
rect -16773 76282 -16738 76334
rect -16859 76270 -16738 76282
rect -16859 76218 -16825 76270
rect -16773 76218 -16738 76270
rect -16859 76206 -16738 76218
rect -16859 76154 -16825 76206
rect -16773 76154 -16738 76206
rect -16859 76142 -16738 76154
rect -16859 76090 -16825 76142
rect -16773 76090 -16738 76142
rect -16859 76078 -16738 76090
rect -16859 76026 -16825 76078
rect -16773 76026 -16738 76078
rect -16859 76014 -16738 76026
rect -16859 75962 -16825 76014
rect -16773 75962 -16738 76014
rect -16859 75950 -16738 75962
rect -16859 75898 -16825 75950
rect -16773 75898 -16738 75950
rect -16859 75886 -16738 75898
rect -16859 75834 -16825 75886
rect -16773 75834 -16738 75886
rect -16859 75822 -16738 75834
rect -16859 75770 -16825 75822
rect -16773 75770 -16738 75822
rect -16859 75758 -16738 75770
rect -16859 75706 -16825 75758
rect -16773 75706 -16738 75758
rect -16859 75694 -16738 75706
rect -16859 75642 -16825 75694
rect -16773 75642 -16738 75694
rect -16859 75630 -16738 75642
rect -16859 75578 -16825 75630
rect -16773 75578 -16738 75630
rect -16859 75566 -16738 75578
rect -16859 75514 -16825 75566
rect -16773 75514 -16738 75566
rect -16859 75502 -16738 75514
rect -16859 75450 -16825 75502
rect -16773 75450 -16738 75502
rect -16859 75438 -16738 75450
rect -16859 75386 -16825 75438
rect -16773 75386 -16738 75438
rect -16859 75374 -16738 75386
rect -16859 75322 -16825 75374
rect -16773 75322 -16738 75374
rect -16859 75310 -16738 75322
rect -16859 75258 -16825 75310
rect -16773 75258 -16738 75310
rect -16859 75246 -16738 75258
rect -15353 75255 -15225 77904
rect 12596 77903 12634 78083
rect 12814 77903 12852 78083
rect 12596 77875 12852 77903
rect 24646 78084 24902 78112
rect 24646 77904 24684 78084
rect 24864 77904 24902 78084
rect 24646 77876 24902 77904
rect 11177 76732 11367 76806
rect -13858 76724 -13737 76729
rect -13858 76672 -13824 76724
rect -13772 76672 -13737 76724
rect -13858 76660 -13737 76672
rect -13858 76608 -13824 76660
rect -13772 76608 -13737 76660
rect -13858 76596 -13737 76608
rect -13858 76544 -13824 76596
rect -13772 76544 -13737 76596
rect -13858 76532 -13737 76544
rect -13858 76480 -13824 76532
rect -13772 76480 -13737 76532
rect -13858 76468 -13737 76480
rect -13858 76416 -13824 76468
rect -13772 76416 -13737 76468
rect -13858 76404 -13737 76416
rect -13858 76352 -13824 76404
rect -13772 76352 -13737 76404
rect -13858 76340 -13737 76352
rect -13858 76288 -13824 76340
rect -13772 76288 -13737 76340
rect -13858 76276 -13737 76288
rect -13858 76224 -13824 76276
rect -13772 76224 -13737 76276
rect -13858 76212 -13737 76224
rect -13858 76160 -13824 76212
rect -13772 76160 -13737 76212
rect -13858 76148 -13737 76160
rect -13858 76096 -13824 76148
rect -13772 76096 -13737 76148
rect -13858 76084 -13737 76096
rect -13858 76032 -13824 76084
rect -13772 76032 -13737 76084
rect -13858 76020 -13737 76032
rect -13858 75968 -13824 76020
rect -13772 75968 -13737 76020
rect -13858 75956 -13737 75968
rect -13858 75904 -13824 75956
rect -13772 75904 -13737 75956
rect -13858 75892 -13737 75904
rect -13858 75840 -13824 75892
rect -13772 75840 -13737 75892
rect -13858 75828 -13737 75840
rect -13858 75776 -13824 75828
rect -13772 75776 -13737 75828
rect -13858 75764 -13737 75776
rect -13858 75712 -13824 75764
rect -13772 75712 -13737 75764
rect -13858 75700 -13737 75712
rect -13858 75648 -13824 75700
rect -13772 75648 -13737 75700
rect -13858 75636 -13737 75648
rect -13858 75584 -13824 75636
rect -13772 75584 -13737 75636
rect -13858 75572 -13737 75584
rect -13858 75520 -13824 75572
rect -13772 75520 -13737 75572
rect -13858 75508 -13737 75520
rect -13858 75456 -13824 75508
rect -13772 75456 -13737 75508
rect -13858 75444 -13737 75456
rect -13858 75392 -13824 75444
rect -13772 75392 -13737 75444
rect -13858 75380 -13737 75392
rect -13858 75328 -13824 75380
rect -13772 75328 -13737 75380
rect -13858 75316 -13737 75328
rect -13858 75264 -13824 75316
rect -13772 75264 -13737 75316
rect -16859 75194 -16825 75246
rect -16773 75194 -16738 75246
rect -16859 75182 -16738 75194
rect -16859 75130 -16825 75182
rect -16773 75130 -16738 75182
rect -16859 75118 -16738 75130
rect -16859 75066 -16825 75118
rect -16773 75066 -16738 75118
rect -16859 75054 -16738 75066
rect -16859 75002 -16825 75054
rect -16773 75002 -16738 75054
rect -16859 74990 -16738 75002
rect -16859 74938 -16825 74990
rect -16773 74938 -16738 74990
rect -16859 74926 -16738 74938
rect -16859 74874 -16825 74926
rect -16773 74874 -16738 74926
rect -16859 74862 -16738 74874
rect -16859 74810 -16825 74862
rect -16773 74810 -16738 74862
rect -16859 74798 -16738 74810
rect -13858 75252 -13737 75264
rect -13858 75200 -13824 75252
rect -13772 75200 -13737 75252
rect -13858 75188 -13737 75200
rect -13858 75136 -13824 75188
rect -13772 75136 -13737 75188
rect -13858 75124 -13737 75136
rect -13858 75072 -13824 75124
rect -13772 75072 -13737 75124
rect -13858 75060 -13737 75072
rect -13858 75008 -13824 75060
rect -13772 75008 -13737 75060
rect -13858 74996 -13737 75008
rect -13858 74944 -13824 74996
rect -13772 74944 -13737 74996
rect -13858 74932 -13737 74944
rect -13858 74880 -13824 74932
rect -13772 74880 -13737 74932
rect -13858 74868 -13737 74880
rect -13858 74816 -13824 74868
rect -13772 74816 -13737 74868
rect -13858 74804 -13737 74816
rect -16859 74746 -16825 74798
rect -16773 74746 -16738 74798
rect -16859 74734 -16738 74746
rect -16859 74682 -16825 74734
rect -16773 74682 -16738 74734
rect -16859 74670 -16738 74682
rect -16859 74618 -16825 74670
rect -16773 74618 -16738 74670
rect -16859 74606 -16738 74618
rect -16859 74554 -16825 74606
rect -16773 74554 -16738 74606
rect -16859 74542 -16738 74554
rect -16859 74490 -16825 74542
rect -16773 74490 -16738 74542
rect -16859 74478 -16738 74490
rect -16859 74426 -16825 74478
rect -16773 74426 -16738 74478
rect -16859 74414 -16738 74426
rect -16859 74362 -16825 74414
rect -16773 74362 -16738 74414
rect -16859 74350 -16738 74362
rect -16859 74298 -16825 74350
rect -16773 74298 -16738 74350
rect -16859 74286 -16738 74298
rect -16859 74234 -16825 74286
rect -16773 74234 -16738 74286
rect -16859 74222 -16738 74234
rect -16859 74170 -16825 74222
rect -16773 74170 -16738 74222
rect -16859 74158 -16738 74170
rect -16859 74106 -16825 74158
rect -16773 74106 -16738 74158
rect -16859 74094 -16738 74106
rect -16859 74042 -16825 74094
rect -16773 74042 -16738 74094
rect -16859 74030 -16738 74042
rect -16859 73978 -16825 74030
rect -16773 73978 -16738 74030
rect -16859 73966 -16738 73978
rect -16859 73914 -16825 73966
rect -16773 73914 -16738 73966
rect -16859 73902 -16738 73914
rect -16859 73850 -16825 73902
rect -16773 73850 -16738 73902
rect -16859 73838 -16738 73850
rect -16859 73786 -16825 73838
rect -16773 73786 -16738 73838
rect -16859 73774 -16738 73786
rect -16859 73722 -16825 73774
rect -16773 73722 -16738 73774
rect -16859 73710 -16738 73722
rect -16859 73658 -16825 73710
rect -16773 73658 -16738 73710
rect -16859 73646 -16738 73658
rect -16859 73594 -16825 73646
rect -16773 73594 -16738 73646
rect -16859 73582 -16738 73594
rect -16859 73530 -16825 73582
rect -16773 73530 -16738 73582
rect -16859 73518 -16738 73530
rect -16859 73466 -16825 73518
rect -16773 73466 -16738 73518
rect -16859 73454 -16738 73466
rect -16859 73402 -16825 73454
rect -16773 73402 -16738 73454
rect -16859 73398 -16738 73402
rect -15353 71958 -15225 74801
rect -13858 74752 -13824 74804
rect -13772 74752 -13737 74804
rect -13858 74740 -13737 74752
rect -13858 74688 -13824 74740
rect -13772 74688 -13737 74740
rect -13858 74676 -13737 74688
rect -13858 74624 -13824 74676
rect -13772 74624 -13737 74676
rect -13858 74612 -13737 74624
rect -13858 74560 -13824 74612
rect -13772 74560 -13737 74612
rect -13858 74548 -13737 74560
rect -13858 74496 -13824 74548
rect -13772 74496 -13737 74548
rect -13858 74484 -13737 74496
rect -13858 74432 -13824 74484
rect -13772 74432 -13737 74484
rect -13858 74420 -13737 74432
rect -13858 74368 -13824 74420
rect -13772 74368 -13737 74420
rect -13858 74356 -13737 74368
rect -13858 74304 -13824 74356
rect -13772 74304 -13737 74356
rect -13858 74292 -13737 74304
rect -13858 74240 -13824 74292
rect -13772 74240 -13737 74292
rect -13858 74228 -13737 74240
rect -13858 74176 -13824 74228
rect -13772 74176 -13737 74228
rect -13858 74164 -13737 74176
rect -13858 74112 -13824 74164
rect -13772 74112 -13737 74164
rect -13858 74100 -13737 74112
rect -13858 74048 -13824 74100
rect -13772 74048 -13737 74100
rect -13858 74036 -13737 74048
rect -13858 73984 -13824 74036
rect -13772 73984 -13737 74036
rect -13858 73972 -13737 73984
rect -13858 73920 -13824 73972
rect -13772 73920 -13737 73972
rect -13858 73908 -13737 73920
rect -13858 73856 -13824 73908
rect -13772 73856 -13737 73908
rect -13858 73844 -13737 73856
rect -13858 73792 -13824 73844
rect -13772 73792 -13737 73844
rect -13858 73780 -13737 73792
rect -13858 73728 -13824 73780
rect -13772 73728 -13737 73780
rect -13858 73716 -13737 73728
rect -13858 73664 -13824 73716
rect -13772 73664 -13737 73716
rect -13858 73652 -13737 73664
rect -13858 73600 -13824 73652
rect -13772 73600 -13737 73652
rect -13858 73588 -13737 73600
rect -13858 73536 -13824 73588
rect -13772 73536 -13737 73588
rect -13858 73524 -13737 73536
rect -13858 73472 -13824 73524
rect -13772 73472 -13737 73524
rect -13858 73460 -13737 73472
rect -13858 73408 -13824 73460
rect -13772 73408 -13737 73460
rect -13858 73404 -13737 73408
rect 11133 76720 11367 76732
rect 11133 73404 11149 76720
rect 11265 73404 11367 76720
rect 11133 73392 11367 73404
rect 11177 73320 11367 73392
rect 12660 73019 12778 77875
rect 14134 76733 14282 76745
rect 14134 73417 14150 76733
rect 14266 73417 14282 76733
rect 14134 73405 14282 73417
rect -16674 71796 -16590 71802
rect -15279 71799 -15195 71805
rect -16674 71744 -16658 71796
rect -16606 71744 -16590 71796
rect -16674 71738 -16590 71744
rect -15496 71792 -15412 71798
rect -15496 71740 -15480 71792
rect -15428 71740 -15412 71792
rect -15279 71747 -15263 71799
rect -15211 71747 -15195 71799
rect -15279 71741 -15195 71747
rect -14145 71796 -14061 71802
rect -14145 71744 -14129 71796
rect -14077 71744 -14061 71796
rect -15496 71734 -15412 71740
rect -14145 71738 -14061 71744
rect -16564 70292 -16480 70298
rect -16564 70240 -16548 70292
rect -16496 70240 -16480 70292
rect -16564 70234 -16480 70240
rect -15450 70278 -15366 70284
rect -15450 70226 -15434 70278
rect -15382 70226 -15366 70278
rect -15450 70220 -15366 70226
rect -15237 70279 -15153 70285
rect -15237 70227 -15221 70279
rect -15169 70227 -15153 70279
rect -15237 70221 -15153 70227
rect -14073 70279 -13989 70285
rect -14073 70227 -14057 70279
rect -14005 70227 -13989 70279
rect -14073 70221 -13989 70227
rect -15432 68494 -15348 68515
rect -15432 68442 -15416 68494
rect -15364 68442 -15348 68494
rect -15432 68430 -15348 68442
rect -15432 68378 -15416 68430
rect -15364 68378 -15348 68430
rect -15432 68366 -15348 68378
rect -15432 68314 -15416 68366
rect -15364 68314 -15348 68366
rect -15432 68302 -15348 68314
rect -15973 68241 -15880 68261
rect -15973 68189 -15953 68241
rect -15901 68189 -15880 68241
rect -15973 68177 -15880 68189
rect -15973 68125 -15953 68177
rect -15901 68125 -15880 68177
rect -15432 68250 -15416 68302
rect -15364 68250 -15348 68302
rect -15432 68238 -15348 68250
rect -15432 68186 -15416 68238
rect -15364 68186 -15348 68238
rect -15432 68166 -15348 68186
rect -14889 68244 -14796 68264
rect -14889 68192 -14869 68244
rect -14817 68192 -14796 68244
rect -14889 68180 -14796 68192
rect -15973 68105 -15880 68125
rect -14889 68128 -14869 68180
rect -14817 68128 -14796 68180
rect -14889 68108 -14796 68128
rect -16587 67607 -16503 67613
rect -14314 67612 -14230 67618
rect -16587 67555 -16571 67607
rect -16519 67555 -16503 67607
rect -16587 67549 -16503 67555
rect -15432 67601 -15348 67607
rect -15432 67549 -15416 67601
rect -15364 67549 -15348 67601
rect -14314 67560 -14298 67612
rect -14246 67560 -14230 67612
rect -14314 67554 -14230 67560
rect -15432 67543 -15348 67549
rect -16123 52998 -15995 66326
rect -14782 53600 -14654 66338
rect -9894 63396 -9432 63402
rect -9894 63344 -9881 63396
rect -9829 63344 -9817 63396
rect -9765 63344 -9753 63396
rect -9701 63344 -9689 63396
rect -9637 63344 -9625 63396
rect -9573 63344 -9561 63396
rect -9509 63344 -9497 63396
rect -9445 63344 -9432 63396
rect -9894 63338 -9432 63344
rect -9237 63338 -8980 63402
rect -8083 63398 -7621 63404
rect -8083 63346 -8070 63398
rect -8018 63346 -8006 63398
rect -7954 63346 -7942 63398
rect -7890 63346 -7878 63398
rect -7826 63346 -7814 63398
rect -7762 63346 -7750 63398
rect -7698 63346 -7686 63398
rect -7634 63346 -7621 63398
rect -8083 63340 -7621 63346
rect -9136 62888 -9072 63338
rect -7427 63332 -7188 63396
rect -6288 63394 -5826 63400
rect -6288 63342 -6275 63394
rect -6223 63342 -6211 63394
rect -6159 63342 -6147 63394
rect -6095 63342 -6083 63394
rect -6031 63342 -6019 63394
rect -5967 63342 -5955 63394
rect -5903 63342 -5891 63394
rect -5839 63342 -5826 63394
rect -6288 63336 -5826 63342
rect -5623 63337 -5392 63401
rect -4489 63392 -4027 63398
rect -4489 63340 -4476 63392
rect -4424 63340 -4412 63392
rect -4360 63340 -4348 63392
rect -4296 63340 -4284 63392
rect -4232 63340 -4220 63392
rect -4168 63340 -4156 63392
rect -4104 63340 -4092 63392
rect -4040 63340 -4027 63392
rect -7341 62888 -7277 63332
rect -6949 63176 -6689 63206
rect -6949 62996 -6909 63176
rect -6729 62996 -6689 63176
rect -6949 62966 -6689 62996
rect -6857 62888 -6793 62966
rect -5541 62888 -5477 63337
rect -4489 63334 -4027 63340
rect -3832 63335 -3572 63399
rect -2698 63396 -2236 63402
rect -2698 63344 -2685 63396
rect -2633 63344 -2621 63396
rect -2569 63344 -2557 63396
rect -2505 63344 -2493 63396
rect -2441 63344 -2429 63396
rect -2377 63344 -2365 63396
rect -2313 63344 -2301 63396
rect -2249 63344 -2236 63396
rect -2698 63338 -2236 63344
rect -2029 63339 -1794 63403
rect -896 63392 -434 63398
rect -896 63340 -883 63392
rect -831 63340 -819 63392
rect -767 63340 -755 63392
rect -703 63340 -691 63392
rect -639 63340 -627 63392
rect -575 63340 -563 63392
rect -511 63340 -499 63392
rect -447 63340 -434 63392
rect -3738 62888 -3674 63335
rect -1934 62888 -1870 63339
rect -896 63334 -434 63340
rect -221 63338 -2 63402
rect -138 63141 -74 63338
rect 747 63202 1297 63232
rect 747 63141 772 63202
rect -138 63077 772 63141
rect -138 62888 -74 63077
rect 747 63022 772 63077
rect 1272 63022 1297 63202
rect 747 62992 1297 63022
rect -9136 62824 -74 62888
rect 337 60808 529 60827
rect -6867 54596 -6803 54597
rect -8567 54589 -8483 54595
rect -8567 54537 -8551 54589
rect -8499 54537 -8483 54589
rect -8567 54531 -8483 54537
rect -6876 54590 -6792 54596
rect -6876 54538 -6860 54590
rect -6808 54538 -6792 54590
rect -6876 54532 -6792 54538
rect -5171 54589 -5087 54595
rect -5171 54537 -5155 54589
rect -5103 54537 -5087 54589
rect -9714 54397 -9452 54403
rect -8557 54401 -8493 54531
rect -6867 54403 -6803 54532
rect -5171 54531 -5087 54537
rect -3375 54589 -3291 54595
rect -3375 54537 -3359 54589
rect -3307 54537 -3291 54589
rect -3375 54531 -3291 54537
rect -1546 54589 -1462 54595
rect -1546 54537 -1530 54589
rect -1478 54537 -1462 54589
rect -1546 54531 -1462 54537
rect -9714 54345 -9673 54397
rect -9621 54345 -9609 54397
rect -9557 54345 -9545 54397
rect -9493 54345 -9452 54397
rect -9714 54339 -9452 54345
rect -9230 54337 -8491 54401
rect -7919 54396 -7657 54402
rect -7919 54344 -7878 54396
rect -7826 54344 -7814 54396
rect -7762 54344 -7750 54396
rect -7698 54344 -7657 54396
rect -7919 54338 -7657 54344
rect -7435 54339 -6803 54403
rect -6119 54398 -5857 54404
rect -5161 54403 -5097 54531
rect -6119 54346 -6078 54398
rect -6026 54346 -6014 54398
rect -5962 54346 -5950 54398
rect -5898 54346 -5857 54398
rect -6119 54340 -5857 54346
rect -5632 54339 -5097 54403
rect -4321 54397 -4059 54403
rect -3365 54401 -3301 54531
rect -4321 54345 -4280 54397
rect -4228 54345 -4216 54397
rect -4164 54345 -4152 54397
rect -4100 54345 -4059 54397
rect -4321 54339 -4059 54345
rect -3832 54339 -3301 54401
rect -2523 54398 -2261 54404
rect -1536 54402 -1472 54531
rect -2523 54346 -2482 54398
rect -2430 54346 -2418 54398
rect -2366 54346 -2354 54398
rect -2302 54346 -2261 54398
rect -2523 54340 -2261 54346
rect -2027 54338 -1472 54402
rect -720 54397 -458 54403
rect -720 54345 -679 54397
rect -627 54345 -615 54397
rect -563 54345 -551 54397
rect -499 54345 -458 54397
rect -720 54339 -458 54345
rect -225 54398 250 54404
rect -225 54346 182 54398
rect 234 54346 250 54398
rect -225 54340 250 54346
rect -14793 53594 -14645 53600
rect -14793 53542 -14777 53594
rect -14725 53542 -14713 53594
rect -14661 53542 -14645 53594
rect -14793 53536 -14645 53542
rect -7560 53594 -7476 53600
rect -7560 53542 -7544 53594
rect -7492 53542 -7476 53594
rect -7560 53536 -7476 53542
rect -6999 53594 -6851 53600
rect -6999 53542 -6983 53594
rect -6931 53542 -6919 53594
rect -6867 53542 -6851 53594
rect -6999 53536 -6851 53542
rect -14782 53520 -14654 53536
rect 337 53140 375 60808
rect 491 53140 529 60808
rect 337 53121 529 53140
rect 10167 60812 10561 60836
rect -16123 52986 -9120 52998
rect -16123 52934 -9392 52986
rect -9340 52934 -9328 52986
rect -9276 52934 -9120 52986
rect -16123 52923 -9120 52934
rect -8864 51221 -8760 51249
rect -8864 51169 -8838 51221
rect -8786 51169 -8760 51221
rect -8864 51157 -8760 51169
rect -8864 51105 -8838 51157
rect -8786 51105 -8760 51157
rect -8864 51093 -8760 51105
rect -8864 51041 -8838 51093
rect -8786 51041 -8760 51093
rect -8864 51014 -8760 51041
rect -5698 51064 -3878 51066
rect -9408 50931 -8690 50937
rect -9408 50879 -9392 50931
rect -9340 50879 -9328 50931
rect -9276 50879 -8690 50931
rect -9408 50873 -8690 50879
rect -7544 50929 -6851 50935
rect -7544 50877 -6983 50929
rect -6931 50877 -6919 50929
rect -6867 50877 -6851 50929
rect -5698 50884 -5678 51064
rect -3898 51024 -3878 51064
rect -3372 51043 -2526 51074
rect -3372 51024 -3359 51043
rect -3898 50988 -3359 51024
rect -2539 51024 -2526 51043
rect -1665 51033 -755 51064
rect -1665 51024 -1652 51033
rect -2539 50988 -1652 51024
rect -768 51024 -755 51033
rect -768 50988 -143 51024
rect -3898 50954 -3879 50988
rect -3845 50954 -3807 50988
rect -3773 50954 -3735 50988
rect -3701 50954 -3663 50988
rect -3629 50954 -3591 50988
rect -3557 50954 -3519 50988
rect -3485 50954 -3447 50988
rect -3413 50954 -3375 50988
rect -2539 50954 -2511 50988
rect -2477 50954 -2439 50988
rect -2405 50954 -2367 50988
rect -2333 50954 -2295 50988
rect -2261 50954 -2223 50988
rect -2189 50954 -2151 50988
rect -2117 50954 -2079 50988
rect -2045 50954 -2007 50988
rect -1973 50954 -1935 50988
rect -1901 50954 -1863 50988
rect -1829 50954 -1791 50988
rect -1757 50954 -1719 50988
rect -1685 50954 -1652 50988
rect -749 50954 -711 50988
rect -677 50954 -639 50988
rect -605 50954 -567 50988
rect -533 50954 -495 50988
rect -461 50954 -423 50988
rect -389 50954 -351 50988
rect -317 50954 -279 50988
rect -245 50954 -207 50988
rect -173 50954 -143 50988
rect -3898 50927 -3359 50954
rect -2539 50927 -1652 50954
rect -3898 50919 -1652 50927
rect -3898 50884 -3878 50919
rect -3372 50896 -2526 50919
rect -1665 50917 -1652 50919
rect -768 50919 -143 50954
rect -768 50917 -755 50919
rect -1665 50886 -755 50917
rect -5698 50883 -3878 50884
rect -7544 50871 -6851 50877
rect -8884 50770 -8770 50791
rect -8884 50718 -8853 50770
rect -8801 50718 -8770 50770
rect -88 50761 131 50774
rect -8884 50706 -8770 50718
rect -8884 50654 -8853 50706
rect -8801 50654 -8770 50706
rect -8884 50642 -8770 50654
rect -8884 50590 -8853 50642
rect -8801 50590 -8770 50642
rect -8884 50578 -8770 50590
rect -8884 50526 -8853 50578
rect -8801 50526 -8770 50578
rect -8884 50514 -8770 50526
rect -8884 50462 -8853 50514
rect -8801 50462 -8770 50514
rect -8884 50450 -8770 50462
rect -8884 50398 -8853 50450
rect -8801 50398 -8770 50450
rect -8884 50378 -8770 50398
rect -5942 50714 -5738 50720
rect -27080 49714 -26716 49720
rect -27080 49662 -27052 49714
rect -27000 49662 -26988 49714
rect -26936 49662 -26924 49714
rect -26872 49662 -26860 49714
rect -26808 49662 -26796 49714
rect -26744 49662 -26716 49714
rect -27080 49656 -26716 49662
rect -26059 49447 -26001 49468
rect -26059 49424 -26047 49447
rect -26070 49418 -26047 49424
rect -26013 49424 -26001 49447
rect -26013 49418 -25986 49424
rect -26418 49407 -26147 49413
rect -26418 49355 -26405 49407
rect -26353 49398 -26341 49407
rect -26289 49398 -26277 49407
rect -26225 49398 -26213 49407
rect -26343 49364 -26341 49398
rect -26353 49355 -26341 49364
rect -26289 49355 -26277 49364
rect -26225 49355 -26213 49364
rect -26161 49355 -26147 49407
rect -26070 49366 -26054 49418
rect -26002 49366 -25986 49418
rect -26070 49361 -25986 49366
rect -26070 49360 -26047 49361
rect -26418 49349 -26147 49355
rect -26059 49327 -26047 49360
rect -26013 49360 -25986 49361
rect -26013 49327 -26001 49360
rect -26059 49295 -26001 49327
rect -25994 49172 -25630 49178
rect -25994 49120 -25966 49172
rect -25914 49120 -25902 49172
rect -25850 49120 -25838 49172
rect -25786 49120 -25774 49172
rect -25722 49120 -25710 49172
rect -25658 49120 -25630 49172
rect -25994 49114 -25630 49120
rect -5942 47782 -5930 50714
rect -5750 47782 -5738 50714
rect -5942 47776 -5738 47782
rect -88 47765 -69 50761
rect 111 47765 131 50761
rect -88 47752 131 47765
rect 10167 47640 10178 60812
rect 10550 47640 10561 60812
rect 10167 47617 10561 47640
rect -5934 46272 -5712 46274
rect -27097 43296 -26980 43313
rect -27097 43244 -27065 43296
rect -27013 43244 -26980 43296
rect -27097 43232 -26980 43244
rect -27097 43180 -27065 43232
rect -27013 43180 -26980 43232
rect -27097 43168 -26980 43180
rect -27097 43116 -27065 43168
rect -27013 43116 -26980 43168
rect -27097 43104 -26980 43116
rect -27097 43052 -27065 43104
rect -27013 43052 -26980 43104
rect -27097 43040 -26980 43052
rect -27097 42988 -27065 43040
rect -27013 42988 -26980 43040
rect -13479 43055 -13395 43061
rect -13479 43003 -13463 43055
rect -13411 43003 -13395 43055
rect -13479 42997 -13395 43003
rect -27097 42976 -26980 42988
rect -27097 42924 -27065 42976
rect -27013 42924 -26980 42976
rect -27097 42912 -26980 42924
rect -27097 42860 -27065 42912
rect -27013 42860 -26980 42912
rect -27097 42848 -26980 42860
rect -27097 42796 -27065 42848
rect -27013 42796 -26980 42848
rect -27097 42779 -26980 42796
rect -27092 42155 -26985 42169
rect -27092 42103 -27065 42155
rect -27013 42103 -26985 42155
rect -27092 42091 -26985 42103
rect -27092 42039 -27065 42091
rect -27013 42039 -26985 42091
rect -27092 42027 -26985 42039
rect -27092 41975 -27065 42027
rect -27013 41975 -26985 42027
rect -27092 41963 -26985 41975
rect -27092 41911 -27065 41963
rect -27013 41911 -26985 41963
rect -27092 41899 -26985 41911
rect -27092 41847 -27065 41899
rect -27013 41847 -26985 41899
rect -27092 41835 -26985 41847
rect -27092 41783 -27065 41835
rect -27013 41783 -26985 41835
rect -27092 41771 -26985 41783
rect -27092 41719 -27065 41771
rect -27013 41719 -26985 41771
rect -27092 41707 -26985 41719
rect -27092 41655 -27065 41707
rect -27013 41655 -26985 41707
rect -27092 41643 -26985 41655
rect -27092 41591 -27065 41643
rect -27013 41591 -26985 41643
rect -27092 41579 -26985 41591
rect -27092 41527 -27065 41579
rect -27013 41527 -26985 41579
rect -27092 41515 -26985 41527
rect -27092 41463 -27065 41515
rect -27013 41463 -26985 41515
rect -27092 41451 -26985 41463
rect -27092 41399 -27065 41451
rect -27013 41399 -26985 41451
rect -27092 41387 -26985 41399
rect -27092 41335 -27065 41387
rect -27013 41335 -26985 41387
rect -27092 41323 -26985 41335
rect -27092 41271 -27065 41323
rect -27013 41271 -26985 41323
rect -27092 41259 -26985 41271
rect -27092 41207 -27065 41259
rect -27013 41207 -26985 41259
rect -27092 41195 -26985 41207
rect -27092 41143 -27065 41195
rect -27013 41143 -26985 41195
rect -27092 41131 -26985 41143
rect -27092 41079 -27065 41131
rect -27013 41079 -26985 41131
rect -27092 41067 -26985 41079
rect -27092 41015 -27065 41067
rect -27013 41015 -26985 41067
rect -27092 41002 -26985 41015
rect -27087 40629 -26980 40643
rect -27087 40577 -27060 40629
rect -27008 40577 -26980 40629
rect -27087 40565 -26980 40577
rect -27087 40513 -27060 40565
rect -27008 40513 -26980 40565
rect -27087 40501 -26980 40513
rect -27087 40449 -27060 40501
rect -27008 40449 -26980 40501
rect -27087 40437 -26980 40449
rect -27087 40385 -27060 40437
rect -27008 40385 -26980 40437
rect -27087 40373 -26980 40385
rect -27087 40321 -27060 40373
rect -27008 40321 -26980 40373
rect -27087 40309 -26980 40321
rect -27087 40257 -27060 40309
rect -27008 40257 -26980 40309
rect -27087 40245 -26980 40257
rect -27087 40193 -27060 40245
rect -27008 40193 -26980 40245
rect -27087 40181 -26980 40193
rect -27087 40129 -27060 40181
rect -27008 40129 -26980 40181
rect -27087 40117 -26980 40129
rect -27087 40065 -27060 40117
rect -27008 40065 -26980 40117
rect -27087 40053 -26980 40065
rect -27087 40001 -27060 40053
rect -27008 40001 -26980 40053
rect -27087 39989 -26980 40001
rect -27087 39937 -27060 39989
rect -27008 39937 -26980 39989
rect -27087 39925 -26980 39937
rect -27087 39873 -27060 39925
rect -27008 39873 -26980 39925
rect -27087 39861 -26980 39873
rect -27087 39809 -27060 39861
rect -27008 39809 -26980 39861
rect -27087 39797 -26980 39809
rect -27087 39745 -27060 39797
rect -27008 39745 -26980 39797
rect -27087 39733 -26980 39745
rect -27087 39681 -27060 39733
rect -27008 39681 -26980 39733
rect -27087 39669 -26980 39681
rect -27087 39617 -27060 39669
rect -27008 39617 -26980 39669
rect -27087 39605 -26980 39617
rect -27087 39553 -27060 39605
rect -27008 39553 -26980 39605
rect -27087 39541 -26980 39553
rect -27087 39489 -27060 39541
rect -27008 39489 -26980 39541
rect -27087 39476 -26980 39489
rect -18893 39520 -18797 39537
rect -18893 39468 -18871 39520
rect -18819 39468 -18797 39520
rect -18893 39456 -18797 39468
rect -18893 39404 -18871 39456
rect -18819 39404 -18797 39456
rect -18893 39392 -18797 39404
rect -18893 39340 -18871 39392
rect -18819 39340 -18797 39392
rect -18893 39328 -18797 39340
rect -18893 39276 -18871 39328
rect -18819 39276 -18797 39328
rect -18893 39264 -18797 39276
rect -18893 39212 -18871 39264
rect -18819 39212 -18797 39264
rect -18893 39200 -18797 39212
rect -31822 39150 -31738 39166
rect -31822 39098 -31806 39150
rect -31754 39098 -31738 39150
rect -18893 39148 -18871 39200
rect -18819 39148 -18797 39200
rect -31146 39126 -31082 39141
rect -31822 39086 -31795 39098
rect -31761 39086 -31738 39098
rect -31549 39092 -31082 39126
rect -18893 39136 -18797 39148
rect -31822 39034 -31806 39086
rect -31754 39034 -31738 39086
rect -31822 39022 -31795 39034
rect -31761 39022 -31738 39034
rect -31822 39007 -31806 39022
rect -31831 38973 -31806 39007
rect -31822 38970 -31806 38973
rect -31754 39007 -31738 39022
rect -31754 38973 -31710 39007
rect -31754 38970 -31738 38973
rect -31822 38958 -31795 38970
rect -31761 38958 -31738 38970
rect -31822 38906 -31806 38958
rect -31754 38906 -31738 38958
rect -31822 38898 -31738 38906
rect -31822 38894 -31795 38898
rect -31761 38894 -31738 38898
rect -31822 38842 -31806 38894
rect -31754 38842 -31738 38894
rect -31146 38886 -31082 39092
rect -31553 38852 -31082 38886
rect -31822 38827 -31738 38842
rect -31821 38595 -31737 38613
rect -31821 38543 -31805 38595
rect -31753 38543 -31737 38595
rect -31146 38570 -31082 38852
rect -31821 38531 -31795 38543
rect -31761 38531 -31737 38543
rect -31553 38536 -31082 38570
rect -31821 38479 -31805 38531
rect -31753 38479 -31737 38531
rect -31821 38478 -31737 38479
rect -31821 38467 -31795 38478
rect -31761 38467 -31737 38478
rect -31821 38415 -31805 38467
rect -31753 38415 -31737 38467
rect -31821 38407 -31737 38415
rect -31831 38406 -31734 38407
rect -31831 38403 -31795 38406
rect -31761 38403 -31734 38406
rect -31831 38373 -31805 38403
rect -31821 38351 -31805 38373
rect -31753 38373 -31734 38403
rect -31753 38351 -31737 38373
rect -31821 38339 -31737 38351
rect -31821 38287 -31805 38339
rect -31753 38287 -31737 38339
rect -31821 38275 -31737 38287
rect -31821 38223 -31805 38275
rect -31753 38223 -31737 38275
rect -31146 38256 -31082 38536
rect -27092 39118 -26988 39120
rect -27092 39066 -27066 39118
rect -27014 39066 -26988 39118
rect -27092 39054 -26988 39066
rect -27092 39002 -27066 39054
rect -27014 39002 -26988 39054
rect -27092 38990 -26988 39002
rect -27092 38938 -27066 38990
rect -27014 38938 -26988 38990
rect -27092 38926 -26988 38938
rect -27092 38874 -27066 38926
rect -27014 38874 -26988 38926
rect -27092 38862 -26988 38874
rect -27092 38810 -27066 38862
rect -27014 38810 -26988 38862
rect -27092 38798 -26988 38810
rect -27092 38746 -27066 38798
rect -27014 38746 -26988 38798
rect -27092 38734 -26988 38746
rect -27092 38682 -27066 38734
rect -27014 38682 -26988 38734
rect -27092 38670 -26988 38682
rect -27092 38618 -27066 38670
rect -27014 38618 -26988 38670
rect -27092 38606 -26988 38618
rect -27092 38554 -27066 38606
rect -27014 38554 -26988 38606
rect -27092 38542 -26988 38554
rect -27092 38490 -27066 38542
rect -27014 38490 -26988 38542
rect -27092 38478 -26988 38490
rect -27092 38426 -27066 38478
rect -27014 38426 -26988 38478
rect -27092 38414 -26988 38426
rect -29624 38407 -29140 38413
rect -29624 38355 -29600 38407
rect -29548 38355 -29536 38407
rect -29484 38355 -29472 38407
rect -29420 38355 -29408 38407
rect -29356 38355 -29344 38407
rect -29292 38355 -29280 38407
rect -29228 38355 -29216 38407
rect -29164 38355 -29140 38407
rect -29624 38349 -29140 38355
rect -27092 38362 -27066 38414
rect -27014 38362 -26988 38414
rect -27092 38350 -26988 38362
rect -27092 38298 -27066 38350
rect -27014 38298 -26988 38350
rect -27092 38286 -26988 38298
rect -31159 38250 -29704 38256
rect -31159 38242 -31024 38250
rect -31821 38211 -31737 38223
rect -31821 38159 -31805 38211
rect -31753 38159 -31737 38211
rect -31553 38208 -31024 38242
rect -31159 38198 -31024 38208
rect -30972 38198 -30960 38250
rect -30908 38198 -29704 38250
rect -27092 38234 -27066 38286
rect -27014 38234 -26988 38286
rect -27092 38232 -26988 38234
rect -18893 39084 -18871 39136
rect -18819 39084 -18797 39136
rect -18893 39072 -18797 39084
rect -18893 39020 -18871 39072
rect -18819 39020 -18797 39072
rect -18893 39008 -18797 39020
rect -18893 38956 -18871 39008
rect -18819 38956 -18797 39008
rect -18893 38944 -18797 38956
rect -18893 38892 -18871 38944
rect -18819 38892 -18797 38944
rect -18893 38880 -18797 38892
rect -18893 38828 -18871 38880
rect -18819 38828 -18797 38880
rect -18893 38816 -18797 38828
rect -18893 38764 -18871 38816
rect -18819 38764 -18797 38816
rect -18893 38752 -18797 38764
rect -18893 38700 -18871 38752
rect -18819 38700 -18797 38752
rect -18893 38688 -18797 38700
rect -18893 38636 -18871 38688
rect -18819 38636 -18797 38688
rect -18893 38624 -18797 38636
rect -18893 38572 -18871 38624
rect -18819 38572 -18797 38624
rect -18893 38560 -18797 38572
rect -18893 38508 -18871 38560
rect -18819 38508 -18797 38560
rect -18893 38496 -18797 38508
rect -18893 38444 -18871 38496
rect -18819 38444 -18797 38496
rect -18893 38432 -18797 38444
rect -18893 38380 -18871 38432
rect -18819 38380 -18797 38432
rect -18893 38368 -18797 38380
rect -18893 38316 -18871 38368
rect -18819 38316 -18797 38368
rect -18893 38304 -18797 38316
rect -18893 38252 -18871 38304
rect -18819 38252 -18797 38304
rect -18893 38240 -18797 38252
rect -31159 38192 -29704 38198
rect -31821 38141 -31737 38159
rect -18893 38188 -18871 38240
rect -18819 38188 -18797 38240
rect -18893 38176 -18797 38188
rect -18893 38124 -18871 38176
rect -18819 38124 -18797 38176
rect -18893 38112 -18797 38124
rect -18893 38060 -18871 38112
rect -18819 38060 -18797 38112
rect -18893 38048 -18797 38060
rect -18893 37996 -18871 38048
rect -18819 37996 -18797 38048
rect -18893 37984 -18797 37996
rect -18893 37932 -18871 37984
rect -18819 37932 -18797 37984
rect -18893 37920 -18797 37932
rect -18893 37868 -18871 37920
rect -18819 37868 -18797 37920
rect -18893 37856 -18797 37868
rect -18893 37804 -18871 37856
rect -18819 37804 -18797 37856
rect -18893 37792 -18797 37804
rect -18893 37740 -18871 37792
rect -18819 37740 -18797 37792
rect -18893 37728 -18797 37740
rect -18893 37676 -18871 37728
rect -18819 37676 -18797 37728
rect -18893 37664 -18797 37676
rect -18893 37612 -18871 37664
rect -18819 37612 -18797 37664
rect -18893 37600 -18797 37612
rect -35528 37540 -35272 37568
rect -35528 37360 -35490 37540
rect -35310 37475 -35272 37540
rect -18893 37548 -18871 37600
rect -18819 37548 -18797 37600
rect -18893 37536 -18797 37548
rect -18893 37484 -18871 37536
rect -18819 37484 -18797 37536
rect -35310 37469 -29696 37475
rect -35310 37417 -30193 37469
rect -30141 37417 -30129 37469
rect -30077 37417 -29696 37469
rect -35310 37411 -29696 37417
rect -18893 37472 -18797 37484
rect -18893 37420 -18871 37472
rect -18819 37420 -18797 37472
rect -35310 37360 -35272 37411
rect -35528 37332 -35272 37360
rect -18893 37408 -18797 37420
rect -18893 37356 -18871 37408
rect -18819 37356 -18797 37408
rect -27089 37351 -26985 37353
rect -29662 37317 -29133 37323
rect -29662 37265 -29648 37317
rect -29596 37265 -29584 37317
rect -29532 37265 -29520 37317
rect -29468 37265 -29456 37317
rect -29404 37265 -29392 37317
rect -29340 37265 -29328 37317
rect -29276 37265 -29264 37317
rect -29212 37265 -29200 37317
rect -29148 37265 -29133 37317
rect -29662 37259 -29133 37265
rect -27089 37299 -27063 37351
rect -27011 37299 -26985 37351
rect -27089 37287 -26985 37299
rect -27089 37235 -27063 37287
rect -27011 37235 -26985 37287
rect -27089 37223 -26985 37235
rect -27089 37171 -27063 37223
rect -27011 37171 -26985 37223
rect -27089 37159 -26985 37171
rect -27089 37107 -27063 37159
rect -27011 37107 -26985 37159
rect -27089 37095 -26985 37107
rect -27089 37043 -27063 37095
rect -27011 37043 -26985 37095
rect -27089 37031 -26985 37043
rect -27089 36979 -27063 37031
rect -27011 36979 -26985 37031
rect -27089 36967 -26985 36979
rect -27089 36915 -27063 36967
rect -27011 36915 -26985 36967
rect -27089 36903 -26985 36915
rect -27089 36851 -27063 36903
rect -27011 36851 -26985 36903
rect -27089 36839 -26985 36851
rect -27089 36787 -27063 36839
rect -27011 36787 -26985 36839
rect -27089 36775 -26985 36787
rect -27089 36723 -27063 36775
rect -27011 36723 -26985 36775
rect -27089 36711 -26985 36723
rect -27089 36659 -27063 36711
rect -27011 36659 -26985 36711
rect -27089 36647 -26985 36659
rect -27089 36595 -27063 36647
rect -27011 36595 -26985 36647
rect -27089 36583 -26985 36595
rect -27089 36531 -27063 36583
rect -27011 36531 -26985 36583
rect -27089 36519 -26985 36531
rect -27089 36467 -27063 36519
rect -27011 36467 -26985 36519
rect -27089 36465 -26985 36467
rect -18893 37344 -18797 37356
rect -18893 37292 -18871 37344
rect -18819 37292 -18797 37344
rect -18893 37280 -18797 37292
rect -18893 37228 -18871 37280
rect -18819 37228 -18797 37280
rect -18893 37216 -18797 37228
rect -18893 37164 -18871 37216
rect -18819 37164 -18797 37216
rect -18893 37152 -18797 37164
rect -18893 37100 -18871 37152
rect -18819 37100 -18797 37152
rect -18893 37088 -18797 37100
rect -18893 37036 -18871 37088
rect -18819 37036 -18797 37088
rect -18893 37024 -18797 37036
rect -18893 36972 -18871 37024
rect -18819 36972 -18797 37024
rect -18893 36960 -18797 36972
rect -18893 36908 -18871 36960
rect -18819 36908 -18797 36960
rect -18893 36896 -18797 36908
rect -18893 36844 -18871 36896
rect -18819 36844 -18797 36896
rect -18893 36832 -18797 36844
rect -18893 36780 -18871 36832
rect -18819 36780 -18797 36832
rect -18893 36768 -18797 36780
rect -18893 36716 -18871 36768
rect -18819 36716 -18797 36768
rect -18893 36704 -18797 36716
rect -18893 36652 -18871 36704
rect -18819 36652 -18797 36704
rect -18893 36640 -18797 36652
rect -18893 36588 -18871 36640
rect -18819 36588 -18797 36640
rect -18893 36576 -18797 36588
rect -18893 36524 -18871 36576
rect -18819 36524 -18797 36576
rect -18893 36512 -18797 36524
rect -18893 36460 -18871 36512
rect -18819 36460 -18797 36512
rect -18893 36448 -18797 36460
rect -18893 36396 -18871 36448
rect -18819 36396 -18797 36448
rect -18893 36384 -18797 36396
rect -18893 36332 -18871 36384
rect -18819 36332 -18797 36384
rect -18893 36320 -18797 36332
rect -18893 36268 -18871 36320
rect -18819 36268 -18797 36320
rect -18893 36256 -18797 36268
rect -18893 36204 -18871 36256
rect -18819 36204 -18797 36256
rect -18893 36192 -18797 36204
rect -27087 36142 -26986 36160
rect -27087 36090 -27063 36142
rect -27011 36090 -26986 36142
rect -18893 36140 -18871 36192
rect -18819 36140 -18797 36192
rect -18893 36124 -18797 36140
rect -27087 36078 -26986 36090
rect -27087 36026 -27063 36078
rect -27011 36026 -26986 36078
rect -27087 36014 -26986 36026
rect -27087 35962 -27063 36014
rect -27011 35962 -26986 36014
rect -27087 35950 -26986 35962
rect -27087 35898 -27063 35950
rect -27011 35898 -26986 35950
rect -27087 35886 -26986 35898
rect -27087 35834 -27063 35886
rect -27011 35834 -26986 35886
rect -27087 35822 -26986 35834
rect -27087 35770 -27063 35822
rect -27011 35770 -26986 35822
rect -27087 35758 -26986 35770
rect -27087 35706 -27063 35758
rect -27011 35706 -26986 35758
rect -27087 35694 -26986 35706
rect -27087 35642 -27063 35694
rect -27011 35642 -26986 35694
rect -27087 35630 -26986 35642
rect -27087 35578 -27063 35630
rect -27011 35578 -26986 35630
rect -27087 35566 -26986 35578
rect -27087 35514 -27063 35566
rect -27011 35514 -26986 35566
rect -27087 35502 -26986 35514
rect -27087 35450 -27063 35502
rect -27011 35450 -26986 35502
rect -27087 35438 -26986 35450
rect -27087 35386 -27063 35438
rect -27011 35386 -26986 35438
rect -27087 35374 -26986 35386
rect -27087 35322 -27063 35374
rect -27011 35322 -26986 35374
rect -27087 35310 -26986 35322
rect -27087 35258 -27063 35310
rect -27011 35258 -26986 35310
rect -27087 35246 -26986 35258
rect -27087 35194 -27063 35246
rect -27011 35194 -26986 35246
rect -27087 35182 -26986 35194
rect -27087 35130 -27063 35182
rect -27011 35130 -26986 35182
rect -27087 35118 -26986 35130
rect -27087 35066 -27063 35118
rect -27011 35066 -26986 35118
rect -27087 35054 -26986 35066
rect -27087 35002 -27063 35054
rect -27011 35002 -26986 35054
rect -27087 34985 -26986 35002
rect -27089 34664 -26990 34691
rect -27089 34612 -27066 34664
rect -27014 34612 -26990 34664
rect -27089 34600 -26990 34612
rect -27089 34548 -27066 34600
rect -27014 34548 -26990 34600
rect -27089 34536 -26990 34548
rect -27089 34484 -27066 34536
rect -27014 34484 -26990 34536
rect -27089 34472 -26990 34484
rect -27089 34420 -27066 34472
rect -27014 34420 -26990 34472
rect -27089 34408 -26990 34420
rect -27089 34356 -27066 34408
rect -27014 34356 -26990 34408
rect -27089 34344 -26990 34356
rect -27089 34292 -27066 34344
rect -27014 34292 -26990 34344
rect -27089 34280 -26990 34292
rect -27089 34228 -27066 34280
rect -27014 34228 -26990 34280
rect -27089 34216 -26990 34228
rect -27089 34164 -27066 34216
rect -27014 34164 -26990 34216
rect -27089 34152 -26990 34164
rect -27089 34100 -27066 34152
rect -27014 34100 -26990 34152
rect -27089 34088 -26990 34100
rect -27089 34036 -27066 34088
rect -27014 34036 -26990 34088
rect -27089 34024 -26990 34036
rect -27089 33972 -27066 34024
rect -27014 33972 -26990 34024
rect -27089 33960 -26990 33972
rect -27089 33908 -27066 33960
rect -27014 33908 -26990 33960
rect -27089 33896 -26990 33908
rect -27089 33844 -27066 33896
rect -27014 33844 -26990 33896
rect -27089 33832 -26990 33844
rect -27089 33780 -27066 33832
rect -27014 33780 -26990 33832
rect -27089 33768 -26990 33780
rect -27089 33716 -27066 33768
rect -27014 33716 -26990 33768
rect -27089 33704 -26990 33716
rect -27089 33652 -27066 33704
rect -27014 33652 -26990 33704
rect -27089 33640 -26990 33652
rect -27089 33588 -27066 33640
rect -27014 33588 -26990 33640
rect -27089 33576 -26990 33588
rect -27089 33524 -27066 33576
rect -27014 33524 -26990 33576
rect -27089 33498 -26990 33524
rect -27094 32882 -26995 32899
rect -27094 32830 -27071 32882
rect -27019 32830 -26995 32882
rect -27094 32818 -26995 32830
rect -27094 32766 -27071 32818
rect -27019 32766 -26995 32818
rect -27094 32754 -26995 32766
rect -27094 32702 -27071 32754
rect -27019 32702 -26995 32754
rect -27094 32690 -26995 32702
rect -27094 32638 -27071 32690
rect -27019 32638 -26995 32690
rect -27094 32626 -26995 32638
rect -27094 32574 -27071 32626
rect -27019 32574 -26995 32626
rect -27094 32562 -26995 32574
rect -27094 32510 -27071 32562
rect -27019 32510 -26995 32562
rect -27094 32498 -26995 32510
rect -27094 32446 -27071 32498
rect -27019 32446 -26995 32498
rect -27094 32434 -26995 32446
rect -27094 32382 -27071 32434
rect -27019 32382 -26995 32434
rect -27094 32365 -26995 32382
rect -13469 29329 -13405 42997
rect -12703 42392 -12619 42398
rect -12703 42340 -12687 42392
rect -12635 42340 -12619 42392
rect -12703 42334 -12619 42340
rect -12693 29752 -12629 42334
rect -5934 39820 -5913 46272
rect -5733 39820 -5712 46272
rect 10170 46127 10561 46128
rect 334 45843 568 45844
rect 93 45365 157 45366
rect -569 45313 157 45365
rect -5934 39819 -5712 39820
rect -6989 39805 -6861 39806
rect -9408 39799 -9260 39805
rect -9408 39747 -9392 39799
rect -9340 39747 -9328 39799
rect -9276 39747 -9260 39799
rect -9408 39741 -9260 39747
rect -6999 39799 -6851 39805
rect -6999 39747 -6983 39799
rect -6931 39747 -6919 39799
rect -6867 39747 -6851 39799
rect -6999 39741 -6851 39747
rect -9398 34670 -9270 39741
rect -9398 34618 -9363 34670
rect -9311 34618 -9270 34670
rect -9398 30305 -9270 34618
rect -6989 33173 -6861 39741
rect -5694 39666 -5662 39846
rect -170 39666 -138 39846
rect 93 38566 157 45313
rect 334 44319 361 45843
rect 541 44319 568 45843
rect 334 44318 568 44319
rect 342 41381 522 41383
rect 342 39857 374 41381
rect 490 39857 522 41381
rect 7082 41306 7200 43012
rect 342 39855 522 39857
rect 2503 38851 2605 38881
rect 2503 38799 2528 38851
rect 2580 38799 2605 38851
rect 2503 38787 2605 38799
rect 2503 38735 2528 38787
rect 2580 38735 2605 38787
rect 2503 38723 2605 38735
rect 2503 38671 2528 38723
rect 2580 38671 2605 38723
rect 2503 38642 2605 38671
rect 5361 38568 5425 40438
rect 83 38560 167 38566
rect 83 38508 99 38560
rect 151 38508 167 38560
rect 83 38502 167 38508
rect 1220 38560 1304 38566
rect 1220 38508 1236 38560
rect 1288 38508 1304 38560
rect 1220 38502 1304 38508
rect 2439 38562 2700 38568
rect 2439 38510 2632 38562
rect 2684 38510 2700 38562
rect 2439 38504 2700 38510
rect 5351 38562 5435 38568
rect 5351 38510 5367 38562
rect 5419 38510 5435 38562
rect 5351 38504 5435 38510
rect 93 37651 157 38502
rect 2505 38394 2624 38420
rect 2505 38342 2538 38394
rect 2590 38342 2624 38394
rect 2505 38330 2624 38342
rect 2505 38278 2538 38330
rect 2590 38278 2624 38330
rect 2505 38266 2624 38278
rect 2505 38214 2538 38266
rect 2590 38214 2624 38266
rect 2505 38202 2624 38214
rect 2505 38150 2538 38202
rect 2590 38150 2624 38202
rect 5361 38155 5425 38504
rect 2505 38138 2624 38150
rect 2505 38086 2538 38138
rect 2590 38086 2624 38138
rect 5351 38149 5435 38155
rect 5351 38097 5367 38149
rect 5419 38097 5435 38149
rect 5351 38091 5435 38097
rect 2505 38074 2624 38086
rect 2505 38022 2538 38074
rect 2590 38022 2624 38074
rect 2505 37996 2624 38022
rect 83 37645 167 37651
rect 83 37593 99 37645
rect 151 37593 167 37645
rect 83 37587 167 37593
rect 3417 37645 3501 37651
rect 3417 37593 3433 37645
rect 3485 37593 3501 37645
rect 3417 37587 3501 37593
rect 93 36816 157 37587
rect 2634 37201 2718 37207
rect 2634 37149 2650 37201
rect 2702 37149 2718 37201
rect 2158 37145 2242 37149
rect 2158 37093 2174 37145
rect 2226 37093 2242 37145
rect 2634 37143 2718 37149
rect 2158 37081 2242 37093
rect 2158 37029 2174 37081
rect 2226 37029 2242 37081
rect 2158 37017 2242 37029
rect 2158 36965 2174 37017
rect 2226 36965 2242 37017
rect 2158 36953 2242 36965
rect 2158 36901 2174 36953
rect 2226 36901 2242 36953
rect 2158 36898 2242 36901
rect 2644 36816 2708 37143
rect 83 36810 167 36816
rect 83 36758 99 36810
rect 151 36758 167 36810
rect 83 36752 167 36758
rect 873 36810 957 36816
rect 873 36758 889 36810
rect 941 36758 957 36810
rect 873 36752 957 36758
rect 2240 36752 2708 36816
rect 93 36750 157 36752
rect 2159 36645 2243 36668
rect 2159 36593 2175 36645
rect 2227 36593 2243 36645
rect 2159 36581 2243 36593
rect 2159 36529 2175 36581
rect 2227 36529 2243 36581
rect 2159 36517 2243 36529
rect 2159 36465 2175 36517
rect 2227 36465 2243 36517
rect 2159 36453 2243 36465
rect 2159 36401 2175 36453
rect 2227 36401 2243 36453
rect 2159 36389 2243 36401
rect 2159 36337 2175 36389
rect 2227 36337 2243 36389
rect 2159 36325 2243 36337
rect 2159 36273 2175 36325
rect 2227 36273 2243 36325
rect 2159 36250 2243 36273
rect 2928 36085 3353 36088
rect 2928 36033 2954 36085
rect 3006 36033 3018 36085
rect 3070 36033 3082 36085
rect 3134 36033 3146 36085
rect 3198 36033 3210 36085
rect 3262 36033 3274 36085
rect 3326 36033 3353 36085
rect 2928 36030 3353 36033
rect 3427 35950 3491 37587
rect 6701 37207 6765 40449
rect 7082 39210 7318 41306
rect 10170 39867 10211 46127
rect 10519 39867 10561 46127
rect 12542 39210 12778 73019
rect 24656 66701 24892 77876
rect 24750 65741 24796 66701
rect 17420 64738 17506 64743
rect 17420 64686 17437 64738
rect 17489 64686 17506 64738
rect 17420 64674 17506 64686
rect 17420 64622 17437 64674
rect 17489 64622 17506 64674
rect 17420 64610 17506 64622
rect 17420 64558 17437 64610
rect 17489 64558 17506 64610
rect 17420 64546 17506 64558
rect 17420 64494 17437 64546
rect 17489 64494 17506 64546
rect 17420 64482 17506 64494
rect 17420 64430 17437 64482
rect 17489 64430 17506 64482
rect 17420 64418 17506 64430
rect 17420 64366 17437 64418
rect 17489 64366 17506 64418
rect 17420 64354 17506 64366
rect 17420 64302 17437 64354
rect 17489 64302 17506 64354
rect 17420 64290 17506 64302
rect 17420 64238 17437 64290
rect 17489 64238 17506 64290
rect 17420 64226 17506 64238
rect 17420 64174 17437 64226
rect 17489 64174 17506 64226
rect 17420 64169 17506 64174
rect 23948 64738 24034 64743
rect 23948 64686 23965 64738
rect 24017 64686 24034 64738
rect 23948 64674 24034 64686
rect 23948 64622 23965 64674
rect 24017 64622 24034 64674
rect 23948 64610 24034 64622
rect 23948 64558 23965 64610
rect 24017 64558 24034 64610
rect 23948 64546 24034 64558
rect 23948 64494 23965 64546
rect 24017 64494 24034 64546
rect 23948 64482 24034 64494
rect 23948 64430 23965 64482
rect 24017 64430 24034 64482
rect 23948 64418 24034 64430
rect 23948 64366 23965 64418
rect 24017 64366 24034 64418
rect 23948 64354 24034 64366
rect 23948 64302 23965 64354
rect 24017 64302 24034 64354
rect 23948 64290 24034 64302
rect 23948 64238 23965 64290
rect 24017 64238 24034 64290
rect 23948 64226 24034 64238
rect 23948 64174 23965 64226
rect 24017 64174 24034 64226
rect 23948 64169 24034 64174
rect 31564 64738 31650 64743
rect 31564 64686 31581 64738
rect 31633 64686 31650 64738
rect 31564 64674 31650 64686
rect 31564 64622 31581 64674
rect 31633 64622 31650 64674
rect 31564 64610 31650 64622
rect 31564 64558 31581 64610
rect 31633 64558 31650 64610
rect 31564 64546 31650 64558
rect 31564 64494 31581 64546
rect 31633 64494 31650 64546
rect 31564 64482 31650 64494
rect 31564 64430 31581 64482
rect 31633 64430 31650 64482
rect 31564 64418 31650 64430
rect 31564 64366 31581 64418
rect 31633 64366 31650 64418
rect 31564 64354 31650 64366
rect 31564 64302 31581 64354
rect 31633 64302 31650 64354
rect 31564 64290 31650 64302
rect 31564 64238 31581 64290
rect 31633 64238 31650 64290
rect 31564 64226 31650 64238
rect 31564 64174 31581 64226
rect 31633 64174 31650 64226
rect 31564 64169 31650 64174
rect 17965 62735 18051 62740
rect 17965 62683 17982 62735
rect 18034 62683 18051 62735
rect 17965 62671 18051 62683
rect 17965 62619 17982 62671
rect 18034 62619 18051 62671
rect 17965 62607 18051 62619
rect 17965 62555 17982 62607
rect 18034 62555 18051 62607
rect 17965 62543 18051 62555
rect 17965 62491 17982 62543
rect 18034 62491 18051 62543
rect 17965 62479 18051 62491
rect 17965 62427 17982 62479
rect 18034 62427 18051 62479
rect 17965 62415 18051 62427
rect 17965 62363 17982 62415
rect 18034 62363 18051 62415
rect 17965 62351 18051 62363
rect 17965 62299 17982 62351
rect 18034 62299 18051 62351
rect 17965 62287 18051 62299
rect 17965 62235 17982 62287
rect 18034 62235 18051 62287
rect 17965 62223 18051 62235
rect 17965 62171 17982 62223
rect 18034 62171 18051 62223
rect 17965 62166 18051 62171
rect 19053 62735 19139 62740
rect 19053 62683 19070 62735
rect 19122 62683 19139 62735
rect 19053 62671 19139 62683
rect 19053 62619 19070 62671
rect 19122 62619 19139 62671
rect 19053 62607 19139 62619
rect 19053 62555 19070 62607
rect 19122 62555 19139 62607
rect 19053 62543 19139 62555
rect 19053 62491 19070 62543
rect 19122 62491 19139 62543
rect 19053 62479 19139 62491
rect 19053 62427 19070 62479
rect 19122 62427 19139 62479
rect 19053 62415 19139 62427
rect 19053 62363 19070 62415
rect 19122 62363 19139 62415
rect 19053 62351 19139 62363
rect 19053 62299 19070 62351
rect 19122 62299 19139 62351
rect 19053 62287 19139 62299
rect 19053 62235 19070 62287
rect 19122 62235 19139 62287
rect 19053 62223 19139 62235
rect 19053 62171 19070 62223
rect 19122 62171 19139 62223
rect 19053 62166 19139 62171
rect 21229 62735 21315 62740
rect 21229 62683 21246 62735
rect 21298 62683 21315 62735
rect 21229 62671 21315 62683
rect 21229 62619 21246 62671
rect 21298 62619 21315 62671
rect 21229 62607 21315 62619
rect 21229 62555 21246 62607
rect 21298 62555 21315 62607
rect 21229 62543 21315 62555
rect 21229 62491 21246 62543
rect 21298 62491 21315 62543
rect 21229 62479 21315 62491
rect 21229 62427 21246 62479
rect 21298 62427 21315 62479
rect 21229 62415 21315 62427
rect 21229 62363 21246 62415
rect 21298 62363 21315 62415
rect 21229 62351 21315 62363
rect 21229 62299 21246 62351
rect 21298 62299 21315 62351
rect 21229 62287 21315 62299
rect 21229 62235 21246 62287
rect 21298 62235 21315 62287
rect 21229 62223 21315 62235
rect 21229 62171 21246 62223
rect 21298 62171 21315 62223
rect 21229 62166 21315 62171
rect 22317 62735 22403 62740
rect 22317 62683 22334 62735
rect 22386 62683 22403 62735
rect 22317 62671 22403 62683
rect 22317 62619 22334 62671
rect 22386 62619 22403 62671
rect 22317 62607 22403 62619
rect 22317 62555 22334 62607
rect 22386 62555 22403 62607
rect 22317 62543 22403 62555
rect 22317 62491 22334 62543
rect 22386 62491 22403 62543
rect 22317 62479 22403 62491
rect 22317 62427 22334 62479
rect 22386 62427 22403 62479
rect 22317 62415 22403 62427
rect 22317 62363 22334 62415
rect 22386 62363 22403 62415
rect 22317 62351 22403 62363
rect 22317 62299 22334 62351
rect 22386 62299 22403 62351
rect 22317 62287 22403 62299
rect 22317 62235 22334 62287
rect 22386 62235 22403 62287
rect 22317 62223 22403 62235
rect 22317 62171 22334 62223
rect 22386 62171 22403 62223
rect 22317 62166 22403 62171
rect 23405 62735 23491 62740
rect 23405 62683 23422 62735
rect 23474 62683 23491 62735
rect 23405 62671 23491 62683
rect 23405 62619 23422 62671
rect 23474 62619 23491 62671
rect 23405 62607 23491 62619
rect 23405 62555 23422 62607
rect 23474 62555 23491 62607
rect 23405 62543 23491 62555
rect 23405 62491 23422 62543
rect 23474 62491 23491 62543
rect 23405 62479 23491 62491
rect 23405 62427 23422 62479
rect 23474 62427 23491 62479
rect 23405 62415 23491 62427
rect 23405 62363 23422 62415
rect 23474 62363 23491 62415
rect 23405 62351 23491 62363
rect 23405 62299 23422 62351
rect 23474 62299 23491 62351
rect 23405 62287 23491 62299
rect 23405 62235 23422 62287
rect 23474 62235 23491 62287
rect 23405 62223 23491 62235
rect 23405 62171 23422 62223
rect 23474 62171 23491 62223
rect 23405 62166 23491 62171
rect 24493 62735 24579 62740
rect 24493 62683 24510 62735
rect 24562 62683 24579 62735
rect 24493 62671 24579 62683
rect 24493 62619 24510 62671
rect 24562 62619 24579 62671
rect 24493 62607 24579 62619
rect 24493 62555 24510 62607
rect 24562 62555 24579 62607
rect 24493 62543 24579 62555
rect 24493 62491 24510 62543
rect 24562 62491 24579 62543
rect 24493 62479 24579 62491
rect 24493 62427 24510 62479
rect 24562 62427 24579 62479
rect 24493 62415 24579 62427
rect 24493 62363 24510 62415
rect 24562 62363 24579 62415
rect 24493 62351 24579 62363
rect 24493 62299 24510 62351
rect 24562 62299 24579 62351
rect 24493 62287 24579 62299
rect 24493 62235 24510 62287
rect 24562 62235 24579 62287
rect 24493 62223 24579 62235
rect 24493 62171 24510 62223
rect 24562 62171 24579 62223
rect 24493 62166 24579 62171
rect 25581 62735 25667 62740
rect 25581 62683 25598 62735
rect 25650 62683 25667 62735
rect 25581 62671 25667 62683
rect 25581 62619 25598 62671
rect 25650 62619 25667 62671
rect 25581 62607 25667 62619
rect 25581 62555 25598 62607
rect 25650 62555 25667 62607
rect 25581 62543 25667 62555
rect 25581 62491 25598 62543
rect 25650 62491 25667 62543
rect 25581 62479 25667 62491
rect 25581 62427 25598 62479
rect 25650 62427 25667 62479
rect 25581 62415 25667 62427
rect 25581 62363 25598 62415
rect 25650 62363 25667 62415
rect 25581 62351 25667 62363
rect 25581 62299 25598 62351
rect 25650 62299 25667 62351
rect 25581 62287 25667 62299
rect 25581 62235 25598 62287
rect 25650 62235 25667 62287
rect 25581 62223 25667 62235
rect 25581 62171 25598 62223
rect 25650 62171 25667 62223
rect 25581 62166 25667 62171
rect 26669 62735 26755 62740
rect 26669 62683 26686 62735
rect 26738 62683 26755 62735
rect 26669 62671 26755 62683
rect 26669 62619 26686 62671
rect 26738 62619 26755 62671
rect 26669 62607 26755 62619
rect 26669 62555 26686 62607
rect 26738 62555 26755 62607
rect 26669 62543 26755 62555
rect 26669 62491 26686 62543
rect 26738 62491 26755 62543
rect 26669 62479 26755 62491
rect 26669 62427 26686 62479
rect 26738 62427 26755 62479
rect 26669 62415 26755 62427
rect 26669 62363 26686 62415
rect 26738 62363 26755 62415
rect 26669 62351 26755 62363
rect 26669 62299 26686 62351
rect 26738 62299 26755 62351
rect 26669 62287 26755 62299
rect 26669 62235 26686 62287
rect 26738 62235 26755 62287
rect 26669 62223 26755 62235
rect 26669 62171 26686 62223
rect 26738 62171 26755 62223
rect 26669 62166 26755 62171
rect 28845 62735 28931 62740
rect 28845 62683 28862 62735
rect 28914 62683 28931 62735
rect 28845 62671 28931 62683
rect 28845 62619 28862 62671
rect 28914 62619 28931 62671
rect 28845 62607 28931 62619
rect 28845 62555 28862 62607
rect 28914 62555 28931 62607
rect 28845 62543 28931 62555
rect 28845 62491 28862 62543
rect 28914 62491 28931 62543
rect 28845 62479 28931 62491
rect 28845 62427 28862 62479
rect 28914 62427 28931 62479
rect 28845 62415 28931 62427
rect 28845 62363 28862 62415
rect 28914 62363 28931 62415
rect 28845 62351 28931 62363
rect 28845 62299 28862 62351
rect 28914 62299 28931 62351
rect 28845 62287 28931 62299
rect 28845 62235 28862 62287
rect 28914 62235 28931 62287
rect 28845 62223 28931 62235
rect 28845 62171 28862 62223
rect 28914 62171 28931 62223
rect 28845 62166 28931 62171
rect 29933 62735 30019 62740
rect 29933 62683 29950 62735
rect 30002 62683 30019 62735
rect 29933 62671 30019 62683
rect 29933 62619 29950 62671
rect 30002 62619 30019 62671
rect 29933 62607 30019 62619
rect 29933 62555 29950 62607
rect 30002 62555 30019 62607
rect 29933 62543 30019 62555
rect 29933 62491 29950 62543
rect 30002 62491 30019 62543
rect 29933 62479 30019 62491
rect 29933 62427 29950 62479
rect 30002 62427 30019 62479
rect 29933 62415 30019 62427
rect 29933 62363 29950 62415
rect 30002 62363 30019 62415
rect 29933 62351 30019 62363
rect 29933 62299 29950 62351
rect 30002 62299 30019 62351
rect 29933 62287 30019 62299
rect 29933 62235 29950 62287
rect 30002 62235 30019 62287
rect 29933 62223 30019 62235
rect 29933 62171 29950 62223
rect 30002 62171 30019 62223
rect 29933 62166 30019 62171
rect 31021 62735 31107 62740
rect 31021 62683 31038 62735
rect 31090 62683 31107 62735
rect 31021 62671 31107 62683
rect 31021 62619 31038 62671
rect 31090 62619 31107 62671
rect 31021 62607 31107 62619
rect 31021 62555 31038 62607
rect 31090 62555 31107 62607
rect 31021 62543 31107 62555
rect 31021 62491 31038 62543
rect 31090 62491 31107 62543
rect 31021 62479 31107 62491
rect 31021 62427 31038 62479
rect 31090 62427 31107 62479
rect 31021 62415 31107 62427
rect 31021 62363 31038 62415
rect 31090 62363 31107 62415
rect 31021 62351 31107 62363
rect 31021 62299 31038 62351
rect 31090 62299 31107 62351
rect 31021 62287 31107 62299
rect 31021 62235 31038 62287
rect 31090 62235 31107 62287
rect 31021 62223 31107 62235
rect 31021 62171 31038 62223
rect 31090 62171 31107 62223
rect 31021 62166 31107 62171
rect 17420 60738 17506 60743
rect 17420 60686 17437 60738
rect 17489 60686 17506 60738
rect 17420 60674 17506 60686
rect 17420 60622 17437 60674
rect 17489 60622 17506 60674
rect 17420 60610 17506 60622
rect 17420 60558 17437 60610
rect 17489 60558 17506 60610
rect 17420 60546 17506 60558
rect 17420 60494 17437 60546
rect 17489 60494 17506 60546
rect 17420 60482 17506 60494
rect 17420 60430 17437 60482
rect 17489 60430 17506 60482
rect 17420 60418 17506 60430
rect 17420 60366 17437 60418
rect 17489 60366 17506 60418
rect 17420 60354 17506 60366
rect 17420 60302 17437 60354
rect 17489 60302 17506 60354
rect 17420 60290 17506 60302
rect 17420 60238 17437 60290
rect 17489 60238 17506 60290
rect 17420 60226 17506 60238
rect 17420 60174 17437 60226
rect 17489 60174 17506 60226
rect 17420 60169 17506 60174
rect 18508 60738 18594 60743
rect 18508 60686 18525 60738
rect 18577 60686 18594 60738
rect 18508 60674 18594 60686
rect 18508 60622 18525 60674
rect 18577 60622 18594 60674
rect 18508 60610 18594 60622
rect 18508 60558 18525 60610
rect 18577 60558 18594 60610
rect 18508 60546 18594 60558
rect 18508 60494 18525 60546
rect 18577 60494 18594 60546
rect 18508 60482 18594 60494
rect 18508 60430 18525 60482
rect 18577 60430 18594 60482
rect 18508 60418 18594 60430
rect 18508 60366 18525 60418
rect 18577 60366 18594 60418
rect 18508 60354 18594 60366
rect 18508 60302 18525 60354
rect 18577 60302 18594 60354
rect 18508 60290 18594 60302
rect 18508 60238 18525 60290
rect 18577 60238 18594 60290
rect 18508 60226 18594 60238
rect 18508 60174 18525 60226
rect 18577 60174 18594 60226
rect 18508 60169 18594 60174
rect 19596 60738 19682 60743
rect 19596 60686 19613 60738
rect 19665 60686 19682 60738
rect 19596 60674 19682 60686
rect 19596 60622 19613 60674
rect 19665 60622 19682 60674
rect 19596 60610 19682 60622
rect 19596 60558 19613 60610
rect 19665 60558 19682 60610
rect 19596 60546 19682 60558
rect 19596 60494 19613 60546
rect 19665 60494 19682 60546
rect 19596 60482 19682 60494
rect 19596 60430 19613 60482
rect 19665 60430 19682 60482
rect 19596 60418 19682 60430
rect 19596 60366 19613 60418
rect 19665 60366 19682 60418
rect 19596 60354 19682 60366
rect 19596 60302 19613 60354
rect 19665 60302 19682 60354
rect 19596 60290 19682 60302
rect 19596 60238 19613 60290
rect 19665 60238 19682 60290
rect 19596 60226 19682 60238
rect 19596 60174 19613 60226
rect 19665 60174 19682 60226
rect 19596 60169 19682 60174
rect 20684 60738 20770 60743
rect 20684 60686 20701 60738
rect 20753 60686 20770 60738
rect 20684 60674 20770 60686
rect 20684 60622 20701 60674
rect 20753 60622 20770 60674
rect 20684 60610 20770 60622
rect 20684 60558 20701 60610
rect 20753 60558 20770 60610
rect 20684 60546 20770 60558
rect 20684 60494 20701 60546
rect 20753 60494 20770 60546
rect 20684 60482 20770 60494
rect 20684 60430 20701 60482
rect 20753 60430 20770 60482
rect 20684 60418 20770 60430
rect 20684 60366 20701 60418
rect 20753 60366 20770 60418
rect 20684 60354 20770 60366
rect 20684 60302 20701 60354
rect 20753 60302 20770 60354
rect 20684 60290 20770 60302
rect 20684 60238 20701 60290
rect 20753 60238 20770 60290
rect 20684 60226 20770 60238
rect 20684 60174 20701 60226
rect 20753 60174 20770 60226
rect 20684 60169 20770 60174
rect 21772 60738 21858 60743
rect 21772 60686 21789 60738
rect 21841 60686 21858 60738
rect 21772 60674 21858 60686
rect 21772 60622 21789 60674
rect 21841 60622 21858 60674
rect 21772 60610 21858 60622
rect 21772 60558 21789 60610
rect 21841 60558 21858 60610
rect 21772 60546 21858 60558
rect 21772 60494 21789 60546
rect 21841 60494 21858 60546
rect 21772 60482 21858 60494
rect 21772 60430 21789 60482
rect 21841 60430 21858 60482
rect 21772 60418 21858 60430
rect 21772 60366 21789 60418
rect 21841 60366 21858 60418
rect 21772 60354 21858 60366
rect 21772 60302 21789 60354
rect 21841 60302 21858 60354
rect 21772 60290 21858 60302
rect 21772 60238 21789 60290
rect 21841 60238 21858 60290
rect 21772 60226 21858 60238
rect 21772 60174 21789 60226
rect 21841 60174 21858 60226
rect 21772 60169 21858 60174
rect 22860 60738 22946 60743
rect 22860 60686 22877 60738
rect 22929 60686 22946 60738
rect 22860 60674 22946 60686
rect 22860 60622 22877 60674
rect 22929 60622 22946 60674
rect 22860 60610 22946 60622
rect 22860 60558 22877 60610
rect 22929 60558 22946 60610
rect 22860 60546 22946 60558
rect 22860 60494 22877 60546
rect 22929 60494 22946 60546
rect 22860 60482 22946 60494
rect 22860 60430 22877 60482
rect 22929 60430 22946 60482
rect 22860 60418 22946 60430
rect 22860 60366 22877 60418
rect 22929 60366 22946 60418
rect 22860 60354 22946 60366
rect 22860 60302 22877 60354
rect 22929 60302 22946 60354
rect 22860 60290 22946 60302
rect 22860 60238 22877 60290
rect 22929 60238 22946 60290
rect 22860 60226 22946 60238
rect 22860 60174 22877 60226
rect 22929 60174 22946 60226
rect 22860 60169 22946 60174
rect 23948 60738 24034 60743
rect 23948 60686 23965 60738
rect 24017 60686 24034 60738
rect 23948 60674 24034 60686
rect 23948 60622 23965 60674
rect 24017 60622 24034 60674
rect 23948 60610 24034 60622
rect 23948 60558 23965 60610
rect 24017 60558 24034 60610
rect 23948 60546 24034 60558
rect 23948 60494 23965 60546
rect 24017 60494 24034 60546
rect 23948 60482 24034 60494
rect 23948 60430 23965 60482
rect 24017 60430 24034 60482
rect 23948 60418 24034 60430
rect 23948 60366 23965 60418
rect 24017 60366 24034 60418
rect 23948 60354 24034 60366
rect 23948 60302 23965 60354
rect 24017 60302 24034 60354
rect 23948 60290 24034 60302
rect 23948 60238 23965 60290
rect 24017 60238 24034 60290
rect 23948 60226 24034 60238
rect 23948 60174 23965 60226
rect 24017 60174 24034 60226
rect 23948 60169 24034 60174
rect 25036 60738 25122 60743
rect 25036 60686 25053 60738
rect 25105 60686 25122 60738
rect 25036 60674 25122 60686
rect 25036 60622 25053 60674
rect 25105 60622 25122 60674
rect 25036 60610 25122 60622
rect 25036 60558 25053 60610
rect 25105 60558 25122 60610
rect 25036 60546 25122 60558
rect 25036 60494 25053 60546
rect 25105 60494 25122 60546
rect 25036 60482 25122 60494
rect 25036 60430 25053 60482
rect 25105 60430 25122 60482
rect 25036 60418 25122 60430
rect 25036 60366 25053 60418
rect 25105 60366 25122 60418
rect 25036 60354 25122 60366
rect 25036 60302 25053 60354
rect 25105 60302 25122 60354
rect 25036 60290 25122 60302
rect 25036 60238 25053 60290
rect 25105 60238 25122 60290
rect 25036 60226 25122 60238
rect 25036 60174 25053 60226
rect 25105 60174 25122 60226
rect 25036 60169 25122 60174
rect 26124 60738 26210 60743
rect 26124 60686 26141 60738
rect 26193 60686 26210 60738
rect 26124 60674 26210 60686
rect 26124 60622 26141 60674
rect 26193 60622 26210 60674
rect 26124 60610 26210 60622
rect 26124 60558 26141 60610
rect 26193 60558 26210 60610
rect 26124 60546 26210 60558
rect 26124 60494 26141 60546
rect 26193 60494 26210 60546
rect 26124 60482 26210 60494
rect 26124 60430 26141 60482
rect 26193 60430 26210 60482
rect 26124 60418 26210 60430
rect 26124 60366 26141 60418
rect 26193 60366 26210 60418
rect 26124 60354 26210 60366
rect 26124 60302 26141 60354
rect 26193 60302 26210 60354
rect 26124 60290 26210 60302
rect 26124 60238 26141 60290
rect 26193 60238 26210 60290
rect 26124 60226 26210 60238
rect 26124 60174 26141 60226
rect 26193 60174 26210 60226
rect 26124 60169 26210 60174
rect 27212 60738 27298 60743
rect 27212 60686 27229 60738
rect 27281 60686 27298 60738
rect 27212 60674 27298 60686
rect 27212 60622 27229 60674
rect 27281 60622 27298 60674
rect 27212 60610 27298 60622
rect 27212 60558 27229 60610
rect 27281 60558 27298 60610
rect 27212 60546 27298 60558
rect 27212 60494 27229 60546
rect 27281 60494 27298 60546
rect 27212 60482 27298 60494
rect 27212 60430 27229 60482
rect 27281 60430 27298 60482
rect 27212 60418 27298 60430
rect 27212 60366 27229 60418
rect 27281 60366 27298 60418
rect 27212 60354 27298 60366
rect 27212 60302 27229 60354
rect 27281 60302 27298 60354
rect 27212 60290 27298 60302
rect 27212 60238 27229 60290
rect 27281 60238 27298 60290
rect 27212 60226 27298 60238
rect 27212 60174 27229 60226
rect 27281 60174 27298 60226
rect 27212 60169 27298 60174
rect 28300 60738 28386 60743
rect 28300 60686 28317 60738
rect 28369 60686 28386 60738
rect 28300 60674 28386 60686
rect 28300 60622 28317 60674
rect 28369 60622 28386 60674
rect 28300 60610 28386 60622
rect 28300 60558 28317 60610
rect 28369 60558 28386 60610
rect 28300 60546 28386 60558
rect 28300 60494 28317 60546
rect 28369 60494 28386 60546
rect 28300 60482 28386 60494
rect 28300 60430 28317 60482
rect 28369 60430 28386 60482
rect 28300 60418 28386 60430
rect 28300 60366 28317 60418
rect 28369 60366 28386 60418
rect 28300 60354 28386 60366
rect 28300 60302 28317 60354
rect 28369 60302 28386 60354
rect 28300 60290 28386 60302
rect 28300 60238 28317 60290
rect 28369 60238 28386 60290
rect 28300 60226 28386 60238
rect 28300 60174 28317 60226
rect 28369 60174 28386 60226
rect 28300 60169 28386 60174
rect 29388 60738 29474 60743
rect 29388 60686 29405 60738
rect 29457 60686 29474 60738
rect 29388 60674 29474 60686
rect 29388 60622 29405 60674
rect 29457 60622 29474 60674
rect 29388 60610 29474 60622
rect 29388 60558 29405 60610
rect 29457 60558 29474 60610
rect 29388 60546 29474 60558
rect 29388 60494 29405 60546
rect 29457 60494 29474 60546
rect 29388 60482 29474 60494
rect 29388 60430 29405 60482
rect 29457 60430 29474 60482
rect 29388 60418 29474 60430
rect 29388 60366 29405 60418
rect 29457 60366 29474 60418
rect 29388 60354 29474 60366
rect 29388 60302 29405 60354
rect 29457 60302 29474 60354
rect 29388 60290 29474 60302
rect 29388 60238 29405 60290
rect 29457 60238 29474 60290
rect 29388 60226 29474 60238
rect 29388 60174 29405 60226
rect 29457 60174 29474 60226
rect 29388 60169 29474 60174
rect 30476 60738 30562 60743
rect 30476 60686 30493 60738
rect 30545 60686 30562 60738
rect 30476 60674 30562 60686
rect 30476 60622 30493 60674
rect 30545 60622 30562 60674
rect 30476 60610 30562 60622
rect 30476 60558 30493 60610
rect 30545 60558 30562 60610
rect 30476 60546 30562 60558
rect 30476 60494 30493 60546
rect 30545 60494 30562 60546
rect 30476 60482 30562 60494
rect 30476 60430 30493 60482
rect 30545 60430 30562 60482
rect 30476 60418 30562 60430
rect 30476 60366 30493 60418
rect 30545 60366 30562 60418
rect 30476 60354 30562 60366
rect 30476 60302 30493 60354
rect 30545 60302 30562 60354
rect 30476 60290 30562 60302
rect 30476 60238 30493 60290
rect 30545 60238 30562 60290
rect 30476 60226 30562 60238
rect 30476 60174 30493 60226
rect 30545 60174 30562 60226
rect 30476 60169 30562 60174
rect 31564 60738 31650 60743
rect 31564 60686 31581 60738
rect 31633 60686 31650 60738
rect 31564 60674 31650 60686
rect 31564 60622 31581 60674
rect 31633 60622 31650 60674
rect 31564 60610 31650 60622
rect 31564 60558 31581 60610
rect 31633 60558 31650 60610
rect 31564 60546 31650 60558
rect 31564 60494 31581 60546
rect 31633 60494 31650 60546
rect 31564 60482 31650 60494
rect 31564 60430 31581 60482
rect 31633 60430 31650 60482
rect 31564 60418 31650 60430
rect 31564 60366 31581 60418
rect 31633 60366 31650 60418
rect 31564 60354 31650 60366
rect 31564 60302 31581 60354
rect 31633 60302 31650 60354
rect 31564 60290 31650 60302
rect 31564 60238 31581 60290
rect 31633 60238 31650 60290
rect 31564 60226 31650 60238
rect 31564 60174 31581 60226
rect 31633 60174 31650 60226
rect 31564 60169 31650 60174
rect 17965 58735 18051 58740
rect 17965 58683 17982 58735
rect 18034 58683 18051 58735
rect 17965 58671 18051 58683
rect 17965 58619 17982 58671
rect 18034 58619 18051 58671
rect 17965 58607 18051 58619
rect 17965 58555 17982 58607
rect 18034 58555 18051 58607
rect 17965 58543 18051 58555
rect 17965 58491 17982 58543
rect 18034 58491 18051 58543
rect 17965 58479 18051 58491
rect 17965 58427 17982 58479
rect 18034 58427 18051 58479
rect 17965 58415 18051 58427
rect 17965 58363 17982 58415
rect 18034 58363 18051 58415
rect 17965 58351 18051 58363
rect 17965 58299 17982 58351
rect 18034 58299 18051 58351
rect 17965 58287 18051 58299
rect 17965 58235 17982 58287
rect 18034 58235 18051 58287
rect 17965 58223 18051 58235
rect 17965 58171 17982 58223
rect 18034 58171 18051 58223
rect 17965 58166 18051 58171
rect 19053 58735 19139 58740
rect 19053 58683 19070 58735
rect 19122 58683 19139 58735
rect 19053 58671 19139 58683
rect 19053 58619 19070 58671
rect 19122 58619 19139 58671
rect 19053 58607 19139 58619
rect 19053 58555 19070 58607
rect 19122 58555 19139 58607
rect 19053 58543 19139 58555
rect 19053 58491 19070 58543
rect 19122 58491 19139 58543
rect 19053 58479 19139 58491
rect 19053 58427 19070 58479
rect 19122 58427 19139 58479
rect 19053 58415 19139 58427
rect 19053 58363 19070 58415
rect 19122 58363 19139 58415
rect 19053 58351 19139 58363
rect 19053 58299 19070 58351
rect 19122 58299 19139 58351
rect 19053 58287 19139 58299
rect 19053 58235 19070 58287
rect 19122 58235 19139 58287
rect 19053 58223 19139 58235
rect 19053 58171 19070 58223
rect 19122 58171 19139 58223
rect 19053 58166 19139 58171
rect 20141 58735 20227 58740
rect 20141 58683 20158 58735
rect 20210 58683 20227 58735
rect 20141 58671 20227 58683
rect 20141 58619 20158 58671
rect 20210 58619 20227 58671
rect 20141 58607 20227 58619
rect 20141 58555 20158 58607
rect 20210 58555 20227 58607
rect 20141 58543 20227 58555
rect 20141 58491 20158 58543
rect 20210 58491 20227 58543
rect 20141 58479 20227 58491
rect 20141 58427 20158 58479
rect 20210 58427 20227 58479
rect 20141 58415 20227 58427
rect 20141 58363 20158 58415
rect 20210 58363 20227 58415
rect 20141 58351 20227 58363
rect 20141 58299 20158 58351
rect 20210 58299 20227 58351
rect 20141 58287 20227 58299
rect 20141 58235 20158 58287
rect 20210 58235 20227 58287
rect 20141 58223 20227 58235
rect 20141 58171 20158 58223
rect 20210 58171 20227 58223
rect 20141 58166 20227 58171
rect 21229 58735 21315 58740
rect 21229 58683 21246 58735
rect 21298 58683 21315 58735
rect 21229 58671 21315 58683
rect 21229 58619 21246 58671
rect 21298 58619 21315 58671
rect 21229 58607 21315 58619
rect 21229 58555 21246 58607
rect 21298 58555 21315 58607
rect 21229 58543 21315 58555
rect 21229 58491 21246 58543
rect 21298 58491 21315 58543
rect 21229 58479 21315 58491
rect 21229 58427 21246 58479
rect 21298 58427 21315 58479
rect 21229 58415 21315 58427
rect 21229 58363 21246 58415
rect 21298 58363 21315 58415
rect 21229 58351 21315 58363
rect 21229 58299 21246 58351
rect 21298 58299 21315 58351
rect 21229 58287 21315 58299
rect 21229 58235 21246 58287
rect 21298 58235 21315 58287
rect 21229 58223 21315 58235
rect 21229 58171 21246 58223
rect 21298 58171 21315 58223
rect 21229 58166 21315 58171
rect 22317 58735 22403 58740
rect 22317 58683 22334 58735
rect 22386 58683 22403 58735
rect 22317 58671 22403 58683
rect 22317 58619 22334 58671
rect 22386 58619 22403 58671
rect 22317 58607 22403 58619
rect 22317 58555 22334 58607
rect 22386 58555 22403 58607
rect 22317 58543 22403 58555
rect 22317 58491 22334 58543
rect 22386 58491 22403 58543
rect 22317 58479 22403 58491
rect 22317 58427 22334 58479
rect 22386 58427 22403 58479
rect 22317 58415 22403 58427
rect 22317 58363 22334 58415
rect 22386 58363 22403 58415
rect 22317 58351 22403 58363
rect 22317 58299 22334 58351
rect 22386 58299 22403 58351
rect 22317 58287 22403 58299
rect 22317 58235 22334 58287
rect 22386 58235 22403 58287
rect 22317 58223 22403 58235
rect 22317 58171 22334 58223
rect 22386 58171 22403 58223
rect 22317 58166 22403 58171
rect 23405 58735 23491 58740
rect 23405 58683 23422 58735
rect 23474 58683 23491 58735
rect 23405 58671 23491 58683
rect 23405 58619 23422 58671
rect 23474 58619 23491 58671
rect 23405 58607 23491 58619
rect 23405 58555 23422 58607
rect 23474 58555 23491 58607
rect 23405 58543 23491 58555
rect 23405 58491 23422 58543
rect 23474 58491 23491 58543
rect 23405 58479 23491 58491
rect 23405 58427 23422 58479
rect 23474 58427 23491 58479
rect 23405 58415 23491 58427
rect 23405 58363 23422 58415
rect 23474 58363 23491 58415
rect 23405 58351 23491 58363
rect 23405 58299 23422 58351
rect 23474 58299 23491 58351
rect 23405 58287 23491 58299
rect 23405 58235 23422 58287
rect 23474 58235 23491 58287
rect 23405 58223 23491 58235
rect 23405 58171 23422 58223
rect 23474 58171 23491 58223
rect 23405 58166 23491 58171
rect 24493 58735 24579 58740
rect 24493 58683 24510 58735
rect 24562 58683 24579 58735
rect 24493 58671 24579 58683
rect 24493 58619 24510 58671
rect 24562 58619 24579 58671
rect 24493 58607 24579 58619
rect 24493 58555 24510 58607
rect 24562 58555 24579 58607
rect 24493 58543 24579 58555
rect 24493 58491 24510 58543
rect 24562 58491 24579 58543
rect 24493 58479 24579 58491
rect 24493 58427 24510 58479
rect 24562 58427 24579 58479
rect 24493 58415 24579 58427
rect 24493 58363 24510 58415
rect 24562 58363 24579 58415
rect 24493 58351 24579 58363
rect 24493 58299 24510 58351
rect 24562 58299 24579 58351
rect 24493 58287 24579 58299
rect 24493 58235 24510 58287
rect 24562 58235 24579 58287
rect 24493 58223 24579 58235
rect 24493 58171 24510 58223
rect 24562 58171 24579 58223
rect 24493 58166 24579 58171
rect 25581 58735 25667 58740
rect 25581 58683 25598 58735
rect 25650 58683 25667 58735
rect 25581 58671 25667 58683
rect 25581 58619 25598 58671
rect 25650 58619 25667 58671
rect 25581 58607 25667 58619
rect 25581 58555 25598 58607
rect 25650 58555 25667 58607
rect 25581 58543 25667 58555
rect 25581 58491 25598 58543
rect 25650 58491 25667 58543
rect 25581 58479 25667 58491
rect 25581 58427 25598 58479
rect 25650 58427 25667 58479
rect 25581 58415 25667 58427
rect 25581 58363 25598 58415
rect 25650 58363 25667 58415
rect 25581 58351 25667 58363
rect 25581 58299 25598 58351
rect 25650 58299 25667 58351
rect 25581 58287 25667 58299
rect 25581 58235 25598 58287
rect 25650 58235 25667 58287
rect 25581 58223 25667 58235
rect 25581 58171 25598 58223
rect 25650 58171 25667 58223
rect 25581 58166 25667 58171
rect 26669 58735 26755 58740
rect 26669 58683 26686 58735
rect 26738 58683 26755 58735
rect 26669 58671 26755 58683
rect 26669 58619 26686 58671
rect 26738 58619 26755 58671
rect 26669 58607 26755 58619
rect 26669 58555 26686 58607
rect 26738 58555 26755 58607
rect 26669 58543 26755 58555
rect 26669 58491 26686 58543
rect 26738 58491 26755 58543
rect 26669 58479 26755 58491
rect 26669 58427 26686 58479
rect 26738 58427 26755 58479
rect 26669 58415 26755 58427
rect 26669 58363 26686 58415
rect 26738 58363 26755 58415
rect 26669 58351 26755 58363
rect 26669 58299 26686 58351
rect 26738 58299 26755 58351
rect 26669 58287 26755 58299
rect 26669 58235 26686 58287
rect 26738 58235 26755 58287
rect 26669 58223 26755 58235
rect 26669 58171 26686 58223
rect 26738 58171 26755 58223
rect 26669 58166 26755 58171
rect 27757 58735 27843 58740
rect 27757 58683 27774 58735
rect 27826 58683 27843 58735
rect 27757 58671 27843 58683
rect 27757 58619 27774 58671
rect 27826 58619 27843 58671
rect 27757 58607 27843 58619
rect 27757 58555 27774 58607
rect 27826 58555 27843 58607
rect 27757 58543 27843 58555
rect 27757 58491 27774 58543
rect 27826 58491 27843 58543
rect 27757 58479 27843 58491
rect 27757 58427 27774 58479
rect 27826 58427 27843 58479
rect 27757 58415 27843 58427
rect 27757 58363 27774 58415
rect 27826 58363 27843 58415
rect 27757 58351 27843 58363
rect 27757 58299 27774 58351
rect 27826 58299 27843 58351
rect 27757 58287 27843 58299
rect 27757 58235 27774 58287
rect 27826 58235 27843 58287
rect 27757 58223 27843 58235
rect 27757 58171 27774 58223
rect 27826 58171 27843 58223
rect 27757 58166 27843 58171
rect 28845 58735 28931 58740
rect 28845 58683 28862 58735
rect 28914 58683 28931 58735
rect 28845 58671 28931 58683
rect 28845 58619 28862 58671
rect 28914 58619 28931 58671
rect 28845 58607 28931 58619
rect 28845 58555 28862 58607
rect 28914 58555 28931 58607
rect 28845 58543 28931 58555
rect 28845 58491 28862 58543
rect 28914 58491 28931 58543
rect 28845 58479 28931 58491
rect 28845 58427 28862 58479
rect 28914 58427 28931 58479
rect 28845 58415 28931 58427
rect 28845 58363 28862 58415
rect 28914 58363 28931 58415
rect 28845 58351 28931 58363
rect 28845 58299 28862 58351
rect 28914 58299 28931 58351
rect 28845 58287 28931 58299
rect 28845 58235 28862 58287
rect 28914 58235 28931 58287
rect 28845 58223 28931 58235
rect 28845 58171 28862 58223
rect 28914 58171 28931 58223
rect 28845 58166 28931 58171
rect 29933 58735 30019 58740
rect 29933 58683 29950 58735
rect 30002 58683 30019 58735
rect 29933 58671 30019 58683
rect 29933 58619 29950 58671
rect 30002 58619 30019 58671
rect 29933 58607 30019 58619
rect 29933 58555 29950 58607
rect 30002 58555 30019 58607
rect 29933 58543 30019 58555
rect 29933 58491 29950 58543
rect 30002 58491 30019 58543
rect 29933 58479 30019 58491
rect 29933 58427 29950 58479
rect 30002 58427 30019 58479
rect 29933 58415 30019 58427
rect 29933 58363 29950 58415
rect 30002 58363 30019 58415
rect 29933 58351 30019 58363
rect 29933 58299 29950 58351
rect 30002 58299 30019 58351
rect 29933 58287 30019 58299
rect 29933 58235 29950 58287
rect 30002 58235 30019 58287
rect 29933 58223 30019 58235
rect 29933 58171 29950 58223
rect 30002 58171 30019 58223
rect 29933 58166 30019 58171
rect 31021 58735 31107 58740
rect 31021 58683 31038 58735
rect 31090 58683 31107 58735
rect 31021 58671 31107 58683
rect 31021 58619 31038 58671
rect 31090 58619 31107 58671
rect 31021 58607 31107 58619
rect 31021 58555 31038 58607
rect 31090 58555 31107 58607
rect 31021 58543 31107 58555
rect 31021 58491 31038 58543
rect 31090 58491 31107 58543
rect 31021 58479 31107 58491
rect 31021 58427 31038 58479
rect 31090 58427 31107 58479
rect 31021 58415 31107 58427
rect 31021 58363 31038 58415
rect 31090 58363 31107 58415
rect 31021 58351 31107 58363
rect 31021 58299 31038 58351
rect 31090 58299 31107 58351
rect 31021 58287 31107 58299
rect 31021 58235 31038 58287
rect 31090 58235 31107 58287
rect 31021 58223 31107 58235
rect 31021 58171 31038 58223
rect 31090 58171 31107 58223
rect 31021 58166 31107 58171
rect 17420 56738 17506 56743
rect 17420 56686 17437 56738
rect 17489 56686 17506 56738
rect 17420 56674 17506 56686
rect 17420 56622 17437 56674
rect 17489 56622 17506 56674
rect 17420 56610 17506 56622
rect 17420 56558 17437 56610
rect 17489 56558 17506 56610
rect 17420 56546 17506 56558
rect 17420 56494 17437 56546
rect 17489 56494 17506 56546
rect 17420 56482 17506 56494
rect 17420 56430 17437 56482
rect 17489 56430 17506 56482
rect 17420 56418 17506 56430
rect 17420 56366 17437 56418
rect 17489 56366 17506 56418
rect 17420 56354 17506 56366
rect 17420 56302 17437 56354
rect 17489 56302 17506 56354
rect 17420 56290 17506 56302
rect 17420 56238 17437 56290
rect 17489 56238 17506 56290
rect 17420 56226 17506 56238
rect 17420 56174 17437 56226
rect 17489 56174 17506 56226
rect 17420 56169 17506 56174
rect 18508 56738 18594 56743
rect 18508 56686 18525 56738
rect 18577 56686 18594 56738
rect 18508 56674 18594 56686
rect 18508 56622 18525 56674
rect 18577 56622 18594 56674
rect 18508 56610 18594 56622
rect 18508 56558 18525 56610
rect 18577 56558 18594 56610
rect 18508 56546 18594 56558
rect 18508 56494 18525 56546
rect 18577 56494 18594 56546
rect 18508 56482 18594 56494
rect 18508 56430 18525 56482
rect 18577 56430 18594 56482
rect 18508 56418 18594 56430
rect 18508 56366 18525 56418
rect 18577 56366 18594 56418
rect 18508 56354 18594 56366
rect 18508 56302 18525 56354
rect 18577 56302 18594 56354
rect 18508 56290 18594 56302
rect 18508 56238 18525 56290
rect 18577 56238 18594 56290
rect 18508 56226 18594 56238
rect 18508 56174 18525 56226
rect 18577 56174 18594 56226
rect 18508 56169 18594 56174
rect 19596 56738 19682 56743
rect 19596 56686 19613 56738
rect 19665 56686 19682 56738
rect 19596 56674 19682 56686
rect 19596 56622 19613 56674
rect 19665 56622 19682 56674
rect 19596 56610 19682 56622
rect 19596 56558 19613 56610
rect 19665 56558 19682 56610
rect 19596 56546 19682 56558
rect 19596 56494 19613 56546
rect 19665 56494 19682 56546
rect 19596 56482 19682 56494
rect 19596 56430 19613 56482
rect 19665 56430 19682 56482
rect 19596 56418 19682 56430
rect 19596 56366 19613 56418
rect 19665 56366 19682 56418
rect 19596 56354 19682 56366
rect 19596 56302 19613 56354
rect 19665 56302 19682 56354
rect 19596 56290 19682 56302
rect 19596 56238 19613 56290
rect 19665 56238 19682 56290
rect 19596 56226 19682 56238
rect 19596 56174 19613 56226
rect 19665 56174 19682 56226
rect 19596 56169 19682 56174
rect 20684 56738 20770 56743
rect 20684 56686 20701 56738
rect 20753 56686 20770 56738
rect 20684 56674 20770 56686
rect 20684 56622 20701 56674
rect 20753 56622 20770 56674
rect 20684 56610 20770 56622
rect 20684 56558 20701 56610
rect 20753 56558 20770 56610
rect 20684 56546 20770 56558
rect 20684 56494 20701 56546
rect 20753 56494 20770 56546
rect 20684 56482 20770 56494
rect 20684 56430 20701 56482
rect 20753 56430 20770 56482
rect 20684 56418 20770 56430
rect 20684 56366 20701 56418
rect 20753 56366 20770 56418
rect 20684 56354 20770 56366
rect 20684 56302 20701 56354
rect 20753 56302 20770 56354
rect 20684 56290 20770 56302
rect 20684 56238 20701 56290
rect 20753 56238 20770 56290
rect 20684 56226 20770 56238
rect 20684 56174 20701 56226
rect 20753 56174 20770 56226
rect 20684 56169 20770 56174
rect 21772 56738 21858 56743
rect 21772 56686 21789 56738
rect 21841 56686 21858 56738
rect 21772 56674 21858 56686
rect 21772 56622 21789 56674
rect 21841 56622 21858 56674
rect 21772 56610 21858 56622
rect 21772 56558 21789 56610
rect 21841 56558 21858 56610
rect 21772 56546 21858 56558
rect 21772 56494 21789 56546
rect 21841 56494 21858 56546
rect 21772 56482 21858 56494
rect 21772 56430 21789 56482
rect 21841 56430 21858 56482
rect 21772 56418 21858 56430
rect 21772 56366 21789 56418
rect 21841 56366 21858 56418
rect 21772 56354 21858 56366
rect 21772 56302 21789 56354
rect 21841 56302 21858 56354
rect 21772 56290 21858 56302
rect 21772 56238 21789 56290
rect 21841 56238 21858 56290
rect 21772 56226 21858 56238
rect 21772 56174 21789 56226
rect 21841 56174 21858 56226
rect 21772 56169 21858 56174
rect 22860 56738 22946 56743
rect 22860 56686 22877 56738
rect 22929 56686 22946 56738
rect 22860 56674 22946 56686
rect 22860 56622 22877 56674
rect 22929 56622 22946 56674
rect 22860 56610 22946 56622
rect 22860 56558 22877 56610
rect 22929 56558 22946 56610
rect 22860 56546 22946 56558
rect 22860 56494 22877 56546
rect 22929 56494 22946 56546
rect 22860 56482 22946 56494
rect 22860 56430 22877 56482
rect 22929 56430 22946 56482
rect 22860 56418 22946 56430
rect 22860 56366 22877 56418
rect 22929 56366 22946 56418
rect 22860 56354 22946 56366
rect 22860 56302 22877 56354
rect 22929 56302 22946 56354
rect 22860 56290 22946 56302
rect 22860 56238 22877 56290
rect 22929 56238 22946 56290
rect 22860 56226 22946 56238
rect 22860 56174 22877 56226
rect 22929 56174 22946 56226
rect 22860 56169 22946 56174
rect 23948 56738 24034 56743
rect 23948 56686 23965 56738
rect 24017 56686 24034 56738
rect 23948 56674 24034 56686
rect 23948 56622 23965 56674
rect 24017 56622 24034 56674
rect 23948 56610 24034 56622
rect 23948 56558 23965 56610
rect 24017 56558 24034 56610
rect 23948 56546 24034 56558
rect 23948 56494 23965 56546
rect 24017 56494 24034 56546
rect 23948 56482 24034 56494
rect 23948 56430 23965 56482
rect 24017 56430 24034 56482
rect 23948 56418 24034 56430
rect 23948 56366 23965 56418
rect 24017 56366 24034 56418
rect 23948 56354 24034 56366
rect 23948 56302 23965 56354
rect 24017 56302 24034 56354
rect 23948 56290 24034 56302
rect 23948 56238 23965 56290
rect 24017 56238 24034 56290
rect 23948 56226 24034 56238
rect 23948 56174 23965 56226
rect 24017 56174 24034 56226
rect 23948 56169 24034 56174
rect 25036 56738 25122 56743
rect 25036 56686 25053 56738
rect 25105 56686 25122 56738
rect 25036 56674 25122 56686
rect 25036 56622 25053 56674
rect 25105 56622 25122 56674
rect 25036 56610 25122 56622
rect 25036 56558 25053 56610
rect 25105 56558 25122 56610
rect 25036 56546 25122 56558
rect 25036 56494 25053 56546
rect 25105 56494 25122 56546
rect 25036 56482 25122 56494
rect 25036 56430 25053 56482
rect 25105 56430 25122 56482
rect 25036 56418 25122 56430
rect 25036 56366 25053 56418
rect 25105 56366 25122 56418
rect 25036 56354 25122 56366
rect 25036 56302 25053 56354
rect 25105 56302 25122 56354
rect 25036 56290 25122 56302
rect 25036 56238 25053 56290
rect 25105 56238 25122 56290
rect 25036 56226 25122 56238
rect 25036 56174 25053 56226
rect 25105 56174 25122 56226
rect 25036 56169 25122 56174
rect 26124 56738 26210 56743
rect 26124 56686 26141 56738
rect 26193 56686 26210 56738
rect 26124 56674 26210 56686
rect 26124 56622 26141 56674
rect 26193 56622 26210 56674
rect 26124 56610 26210 56622
rect 26124 56558 26141 56610
rect 26193 56558 26210 56610
rect 26124 56546 26210 56558
rect 26124 56494 26141 56546
rect 26193 56494 26210 56546
rect 26124 56482 26210 56494
rect 26124 56430 26141 56482
rect 26193 56430 26210 56482
rect 26124 56418 26210 56430
rect 26124 56366 26141 56418
rect 26193 56366 26210 56418
rect 26124 56354 26210 56366
rect 26124 56302 26141 56354
rect 26193 56302 26210 56354
rect 26124 56290 26210 56302
rect 26124 56238 26141 56290
rect 26193 56238 26210 56290
rect 26124 56226 26210 56238
rect 26124 56174 26141 56226
rect 26193 56174 26210 56226
rect 26124 56169 26210 56174
rect 27212 56738 27298 56743
rect 27212 56686 27229 56738
rect 27281 56686 27298 56738
rect 27212 56674 27298 56686
rect 27212 56622 27229 56674
rect 27281 56622 27298 56674
rect 27212 56610 27298 56622
rect 27212 56558 27229 56610
rect 27281 56558 27298 56610
rect 27212 56546 27298 56558
rect 27212 56494 27229 56546
rect 27281 56494 27298 56546
rect 27212 56482 27298 56494
rect 27212 56430 27229 56482
rect 27281 56430 27298 56482
rect 27212 56418 27298 56430
rect 27212 56366 27229 56418
rect 27281 56366 27298 56418
rect 27212 56354 27298 56366
rect 27212 56302 27229 56354
rect 27281 56302 27298 56354
rect 27212 56290 27298 56302
rect 27212 56238 27229 56290
rect 27281 56238 27298 56290
rect 27212 56226 27298 56238
rect 27212 56174 27229 56226
rect 27281 56174 27298 56226
rect 27212 56169 27298 56174
rect 28300 56738 28386 56743
rect 28300 56686 28317 56738
rect 28369 56686 28386 56738
rect 28300 56674 28386 56686
rect 28300 56622 28317 56674
rect 28369 56622 28386 56674
rect 28300 56610 28386 56622
rect 28300 56558 28317 56610
rect 28369 56558 28386 56610
rect 28300 56546 28386 56558
rect 28300 56494 28317 56546
rect 28369 56494 28386 56546
rect 28300 56482 28386 56494
rect 28300 56430 28317 56482
rect 28369 56430 28386 56482
rect 28300 56418 28386 56430
rect 28300 56366 28317 56418
rect 28369 56366 28386 56418
rect 28300 56354 28386 56366
rect 28300 56302 28317 56354
rect 28369 56302 28386 56354
rect 28300 56290 28386 56302
rect 28300 56238 28317 56290
rect 28369 56238 28386 56290
rect 28300 56226 28386 56238
rect 28300 56174 28317 56226
rect 28369 56174 28386 56226
rect 28300 56169 28386 56174
rect 29388 56738 29474 56743
rect 29388 56686 29405 56738
rect 29457 56686 29474 56738
rect 29388 56674 29474 56686
rect 29388 56622 29405 56674
rect 29457 56622 29474 56674
rect 29388 56610 29474 56622
rect 29388 56558 29405 56610
rect 29457 56558 29474 56610
rect 29388 56546 29474 56558
rect 29388 56494 29405 56546
rect 29457 56494 29474 56546
rect 29388 56482 29474 56494
rect 29388 56430 29405 56482
rect 29457 56430 29474 56482
rect 29388 56418 29474 56430
rect 29388 56366 29405 56418
rect 29457 56366 29474 56418
rect 29388 56354 29474 56366
rect 29388 56302 29405 56354
rect 29457 56302 29474 56354
rect 29388 56290 29474 56302
rect 29388 56238 29405 56290
rect 29457 56238 29474 56290
rect 29388 56226 29474 56238
rect 29388 56174 29405 56226
rect 29457 56174 29474 56226
rect 29388 56169 29474 56174
rect 30476 56738 30562 56743
rect 30476 56686 30493 56738
rect 30545 56686 30562 56738
rect 30476 56674 30562 56686
rect 30476 56622 30493 56674
rect 30545 56622 30562 56674
rect 30476 56610 30562 56622
rect 30476 56558 30493 56610
rect 30545 56558 30562 56610
rect 30476 56546 30562 56558
rect 30476 56494 30493 56546
rect 30545 56494 30562 56546
rect 30476 56482 30562 56494
rect 30476 56430 30493 56482
rect 30545 56430 30562 56482
rect 30476 56418 30562 56430
rect 30476 56366 30493 56418
rect 30545 56366 30562 56418
rect 30476 56354 30562 56366
rect 30476 56302 30493 56354
rect 30545 56302 30562 56354
rect 30476 56290 30562 56302
rect 30476 56238 30493 56290
rect 30545 56238 30562 56290
rect 30476 56226 30562 56238
rect 30476 56174 30493 56226
rect 30545 56174 30562 56226
rect 30476 56169 30562 56174
rect 31564 56738 31650 56743
rect 31564 56686 31581 56738
rect 31633 56686 31650 56738
rect 31564 56674 31650 56686
rect 31564 56622 31581 56674
rect 31633 56622 31650 56674
rect 31564 56610 31650 56622
rect 31564 56558 31581 56610
rect 31633 56558 31650 56610
rect 31564 56546 31650 56558
rect 31564 56494 31581 56546
rect 31633 56494 31650 56546
rect 31564 56482 31650 56494
rect 31564 56430 31581 56482
rect 31633 56430 31650 56482
rect 31564 56418 31650 56430
rect 31564 56366 31581 56418
rect 31633 56366 31650 56418
rect 31564 56354 31650 56366
rect 31564 56302 31581 56354
rect 31633 56302 31650 56354
rect 31564 56290 31650 56302
rect 31564 56238 31581 56290
rect 31633 56238 31650 56290
rect 31564 56226 31650 56238
rect 31564 56174 31581 56226
rect 31633 56174 31650 56226
rect 31564 56169 31650 56174
rect 17965 54735 18051 54740
rect 17965 54683 17982 54735
rect 18034 54683 18051 54735
rect 17965 54671 18051 54683
rect 17965 54619 17982 54671
rect 18034 54619 18051 54671
rect 17965 54607 18051 54619
rect 17965 54555 17982 54607
rect 18034 54555 18051 54607
rect 17965 54543 18051 54555
rect 17965 54491 17982 54543
rect 18034 54491 18051 54543
rect 17965 54479 18051 54491
rect 17965 54427 17982 54479
rect 18034 54427 18051 54479
rect 17965 54415 18051 54427
rect 17965 54363 17982 54415
rect 18034 54363 18051 54415
rect 17965 54351 18051 54363
rect 17965 54299 17982 54351
rect 18034 54299 18051 54351
rect 17965 54287 18051 54299
rect 17965 54235 17982 54287
rect 18034 54235 18051 54287
rect 17965 54223 18051 54235
rect 17965 54171 17982 54223
rect 18034 54171 18051 54223
rect 17965 54166 18051 54171
rect 19053 54735 19139 54740
rect 19053 54683 19070 54735
rect 19122 54683 19139 54735
rect 19053 54671 19139 54683
rect 19053 54619 19070 54671
rect 19122 54619 19139 54671
rect 19053 54607 19139 54619
rect 19053 54555 19070 54607
rect 19122 54555 19139 54607
rect 19053 54543 19139 54555
rect 19053 54491 19070 54543
rect 19122 54491 19139 54543
rect 19053 54479 19139 54491
rect 19053 54427 19070 54479
rect 19122 54427 19139 54479
rect 19053 54415 19139 54427
rect 19053 54363 19070 54415
rect 19122 54363 19139 54415
rect 19053 54351 19139 54363
rect 19053 54299 19070 54351
rect 19122 54299 19139 54351
rect 19053 54287 19139 54299
rect 19053 54235 19070 54287
rect 19122 54235 19139 54287
rect 19053 54223 19139 54235
rect 19053 54171 19070 54223
rect 19122 54171 19139 54223
rect 19053 54166 19139 54171
rect 20141 54735 20227 54740
rect 20141 54683 20158 54735
rect 20210 54683 20227 54735
rect 20141 54671 20227 54683
rect 20141 54619 20158 54671
rect 20210 54619 20227 54671
rect 20141 54607 20227 54619
rect 20141 54555 20158 54607
rect 20210 54555 20227 54607
rect 20141 54543 20227 54555
rect 20141 54491 20158 54543
rect 20210 54491 20227 54543
rect 20141 54479 20227 54491
rect 20141 54427 20158 54479
rect 20210 54427 20227 54479
rect 20141 54415 20227 54427
rect 20141 54363 20158 54415
rect 20210 54363 20227 54415
rect 20141 54351 20227 54363
rect 20141 54299 20158 54351
rect 20210 54299 20227 54351
rect 20141 54287 20227 54299
rect 20141 54235 20158 54287
rect 20210 54235 20227 54287
rect 20141 54223 20227 54235
rect 20141 54171 20158 54223
rect 20210 54171 20227 54223
rect 20141 54166 20227 54171
rect 21229 54735 21315 54740
rect 21229 54683 21246 54735
rect 21298 54683 21315 54735
rect 21229 54671 21315 54683
rect 21229 54619 21246 54671
rect 21298 54619 21315 54671
rect 21229 54607 21315 54619
rect 21229 54555 21246 54607
rect 21298 54555 21315 54607
rect 21229 54543 21315 54555
rect 21229 54491 21246 54543
rect 21298 54491 21315 54543
rect 21229 54479 21315 54491
rect 21229 54427 21246 54479
rect 21298 54427 21315 54479
rect 21229 54415 21315 54427
rect 21229 54363 21246 54415
rect 21298 54363 21315 54415
rect 21229 54351 21315 54363
rect 21229 54299 21246 54351
rect 21298 54299 21315 54351
rect 21229 54287 21315 54299
rect 21229 54235 21246 54287
rect 21298 54235 21315 54287
rect 21229 54223 21315 54235
rect 21229 54171 21246 54223
rect 21298 54171 21315 54223
rect 21229 54166 21315 54171
rect 22317 54735 22403 54740
rect 22317 54683 22334 54735
rect 22386 54683 22403 54735
rect 22317 54671 22403 54683
rect 22317 54619 22334 54671
rect 22386 54619 22403 54671
rect 22317 54607 22403 54619
rect 22317 54555 22334 54607
rect 22386 54555 22403 54607
rect 22317 54543 22403 54555
rect 22317 54491 22334 54543
rect 22386 54491 22403 54543
rect 22317 54479 22403 54491
rect 22317 54427 22334 54479
rect 22386 54427 22403 54479
rect 22317 54415 22403 54427
rect 22317 54363 22334 54415
rect 22386 54363 22403 54415
rect 22317 54351 22403 54363
rect 22317 54299 22334 54351
rect 22386 54299 22403 54351
rect 22317 54287 22403 54299
rect 22317 54235 22334 54287
rect 22386 54235 22403 54287
rect 22317 54223 22403 54235
rect 22317 54171 22334 54223
rect 22386 54171 22403 54223
rect 22317 54166 22403 54171
rect 23405 54735 23491 54740
rect 23405 54683 23422 54735
rect 23474 54683 23491 54735
rect 23405 54671 23491 54683
rect 23405 54619 23422 54671
rect 23474 54619 23491 54671
rect 23405 54607 23491 54619
rect 23405 54555 23422 54607
rect 23474 54555 23491 54607
rect 23405 54543 23491 54555
rect 23405 54491 23422 54543
rect 23474 54491 23491 54543
rect 23405 54479 23491 54491
rect 23405 54427 23422 54479
rect 23474 54427 23491 54479
rect 23405 54415 23491 54427
rect 23405 54363 23422 54415
rect 23474 54363 23491 54415
rect 23405 54351 23491 54363
rect 23405 54299 23422 54351
rect 23474 54299 23491 54351
rect 23405 54287 23491 54299
rect 23405 54235 23422 54287
rect 23474 54235 23491 54287
rect 23405 54223 23491 54235
rect 23405 54171 23422 54223
rect 23474 54171 23491 54223
rect 23405 54166 23491 54171
rect 24493 54735 24579 54740
rect 24493 54683 24510 54735
rect 24562 54683 24579 54735
rect 24493 54671 24579 54683
rect 24493 54619 24510 54671
rect 24562 54619 24579 54671
rect 24493 54607 24579 54619
rect 24493 54555 24510 54607
rect 24562 54555 24579 54607
rect 24493 54543 24579 54555
rect 24493 54491 24510 54543
rect 24562 54491 24579 54543
rect 24493 54479 24579 54491
rect 24493 54427 24510 54479
rect 24562 54427 24579 54479
rect 24493 54415 24579 54427
rect 24493 54363 24510 54415
rect 24562 54363 24579 54415
rect 24493 54351 24579 54363
rect 24493 54299 24510 54351
rect 24562 54299 24579 54351
rect 24493 54287 24579 54299
rect 24493 54235 24510 54287
rect 24562 54235 24579 54287
rect 24493 54223 24579 54235
rect 24493 54171 24510 54223
rect 24562 54171 24579 54223
rect 24493 54166 24579 54171
rect 25581 54735 25667 54740
rect 25581 54683 25598 54735
rect 25650 54683 25667 54735
rect 25581 54671 25667 54683
rect 25581 54619 25598 54671
rect 25650 54619 25667 54671
rect 25581 54607 25667 54619
rect 25581 54555 25598 54607
rect 25650 54555 25667 54607
rect 25581 54543 25667 54555
rect 25581 54491 25598 54543
rect 25650 54491 25667 54543
rect 25581 54479 25667 54491
rect 25581 54427 25598 54479
rect 25650 54427 25667 54479
rect 25581 54415 25667 54427
rect 25581 54363 25598 54415
rect 25650 54363 25667 54415
rect 25581 54351 25667 54363
rect 25581 54299 25598 54351
rect 25650 54299 25667 54351
rect 25581 54287 25667 54299
rect 25581 54235 25598 54287
rect 25650 54235 25667 54287
rect 25581 54223 25667 54235
rect 25581 54171 25598 54223
rect 25650 54171 25667 54223
rect 25581 54166 25667 54171
rect 26669 54735 26755 54740
rect 26669 54683 26686 54735
rect 26738 54683 26755 54735
rect 26669 54671 26755 54683
rect 26669 54619 26686 54671
rect 26738 54619 26755 54671
rect 26669 54607 26755 54619
rect 26669 54555 26686 54607
rect 26738 54555 26755 54607
rect 26669 54543 26755 54555
rect 26669 54491 26686 54543
rect 26738 54491 26755 54543
rect 26669 54479 26755 54491
rect 26669 54427 26686 54479
rect 26738 54427 26755 54479
rect 26669 54415 26755 54427
rect 26669 54363 26686 54415
rect 26738 54363 26755 54415
rect 26669 54351 26755 54363
rect 26669 54299 26686 54351
rect 26738 54299 26755 54351
rect 26669 54287 26755 54299
rect 26669 54235 26686 54287
rect 26738 54235 26755 54287
rect 26669 54223 26755 54235
rect 26669 54171 26686 54223
rect 26738 54171 26755 54223
rect 26669 54166 26755 54171
rect 27757 54735 27843 54740
rect 27757 54683 27774 54735
rect 27826 54683 27843 54735
rect 27757 54671 27843 54683
rect 27757 54619 27774 54671
rect 27826 54619 27843 54671
rect 27757 54607 27843 54619
rect 27757 54555 27774 54607
rect 27826 54555 27843 54607
rect 27757 54543 27843 54555
rect 27757 54491 27774 54543
rect 27826 54491 27843 54543
rect 27757 54479 27843 54491
rect 27757 54427 27774 54479
rect 27826 54427 27843 54479
rect 27757 54415 27843 54427
rect 27757 54363 27774 54415
rect 27826 54363 27843 54415
rect 27757 54351 27843 54363
rect 27757 54299 27774 54351
rect 27826 54299 27843 54351
rect 27757 54287 27843 54299
rect 27757 54235 27774 54287
rect 27826 54235 27843 54287
rect 27757 54223 27843 54235
rect 27757 54171 27774 54223
rect 27826 54171 27843 54223
rect 27757 54166 27843 54171
rect 28845 54735 28931 54740
rect 28845 54683 28862 54735
rect 28914 54683 28931 54735
rect 28845 54671 28931 54683
rect 28845 54619 28862 54671
rect 28914 54619 28931 54671
rect 28845 54607 28931 54619
rect 28845 54555 28862 54607
rect 28914 54555 28931 54607
rect 28845 54543 28931 54555
rect 28845 54491 28862 54543
rect 28914 54491 28931 54543
rect 28845 54479 28931 54491
rect 28845 54427 28862 54479
rect 28914 54427 28931 54479
rect 28845 54415 28931 54427
rect 28845 54363 28862 54415
rect 28914 54363 28931 54415
rect 28845 54351 28931 54363
rect 28845 54299 28862 54351
rect 28914 54299 28931 54351
rect 28845 54287 28931 54299
rect 28845 54235 28862 54287
rect 28914 54235 28931 54287
rect 28845 54223 28931 54235
rect 28845 54171 28862 54223
rect 28914 54171 28931 54223
rect 28845 54166 28931 54171
rect 29933 54735 30019 54740
rect 29933 54683 29950 54735
rect 30002 54683 30019 54735
rect 29933 54671 30019 54683
rect 29933 54619 29950 54671
rect 30002 54619 30019 54671
rect 29933 54607 30019 54619
rect 29933 54555 29950 54607
rect 30002 54555 30019 54607
rect 29933 54543 30019 54555
rect 29933 54491 29950 54543
rect 30002 54491 30019 54543
rect 29933 54479 30019 54491
rect 29933 54427 29950 54479
rect 30002 54427 30019 54479
rect 29933 54415 30019 54427
rect 29933 54363 29950 54415
rect 30002 54363 30019 54415
rect 29933 54351 30019 54363
rect 29933 54299 29950 54351
rect 30002 54299 30019 54351
rect 29933 54287 30019 54299
rect 29933 54235 29950 54287
rect 30002 54235 30019 54287
rect 29933 54223 30019 54235
rect 29933 54171 29950 54223
rect 30002 54171 30019 54223
rect 29933 54166 30019 54171
rect 31021 54735 31107 54740
rect 31021 54683 31038 54735
rect 31090 54683 31107 54735
rect 31021 54671 31107 54683
rect 31021 54619 31038 54671
rect 31090 54619 31107 54671
rect 31021 54607 31107 54619
rect 31021 54555 31038 54607
rect 31090 54555 31107 54607
rect 31021 54543 31107 54555
rect 31021 54491 31038 54543
rect 31090 54491 31107 54543
rect 31021 54479 31107 54491
rect 31021 54427 31038 54479
rect 31090 54427 31107 54479
rect 31021 54415 31107 54427
rect 31021 54363 31038 54415
rect 31090 54363 31107 54415
rect 31021 54351 31107 54363
rect 31021 54299 31038 54351
rect 31090 54299 31107 54351
rect 31021 54287 31107 54299
rect 31021 54235 31038 54287
rect 31090 54235 31107 54287
rect 31021 54223 31107 54235
rect 31021 54171 31038 54223
rect 31090 54171 31107 54223
rect 31021 54166 31107 54171
rect 17420 52738 17506 52743
rect 17420 52686 17437 52738
rect 17489 52686 17506 52738
rect 17420 52674 17506 52686
rect 17420 52622 17437 52674
rect 17489 52622 17506 52674
rect 17420 52610 17506 52622
rect 17420 52558 17437 52610
rect 17489 52558 17506 52610
rect 17420 52546 17506 52558
rect 17420 52494 17437 52546
rect 17489 52494 17506 52546
rect 17420 52482 17506 52494
rect 17420 52430 17437 52482
rect 17489 52430 17506 52482
rect 17420 52418 17506 52430
rect 17420 52366 17437 52418
rect 17489 52366 17506 52418
rect 17420 52354 17506 52366
rect 17420 52302 17437 52354
rect 17489 52302 17506 52354
rect 17420 52290 17506 52302
rect 17420 52238 17437 52290
rect 17489 52238 17506 52290
rect 17420 52226 17506 52238
rect 17420 52174 17437 52226
rect 17489 52174 17506 52226
rect 17420 52169 17506 52174
rect 18508 52738 18594 52743
rect 18508 52686 18525 52738
rect 18577 52686 18594 52738
rect 18508 52674 18594 52686
rect 18508 52622 18525 52674
rect 18577 52622 18594 52674
rect 18508 52610 18594 52622
rect 18508 52558 18525 52610
rect 18577 52558 18594 52610
rect 18508 52546 18594 52558
rect 18508 52494 18525 52546
rect 18577 52494 18594 52546
rect 18508 52482 18594 52494
rect 18508 52430 18525 52482
rect 18577 52430 18594 52482
rect 18508 52418 18594 52430
rect 18508 52366 18525 52418
rect 18577 52366 18594 52418
rect 18508 52354 18594 52366
rect 18508 52302 18525 52354
rect 18577 52302 18594 52354
rect 18508 52290 18594 52302
rect 18508 52238 18525 52290
rect 18577 52238 18594 52290
rect 18508 52226 18594 52238
rect 18508 52174 18525 52226
rect 18577 52174 18594 52226
rect 18508 52169 18594 52174
rect 19596 52738 19682 52743
rect 19596 52686 19613 52738
rect 19665 52686 19682 52738
rect 19596 52674 19682 52686
rect 19596 52622 19613 52674
rect 19665 52622 19682 52674
rect 19596 52610 19682 52622
rect 19596 52558 19613 52610
rect 19665 52558 19682 52610
rect 19596 52546 19682 52558
rect 19596 52494 19613 52546
rect 19665 52494 19682 52546
rect 19596 52482 19682 52494
rect 19596 52430 19613 52482
rect 19665 52430 19682 52482
rect 19596 52418 19682 52430
rect 19596 52366 19613 52418
rect 19665 52366 19682 52418
rect 19596 52354 19682 52366
rect 19596 52302 19613 52354
rect 19665 52302 19682 52354
rect 19596 52290 19682 52302
rect 19596 52238 19613 52290
rect 19665 52238 19682 52290
rect 19596 52226 19682 52238
rect 19596 52174 19613 52226
rect 19665 52174 19682 52226
rect 19596 52169 19682 52174
rect 20684 52738 20770 52743
rect 20684 52686 20701 52738
rect 20753 52686 20770 52738
rect 20684 52674 20770 52686
rect 20684 52622 20701 52674
rect 20753 52622 20770 52674
rect 20684 52610 20770 52622
rect 20684 52558 20701 52610
rect 20753 52558 20770 52610
rect 20684 52546 20770 52558
rect 20684 52494 20701 52546
rect 20753 52494 20770 52546
rect 20684 52482 20770 52494
rect 20684 52430 20701 52482
rect 20753 52430 20770 52482
rect 20684 52418 20770 52430
rect 20684 52366 20701 52418
rect 20753 52366 20770 52418
rect 20684 52354 20770 52366
rect 20684 52302 20701 52354
rect 20753 52302 20770 52354
rect 20684 52290 20770 52302
rect 20684 52238 20701 52290
rect 20753 52238 20770 52290
rect 20684 52226 20770 52238
rect 20684 52174 20701 52226
rect 20753 52174 20770 52226
rect 20684 52169 20770 52174
rect 21772 52738 21858 52743
rect 21772 52686 21789 52738
rect 21841 52686 21858 52738
rect 21772 52674 21858 52686
rect 21772 52622 21789 52674
rect 21841 52622 21858 52674
rect 21772 52610 21858 52622
rect 21772 52558 21789 52610
rect 21841 52558 21858 52610
rect 21772 52546 21858 52558
rect 21772 52494 21789 52546
rect 21841 52494 21858 52546
rect 21772 52482 21858 52494
rect 21772 52430 21789 52482
rect 21841 52430 21858 52482
rect 21772 52418 21858 52430
rect 21772 52366 21789 52418
rect 21841 52366 21858 52418
rect 21772 52354 21858 52366
rect 21772 52302 21789 52354
rect 21841 52302 21858 52354
rect 21772 52290 21858 52302
rect 21772 52238 21789 52290
rect 21841 52238 21858 52290
rect 21772 52226 21858 52238
rect 21772 52174 21789 52226
rect 21841 52174 21858 52226
rect 21772 52169 21858 52174
rect 22860 52738 22946 52743
rect 22860 52686 22877 52738
rect 22929 52686 22946 52738
rect 22860 52674 22946 52686
rect 22860 52622 22877 52674
rect 22929 52622 22946 52674
rect 22860 52610 22946 52622
rect 22860 52558 22877 52610
rect 22929 52558 22946 52610
rect 22860 52546 22946 52558
rect 22860 52494 22877 52546
rect 22929 52494 22946 52546
rect 22860 52482 22946 52494
rect 22860 52430 22877 52482
rect 22929 52430 22946 52482
rect 22860 52418 22946 52430
rect 22860 52366 22877 52418
rect 22929 52366 22946 52418
rect 22860 52354 22946 52366
rect 22860 52302 22877 52354
rect 22929 52302 22946 52354
rect 22860 52290 22946 52302
rect 22860 52238 22877 52290
rect 22929 52238 22946 52290
rect 22860 52226 22946 52238
rect 22860 52174 22877 52226
rect 22929 52174 22946 52226
rect 22860 52169 22946 52174
rect 23948 52738 24034 52743
rect 23948 52686 23965 52738
rect 24017 52686 24034 52738
rect 23948 52674 24034 52686
rect 23948 52622 23965 52674
rect 24017 52622 24034 52674
rect 23948 52610 24034 52622
rect 23948 52558 23965 52610
rect 24017 52558 24034 52610
rect 23948 52546 24034 52558
rect 23948 52494 23965 52546
rect 24017 52494 24034 52546
rect 23948 52482 24034 52494
rect 23948 52430 23965 52482
rect 24017 52430 24034 52482
rect 23948 52418 24034 52430
rect 23948 52366 23965 52418
rect 24017 52366 24034 52418
rect 23948 52354 24034 52366
rect 23948 52302 23965 52354
rect 24017 52302 24034 52354
rect 23948 52290 24034 52302
rect 23948 52238 23965 52290
rect 24017 52238 24034 52290
rect 23948 52226 24034 52238
rect 23948 52174 23965 52226
rect 24017 52174 24034 52226
rect 23948 52169 24034 52174
rect 25036 52738 25122 52743
rect 25036 52686 25053 52738
rect 25105 52686 25122 52738
rect 25036 52674 25122 52686
rect 25036 52622 25053 52674
rect 25105 52622 25122 52674
rect 25036 52610 25122 52622
rect 25036 52558 25053 52610
rect 25105 52558 25122 52610
rect 25036 52546 25122 52558
rect 25036 52494 25053 52546
rect 25105 52494 25122 52546
rect 25036 52482 25122 52494
rect 25036 52430 25053 52482
rect 25105 52430 25122 52482
rect 25036 52418 25122 52430
rect 25036 52366 25053 52418
rect 25105 52366 25122 52418
rect 25036 52354 25122 52366
rect 25036 52302 25053 52354
rect 25105 52302 25122 52354
rect 25036 52290 25122 52302
rect 25036 52238 25053 52290
rect 25105 52238 25122 52290
rect 25036 52226 25122 52238
rect 25036 52174 25053 52226
rect 25105 52174 25122 52226
rect 25036 52169 25122 52174
rect 26124 52738 26210 52743
rect 26124 52686 26141 52738
rect 26193 52686 26210 52738
rect 26124 52674 26210 52686
rect 26124 52622 26141 52674
rect 26193 52622 26210 52674
rect 26124 52610 26210 52622
rect 26124 52558 26141 52610
rect 26193 52558 26210 52610
rect 26124 52546 26210 52558
rect 26124 52494 26141 52546
rect 26193 52494 26210 52546
rect 26124 52482 26210 52494
rect 26124 52430 26141 52482
rect 26193 52430 26210 52482
rect 26124 52418 26210 52430
rect 26124 52366 26141 52418
rect 26193 52366 26210 52418
rect 26124 52354 26210 52366
rect 26124 52302 26141 52354
rect 26193 52302 26210 52354
rect 26124 52290 26210 52302
rect 26124 52238 26141 52290
rect 26193 52238 26210 52290
rect 26124 52226 26210 52238
rect 26124 52174 26141 52226
rect 26193 52174 26210 52226
rect 26124 52169 26210 52174
rect 27212 52738 27298 52743
rect 27212 52686 27229 52738
rect 27281 52686 27298 52738
rect 27212 52674 27298 52686
rect 27212 52622 27229 52674
rect 27281 52622 27298 52674
rect 27212 52610 27298 52622
rect 27212 52558 27229 52610
rect 27281 52558 27298 52610
rect 27212 52546 27298 52558
rect 27212 52494 27229 52546
rect 27281 52494 27298 52546
rect 27212 52482 27298 52494
rect 27212 52430 27229 52482
rect 27281 52430 27298 52482
rect 27212 52418 27298 52430
rect 27212 52366 27229 52418
rect 27281 52366 27298 52418
rect 27212 52354 27298 52366
rect 27212 52302 27229 52354
rect 27281 52302 27298 52354
rect 27212 52290 27298 52302
rect 27212 52238 27229 52290
rect 27281 52238 27298 52290
rect 27212 52226 27298 52238
rect 27212 52174 27229 52226
rect 27281 52174 27298 52226
rect 27212 52169 27298 52174
rect 28300 52738 28386 52743
rect 28300 52686 28317 52738
rect 28369 52686 28386 52738
rect 28300 52674 28386 52686
rect 28300 52622 28317 52674
rect 28369 52622 28386 52674
rect 28300 52610 28386 52622
rect 28300 52558 28317 52610
rect 28369 52558 28386 52610
rect 28300 52546 28386 52558
rect 28300 52494 28317 52546
rect 28369 52494 28386 52546
rect 28300 52482 28386 52494
rect 28300 52430 28317 52482
rect 28369 52430 28386 52482
rect 28300 52418 28386 52430
rect 28300 52366 28317 52418
rect 28369 52366 28386 52418
rect 28300 52354 28386 52366
rect 28300 52302 28317 52354
rect 28369 52302 28386 52354
rect 28300 52290 28386 52302
rect 28300 52238 28317 52290
rect 28369 52238 28386 52290
rect 28300 52226 28386 52238
rect 28300 52174 28317 52226
rect 28369 52174 28386 52226
rect 28300 52169 28386 52174
rect 29388 52738 29474 52743
rect 29388 52686 29405 52738
rect 29457 52686 29474 52738
rect 29388 52674 29474 52686
rect 29388 52622 29405 52674
rect 29457 52622 29474 52674
rect 29388 52610 29474 52622
rect 29388 52558 29405 52610
rect 29457 52558 29474 52610
rect 29388 52546 29474 52558
rect 29388 52494 29405 52546
rect 29457 52494 29474 52546
rect 29388 52482 29474 52494
rect 29388 52430 29405 52482
rect 29457 52430 29474 52482
rect 29388 52418 29474 52430
rect 29388 52366 29405 52418
rect 29457 52366 29474 52418
rect 29388 52354 29474 52366
rect 29388 52302 29405 52354
rect 29457 52302 29474 52354
rect 29388 52290 29474 52302
rect 29388 52238 29405 52290
rect 29457 52238 29474 52290
rect 29388 52226 29474 52238
rect 29388 52174 29405 52226
rect 29457 52174 29474 52226
rect 29388 52169 29474 52174
rect 30476 52738 30562 52743
rect 30476 52686 30493 52738
rect 30545 52686 30562 52738
rect 30476 52674 30562 52686
rect 30476 52622 30493 52674
rect 30545 52622 30562 52674
rect 30476 52610 30562 52622
rect 30476 52558 30493 52610
rect 30545 52558 30562 52610
rect 30476 52546 30562 52558
rect 30476 52494 30493 52546
rect 30545 52494 30562 52546
rect 30476 52482 30562 52494
rect 30476 52430 30493 52482
rect 30545 52430 30562 52482
rect 30476 52418 30562 52430
rect 30476 52366 30493 52418
rect 30545 52366 30562 52418
rect 30476 52354 30562 52366
rect 30476 52302 30493 52354
rect 30545 52302 30562 52354
rect 30476 52290 30562 52302
rect 30476 52238 30493 52290
rect 30545 52238 30562 52290
rect 30476 52226 30562 52238
rect 30476 52174 30493 52226
rect 30545 52174 30562 52226
rect 30476 52169 30562 52174
rect 31564 52738 31650 52743
rect 31564 52686 31581 52738
rect 31633 52686 31650 52738
rect 31564 52674 31650 52686
rect 31564 52622 31581 52674
rect 31633 52622 31650 52674
rect 31564 52610 31650 52622
rect 31564 52558 31581 52610
rect 31633 52558 31650 52610
rect 31564 52546 31650 52558
rect 31564 52494 31581 52546
rect 31633 52494 31650 52546
rect 31564 52482 31650 52494
rect 31564 52430 31581 52482
rect 31633 52430 31650 52482
rect 31564 52418 31650 52430
rect 31564 52366 31581 52418
rect 31633 52366 31650 52418
rect 31564 52354 31650 52366
rect 31564 52302 31581 52354
rect 31633 52302 31650 52354
rect 31564 52290 31650 52302
rect 31564 52238 31581 52290
rect 31633 52238 31650 52290
rect 31564 52226 31650 52238
rect 31564 52174 31581 52226
rect 31633 52174 31650 52226
rect 31564 52169 31650 52174
rect 17965 50735 18051 50740
rect 17965 50683 17982 50735
rect 18034 50683 18051 50735
rect 17965 50671 18051 50683
rect 17965 50619 17982 50671
rect 18034 50619 18051 50671
rect 17965 50607 18051 50619
rect 17965 50555 17982 50607
rect 18034 50555 18051 50607
rect 17965 50543 18051 50555
rect 17965 50491 17982 50543
rect 18034 50491 18051 50543
rect 17965 50479 18051 50491
rect 17965 50427 17982 50479
rect 18034 50427 18051 50479
rect 17965 50415 18051 50427
rect 17965 50363 17982 50415
rect 18034 50363 18051 50415
rect 17965 50351 18051 50363
rect 17965 50299 17982 50351
rect 18034 50299 18051 50351
rect 17965 50287 18051 50299
rect 17965 50235 17982 50287
rect 18034 50235 18051 50287
rect 17965 50223 18051 50235
rect 17965 50171 17982 50223
rect 18034 50171 18051 50223
rect 17965 50166 18051 50171
rect 20141 50735 20227 50740
rect 20141 50683 20158 50735
rect 20210 50683 20227 50735
rect 20141 50671 20227 50683
rect 20141 50619 20158 50671
rect 20210 50619 20227 50671
rect 20141 50607 20227 50619
rect 20141 50555 20158 50607
rect 20210 50555 20227 50607
rect 20141 50543 20227 50555
rect 20141 50491 20158 50543
rect 20210 50491 20227 50543
rect 20141 50479 20227 50491
rect 20141 50427 20158 50479
rect 20210 50427 20227 50479
rect 20141 50415 20227 50427
rect 20141 50363 20158 50415
rect 20210 50363 20227 50415
rect 20141 50351 20227 50363
rect 20141 50299 20158 50351
rect 20210 50299 20227 50351
rect 20141 50287 20227 50299
rect 20141 50235 20158 50287
rect 20210 50235 20227 50287
rect 20141 50223 20227 50235
rect 20141 50171 20158 50223
rect 20210 50171 20227 50223
rect 20141 50166 20227 50171
rect 21229 50735 21315 50740
rect 21229 50683 21246 50735
rect 21298 50683 21315 50735
rect 21229 50671 21315 50683
rect 21229 50619 21246 50671
rect 21298 50619 21315 50671
rect 21229 50607 21315 50619
rect 21229 50555 21246 50607
rect 21298 50555 21315 50607
rect 21229 50543 21315 50555
rect 21229 50491 21246 50543
rect 21298 50491 21315 50543
rect 21229 50479 21315 50491
rect 21229 50427 21246 50479
rect 21298 50427 21315 50479
rect 21229 50415 21315 50427
rect 21229 50363 21246 50415
rect 21298 50363 21315 50415
rect 21229 50351 21315 50363
rect 21229 50299 21246 50351
rect 21298 50299 21315 50351
rect 21229 50287 21315 50299
rect 21229 50235 21246 50287
rect 21298 50235 21315 50287
rect 21229 50223 21315 50235
rect 21229 50171 21246 50223
rect 21298 50171 21315 50223
rect 21229 50166 21315 50171
rect 23405 50735 23491 50740
rect 23405 50683 23422 50735
rect 23474 50683 23491 50735
rect 23405 50671 23491 50683
rect 23405 50619 23422 50671
rect 23474 50619 23491 50671
rect 23405 50607 23491 50619
rect 23405 50555 23422 50607
rect 23474 50555 23491 50607
rect 23405 50543 23491 50555
rect 23405 50491 23422 50543
rect 23474 50491 23491 50543
rect 23405 50479 23491 50491
rect 23405 50427 23422 50479
rect 23474 50427 23491 50479
rect 23405 50415 23491 50427
rect 23405 50363 23422 50415
rect 23474 50363 23491 50415
rect 23405 50351 23491 50363
rect 23405 50299 23422 50351
rect 23474 50299 23491 50351
rect 23405 50287 23491 50299
rect 23405 50235 23422 50287
rect 23474 50235 23491 50287
rect 23405 50223 23491 50235
rect 23405 50171 23422 50223
rect 23474 50171 23491 50223
rect 23405 50166 23491 50171
rect 24493 50735 24579 50740
rect 24493 50683 24510 50735
rect 24562 50683 24579 50735
rect 24493 50671 24579 50683
rect 24493 50619 24510 50671
rect 24562 50619 24579 50671
rect 24493 50607 24579 50619
rect 24493 50555 24510 50607
rect 24562 50555 24579 50607
rect 24493 50543 24579 50555
rect 24493 50491 24510 50543
rect 24562 50491 24579 50543
rect 24493 50479 24579 50491
rect 24493 50427 24510 50479
rect 24562 50427 24579 50479
rect 24493 50415 24579 50427
rect 24493 50363 24510 50415
rect 24562 50363 24579 50415
rect 24493 50351 24579 50363
rect 24493 50299 24510 50351
rect 24562 50299 24579 50351
rect 24493 50287 24579 50299
rect 24493 50235 24510 50287
rect 24562 50235 24579 50287
rect 24493 50223 24579 50235
rect 24493 50171 24510 50223
rect 24562 50171 24579 50223
rect 24493 50166 24579 50171
rect 25581 50735 25667 50740
rect 25581 50683 25598 50735
rect 25650 50683 25667 50735
rect 25581 50671 25667 50683
rect 25581 50619 25598 50671
rect 25650 50619 25667 50671
rect 25581 50607 25667 50619
rect 25581 50555 25598 50607
rect 25650 50555 25667 50607
rect 25581 50543 25667 50555
rect 25581 50491 25598 50543
rect 25650 50491 25667 50543
rect 25581 50479 25667 50491
rect 25581 50427 25598 50479
rect 25650 50427 25667 50479
rect 25581 50415 25667 50427
rect 25581 50363 25598 50415
rect 25650 50363 25667 50415
rect 25581 50351 25667 50363
rect 25581 50299 25598 50351
rect 25650 50299 25667 50351
rect 25581 50287 25667 50299
rect 25581 50235 25598 50287
rect 25650 50235 25667 50287
rect 25581 50223 25667 50235
rect 25581 50171 25598 50223
rect 25650 50171 25667 50223
rect 25581 50166 25667 50171
rect 27757 50735 27843 50740
rect 27757 50683 27774 50735
rect 27826 50683 27843 50735
rect 27757 50671 27843 50683
rect 27757 50619 27774 50671
rect 27826 50619 27843 50671
rect 27757 50607 27843 50619
rect 27757 50555 27774 50607
rect 27826 50555 27843 50607
rect 27757 50543 27843 50555
rect 27757 50491 27774 50543
rect 27826 50491 27843 50543
rect 27757 50479 27843 50491
rect 27757 50427 27774 50479
rect 27826 50427 27843 50479
rect 27757 50415 27843 50427
rect 27757 50363 27774 50415
rect 27826 50363 27843 50415
rect 27757 50351 27843 50363
rect 27757 50299 27774 50351
rect 27826 50299 27843 50351
rect 27757 50287 27843 50299
rect 27757 50235 27774 50287
rect 27826 50235 27843 50287
rect 27757 50223 27843 50235
rect 27757 50171 27774 50223
rect 27826 50171 27843 50223
rect 27757 50166 27843 50171
rect 28845 50735 28931 50740
rect 28845 50683 28862 50735
rect 28914 50683 28931 50735
rect 28845 50671 28931 50683
rect 28845 50619 28862 50671
rect 28914 50619 28931 50671
rect 28845 50607 28931 50619
rect 28845 50555 28862 50607
rect 28914 50555 28931 50607
rect 28845 50543 28931 50555
rect 28845 50491 28862 50543
rect 28914 50491 28931 50543
rect 28845 50479 28931 50491
rect 28845 50427 28862 50479
rect 28914 50427 28931 50479
rect 28845 50415 28931 50427
rect 28845 50363 28862 50415
rect 28914 50363 28931 50415
rect 28845 50351 28931 50363
rect 28845 50299 28862 50351
rect 28914 50299 28931 50351
rect 28845 50287 28931 50299
rect 28845 50235 28862 50287
rect 28914 50235 28931 50287
rect 28845 50223 28931 50235
rect 28845 50171 28862 50223
rect 28914 50171 28931 50223
rect 28845 50166 28931 50171
rect 31021 50735 31107 50740
rect 31021 50683 31038 50735
rect 31090 50683 31107 50735
rect 31021 50671 31107 50683
rect 31021 50619 31038 50671
rect 31090 50619 31107 50671
rect 31021 50607 31107 50619
rect 31021 50555 31038 50607
rect 31090 50555 31107 50607
rect 31021 50543 31107 50555
rect 31021 50491 31038 50543
rect 31090 50491 31107 50543
rect 31021 50479 31107 50491
rect 31021 50427 31038 50479
rect 31090 50427 31107 50479
rect 31021 50415 31107 50427
rect 31021 50363 31038 50415
rect 31090 50363 31107 50415
rect 31021 50351 31107 50363
rect 31021 50299 31038 50351
rect 31090 50299 31107 50351
rect 31021 50287 31107 50299
rect 31021 50235 31038 50287
rect 31090 50235 31107 50287
rect 31021 50223 31107 50235
rect 31021 50171 31038 50223
rect 31090 50171 31107 50223
rect 31021 50166 31107 50171
rect 17420 48738 17506 48743
rect 17420 48686 17437 48738
rect 17489 48686 17506 48738
rect 17420 48674 17506 48686
rect 17420 48622 17437 48674
rect 17489 48622 17506 48674
rect 17420 48610 17506 48622
rect 17420 48558 17437 48610
rect 17489 48558 17506 48610
rect 17420 48546 17506 48558
rect 17420 48494 17437 48546
rect 17489 48494 17506 48546
rect 17420 48482 17506 48494
rect 17420 48430 17437 48482
rect 17489 48430 17506 48482
rect 17420 48418 17506 48430
rect 17420 48366 17437 48418
rect 17489 48366 17506 48418
rect 17420 48354 17506 48366
rect 17420 48302 17437 48354
rect 17489 48302 17506 48354
rect 17420 48290 17506 48302
rect 17420 48238 17437 48290
rect 17489 48238 17506 48290
rect 17420 48226 17506 48238
rect 17420 48174 17437 48226
rect 17489 48174 17506 48226
rect 17420 48169 17506 48174
rect 18508 48738 18594 48743
rect 18508 48686 18525 48738
rect 18577 48686 18594 48738
rect 18508 48674 18594 48686
rect 18508 48622 18525 48674
rect 18577 48622 18594 48674
rect 18508 48610 18594 48622
rect 18508 48558 18525 48610
rect 18577 48558 18594 48610
rect 18508 48546 18594 48558
rect 18508 48494 18525 48546
rect 18577 48494 18594 48546
rect 18508 48482 18594 48494
rect 18508 48430 18525 48482
rect 18577 48430 18594 48482
rect 18508 48418 18594 48430
rect 18508 48366 18525 48418
rect 18577 48366 18594 48418
rect 18508 48354 18594 48366
rect 18508 48302 18525 48354
rect 18577 48302 18594 48354
rect 18508 48290 18594 48302
rect 18508 48238 18525 48290
rect 18577 48238 18594 48290
rect 18508 48226 18594 48238
rect 18508 48174 18525 48226
rect 18577 48174 18594 48226
rect 18508 48169 18594 48174
rect 19596 48738 19682 48743
rect 19596 48686 19613 48738
rect 19665 48686 19682 48738
rect 19596 48674 19682 48686
rect 19596 48622 19613 48674
rect 19665 48622 19682 48674
rect 19596 48610 19682 48622
rect 19596 48558 19613 48610
rect 19665 48558 19682 48610
rect 19596 48546 19682 48558
rect 19596 48494 19613 48546
rect 19665 48494 19682 48546
rect 19596 48482 19682 48494
rect 19596 48430 19613 48482
rect 19665 48430 19682 48482
rect 19596 48418 19682 48430
rect 19596 48366 19613 48418
rect 19665 48366 19682 48418
rect 19596 48354 19682 48366
rect 19596 48302 19613 48354
rect 19665 48302 19682 48354
rect 19596 48290 19682 48302
rect 19596 48238 19613 48290
rect 19665 48238 19682 48290
rect 19596 48226 19682 48238
rect 19596 48174 19613 48226
rect 19665 48174 19682 48226
rect 19596 48169 19682 48174
rect 20684 48738 20770 48743
rect 20684 48686 20701 48738
rect 20753 48686 20770 48738
rect 20684 48674 20770 48686
rect 20684 48622 20701 48674
rect 20753 48622 20770 48674
rect 20684 48610 20770 48622
rect 20684 48558 20701 48610
rect 20753 48558 20770 48610
rect 20684 48546 20770 48558
rect 20684 48494 20701 48546
rect 20753 48494 20770 48546
rect 20684 48482 20770 48494
rect 20684 48430 20701 48482
rect 20753 48430 20770 48482
rect 20684 48418 20770 48430
rect 20684 48366 20701 48418
rect 20753 48366 20770 48418
rect 20684 48354 20770 48366
rect 20684 48302 20701 48354
rect 20753 48302 20770 48354
rect 20684 48290 20770 48302
rect 20684 48238 20701 48290
rect 20753 48238 20770 48290
rect 20684 48226 20770 48238
rect 20684 48174 20701 48226
rect 20753 48174 20770 48226
rect 20684 48169 20770 48174
rect 21772 48738 21858 48743
rect 21772 48686 21789 48738
rect 21841 48686 21858 48738
rect 21772 48674 21858 48686
rect 21772 48622 21789 48674
rect 21841 48622 21858 48674
rect 21772 48610 21858 48622
rect 21772 48558 21789 48610
rect 21841 48558 21858 48610
rect 21772 48546 21858 48558
rect 21772 48494 21789 48546
rect 21841 48494 21858 48546
rect 21772 48482 21858 48494
rect 21772 48430 21789 48482
rect 21841 48430 21858 48482
rect 21772 48418 21858 48430
rect 21772 48366 21789 48418
rect 21841 48366 21858 48418
rect 21772 48354 21858 48366
rect 21772 48302 21789 48354
rect 21841 48302 21858 48354
rect 21772 48290 21858 48302
rect 21772 48238 21789 48290
rect 21841 48238 21858 48290
rect 21772 48226 21858 48238
rect 21772 48174 21789 48226
rect 21841 48174 21858 48226
rect 21772 48169 21858 48174
rect 22860 48738 22946 48743
rect 22860 48686 22877 48738
rect 22929 48686 22946 48738
rect 22860 48674 22946 48686
rect 22860 48622 22877 48674
rect 22929 48622 22946 48674
rect 22860 48610 22946 48622
rect 22860 48558 22877 48610
rect 22929 48558 22946 48610
rect 22860 48546 22946 48558
rect 22860 48494 22877 48546
rect 22929 48494 22946 48546
rect 22860 48482 22946 48494
rect 22860 48430 22877 48482
rect 22929 48430 22946 48482
rect 22860 48418 22946 48430
rect 22860 48366 22877 48418
rect 22929 48366 22946 48418
rect 22860 48354 22946 48366
rect 22860 48302 22877 48354
rect 22929 48302 22946 48354
rect 22860 48290 22946 48302
rect 22860 48238 22877 48290
rect 22929 48238 22946 48290
rect 22860 48226 22946 48238
rect 22860 48174 22877 48226
rect 22929 48174 22946 48226
rect 22860 48169 22946 48174
rect 23948 48738 24034 48743
rect 23948 48686 23965 48738
rect 24017 48686 24034 48738
rect 23948 48674 24034 48686
rect 23948 48622 23965 48674
rect 24017 48622 24034 48674
rect 23948 48610 24034 48622
rect 23948 48558 23965 48610
rect 24017 48558 24034 48610
rect 23948 48546 24034 48558
rect 23948 48494 23965 48546
rect 24017 48494 24034 48546
rect 23948 48482 24034 48494
rect 23948 48430 23965 48482
rect 24017 48430 24034 48482
rect 23948 48418 24034 48430
rect 23948 48366 23965 48418
rect 24017 48366 24034 48418
rect 23948 48354 24034 48366
rect 23948 48302 23965 48354
rect 24017 48302 24034 48354
rect 23948 48290 24034 48302
rect 23948 48238 23965 48290
rect 24017 48238 24034 48290
rect 23948 48226 24034 48238
rect 23948 48174 23965 48226
rect 24017 48174 24034 48226
rect 23948 48169 24034 48174
rect 29388 48738 29474 48743
rect 29388 48686 29405 48738
rect 29457 48686 29474 48738
rect 29388 48674 29474 48686
rect 29388 48622 29405 48674
rect 29457 48622 29474 48674
rect 29388 48610 29474 48622
rect 29388 48558 29405 48610
rect 29457 48558 29474 48610
rect 29388 48546 29474 48558
rect 29388 48494 29405 48546
rect 29457 48494 29474 48546
rect 29388 48482 29474 48494
rect 29388 48430 29405 48482
rect 29457 48430 29474 48482
rect 29388 48418 29474 48430
rect 29388 48366 29405 48418
rect 29457 48366 29474 48418
rect 29388 48354 29474 48366
rect 29388 48302 29405 48354
rect 29457 48302 29474 48354
rect 29388 48290 29474 48302
rect 29388 48238 29405 48290
rect 29457 48238 29474 48290
rect 29388 48226 29474 48238
rect 29388 48174 29405 48226
rect 29457 48174 29474 48226
rect 29388 48169 29474 48174
rect 30476 48738 30562 48743
rect 30476 48686 30493 48738
rect 30545 48686 30562 48738
rect 30476 48674 30562 48686
rect 30476 48622 30493 48674
rect 30545 48622 30562 48674
rect 30476 48610 30562 48622
rect 30476 48558 30493 48610
rect 30545 48558 30562 48610
rect 30476 48546 30562 48558
rect 30476 48494 30493 48546
rect 30545 48494 30562 48546
rect 30476 48482 30562 48494
rect 30476 48430 30493 48482
rect 30545 48430 30562 48482
rect 30476 48418 30562 48430
rect 30476 48366 30493 48418
rect 30545 48366 30562 48418
rect 30476 48354 30562 48366
rect 30476 48302 30493 48354
rect 30545 48302 30562 48354
rect 30476 48290 30562 48302
rect 30476 48238 30493 48290
rect 30545 48238 30562 48290
rect 30476 48226 30562 48238
rect 30476 48174 30493 48226
rect 30545 48174 30562 48226
rect 30476 48169 30562 48174
rect 31564 48738 31650 48743
rect 31564 48686 31581 48738
rect 31633 48686 31650 48738
rect 31564 48674 31650 48686
rect 31564 48622 31581 48674
rect 31633 48622 31650 48674
rect 31564 48610 31650 48622
rect 31564 48558 31581 48610
rect 31633 48558 31650 48610
rect 31564 48546 31650 48558
rect 31564 48494 31581 48546
rect 31633 48494 31650 48546
rect 31564 48482 31650 48494
rect 31564 48430 31581 48482
rect 31633 48430 31650 48482
rect 31564 48418 31650 48430
rect 31564 48366 31581 48418
rect 31633 48366 31650 48418
rect 31564 48354 31650 48366
rect 31564 48302 31581 48354
rect 31633 48302 31650 48354
rect 31564 48290 31650 48302
rect 31564 48238 31581 48290
rect 31633 48238 31650 48290
rect 31564 48226 31650 48238
rect 31564 48174 31581 48226
rect 31633 48174 31650 48226
rect 31564 48169 31650 48174
rect 17965 46735 18051 46740
rect 17965 46683 17982 46735
rect 18034 46683 18051 46735
rect 17965 46671 18051 46683
rect 17965 46619 17982 46671
rect 18034 46619 18051 46671
rect 17965 46607 18051 46619
rect 17965 46555 17982 46607
rect 18034 46555 18051 46607
rect 17965 46543 18051 46555
rect 17965 46491 17982 46543
rect 18034 46491 18051 46543
rect 17965 46479 18051 46491
rect 17965 46427 17982 46479
rect 18034 46427 18051 46479
rect 17965 46415 18051 46427
rect 17965 46363 17982 46415
rect 18034 46363 18051 46415
rect 17965 46351 18051 46363
rect 17965 46299 17982 46351
rect 18034 46299 18051 46351
rect 17965 46287 18051 46299
rect 17965 46235 17982 46287
rect 18034 46235 18051 46287
rect 17965 46223 18051 46235
rect 17965 46171 17982 46223
rect 18034 46171 18051 46223
rect 17965 46166 18051 46171
rect 19053 46735 19139 46740
rect 19053 46683 19070 46735
rect 19122 46683 19139 46735
rect 19053 46671 19139 46683
rect 19053 46619 19070 46671
rect 19122 46619 19139 46671
rect 19053 46607 19139 46619
rect 19053 46555 19070 46607
rect 19122 46555 19139 46607
rect 19053 46543 19139 46555
rect 19053 46491 19070 46543
rect 19122 46491 19139 46543
rect 19053 46479 19139 46491
rect 19053 46427 19070 46479
rect 19122 46427 19139 46479
rect 19053 46415 19139 46427
rect 19053 46363 19070 46415
rect 19122 46363 19139 46415
rect 19053 46351 19139 46363
rect 19053 46299 19070 46351
rect 19122 46299 19139 46351
rect 19053 46287 19139 46299
rect 19053 46235 19070 46287
rect 19122 46235 19139 46287
rect 19053 46223 19139 46235
rect 19053 46171 19070 46223
rect 19122 46171 19139 46223
rect 19053 46166 19139 46171
rect 20141 46735 20227 46740
rect 20141 46683 20158 46735
rect 20210 46683 20227 46735
rect 20141 46671 20227 46683
rect 20141 46619 20158 46671
rect 20210 46619 20227 46671
rect 20141 46607 20227 46619
rect 20141 46555 20158 46607
rect 20210 46555 20227 46607
rect 20141 46543 20227 46555
rect 20141 46491 20158 46543
rect 20210 46491 20227 46543
rect 20141 46479 20227 46491
rect 20141 46427 20158 46479
rect 20210 46427 20227 46479
rect 20141 46415 20227 46427
rect 20141 46363 20158 46415
rect 20210 46363 20227 46415
rect 20141 46351 20227 46363
rect 20141 46299 20158 46351
rect 20210 46299 20227 46351
rect 20141 46287 20227 46299
rect 20141 46235 20158 46287
rect 20210 46235 20227 46287
rect 20141 46223 20227 46235
rect 20141 46171 20158 46223
rect 20210 46171 20227 46223
rect 20141 46166 20227 46171
rect 21229 46735 21315 46740
rect 21229 46683 21246 46735
rect 21298 46683 21315 46735
rect 21229 46671 21315 46683
rect 21229 46619 21246 46671
rect 21298 46619 21315 46671
rect 21229 46607 21315 46619
rect 21229 46555 21246 46607
rect 21298 46555 21315 46607
rect 21229 46543 21315 46555
rect 21229 46491 21246 46543
rect 21298 46491 21315 46543
rect 21229 46479 21315 46491
rect 21229 46427 21246 46479
rect 21298 46427 21315 46479
rect 21229 46415 21315 46427
rect 21229 46363 21246 46415
rect 21298 46363 21315 46415
rect 21229 46351 21315 46363
rect 21229 46299 21246 46351
rect 21298 46299 21315 46351
rect 21229 46287 21315 46299
rect 21229 46235 21246 46287
rect 21298 46235 21315 46287
rect 21229 46223 21315 46235
rect 21229 46171 21246 46223
rect 21298 46171 21315 46223
rect 21229 46166 21315 46171
rect 22317 46735 22403 46740
rect 22317 46683 22334 46735
rect 22386 46683 22403 46735
rect 22317 46671 22403 46683
rect 22317 46619 22334 46671
rect 22386 46619 22403 46671
rect 22317 46607 22403 46619
rect 22317 46555 22334 46607
rect 22386 46555 22403 46607
rect 22317 46543 22403 46555
rect 22317 46491 22334 46543
rect 22386 46491 22403 46543
rect 22317 46479 22403 46491
rect 22317 46427 22334 46479
rect 22386 46427 22403 46479
rect 22317 46415 22403 46427
rect 22317 46363 22334 46415
rect 22386 46363 22403 46415
rect 22317 46351 22403 46363
rect 22317 46299 22334 46351
rect 22386 46299 22403 46351
rect 22317 46287 22403 46299
rect 22317 46235 22334 46287
rect 22386 46235 22403 46287
rect 22317 46223 22403 46235
rect 22317 46171 22334 46223
rect 22386 46171 22403 46223
rect 22317 46166 22403 46171
rect 24493 46735 24579 46740
rect 24493 46683 24510 46735
rect 24562 46683 24579 46735
rect 24493 46671 24579 46683
rect 24493 46619 24510 46671
rect 24562 46619 24579 46671
rect 24493 46607 24579 46619
rect 24493 46555 24510 46607
rect 24562 46555 24579 46607
rect 24493 46543 24579 46555
rect 24493 46491 24510 46543
rect 24562 46491 24579 46543
rect 24493 46479 24579 46491
rect 24493 46427 24510 46479
rect 24562 46427 24579 46479
rect 24493 46415 24579 46427
rect 24493 46363 24510 46415
rect 24562 46363 24579 46415
rect 24493 46351 24579 46363
rect 24493 46299 24510 46351
rect 24562 46299 24579 46351
rect 24493 46287 24579 46299
rect 24493 46235 24510 46287
rect 24562 46235 24579 46287
rect 24493 46223 24579 46235
rect 24493 46171 24510 46223
rect 24562 46171 24579 46223
rect 24493 46166 24579 46171
rect 25581 46735 25667 46740
rect 25581 46683 25598 46735
rect 25650 46683 25667 46735
rect 25581 46671 25667 46683
rect 25581 46619 25598 46671
rect 25650 46619 25667 46671
rect 25581 46607 25667 46619
rect 25581 46555 25598 46607
rect 25650 46555 25667 46607
rect 25581 46543 25667 46555
rect 25581 46491 25598 46543
rect 25650 46491 25667 46543
rect 25581 46479 25667 46491
rect 25581 46427 25598 46479
rect 25650 46427 25667 46479
rect 25581 46415 25667 46427
rect 25581 46363 25598 46415
rect 25650 46363 25667 46415
rect 25581 46351 25667 46363
rect 25581 46299 25598 46351
rect 25650 46299 25667 46351
rect 25581 46287 25667 46299
rect 25581 46235 25598 46287
rect 25650 46235 25667 46287
rect 25581 46223 25667 46235
rect 25581 46171 25598 46223
rect 25650 46171 25667 46223
rect 25581 46166 25667 46171
rect 26669 46735 26755 46740
rect 26669 46683 26686 46735
rect 26738 46683 26755 46735
rect 26669 46671 26755 46683
rect 26669 46619 26686 46671
rect 26738 46619 26755 46671
rect 26669 46607 26755 46619
rect 26669 46555 26686 46607
rect 26738 46555 26755 46607
rect 26669 46543 26755 46555
rect 26669 46491 26686 46543
rect 26738 46491 26755 46543
rect 26669 46479 26755 46491
rect 26669 46427 26686 46479
rect 26738 46427 26755 46479
rect 26669 46415 26755 46427
rect 26669 46363 26686 46415
rect 26738 46363 26755 46415
rect 26669 46351 26755 46363
rect 26669 46299 26686 46351
rect 26738 46299 26755 46351
rect 26669 46287 26755 46299
rect 26669 46235 26686 46287
rect 26738 46235 26755 46287
rect 26669 46223 26755 46235
rect 26669 46171 26686 46223
rect 26738 46171 26755 46223
rect 26669 46166 26755 46171
rect 27757 46735 27843 46740
rect 27757 46683 27774 46735
rect 27826 46683 27843 46735
rect 27757 46671 27843 46683
rect 27757 46619 27774 46671
rect 27826 46619 27843 46671
rect 27757 46607 27843 46619
rect 27757 46555 27774 46607
rect 27826 46555 27843 46607
rect 27757 46543 27843 46555
rect 27757 46491 27774 46543
rect 27826 46491 27843 46543
rect 27757 46479 27843 46491
rect 27757 46427 27774 46479
rect 27826 46427 27843 46479
rect 27757 46415 27843 46427
rect 27757 46363 27774 46415
rect 27826 46363 27843 46415
rect 27757 46351 27843 46363
rect 27757 46299 27774 46351
rect 27826 46299 27843 46351
rect 27757 46287 27843 46299
rect 27757 46235 27774 46287
rect 27826 46235 27843 46287
rect 27757 46223 27843 46235
rect 27757 46171 27774 46223
rect 27826 46171 27843 46223
rect 27757 46166 27843 46171
rect 28845 46735 28931 46740
rect 28845 46683 28862 46735
rect 28914 46683 28931 46735
rect 28845 46671 28931 46683
rect 28845 46619 28862 46671
rect 28914 46619 28931 46671
rect 28845 46607 28931 46619
rect 28845 46555 28862 46607
rect 28914 46555 28931 46607
rect 28845 46543 28931 46555
rect 28845 46491 28862 46543
rect 28914 46491 28931 46543
rect 28845 46479 28931 46491
rect 28845 46427 28862 46479
rect 28914 46427 28931 46479
rect 28845 46415 28931 46427
rect 28845 46363 28862 46415
rect 28914 46363 28931 46415
rect 28845 46351 28931 46363
rect 28845 46299 28862 46351
rect 28914 46299 28931 46351
rect 28845 46287 28931 46299
rect 28845 46235 28862 46287
rect 28914 46235 28931 46287
rect 28845 46223 28931 46235
rect 28845 46171 28862 46223
rect 28914 46171 28931 46223
rect 28845 46166 28931 46171
rect 29933 46735 30019 46740
rect 29933 46683 29950 46735
rect 30002 46683 30019 46735
rect 29933 46671 30019 46683
rect 29933 46619 29950 46671
rect 30002 46619 30019 46671
rect 29933 46607 30019 46619
rect 29933 46555 29950 46607
rect 30002 46555 30019 46607
rect 29933 46543 30019 46555
rect 29933 46491 29950 46543
rect 30002 46491 30019 46543
rect 29933 46479 30019 46491
rect 29933 46427 29950 46479
rect 30002 46427 30019 46479
rect 29933 46415 30019 46427
rect 29933 46363 29950 46415
rect 30002 46363 30019 46415
rect 29933 46351 30019 46363
rect 29933 46299 29950 46351
rect 30002 46299 30019 46351
rect 29933 46287 30019 46299
rect 29933 46235 29950 46287
rect 30002 46235 30019 46287
rect 29933 46223 30019 46235
rect 29933 46171 29950 46223
rect 30002 46171 30019 46223
rect 29933 46166 30019 46171
rect 31021 46735 31107 46740
rect 31021 46683 31038 46735
rect 31090 46683 31107 46735
rect 31021 46671 31107 46683
rect 31021 46619 31038 46671
rect 31090 46619 31107 46671
rect 31021 46607 31107 46619
rect 31021 46555 31038 46607
rect 31090 46555 31107 46607
rect 31021 46543 31107 46555
rect 31021 46491 31038 46543
rect 31090 46491 31107 46543
rect 31021 46479 31107 46491
rect 31021 46427 31038 46479
rect 31090 46427 31107 46479
rect 31021 46415 31107 46427
rect 31021 46363 31038 46415
rect 31090 46363 31107 46415
rect 31021 46351 31107 46363
rect 31021 46299 31038 46351
rect 31090 46299 31107 46351
rect 31021 46287 31107 46299
rect 31021 46235 31038 46287
rect 31090 46235 31107 46287
rect 31021 46223 31107 46235
rect 31021 46171 31038 46223
rect 31090 46171 31107 46223
rect 31021 46166 31107 46171
rect 18235 45742 18319 45748
rect 18235 45690 18251 45742
rect 18303 45690 18319 45742
rect 18235 45684 18319 45690
rect 18781 45742 18865 45748
rect 18781 45690 18797 45742
rect 18849 45690 18865 45742
rect 18781 45684 18865 45690
rect 19327 45733 19411 45739
rect 19327 45681 19343 45733
rect 19395 45681 19411 45733
rect 19327 45675 19411 45681
rect 19872 45732 19956 45738
rect 19872 45680 19888 45732
rect 19940 45680 19956 45732
rect 25853 45732 25937 45738
rect 19872 45674 19956 45680
rect 21503 45720 21587 45726
rect 21503 45668 21519 45720
rect 21571 45668 21587 45720
rect 21503 45662 21587 45668
rect 22046 45717 22130 45723
rect 22046 45665 22062 45717
rect 22114 45665 22130 45717
rect 22046 45659 22130 45665
rect 22588 45716 22672 45722
rect 22588 45664 22604 45716
rect 22656 45664 22672 45716
rect 22588 45658 22672 45664
rect 23135 45721 23219 45727
rect 23135 45669 23151 45721
rect 23203 45669 23219 45721
rect 25853 45680 25869 45732
rect 25921 45680 25937 45732
rect 25853 45674 25937 45680
rect 26396 45736 26480 45742
rect 26396 45684 26412 45736
rect 26464 45684 26480 45736
rect 26396 45678 26480 45684
rect 26938 45730 27022 45736
rect 26938 45678 26954 45730
rect 27006 45678 27022 45730
rect 29119 45732 29203 45738
rect 26938 45672 27022 45678
rect 27495 45721 27579 45727
rect 23135 45663 23219 45669
rect 27495 45669 27511 45721
rect 27563 45669 27579 45721
rect 29119 45680 29135 45732
rect 29187 45680 29203 45732
rect 29119 45674 29203 45680
rect 29663 45725 29747 45731
rect 27495 45663 27579 45669
rect 29663 45673 29679 45725
rect 29731 45673 29747 45725
rect 29663 45667 29747 45673
rect 30213 45729 30297 45735
rect 30213 45677 30229 45729
rect 30281 45677 30297 45729
rect 30213 45671 30297 45677
rect 30746 45729 30830 45735
rect 30746 45677 30762 45729
rect 30814 45677 30830 45729
rect 30746 45671 30830 45677
rect 44744 45066 45316 45074
rect 44744 45014 44780 45066
rect 44832 45014 44844 45066
rect 44896 45014 44908 45066
rect 44960 45014 44972 45066
rect 45024 45014 45036 45066
rect 45088 45014 45100 45066
rect 45152 45014 45164 45066
rect 45216 45014 45228 45066
rect 45280 45014 45316 45066
rect 44744 45007 45316 45014
rect 41802 44927 41848 44948
rect 41802 44893 41808 44927
rect 41842 44893 41848 44927
rect 39547 44885 39631 44891
rect 39547 44833 39563 44885
rect 39615 44861 39631 44885
rect 39615 44833 40018 44861
rect 39547 44827 40018 44833
rect 41802 44855 41848 44893
rect 39972 44823 40018 44827
rect 39972 44817 40030 44823
rect 39972 44783 39984 44817
rect 40018 44783 40030 44817
rect 39972 44777 40030 44783
rect 40585 44778 40595 44830
rect 40647 44778 40657 44830
rect 40591 44776 40649 44778
rect 40985 44767 40995 44819
rect 41047 44767 41057 44819
rect 41142 44771 41152 44823
rect 41204 44771 41214 44823
rect 41802 44821 41808 44855
rect 41842 44821 41848 44855
rect 46284 44911 46540 44939
rect 46284 44853 46322 44911
rect 43269 44836 43327 44842
rect 43441 44836 43499 44842
rect 43613 44836 43671 44842
rect 43785 44836 43843 44842
rect 43957 44836 44015 44842
rect 44162 44836 44220 44842
rect 44339 44836 44397 44842
rect 44511 44836 44569 44842
rect 44683 44836 44741 44842
rect 44855 44836 44913 44842
rect 45027 44836 45085 44842
rect 45199 44836 45257 44842
rect 45864 44836 46322 44853
rect 41802 44783 41848 44821
rect 40116 44736 40174 44742
rect 40116 44702 40128 44736
rect 40162 44702 40174 44736
rect 40884 44710 40894 44762
rect 40946 44710 40956 44762
rect 41802 44749 41808 44783
rect 41842 44753 41848 44783
rect 42997 44786 43044 44830
rect 43269 44802 43281 44836
rect 43315 44802 43453 44836
rect 43487 44802 43625 44836
rect 43659 44802 43797 44836
rect 43831 44802 43969 44836
rect 44003 44802 44174 44836
rect 44208 44802 44351 44836
rect 44385 44802 44523 44836
rect 44557 44802 44695 44836
rect 44729 44802 44867 44836
rect 44901 44802 45039 44836
rect 45073 44802 45211 44836
rect 45245 44802 46322 44836
rect 43269 44796 43327 44802
rect 43441 44796 43499 44802
rect 43613 44796 43671 44802
rect 43785 44796 43843 44802
rect 43957 44796 44015 44802
rect 44162 44796 44220 44802
rect 44339 44796 44397 44802
rect 44511 44796 44569 44802
rect 44683 44796 44741 44802
rect 44855 44796 44913 44802
rect 45027 44796 45085 44802
rect 45199 44796 45257 44802
rect 45864 44789 46322 44802
rect 41842 44749 42948 44753
rect 41802 44747 42948 44749
rect 41802 44713 42539 44747
rect 42573 44713 42611 44747
rect 42645 44713 42683 44747
rect 42717 44713 42755 44747
rect 42789 44713 42827 44747
rect 42861 44713 42899 44747
rect 42933 44713 42948 44747
rect 41802 44711 42948 44713
rect 40116 44701 40174 44702
rect 39547 44696 40174 44701
rect 39547 44695 40162 44696
rect 39547 44643 39563 44695
rect 39615 44667 40162 44695
rect 41802 44677 41808 44711
rect 41842 44708 42948 44711
rect 41842 44677 41848 44708
rect 42525 44707 42948 44708
rect 42997 44752 43003 44786
rect 43037 44756 43044 44786
rect 43037 44752 43507 44756
rect 42997 44750 43507 44752
rect 42997 44716 43277 44750
rect 43311 44716 43349 44750
rect 43383 44716 43507 44750
rect 42997 44714 43507 44716
rect 39615 44643 39631 44667
rect 39547 44637 39631 44643
rect 41802 44639 41848 44677
rect 41802 44605 41808 44639
rect 41842 44605 41848 44639
rect 42997 44680 43003 44714
rect 43037 44710 43507 44714
rect 46284 44731 46322 44789
rect 46502 44731 46540 44911
rect 43037 44680 43044 44710
rect 46284 44703 46540 44731
rect 42997 44636 43044 44680
rect 41802 44584 41848 44605
rect 41506 44520 41884 44527
rect 41506 44468 41541 44520
rect 41593 44468 41605 44520
rect 41657 44468 41669 44520
rect 41721 44468 41733 44520
rect 41785 44468 41797 44520
rect 41849 44468 41884 44520
rect 41506 44462 41884 44468
rect 44756 43915 45303 43925
rect 44756 43863 44779 43915
rect 44831 43863 44843 43915
rect 44895 43863 44907 43915
rect 44959 43863 44971 43915
rect 45023 43863 45035 43915
rect 45087 43863 45099 43915
rect 45151 43863 45163 43915
rect 45215 43863 45227 43915
rect 45279 43863 45303 43915
rect 44756 43854 45303 43863
rect 41802 43777 41848 43798
rect 41802 43743 41808 43777
rect 41842 43743 41848 43777
rect 39547 43735 39631 43741
rect 39547 43683 39563 43735
rect 39615 43711 39631 43735
rect 39615 43683 40018 43711
rect 39547 43677 40018 43683
rect 41802 43705 41848 43743
rect 39972 43673 40018 43677
rect 39972 43667 40030 43673
rect 39972 43633 39984 43667
rect 40018 43633 40030 43667
rect 39972 43627 40030 43633
rect 40585 43628 40595 43680
rect 40647 43628 40657 43680
rect 40591 43626 40649 43628
rect 40985 43617 40995 43669
rect 41047 43617 41057 43669
rect 41142 43621 41152 43673
rect 41204 43621 41214 43673
rect 41802 43671 41808 43705
rect 41842 43671 41848 43705
rect 46272 43760 46528 43788
rect 46272 43703 46310 43760
rect 43269 43686 43327 43692
rect 43441 43686 43499 43692
rect 43613 43686 43671 43692
rect 43785 43686 43843 43692
rect 43957 43686 44015 43692
rect 44162 43686 44220 43692
rect 44339 43686 44397 43692
rect 44511 43686 44569 43692
rect 44683 43686 44741 43692
rect 44855 43686 44913 43692
rect 45027 43686 45085 43692
rect 45199 43686 45257 43692
rect 45864 43686 46310 43703
rect 41802 43633 41848 43671
rect 40116 43586 40174 43592
rect 40116 43552 40128 43586
rect 40162 43552 40174 43586
rect 40884 43560 40894 43612
rect 40946 43560 40956 43612
rect 41802 43599 41808 43633
rect 41842 43603 41848 43633
rect 42997 43636 43044 43680
rect 43269 43652 43281 43686
rect 43315 43652 43453 43686
rect 43487 43652 43625 43686
rect 43659 43652 43797 43686
rect 43831 43652 43969 43686
rect 44003 43652 44174 43686
rect 44208 43652 44351 43686
rect 44385 43652 44523 43686
rect 44557 43652 44695 43686
rect 44729 43652 44867 43686
rect 44901 43652 45039 43686
rect 45073 43652 45211 43686
rect 45245 43652 46310 43686
rect 43269 43646 43327 43652
rect 43441 43646 43499 43652
rect 43613 43646 43671 43652
rect 43785 43646 43843 43652
rect 43957 43646 44015 43652
rect 44162 43646 44220 43652
rect 44339 43646 44397 43652
rect 44511 43646 44569 43652
rect 44683 43646 44741 43652
rect 44855 43646 44913 43652
rect 45027 43646 45085 43652
rect 45199 43646 45257 43652
rect 45864 43639 46310 43652
rect 41842 43599 42948 43603
rect 41802 43597 42948 43599
rect 41802 43563 42539 43597
rect 42573 43563 42611 43597
rect 42645 43563 42683 43597
rect 42717 43563 42755 43597
rect 42789 43563 42827 43597
rect 42861 43563 42899 43597
rect 42933 43563 42948 43597
rect 41802 43561 42948 43563
rect 40116 43551 40174 43552
rect 39547 43546 40174 43551
rect 39547 43545 40162 43546
rect 39547 43493 39563 43545
rect 39615 43517 40162 43545
rect 41802 43527 41808 43561
rect 41842 43558 42948 43561
rect 41842 43527 41848 43558
rect 42525 43557 42948 43558
rect 42997 43602 43003 43636
rect 43037 43606 43044 43636
rect 43037 43602 43507 43606
rect 42997 43600 43507 43602
rect 42997 43566 43277 43600
rect 43311 43566 43349 43600
rect 43383 43566 43507 43600
rect 42997 43564 43507 43566
rect 39615 43493 39631 43517
rect 39547 43487 39631 43493
rect 41802 43489 41848 43527
rect 41802 43455 41808 43489
rect 41842 43455 41848 43489
rect 42997 43530 43003 43564
rect 43037 43560 43507 43564
rect 46272 43580 46310 43639
rect 46490 43580 46528 43760
rect 43037 43530 43044 43560
rect 46272 43552 46528 43580
rect 42997 43486 43044 43530
rect 41802 43434 41848 43455
rect 41504 43370 41882 43377
rect 41504 43318 41539 43370
rect 41591 43318 41603 43370
rect 41655 43318 41667 43370
rect 41719 43318 41731 43370
rect 41783 43318 41795 43370
rect 41847 43318 41882 43370
rect 41504 43312 41882 43318
rect 44746 41373 45293 41383
rect 44746 41321 44769 41373
rect 44821 41321 44833 41373
rect 44885 41321 44897 41373
rect 44949 41321 44961 41373
rect 45013 41321 45025 41373
rect 45077 41321 45089 41373
rect 45141 41321 45153 41373
rect 45205 41321 45217 41373
rect 45269 41321 45293 41373
rect 44746 41312 45293 41321
rect 41802 41237 41848 41258
rect 41802 41203 41808 41237
rect 41842 41203 41848 41237
rect 39547 41195 39631 41201
rect 39547 41143 39563 41195
rect 39615 41171 39631 41195
rect 39615 41143 40018 41171
rect 39547 41137 40018 41143
rect 41802 41165 41848 41203
rect 39972 41133 40018 41137
rect 39972 41127 40030 41133
rect 39972 41093 39984 41127
rect 40018 41093 40030 41127
rect 39972 41087 40030 41093
rect 40585 41088 40595 41140
rect 40647 41088 40657 41140
rect 40591 41086 40649 41088
rect 40985 41077 40995 41129
rect 41047 41077 41057 41129
rect 41142 41081 41152 41133
rect 41204 41081 41214 41133
rect 41802 41131 41808 41165
rect 41842 41131 41848 41165
rect 46130 41228 46386 41256
rect 46130 41162 46168 41228
rect 43269 41146 43327 41152
rect 43441 41146 43499 41152
rect 43613 41146 43671 41152
rect 43785 41146 43843 41152
rect 43957 41146 44015 41152
rect 44162 41146 44220 41152
rect 44339 41146 44397 41152
rect 44511 41146 44569 41152
rect 44683 41146 44741 41152
rect 44855 41146 44913 41152
rect 45027 41146 45085 41152
rect 45199 41146 45257 41152
rect 45864 41146 46168 41162
rect 41802 41093 41848 41131
rect 40116 41046 40174 41052
rect 40116 41012 40128 41046
rect 40162 41012 40174 41046
rect 40884 41020 40894 41072
rect 40946 41020 40956 41072
rect 41802 41059 41808 41093
rect 41842 41063 41848 41093
rect 42997 41096 43044 41140
rect 43269 41112 43281 41146
rect 43315 41112 43453 41146
rect 43487 41112 43625 41146
rect 43659 41112 43797 41146
rect 43831 41112 43969 41146
rect 44003 41112 44174 41146
rect 44208 41112 44351 41146
rect 44385 41112 44523 41146
rect 44557 41112 44695 41146
rect 44729 41112 44867 41146
rect 44901 41112 45039 41146
rect 45073 41112 45211 41146
rect 45245 41112 46168 41146
rect 43269 41106 43327 41112
rect 43441 41106 43499 41112
rect 43613 41106 43671 41112
rect 43785 41106 43843 41112
rect 43957 41106 44015 41112
rect 44162 41106 44220 41112
rect 44339 41106 44397 41112
rect 44511 41106 44569 41112
rect 44683 41106 44741 41112
rect 44855 41106 44913 41112
rect 45027 41106 45085 41112
rect 45199 41106 45257 41112
rect 45864 41098 46168 41112
rect 41842 41059 42948 41063
rect 41802 41057 42948 41059
rect 41802 41023 42539 41057
rect 42573 41023 42611 41057
rect 42645 41023 42683 41057
rect 42717 41023 42755 41057
rect 42789 41023 42827 41057
rect 42861 41023 42899 41057
rect 42933 41023 42948 41057
rect 41802 41021 42948 41023
rect 40116 41011 40174 41012
rect 39547 41006 40174 41011
rect 39547 41005 40162 41006
rect 39547 40953 39563 41005
rect 39615 40977 40162 41005
rect 41802 40987 41808 41021
rect 41842 41018 42948 41021
rect 41842 40987 41848 41018
rect 42525 41017 42948 41018
rect 42997 41062 43003 41096
rect 43037 41066 43044 41096
rect 43037 41062 43507 41066
rect 42997 41060 43507 41062
rect 42997 41026 43277 41060
rect 43311 41026 43349 41060
rect 43383 41026 43507 41060
rect 42997 41024 43507 41026
rect 39615 40953 39631 40977
rect 39547 40947 39631 40953
rect 41802 40949 41848 40987
rect 41802 40915 41808 40949
rect 41842 40915 41848 40949
rect 42997 40990 43003 41024
rect 43037 41020 43507 41024
rect 46130 41048 46168 41098
rect 46348 41048 46386 41228
rect 46130 41020 46386 41048
rect 43037 40990 43044 41020
rect 42997 40946 43044 40990
rect 41802 40894 41848 40915
rect 41422 40829 41800 40836
rect 41422 40777 41457 40829
rect 41509 40777 41521 40829
rect 41573 40777 41585 40829
rect 41637 40777 41649 40829
rect 41701 40777 41713 40829
rect 41765 40777 41800 40829
rect 41422 40771 41800 40777
rect 44746 40103 45293 40113
rect 44746 40051 44769 40103
rect 44821 40051 44833 40103
rect 44885 40051 44897 40103
rect 44949 40051 44961 40103
rect 45013 40051 45025 40103
rect 45077 40051 45089 40103
rect 45141 40051 45153 40103
rect 45205 40051 45217 40103
rect 45269 40051 45293 40103
rect 44746 40042 45293 40051
rect 41802 39967 41848 39988
rect 41802 39933 41808 39967
rect 41842 39933 41848 39967
rect 39547 39925 39631 39931
rect 39547 39873 39563 39925
rect 39615 39901 39631 39925
rect 39615 39873 40018 39901
rect 39547 39867 40018 39873
rect 41802 39895 41848 39933
rect 39972 39863 40018 39867
rect 39972 39857 40030 39863
rect 39972 39823 39984 39857
rect 40018 39823 40030 39857
rect 39972 39817 40030 39823
rect 40585 39818 40595 39870
rect 40647 39818 40657 39870
rect 40591 39816 40649 39818
rect 40985 39807 40995 39859
rect 41047 39807 41057 39859
rect 41142 39811 41152 39863
rect 41204 39811 41214 39863
rect 41802 39861 41808 39895
rect 41842 39861 41848 39895
rect 46101 39938 46357 39966
rect 46101 39892 46139 39938
rect 43269 39876 43327 39882
rect 43441 39876 43499 39882
rect 43613 39876 43671 39882
rect 43785 39876 43843 39882
rect 43957 39876 44015 39882
rect 44162 39876 44220 39882
rect 44339 39876 44397 39882
rect 44511 39876 44569 39882
rect 44683 39876 44741 39882
rect 44855 39876 44913 39882
rect 45027 39876 45085 39882
rect 45199 39876 45257 39882
rect 45864 39876 46139 39892
rect 41802 39823 41848 39861
rect 40116 39776 40174 39782
rect 40116 39742 40128 39776
rect 40162 39742 40174 39776
rect 40884 39750 40894 39802
rect 40946 39750 40956 39802
rect 41802 39789 41808 39823
rect 41842 39793 41848 39823
rect 42997 39826 43044 39870
rect 43269 39842 43281 39876
rect 43315 39842 43453 39876
rect 43487 39842 43625 39876
rect 43659 39842 43797 39876
rect 43831 39842 43969 39876
rect 44003 39842 44174 39876
rect 44208 39842 44351 39876
rect 44385 39842 44523 39876
rect 44557 39842 44695 39876
rect 44729 39842 44867 39876
rect 44901 39842 45039 39876
rect 45073 39842 45211 39876
rect 45245 39842 46139 39876
rect 43269 39836 43327 39842
rect 43441 39836 43499 39842
rect 43613 39836 43671 39842
rect 43785 39836 43843 39842
rect 43957 39836 44015 39842
rect 44162 39836 44220 39842
rect 44339 39836 44397 39842
rect 44511 39836 44569 39842
rect 44683 39836 44741 39842
rect 44855 39836 44913 39842
rect 45027 39836 45085 39842
rect 45199 39836 45257 39842
rect 45864 39828 46139 39842
rect 41842 39789 42948 39793
rect 41802 39787 42948 39789
rect 41802 39753 42539 39787
rect 42573 39753 42611 39787
rect 42645 39753 42683 39787
rect 42717 39753 42755 39787
rect 42789 39753 42827 39787
rect 42861 39753 42899 39787
rect 42933 39753 42948 39787
rect 41802 39751 42948 39753
rect 40116 39741 40174 39742
rect 39547 39736 40174 39741
rect 39547 39735 40162 39736
rect 39547 39683 39563 39735
rect 39615 39707 40162 39735
rect 41802 39717 41808 39751
rect 41842 39748 42948 39751
rect 41842 39717 41848 39748
rect 42525 39747 42948 39748
rect 42997 39792 43003 39826
rect 43037 39796 43044 39826
rect 43037 39792 43507 39796
rect 42997 39790 43507 39792
rect 42997 39756 43277 39790
rect 43311 39756 43349 39790
rect 43383 39756 43507 39790
rect 42997 39754 43507 39756
rect 39615 39683 39631 39707
rect 39547 39677 39631 39683
rect 41802 39679 41848 39717
rect 41802 39645 41808 39679
rect 41842 39645 41848 39679
rect 42997 39720 43003 39754
rect 43037 39750 43507 39754
rect 46101 39758 46139 39828
rect 46319 39758 46357 39938
rect 43037 39720 43044 39750
rect 46101 39730 46357 39758
rect 42997 39676 43044 39720
rect 41802 39624 41848 39645
rect 41420 39560 41798 39567
rect 41420 39508 41455 39560
rect 41507 39508 41519 39560
rect 41571 39508 41583 39560
rect 41635 39508 41647 39560
rect 41699 39508 41711 39560
rect 41763 39508 41798 39560
rect 41420 39502 41798 39508
rect 7072 39182 7328 39210
rect 7072 39002 7110 39182
rect 7290 39002 7328 39182
rect 7072 38974 7328 39002
rect 12532 39182 12788 39210
rect 12532 39002 12570 39182
rect 12750 39002 12788 39182
rect 12532 38974 12788 39002
rect 12660 38964 12778 38974
rect 7236 38155 7300 38168
rect 7226 38149 7310 38155
rect 7226 38097 7242 38149
rect 7294 38097 7310 38149
rect 7226 38091 7310 38097
rect 5419 37201 5503 37207
rect 5419 37149 5435 37201
rect 5487 37149 5503 37201
rect 5419 37143 5503 37149
rect 6691 37201 6775 37207
rect 6691 37149 6707 37201
rect 6759 37149 6775 37201
rect 6691 37143 6775 37149
rect 3572 36088 3821 36094
rect 3572 36036 3606 36088
rect 3658 36036 3670 36088
rect 3722 36036 3734 36088
rect 3786 36036 3821 36088
rect 3572 36030 3821 36036
rect 5045 36087 5361 36104
rect 5045 36035 5081 36087
rect 5133 36035 5145 36087
rect 5197 36035 5209 36087
rect 5261 36035 5273 36087
rect 5325 36035 5361 36087
rect 5045 36018 5361 36035
rect 5429 35945 5493 37143
rect 7236 36107 7300 38091
rect 9418 37645 9502 37651
rect 9418 37593 9434 37645
rect 9486 37593 9502 37645
rect 9418 37587 9502 37593
rect 5564 36088 5811 36097
rect 5564 36036 5597 36088
rect 5649 36036 5661 36088
rect 5713 36036 5725 36088
rect 5777 36036 5811 36088
rect 5564 36027 5811 36036
rect 6926 36080 7167 36089
rect 6926 36028 6956 36080
rect 7008 36028 7020 36080
rect 7072 36028 7084 36080
rect 7136 36028 7167 36080
rect 7373 36087 7691 36094
rect 7373 36035 7410 36087
rect 7462 36035 7474 36087
rect 7526 36035 7538 36087
rect 7590 36035 7602 36087
rect 7654 36035 7691 36087
rect 7373 36028 7691 36035
rect 8911 36086 9358 36093
rect 8911 36034 8948 36086
rect 9000 36034 9012 36086
rect 9064 36034 9076 36086
rect 9128 36034 9140 36086
rect 9192 36034 9204 36086
rect 9256 36034 9268 36086
rect 9320 36034 9358 36086
rect 8911 36028 9358 36034
rect 6926 36020 7167 36028
rect 9428 35940 9492 37587
rect 9565 36083 9812 36091
rect 9565 36031 9598 36083
rect 9650 36031 9662 36083
rect 9714 36031 9726 36083
rect 9778 36031 9812 36083
rect 9565 36023 9812 36031
rect 5420 35014 5504 35020
rect 5420 34962 5436 35014
rect 5488 34962 5504 35014
rect 5420 34956 5504 34962
rect 7232 35012 7316 35018
rect 7232 34960 7248 35012
rect 7300 34960 7316 35012
rect 7232 34954 7316 34960
rect 3866 34780 4878 34844
rect 7854 34781 8873 34845
rect 3745 33850 3797 34654
rect 3735 33798 3745 33850
rect 3797 33798 3807 33850
rect -6989 33121 -6942 33173
rect -6890 33121 -6861 33173
rect -6989 31811 -6861 33121
rect -6999 31805 -6851 31811
rect -6999 31753 -6983 31805
rect -6931 31753 -6919 31805
rect -6867 31753 -6851 31805
rect -6999 31747 -6851 31753
rect -6989 31712 -6861 31747
rect 4354 30432 4418 34780
rect 5420 34419 5504 34425
rect 5420 34367 5436 34419
rect 5488 34367 5504 34419
rect 5420 34361 5504 34367
rect 7232 34419 7316 34425
rect 7232 34367 7248 34419
rect 7300 34367 7316 34419
rect 7232 34361 7316 34367
rect 5430 33561 5494 34361
rect 7242 34328 7306 34361
rect 7242 34264 7492 34328
rect 7428 33569 7492 34264
rect 7418 33563 7502 33569
rect 5420 33555 5504 33561
rect 5420 33503 5436 33555
rect 5488 33503 5504 33555
rect 7418 33511 7434 33563
rect 7486 33511 7502 33563
rect 7418 33505 7502 33511
rect 5420 33497 5504 33503
rect 5430 33480 5494 33497
rect 8328 30437 8392 34781
rect 9745 33850 9797 34662
rect 9735 33798 9745 33850
rect 9797 33798 9807 33850
rect 9745 33795 9797 33798
rect 4344 30426 4428 30432
rect 4344 30374 4360 30426
rect 4412 30374 4428 30426
rect 4344 30368 4428 30374
rect 8318 30431 8402 30437
rect 8318 30379 8334 30431
rect 8386 30379 8402 30431
rect 8318 30373 8402 30379
rect -9407 30299 -9259 30305
rect -9407 30247 -9391 30299
rect -9339 30247 -9327 30299
rect -9275 30247 -9259 30299
rect -9407 30241 -9259 30247
rect -9398 30201 -9270 30241
rect -12703 29746 -12619 29752
rect -12703 29694 -12687 29746
rect -12635 29694 -12619 29746
rect -12703 29688 -12619 29694
rect -13479 29323 -13395 29329
rect -30209 29281 -18384 29288
rect -30209 29165 -30193 29281
rect -30077 29165 -18517 29281
rect -18401 29165 -18384 29281
rect -13479 29271 -13463 29323
rect -13411 29271 -13395 29323
rect -13479 29265 -13395 29271
rect -30209 29159 -18384 29165
rect 7950 28840 8034 28846
rect 1941 28802 2089 28808
rect 1941 28750 1957 28802
rect 2009 28750 2021 28802
rect 2073 28750 2089 28802
rect 7950 28788 7966 28840
rect 8018 28788 8034 28840
rect 7950 28782 8034 28788
rect 1941 28744 2089 28750
rect 1951 28644 2079 28744
rect -11888 28602 2079 28644
rect -11888 28550 -6080 28602
rect -6028 28550 -6016 28602
rect -5964 28550 2079 28602
rect -11888 28516 2079 28550
rect 3368 28589 3496 28627
rect 3368 28537 3405 28589
rect 3457 28537 3496 28589
rect -15722 28089 -15603 28098
rect -15722 28037 -15689 28089
rect -15637 28037 -15603 28089
rect -15722 28025 -15603 28037
rect -15722 27973 -15689 28025
rect -15637 27973 -15603 28025
rect -13993 28014 -13983 28066
rect -13931 28014 -13694 28066
rect -12399 28059 -12306 28076
rect -15722 27961 -15603 27973
rect -31040 27923 -19244 27930
rect -31040 27807 -31024 27923
rect -30908 27807 -19377 27923
rect -19261 27807 -19244 27923
rect -31040 27801 -19244 27807
rect -15722 27909 -15689 27961
rect -15637 27909 -15603 27961
rect -15722 27897 -15603 27909
rect -15722 27845 -15689 27897
rect -15637 27845 -15603 27897
rect -15722 27833 -15603 27845
rect -15722 27781 -15689 27833
rect -15637 27781 -15603 27833
rect -15722 27769 -15603 27781
rect -15722 27717 -15689 27769
rect -15637 27717 -15603 27769
rect -15722 27705 -15603 27717
rect -15722 27653 -15689 27705
rect -15637 27653 -15603 27705
rect -12399 28007 -12379 28059
rect -12327 28007 -12306 28059
rect -12399 27995 -12306 28007
rect -12399 27943 -12379 27995
rect -12327 27943 -12306 27995
rect -12399 27931 -12306 27943
rect -12399 27879 -12379 27931
rect -12327 27879 -12306 27931
rect -12399 27867 -12306 27879
rect -12399 27815 -12379 27867
rect -12327 27815 -12306 27867
rect -12399 27803 -12306 27815
rect -12399 27751 -12379 27803
rect -12327 27751 -12306 27803
rect -12399 27739 -12306 27751
rect -12399 27687 -12379 27739
rect -12327 27687 -12306 27739
rect -12399 27670 -12306 27687
rect -15722 27645 -15603 27653
rect -17645 27638 -17497 27644
rect -18326 27575 -18262 27600
rect -18336 27569 -18252 27575
rect -18336 27517 -18320 27569
rect -18268 27517 -18252 27569
rect -18336 27511 -18252 27517
rect -17645 27522 -17629 27638
rect -17513 27568 -17497 27638
rect -11888 27634 -11760 28516
rect -12206 27579 -11760 27634
rect -17513 27522 -17334 27568
rect -17645 27516 -17334 27522
rect -14916 27519 -14906 27571
rect -14854 27519 -13619 27571
rect -12491 27515 -11760 27579
rect -18326 27098 -18262 27511
rect -12206 27506 -11760 27515
rect -12404 27402 -12287 27427
rect -12404 27350 -12372 27402
rect -12320 27350 -12287 27402
rect -12404 27338 -12287 27350
rect -12404 27286 -12372 27338
rect -12320 27286 -12287 27338
rect -12404 27274 -12287 27286
rect -14414 27207 -14404 27259
rect -14352 27207 -13728 27259
rect -12404 27222 -12372 27274
rect -12320 27222 -12287 27274
rect -12404 27198 -12287 27222
rect -18336 27092 -18252 27098
rect -18336 27040 -18320 27092
rect -18268 27040 -18252 27092
rect -15239 27082 -14906 27083
rect -18336 27034 -18252 27040
rect -18891 26754 -18807 26760
rect -18891 26702 -18875 26754
rect -18823 26702 -18807 26754
rect -18891 26696 -18807 26702
rect -38200 26588 -34846 26611
rect -38200 26536 -38181 26588
rect -38129 26536 -38117 26588
rect -38065 26536 -38053 26588
rect -38001 26536 -37989 26588
rect -37937 26536 -37925 26588
rect -37873 26536 -37861 26588
rect -37809 26536 -37797 26588
rect -37745 26536 -37733 26588
rect -37681 26536 -37669 26588
rect -37617 26536 -37605 26588
rect -37553 26536 -37541 26588
rect -37489 26536 -37477 26588
rect -37425 26536 -37413 26588
rect -37361 26536 -37349 26588
rect -37297 26536 -37285 26588
rect -37233 26536 -37221 26588
rect -37169 26536 -37157 26588
rect -37105 26536 -37093 26588
rect -37041 26536 -37029 26588
rect -36977 26536 -36965 26588
rect -36913 26536 -36901 26588
rect -36849 26536 -36837 26588
rect -36785 26536 -36773 26588
rect -36721 26536 -36709 26588
rect -36657 26536 -36645 26588
rect -36593 26536 -36581 26588
rect -36529 26536 -36517 26588
rect -36465 26536 -36453 26588
rect -36401 26536 -36389 26588
rect -36337 26536 -36325 26588
rect -36273 26536 -36261 26588
rect -36209 26536 -36197 26588
rect -36145 26536 -36133 26588
rect -36081 26536 -36069 26588
rect -36017 26536 -36005 26588
rect -35953 26536 -35941 26588
rect -35889 26536 -35877 26588
rect -35825 26536 -35813 26588
rect -35761 26536 -35749 26588
rect -35697 26536 -35685 26588
rect -35633 26536 -35621 26588
rect -35569 26536 -35557 26588
rect -35505 26536 -35493 26588
rect -35441 26536 -35429 26588
rect -35377 26536 -35365 26588
rect -35313 26536 -35301 26588
rect -35249 26536 -35237 26588
rect -35185 26536 -35173 26588
rect -35121 26536 -35109 26588
rect -35057 26536 -35045 26588
rect -34993 26536 -34981 26588
rect -34929 26536 -34917 26588
rect -34865 26536 -34846 26588
rect -38200 26514 -34846 26536
rect -18881 25977 -18817 26696
rect -18892 25971 -18808 25977
rect -18892 25919 -18876 25971
rect -18824 25919 -18808 25971
rect -18892 25913 -18808 25919
rect -25459 25450 -25359 25482
rect -25459 25398 -25435 25450
rect -25383 25398 -25359 25450
rect -25459 25386 -25359 25398
rect -25459 25334 -25435 25386
rect -25383 25334 -25359 25386
rect -25459 25322 -25359 25334
rect -25459 25270 -25435 25322
rect -25383 25270 -25359 25322
rect -25459 25258 -25359 25270
rect -25459 25206 -25435 25258
rect -25383 25206 -25359 25258
rect -25459 25175 -25359 25206
rect -40603 25143 -40347 25171
rect -40603 24963 -40565 25143
rect -40385 25112 -40347 25143
rect -40385 25106 -26683 25112
rect -40385 24990 -32985 25106
rect -32869 24990 -26683 25106
rect -40385 24984 -26683 24990
rect -25335 24984 -24122 25112
rect -40385 24963 -40347 24984
rect -40603 24935 -40347 24963
rect -25462 24919 -25355 24945
rect -25462 24867 -25435 24919
rect -25383 24867 -25355 24919
rect -25462 24855 -25355 24867
rect -25462 24803 -25435 24855
rect -25383 24803 -25355 24855
rect -25462 24791 -25355 24803
rect -25462 24739 -25435 24791
rect -25383 24739 -25355 24791
rect -25462 24714 -25355 24739
rect -38192 23580 -34842 23605
rect -38192 23528 -38175 23580
rect -38123 23528 -38111 23580
rect -38059 23528 -38047 23580
rect -37995 23528 -37983 23580
rect -37931 23528 -37919 23580
rect -37867 23528 -37855 23580
rect -37803 23528 -37791 23580
rect -37739 23528 -37727 23580
rect -37675 23528 -37663 23580
rect -37611 23528 -37599 23580
rect -37547 23528 -37535 23580
rect -37483 23528 -37471 23580
rect -37419 23528 -37407 23580
rect -37355 23528 -37343 23580
rect -37291 23528 -37279 23580
rect -37227 23528 -37215 23580
rect -37163 23528 -37151 23580
rect -37099 23528 -37087 23580
rect -37035 23528 -37023 23580
rect -36971 23528 -36959 23580
rect -36907 23528 -36895 23580
rect -36843 23528 -36831 23580
rect -36779 23528 -36767 23580
rect -36715 23528 -36703 23580
rect -36651 23528 -36639 23580
rect -36587 23528 -36575 23580
rect -36523 23528 -36511 23580
rect -36459 23528 -36447 23580
rect -36395 23528 -36383 23580
rect -36331 23528 -36319 23580
rect -36267 23528 -36255 23580
rect -36203 23528 -36191 23580
rect -36139 23528 -36127 23580
rect -36075 23528 -36063 23580
rect -36011 23528 -35999 23580
rect -35947 23528 -35935 23580
rect -35883 23528 -35871 23580
rect -35819 23528 -35807 23580
rect -35755 23528 -35743 23580
rect -35691 23528 -35679 23580
rect -35627 23528 -35615 23580
rect -35563 23528 -35551 23580
rect -35499 23528 -35487 23580
rect -35435 23528 -35423 23580
rect -35371 23528 -35359 23580
rect -35307 23528 -35295 23580
rect -35243 23528 -35231 23580
rect -35179 23528 -35167 23580
rect -35115 23528 -35103 23580
rect -35051 23528 -35039 23580
rect -34987 23528 -34975 23580
rect -34923 23528 -34911 23580
rect -34859 23528 -34842 23580
rect -38192 23503 -34842 23528
rect -24250 21702 -24122 24984
rect -18881 24118 -18817 25913
rect -18326 24457 -18262 27034
rect -15242 27031 -14906 27082
rect -14854 27031 -14844 27083
rect -17266 26754 -17182 26760
rect -17266 26702 -17250 26754
rect -17198 26702 -17182 26754
rect -17266 26696 -17182 26702
rect -11912 26582 -9878 26588
rect -11912 26530 -10010 26582
rect -9958 26530 -9946 26582
rect -9894 26530 -9878 26582
rect -11912 26524 -9878 26530
rect -17645 26409 -17334 26415
rect -13993 26414 -13983 26466
rect -13931 26414 -13722 26466
rect -12406 26457 -12291 26486
rect -17645 26293 -17629 26409
rect -17513 26363 -17334 26409
rect -12406 26405 -12375 26457
rect -12323 26405 -12291 26457
rect -12406 26393 -12291 26405
rect -17513 26293 -17497 26363
rect -17645 26287 -17497 26293
rect -12406 26341 -12375 26393
rect -12323 26341 -12291 26393
rect -12406 26329 -12291 26341
rect -15735 26252 -15626 26281
rect -15735 26200 -15707 26252
rect -15655 26200 -15626 26252
rect -15735 26188 -15626 26200
rect -15735 26136 -15707 26188
rect -15655 26136 -15626 26188
rect -15735 26124 -15626 26136
rect -15735 26072 -15707 26124
rect -15655 26072 -15626 26124
rect -15735 26044 -15626 26072
rect -12406 26277 -12375 26329
rect -12323 26277 -12291 26329
rect -12406 26265 -12291 26277
rect -12406 26213 -12375 26265
rect -12323 26213 -12291 26265
rect -12406 26201 -12291 26213
rect -12406 26149 -12375 26201
rect -12323 26149 -12291 26201
rect -12406 26137 -12291 26149
rect -12406 26085 -12375 26137
rect -12323 26085 -12291 26137
rect -12406 26057 -12291 26085
rect -11912 25978 -11848 26524
rect -14916 25915 -14906 25967
rect -14854 25915 -13624 25967
rect -12478 25914 -11848 25978
rect -12394 25803 -12311 25823
rect 1952 25820 2080 25825
rect -12394 25751 -12379 25803
rect -12327 25751 -12311 25803
rect 1942 25814 2090 25820
rect 1942 25762 1958 25814
rect 2010 25762 2022 25814
rect 2074 25762 2090 25814
rect 1942 25756 2090 25762
rect -12394 25739 -12311 25751
rect -12394 25687 -12379 25739
rect -12327 25687 -12311 25739
rect -12394 25675 -12311 25687
rect -14414 25607 -14404 25659
rect -14352 25607 -13741 25659
rect -12394 25623 -12379 25675
rect -12327 25623 -12311 25675
rect -12394 25604 -12311 25623
rect 1952 25448 2080 25756
rect -15737 25418 -15622 25447
rect -15737 25366 -15706 25418
rect -15654 25366 -15622 25418
rect -15737 25354 -15622 25366
rect -15737 25302 -15706 25354
rect -15654 25302 -15622 25354
rect -15737 25290 -15622 25302
rect -15737 25238 -15706 25290
rect -15654 25238 -15622 25290
rect -15737 25226 -15622 25238
rect -15737 25174 -15706 25226
rect -15654 25174 -15622 25226
rect -15737 25162 -15622 25174
rect -15737 25110 -15706 25162
rect -15654 25110 -15622 25162
rect -15737 25098 -15622 25110
rect -15737 25046 -15706 25098
rect -15654 25046 -15622 25098
rect -15737 25018 -15622 25046
rect -11886 25408 2080 25448
rect -11886 25356 -3495 25408
rect -3443 25356 -3431 25408
rect -3379 25356 2080 25408
rect -11886 25320 2080 25356
rect -17645 24996 -17497 25002
rect -17645 24880 -17629 24996
rect -17513 24926 -17497 24996
rect -17513 24880 -17339 24926
rect -17645 24874 -17339 24880
rect -13993 24814 -13983 24866
rect -13931 24814 -13749 24866
rect -12403 24707 -12318 24712
rect -12403 24655 -12387 24707
rect -12335 24655 -12318 24707
rect -12403 24643 -12318 24655
rect -12403 24591 -12387 24643
rect -12335 24591 -12318 24643
rect -12403 24579 -12318 24591
rect -12403 24527 -12387 24579
rect -12335 24527 -12318 24579
rect -12403 24515 -12318 24527
rect -12403 24463 -12387 24515
rect -12335 24463 -12318 24515
rect -12403 24458 -12318 24463
rect -18336 24451 -18252 24457
rect -18336 24399 -18320 24451
rect -18268 24399 -18252 24451
rect -18336 24393 -18252 24399
rect -15202 24389 -14908 24441
rect -14856 24389 -14850 24441
rect -11886 24408 -11758 25320
rect -14908 24369 -14850 24389
rect -12198 24376 -11758 24408
rect -14908 24317 -13620 24369
rect -12469 24312 -11758 24376
rect -12198 24280 -11758 24312
rect -12408 24211 -12306 24239
rect -12408 24159 -12383 24211
rect -12331 24159 -12306 24211
rect -12408 24147 -12306 24159
rect -18891 24112 -18807 24118
rect -18891 24060 -18875 24112
rect -18823 24060 -18807 24112
rect -18891 24054 -18807 24060
rect -17273 24112 -17189 24118
rect -17273 24060 -17257 24112
rect -17205 24060 -17189 24112
rect -17273 24054 -17189 24060
rect -12408 24095 -12383 24147
rect -12331 24095 -12306 24147
rect -12408 24083 -12306 24095
rect -14414 24007 -14404 24059
rect -14352 24007 -13733 24059
rect -12408 24031 -12383 24083
rect -12331 24031 -12306 24083
rect -12408 24003 -12306 24031
rect 3368 24095 3496 28537
rect 7960 25820 8024 28782
rect 9366 28586 9494 28632
rect 9366 28534 9405 28586
rect 9457 28534 9494 28586
rect 7950 25814 8034 25820
rect 7950 25762 7966 25814
rect 8018 25762 8034 25814
rect 7950 25756 8034 25762
rect 5705 24576 5793 24594
rect 5705 24524 5723 24576
rect 5775 24524 5793 24576
rect 5705 24512 5793 24524
rect 5705 24460 5723 24512
rect 5775 24460 5793 24512
rect 5705 24448 5793 24460
rect 5705 24396 5723 24448
rect 5775 24396 5793 24448
rect 5705 24384 5793 24396
rect 5705 24332 5723 24384
rect 5775 24332 5793 24384
rect 5705 24320 5793 24332
rect 5705 24268 5723 24320
rect 5775 24268 5793 24320
rect 5705 24256 5793 24268
rect 5705 24204 5723 24256
rect 5775 24204 5793 24256
rect 5705 24186 5793 24204
rect 3368 24043 3405 24095
rect 3457 24043 3496 24095
rect -17645 23767 -17338 23773
rect -17645 23651 -17629 23767
rect -17513 23721 -17338 23767
rect -17513 23651 -17497 23721
rect -17645 23645 -17497 23651
rect -15735 23611 -15648 23637
rect -15735 23559 -15718 23611
rect -15666 23559 -15648 23611
rect -15735 23547 -15648 23559
rect -15735 23495 -15718 23547
rect -15666 23495 -15648 23547
rect -15735 23483 -15648 23495
rect -15735 23431 -15718 23483
rect -15666 23431 -15648 23483
rect -15735 23405 -15648 23431
rect 3368 23415 3496 24043
rect 5633 24091 5717 24097
rect 5633 24039 5649 24091
rect 5701 24039 5717 24091
rect 5633 24033 5717 24039
rect 7007 24095 7091 24101
rect 7007 24043 7023 24095
rect 7075 24043 7091 24095
rect 7007 24037 7091 24043
rect 9366 24095 9494 28534
rect 9366 24043 9405 24095
rect 9457 24043 9494 24095
rect 42846 24145 46200 24174
rect 42846 24093 42865 24145
rect 42917 24093 42929 24145
rect 42981 24093 42993 24145
rect 43045 24093 43057 24145
rect 43109 24093 43121 24145
rect 43173 24093 43185 24145
rect 43237 24093 43249 24145
rect 43301 24093 43313 24145
rect 43365 24093 43377 24145
rect 43429 24093 43441 24145
rect 43493 24093 43505 24145
rect 43557 24093 43569 24145
rect 43621 24093 43633 24145
rect 43685 24093 43697 24145
rect 43749 24093 43761 24145
rect 43813 24093 43825 24145
rect 43877 24093 43889 24145
rect 43941 24093 43953 24145
rect 44005 24093 44017 24145
rect 44069 24093 44081 24145
rect 44133 24093 44145 24145
rect 44197 24093 44209 24145
rect 44261 24093 44273 24145
rect 44325 24093 44337 24145
rect 44389 24093 44401 24145
rect 44453 24093 44465 24145
rect 44517 24093 44529 24145
rect 44581 24093 44593 24145
rect 44645 24093 44657 24145
rect 44709 24093 44721 24145
rect 44773 24093 44785 24145
rect 44837 24093 44849 24145
rect 44901 24093 44913 24145
rect 44965 24093 44977 24145
rect 45029 24093 45041 24145
rect 45093 24093 45105 24145
rect 45157 24093 45169 24145
rect 45221 24093 45233 24145
rect 45285 24093 45297 24145
rect 45349 24093 45361 24145
rect 45413 24093 45425 24145
rect 45477 24093 45489 24145
rect 45541 24093 45553 24145
rect 45605 24093 45617 24145
rect 45669 24093 45681 24145
rect 45733 24093 45745 24145
rect 45797 24093 45809 24145
rect 45861 24093 45873 24145
rect 45925 24093 45937 24145
rect 45989 24093 46001 24145
rect 46053 24093 46065 24145
rect 46117 24093 46129 24145
rect 46181 24093 46200 24145
rect 42846 24065 46200 24093
rect 5724 23395 5788 23661
rect 9366 23423 9494 24043
rect 35142 23860 35226 23866
rect 35142 23808 35158 23860
rect 35210 23808 35226 23860
rect 35142 23802 35226 23808
rect 39336 23693 39430 23714
rect 39336 23641 39357 23693
rect 39409 23641 39430 23693
rect 39336 23629 39430 23641
rect 37809 23609 37902 23611
rect 37809 23557 37829 23609
rect 37881 23557 37902 23609
rect 37809 23545 37902 23557
rect 37809 23493 37829 23545
rect 37881 23493 37902 23545
rect 39336 23577 39357 23629
rect 39409 23577 39430 23629
rect 39336 23565 39430 23577
rect 39336 23513 39357 23565
rect 39409 23513 39430 23565
rect 39336 23493 39430 23513
rect 37809 23492 37902 23493
rect 2550 23328 2850 23392
rect 3860 23331 9002 23395
rect -13993 23214 -13983 23266
rect -13931 23214 -13709 23266
rect -12399 23253 -12309 23277
rect -12399 23201 -12380 23253
rect -12328 23201 -12309 23253
rect -12399 23189 -12309 23201
rect -12399 23137 -12380 23189
rect -12328 23137 -12309 23189
rect -12399 23125 -12309 23137
rect -12399 23073 -12380 23125
rect -12328 23073 -12309 23125
rect -12399 23061 -12309 23073
rect 2550 23063 2614 23328
rect 8777 23327 8953 23331
rect 8777 23275 8807 23327
rect 8859 23275 8871 23327
rect 8923 23275 8953 23327
rect 10068 23326 10266 23390
rect 8777 23246 8953 23275
rect 10202 23063 10266 23326
rect 11296 23295 33935 23423
rect 39446 23303 39682 23431
rect -12399 23009 -12380 23061
rect -12328 23009 -12309 23061
rect -12399 22997 -12309 23009
rect 2540 23057 2624 23063
rect 2540 23005 2556 23057
rect 2608 23005 2624 23057
rect 2540 22999 2624 23005
rect 10192 23057 10276 23063
rect 10192 23005 10208 23057
rect 10260 23005 10276 23057
rect 10192 22999 10276 23005
rect -12399 22945 -12380 22997
rect -12328 22945 -12309 22997
rect -12399 22933 -12309 22945
rect -12399 22881 -12380 22933
rect -12328 22881 -12309 22933
rect -12399 22857 -12309 22881
rect -12465 22773 -11463 22776
rect -14918 22719 -14908 22771
rect -14856 22719 -13614 22771
rect -12460 22770 -11463 22773
rect -12460 22718 -11595 22770
rect -11543 22718 -11531 22770
rect -11479 22718 -11463 22770
rect -12460 22712 -11463 22718
rect -12401 22601 -12313 22624
rect -12401 22549 -12383 22601
rect -12331 22549 -12313 22601
rect -12401 22537 -12313 22549
rect -12401 22485 -12383 22537
rect -12331 22485 -12313 22537
rect -12401 22473 -12313 22485
rect -14414 22407 -14404 22459
rect -14352 22407 -13740 22459
rect -12401 22421 -12383 22473
rect -12331 22421 -12313 22473
rect -12401 22399 -12313 22421
rect 3395 22101 3459 22106
rect -24250 21665 -5931 21702
rect -24250 21613 -6080 21665
rect -6028 21613 -6016 21665
rect -5964 21613 -5931 21665
rect -24250 21574 -5931 21613
rect -24284 20803 -3339 20842
rect -24284 20751 -3495 20803
rect -3443 20751 -3431 20803
rect -3379 20751 -3339 20803
rect -24284 20714 -3339 20751
rect -38178 19052 -34851 19065
rect -38178 19000 -38141 19052
rect -38089 19000 -38077 19052
rect -38025 19000 -38013 19052
rect -37961 19000 -37949 19052
rect -37897 19000 -37885 19052
rect -37833 19000 -37821 19052
rect -37769 19000 -37757 19052
rect -37705 19000 -37693 19052
rect -37641 19000 -37629 19052
rect -37577 19000 -37565 19052
rect -37513 19000 -37501 19052
rect -37449 19000 -37437 19052
rect -37385 19000 -37373 19052
rect -37321 19000 -37309 19052
rect -37257 19000 -37245 19052
rect -37193 19000 -37181 19052
rect -37129 19000 -37117 19052
rect -37065 19000 -37053 19052
rect -37001 19000 -36989 19052
rect -36937 19000 -36925 19052
rect -36873 19000 -36861 19052
rect -36809 19000 -36797 19052
rect -36745 19000 -36733 19052
rect -36681 19000 -36669 19052
rect -36617 19000 -36605 19052
rect -36553 19000 -36541 19052
rect -36489 19000 -36477 19052
rect -36425 19000 -36413 19052
rect -36361 19000 -36349 19052
rect -36297 19000 -36285 19052
rect -36233 19000 -36221 19052
rect -36169 19000 -36157 19052
rect -36105 19000 -36093 19052
rect -36041 19000 -36029 19052
rect -35977 19000 -35965 19052
rect -35913 19000 -35901 19052
rect -35849 19000 -35837 19052
rect -35785 19000 -35773 19052
rect -35721 19000 -35709 19052
rect -35657 19000 -35645 19052
rect -35593 19000 -35581 19052
rect -35529 19000 -35517 19052
rect -35465 19000 -35453 19052
rect -35401 19000 -35389 19052
rect -35337 19000 -35325 19052
rect -35273 19000 -35261 19052
rect -35209 19000 -35197 19052
rect -35145 19000 -35133 19052
rect -35081 19000 -35069 19052
rect -35017 19000 -35005 19052
rect -34953 19000 -34941 19052
rect -34889 19000 -34851 19052
rect -38178 18987 -34851 19000
rect -25462 17896 -25377 17922
rect -25462 17844 -25446 17896
rect -25394 17844 -25377 17896
rect -25462 17832 -25377 17844
rect -25462 17780 -25446 17832
rect -25394 17780 -25377 17832
rect -25462 17768 -25377 17780
rect -25462 17716 -25446 17768
rect -25394 17716 -25377 17768
rect -25462 17704 -25377 17716
rect -25462 17652 -25446 17704
rect -25394 17652 -25377 17704
rect -40606 17602 -40350 17630
rect -25462 17627 -25377 17652
rect -40606 17422 -40568 17602
rect -40388 17582 -40350 17602
rect -40388 17576 -26675 17582
rect -24284 17579 -24156 20714
rect -454 20103 -370 20109
rect -454 20051 -438 20103
rect -386 20051 -370 20103
rect -454 20039 -370 20051
rect -454 19987 -438 20039
rect -386 19987 -370 20039
rect -454 19981 -370 19987
rect -444 18993 -380 19981
rect 1674 19404 1812 19410
rect 1674 19352 1690 19404
rect 1742 19352 1812 19404
rect 1674 19340 1812 19352
rect 1674 19288 1690 19340
rect 1742 19288 1812 19340
rect 1674 19282 1812 19288
rect 223 17766 307 17772
rect -40388 17460 -31124 17576
rect -31008 17460 -26675 17576
rect -40388 17454 -26675 17460
rect -40388 17422 -40350 17454
rect -25357 17451 -24156 17579
rect -821 17525 -757 17735
rect 223 17714 239 17766
rect 291 17714 307 17766
rect 223 17708 307 17714
rect -831 17519 -747 17525
rect -831 17467 -815 17519
rect -763 17467 -747 17519
rect -831 17461 -747 17467
rect -40606 17394 -40350 17422
rect -25460 17376 -25368 17404
rect -25460 17324 -25440 17376
rect -25388 17324 -25368 17376
rect -25460 17312 -25368 17324
rect -25460 17260 -25440 17312
rect -25388 17260 -25368 17312
rect -25460 17248 -25368 17260
rect -25460 17196 -25440 17248
rect -25388 17196 -25368 17248
rect -445 17221 -381 17690
rect 1684 17221 1812 19282
rect 3361 19340 3489 22101
rect 4387 21985 4397 22037
rect 4449 21985 4459 22037
rect 8218 21985 8228 22037
rect 8280 21985 8290 22037
rect 4397 20945 4449 21985
rect 8228 20945 8280 21985
rect 4387 20893 4397 20945
rect 4449 20893 4459 20945
rect 8218 20893 8228 20945
rect 8280 20893 8290 20945
rect 8228 20883 8280 20893
rect 5384 20103 5468 20109
rect 5384 20051 5400 20103
rect 5452 20051 5468 20103
rect 5384 20039 5468 20051
rect 5384 19987 5400 20039
rect 5452 19987 5468 20039
rect 5384 19981 5468 19987
rect 9363 20103 9491 22105
rect 9363 20051 9400 20103
rect 9452 20051 9491 20103
rect 9363 20039 9491 20051
rect 9363 19987 9400 20039
rect 9452 19987 9491 20039
rect 3361 19288 3401 19340
rect 3453 19288 3489 19340
rect 3051 19100 3135 19106
rect 3051 19048 3067 19100
rect 3119 19048 3135 19100
rect 3361 19072 3489 19288
rect 4847 19158 5204 19173
rect 3051 19042 3135 19048
rect 3883 18987 4359 19051
rect 4847 19042 4871 19158
rect 5179 19042 5204 19158
rect 5394 19098 5458 19981
rect 7384 19404 7468 19410
rect 7384 19352 7400 19404
rect 7452 19352 7468 19404
rect 7384 19340 7468 19352
rect 7384 19288 7400 19340
rect 7452 19288 7468 19340
rect 7384 19282 7468 19288
rect 7075 19100 7159 19106
rect 7394 19103 7458 19282
rect 4847 19027 5204 19042
rect 5882 18991 6291 19055
rect 7075 19048 7091 19100
rect 7143 19048 7159 19100
rect 8971 19100 9055 19106
rect 7075 19042 7159 19048
rect -25460 17169 -25368 17196
rect -455 17215 -371 17221
rect -455 17163 -439 17215
rect -387 17163 -371 17215
rect -455 17151 -371 17163
rect -455 17099 -439 17151
rect -387 17099 -371 17151
rect -455 17093 -371 17099
rect 1674 17215 1812 17221
rect 1674 17163 1690 17215
rect 1742 17163 1812 17215
rect 1674 17151 1812 17163
rect 1674 17099 1690 17151
rect 1742 17099 1812 17151
rect 1674 17093 1812 17099
rect 3393 16866 3457 17769
rect 4295 17289 4359 18987
rect 4285 17283 4369 17289
rect 4285 17231 4301 17283
rect 4353 17231 4369 17283
rect 4285 17225 4369 17231
rect 5393 16866 5457 17768
rect 6227 17289 6291 18991
rect 7877 18989 8344 19053
rect 8971 19048 8987 19100
rect 9039 19048 9055 19100
rect 9363 19074 9491 19987
rect 11296 19412 11424 23295
rect 39325 23198 39431 23200
rect 37809 23192 37915 23194
rect 37809 23140 37836 23192
rect 37888 23140 37915 23192
rect 37809 23128 37915 23140
rect 37809 23076 37836 23128
rect 37888 23076 37915 23128
rect 37809 23064 37915 23076
rect 37809 23012 37836 23064
rect 37888 23012 37915 23064
rect 37809 23000 37915 23012
rect 37809 22948 37836 23000
rect 37888 22948 37915 23000
rect 39325 23146 39352 23198
rect 39404 23146 39431 23198
rect 39325 23134 39431 23146
rect 39325 23082 39352 23134
rect 39404 23082 39431 23134
rect 39325 23070 39431 23082
rect 39325 23018 39352 23070
rect 39404 23018 39431 23070
rect 39325 23006 39431 23018
rect 39325 22954 39352 23006
rect 39404 22954 39431 23006
rect 39325 22952 39431 22954
rect 37809 22946 37915 22948
rect 35090 22610 35100 22790
rect 35280 22610 35290 22790
rect 35750 22725 36031 22730
rect 35750 22673 35768 22725
rect 35820 22673 35832 22725
rect 35884 22673 35896 22725
rect 35948 22673 35960 22725
rect 36012 22673 36031 22725
rect 35750 22668 36031 22673
rect 39554 22677 39682 23303
rect 47546 22706 47802 22734
rect 47546 22677 47584 22706
rect 39554 22549 47584 22677
rect 39336 22367 39430 22388
rect 39336 22315 39357 22367
rect 39409 22315 39430 22367
rect 39336 22303 39430 22315
rect 37816 22273 37906 22280
rect 37816 22221 37835 22273
rect 37887 22221 37906 22273
rect 37816 22209 37906 22221
rect 37816 22157 37835 22209
rect 37887 22157 37906 22209
rect 39336 22251 39357 22303
rect 39409 22251 39430 22303
rect 39336 22239 39430 22251
rect 39336 22187 39357 22239
rect 39409 22187 39430 22239
rect 39336 22167 39430 22187
rect 37816 22151 37906 22157
rect 12373 21996 33915 22124
rect 39556 22107 39684 22549
rect 47546 22526 47584 22549
rect 47764 22526 47802 22706
rect 47546 22498 47802 22526
rect 12373 20111 12501 21996
rect 39464 21979 39684 22107
rect 39331 21832 39437 21834
rect 37804 21812 37909 21823
rect 37804 21760 37830 21812
rect 37882 21760 37909 21812
rect 37804 21748 37909 21760
rect 37804 21696 37830 21748
rect 37882 21696 37909 21748
rect 37804 21684 37909 21696
rect 37804 21632 37830 21684
rect 37882 21632 37909 21684
rect 37804 21621 37909 21632
rect 39331 21780 39358 21832
rect 39410 21780 39437 21832
rect 39331 21768 39437 21780
rect 39331 21716 39358 21768
rect 39410 21716 39437 21768
rect 39331 21704 39437 21716
rect 39331 21652 39358 21704
rect 39410 21652 39437 21704
rect 39331 21640 39437 21652
rect 39331 21588 39358 21640
rect 39410 21588 39437 21640
rect 39331 21586 39437 21588
rect 35142 21579 35226 21585
rect 35142 21527 35158 21579
rect 35210 21527 35226 21579
rect 35142 21521 35226 21527
rect 42844 21149 46198 21178
rect 42844 21097 42863 21149
rect 42915 21097 42927 21149
rect 42979 21097 42991 21149
rect 43043 21097 43055 21149
rect 43107 21097 43119 21149
rect 43171 21097 43183 21149
rect 43235 21097 43247 21149
rect 43299 21097 43311 21149
rect 43363 21097 43375 21149
rect 43427 21097 43439 21149
rect 43491 21097 43503 21149
rect 43555 21097 43567 21149
rect 43619 21097 43631 21149
rect 43683 21097 43695 21149
rect 43747 21097 43759 21149
rect 43811 21097 43823 21149
rect 43875 21097 43887 21149
rect 43939 21097 43951 21149
rect 44003 21097 44015 21149
rect 44067 21097 44079 21149
rect 44131 21097 44143 21149
rect 44195 21097 44207 21149
rect 44259 21097 44271 21149
rect 44323 21097 44335 21149
rect 44387 21097 44399 21149
rect 44451 21097 44463 21149
rect 44515 21097 44527 21149
rect 44579 21097 44591 21149
rect 44643 21097 44655 21149
rect 44707 21097 44719 21149
rect 44771 21097 44783 21149
rect 44835 21097 44847 21149
rect 44899 21097 44911 21149
rect 44963 21097 44975 21149
rect 45027 21097 45039 21149
rect 45091 21097 45103 21149
rect 45155 21097 45167 21149
rect 45219 21097 45231 21149
rect 45283 21097 45295 21149
rect 45347 21097 45359 21149
rect 45411 21097 45423 21149
rect 45475 21097 45487 21149
rect 45539 21097 45551 21149
rect 45603 21097 45615 21149
rect 45667 21097 45679 21149
rect 45731 21097 45743 21149
rect 45795 21097 45807 21149
rect 45859 21097 45871 21149
rect 45923 21097 45935 21149
rect 45987 21097 45999 21149
rect 46051 21097 46063 21149
rect 46115 21097 46127 21149
rect 46179 21097 46198 21149
rect 42844 21069 46198 21097
rect 14678 21021 14762 21027
rect 14678 20969 14694 21021
rect 14746 20969 14762 21021
rect 14678 20963 14762 20969
rect 14688 20497 14752 20963
rect 23660 20210 23744 20216
rect 23660 20158 23676 20210
rect 23728 20158 23744 20210
rect 23660 20152 23744 20158
rect 12363 20105 12511 20111
rect 12363 19989 12379 20105
rect 12495 19989 12511 20105
rect 12363 19983 12511 19989
rect 11285 19406 11433 19412
rect 11285 19290 11301 19406
rect 11417 19290 11433 19406
rect 23679 19376 23763 19382
rect 23679 19324 23695 19376
rect 23747 19324 23763 19376
rect 23679 19318 23763 19324
rect 11285 19284 11433 19290
rect 11296 19261 11424 19284
rect 8971 19042 9055 19048
rect 9877 19052 10306 19058
rect 9877 19000 10238 19052
rect 10290 19000 10306 19052
rect 9877 18994 10306 19000
rect 8280 18718 8344 18989
rect 8270 18712 8354 18718
rect 8270 18660 8286 18712
rect 8338 18660 8354 18712
rect 14667 18688 14701 18743
rect 8270 18654 8354 18660
rect 13564 18682 14728 18688
rect 13564 18630 13580 18682
rect 13632 18630 14728 18682
rect 13564 18624 14728 18630
rect 23648 18422 23732 18428
rect 23648 18370 23664 18422
rect 23716 18370 23732 18422
rect 23648 18364 23732 18370
rect 13877 17983 13961 18047
rect 7393 17359 7457 17775
rect 9396 17359 9460 17774
rect 23679 17546 23763 17552
rect 23679 17494 23695 17546
rect 23747 17494 23763 17546
rect 23679 17488 23763 17494
rect 7383 17353 7467 17359
rect 7383 17301 7399 17353
rect 7451 17301 7467 17353
rect 7383 17289 7467 17301
rect 6217 17283 6301 17289
rect 6217 17231 6233 17283
rect 6285 17231 6301 17283
rect 7383 17237 7399 17289
rect 7451 17237 7467 17289
rect 7383 17231 7467 17237
rect 9386 17353 9470 17359
rect 9386 17301 9402 17353
rect 9454 17301 9470 17353
rect 9386 17289 9470 17301
rect 9386 17237 9402 17289
rect 9454 17237 9470 17289
rect 9386 17231 9470 17237
rect 13875 17353 13959 17359
rect 13875 17301 13891 17353
rect 13943 17301 13959 17353
rect 13875 17289 13959 17301
rect 13875 17237 13891 17289
rect 13943 17237 13959 17289
rect 13875 17231 13959 17237
rect 6217 17225 6301 17231
rect 14680 17077 14764 17083
rect 14680 17025 14696 17077
rect 14748 17025 14764 17077
rect 14680 17019 14764 17025
rect 14690 16894 14754 17019
rect 3383 16860 3467 16866
rect 3383 16808 3399 16860
rect 3451 16808 3467 16860
rect 3383 16796 3467 16808
rect 3383 16744 3399 16796
rect 3451 16744 3467 16796
rect 3383 16738 3467 16744
rect 5383 16860 5467 16866
rect 5383 16808 5399 16860
rect 5451 16808 5467 16860
rect 5383 16796 5467 16808
rect 5383 16744 5399 16796
rect 5451 16744 5467 16796
rect 5383 16738 5467 16744
rect 13267 16860 13351 16866
rect 13267 16808 13283 16860
rect 13335 16808 13351 16860
rect 13267 16796 13351 16808
rect 13267 16744 13283 16796
rect 13335 16744 13351 16796
rect 13267 16738 13351 16744
rect 23062 16656 23727 16720
rect 241 16432 11149 16446
rect -3926 16288 -3862 16297
rect -3936 16282 -3852 16288
rect -3936 16230 -3920 16282
rect -3868 16230 -3852 16282
rect 241 16252 261 16432
rect 11129 16252 11149 16432
rect 241 16238 11149 16252
rect -3936 16224 -3852 16230
rect 18 16160 197 16189
rect -38184 16057 -34842 16075
rect -38184 16005 -38171 16057
rect -38119 16005 -38107 16057
rect -38055 16005 -38043 16057
rect -37991 16005 -37979 16057
rect -37927 16005 -37915 16057
rect -37863 16005 -37851 16057
rect -37799 16005 -37787 16057
rect -37735 16005 -37723 16057
rect -37671 16005 -37659 16057
rect -37607 16005 -37595 16057
rect -37543 16005 -37531 16057
rect -37479 16005 -37467 16057
rect -37415 16005 -37403 16057
rect -37351 16005 -37339 16057
rect -37287 16005 -37275 16057
rect -37223 16005 -37211 16057
rect -37159 16005 -37147 16057
rect -37095 16005 -37083 16057
rect -37031 16005 -37019 16057
rect -36967 16005 -36955 16057
rect -36903 16005 -36891 16057
rect -36839 16005 -36827 16057
rect -36775 16005 -36763 16057
rect -36711 16005 -36699 16057
rect -36647 16005 -36635 16057
rect -36583 16005 -36571 16057
rect -36519 16005 -36507 16057
rect -36455 16005 -36443 16057
rect -36391 16005 -36379 16057
rect -36327 16005 -36315 16057
rect -36263 16005 -36251 16057
rect -36199 16005 -36187 16057
rect -36135 16005 -36123 16057
rect -36071 16005 -36059 16057
rect -36007 16005 -35995 16057
rect -35943 16005 -35931 16057
rect -35879 16005 -35867 16057
rect -35815 16005 -35803 16057
rect -35751 16005 -35739 16057
rect -35687 16005 -35675 16057
rect -35623 16005 -35611 16057
rect -35559 16005 -35547 16057
rect -35495 16005 -35483 16057
rect -35431 16005 -35419 16057
rect -35367 16005 -35355 16057
rect -35303 16005 -35291 16057
rect -35239 16005 -35227 16057
rect -35175 16005 -35163 16057
rect -35111 16005 -35099 16057
rect -35047 16005 -35035 16057
rect -34983 16005 -34971 16057
rect -34919 16005 -34907 16057
rect -34855 16005 -34842 16057
rect -38184 15987 -34842 16005
rect -5787 15708 -3049 15709
rect -5796 15702 -3049 15708
rect -5796 15650 -5780 15702
rect -5728 15650 -3049 15702
rect -5796 15645 -3049 15650
rect -5796 15644 -5712 15645
rect -3113 15543 -3049 15645
rect -3927 15083 -3914 15135
rect -3862 15083 -2971 15135
rect -1824 15084 -678 15136
rect -626 15084 -616 15136
rect -3154 14980 -3051 14998
rect -3154 14928 -3129 14980
rect -3077 14928 -3051 14980
rect -3154 14916 -3051 14928
rect -3154 14864 -3129 14916
rect -3077 14864 -3051 14916
rect -3154 14852 -3051 14864
rect -3154 14800 -3129 14852
rect -3077 14800 -3051 14852
rect -3154 14788 -3051 14800
rect -3154 14736 -3129 14788
rect -3077 14736 -3051 14788
rect -3154 14719 -3051 14736
rect -25527 14423 -25434 14446
rect -25527 14371 -25507 14423
rect -25455 14371 -25434 14423
rect -25527 14359 -25434 14371
rect -25527 14307 -25507 14359
rect -25455 14307 -25434 14359
rect -25527 14295 -25434 14307
rect -25527 14243 -25507 14295
rect -25455 14243 -25434 14295
rect -25527 14231 -25434 14243
rect -4912 14431 -4822 14446
rect -4912 14379 -4893 14431
rect -4841 14379 -4822 14431
rect -4912 14367 -4822 14379
rect -4912 14315 -4893 14367
rect -4841 14315 -4822 14367
rect -4912 14303 -4822 14315
rect -4912 14251 -4893 14303
rect -4841 14251 -4822 14303
rect -4912 14236 -4822 14251
rect -25527 14179 -25507 14231
rect -25455 14179 -25434 14231
rect -25527 14157 -25434 14179
rect -13074 14135 -6287 14141
rect -33001 14096 -26755 14102
rect -33001 13980 -32985 14096
rect -32869 13980 -26755 14096
rect -25361 14073 -18140 14105
rect -13074 14083 -13058 14135
rect -13006 14083 -6538 14135
rect -6486 14083 -6287 14135
rect -4816 14087 -3914 14139
rect -3862 14087 -3852 14139
rect -13074 14077 -6287 14083
rect -25592 14067 -18140 14073
rect -25592 14015 -18217 14067
rect -18165 14015 -18140 14067
rect -25592 14009 -18140 14015
rect -33001 13974 -26755 13980
rect -25361 13977 -18140 14009
rect -4927 13974 -4823 13998
rect -25528 13897 -25436 13925
rect -25528 13845 -25508 13897
rect -25456 13845 -25436 13897
rect -25528 13833 -25436 13845
rect -25528 13781 -25508 13833
rect -25456 13781 -25436 13833
rect -25528 13769 -25436 13781
rect -25528 13717 -25508 13769
rect -25456 13717 -25436 13769
rect -25528 13690 -25436 13717
rect -4927 13922 -4901 13974
rect -4849 13922 -4823 13974
rect -4927 13910 -4823 13922
rect -4927 13858 -4901 13910
rect -4849 13858 -4823 13910
rect -4927 13846 -4823 13858
rect -4927 13794 -4901 13846
rect -4849 13794 -4823 13846
rect -4927 13782 -4823 13794
rect -4927 13730 -4901 13782
rect -4849 13730 -4823 13782
rect -4927 13706 -4823 13730
rect -1818 13115 -1715 13133
rect -1818 13063 -1793 13115
rect -1741 13063 -1715 13115
rect -1818 13051 -1715 13063
rect -1818 12999 -1793 13051
rect -1741 12999 -1715 13051
rect -1818 12987 -1715 12999
rect -1818 12935 -1793 12987
rect -1741 12935 -1715 12987
rect -1818 12923 -1715 12935
rect -6554 12886 -5777 12892
rect -6554 12834 -6538 12886
rect -6486 12834 -5845 12886
rect -5793 12834 -5777 12886
rect -6554 12828 -5777 12834
rect -1818 12871 -1793 12923
rect -1741 12871 -1715 12923
rect -1818 12859 -1715 12871
rect -1818 12807 -1793 12859
rect -1741 12807 -1715 12859
rect -1818 12795 -1715 12807
rect -1818 12743 -1793 12795
rect -1741 12743 -1715 12795
rect -1818 12726 -1715 12743
rect -3914 12635 -3027 12636
rect -3924 12583 -3914 12635
rect -3862 12583 -3027 12635
rect -1725 12585 -279 12637
rect -227 12585 -217 12637
rect -1785 12403 -1424 12409
rect -1785 12351 -1492 12403
rect -1440 12351 -1424 12403
rect -1785 12345 -1424 12351
rect -5861 12213 -5777 12219
rect -5861 12161 -5845 12213
rect -5793 12161 -5777 12213
rect -5861 12155 -5777 12161
rect -1798 11529 -1703 11530
rect -1798 11520 -1683 11529
rect -1798 11468 -1752 11520
rect -1700 11468 -1683 11520
rect -1798 11456 -1683 11468
rect -1798 11404 -1752 11456
rect -1700 11404 -1683 11456
rect -1798 11392 -1683 11404
rect -1798 11340 -1752 11392
rect -1700 11340 -1683 11392
rect -1798 11328 -1683 11340
rect -1798 11276 -1752 11328
rect -1700 11276 -1683 11328
rect -1798 11264 -1683 11276
rect -1798 11212 -1752 11264
rect -1700 11212 -1683 11264
rect -1798 11200 -1683 11212
rect -1798 11148 -1752 11200
rect -1700 11148 -1683 11200
rect -1798 11140 -1683 11148
rect -1798 11139 -1703 11140
rect -3425 10982 -3415 11034
rect -3363 10982 -3032 11034
rect -1724 10983 -279 11035
rect -227 10983 -217 11035
rect -5855 10891 -5845 10943
rect -5793 10891 -5783 10943
rect -6172 10821 -5927 10833
rect -6172 10769 -6140 10821
rect -6088 10769 -6076 10821
rect -6024 10769 -6012 10821
rect -5960 10769 -5927 10821
rect -6172 10758 -5927 10769
rect -5717 10820 -5391 10838
rect -5717 10768 -5676 10820
rect -5624 10768 -5612 10820
rect -5560 10768 -5548 10820
rect -5496 10768 -5484 10820
rect -5432 10768 -5391 10820
rect -5717 10751 -5391 10768
rect -1803 10777 -1424 10783
rect -1803 10725 -1492 10777
rect -1440 10725 -1424 10777
rect -1803 10719 -1424 10725
rect 18 10668 49 16160
rect 165 10668 197 16160
rect 11229 16163 11409 16184
rect 11229 14447 11261 16163
rect 11377 14447 11409 16163
rect 23062 15496 23126 16656
rect 23676 15782 23760 15788
rect 23676 15730 23692 15782
rect 23744 15730 23760 15782
rect 23676 15724 23760 15730
rect 20918 15490 23763 15496
rect 20918 15438 20934 15490
rect 20986 15438 23763 15490
rect 20918 15432 23763 15438
rect 14680 15222 14764 15228
rect 14680 15170 14696 15222
rect 14748 15170 14764 15222
rect 14680 15164 14764 15170
rect 14690 15130 14754 15164
rect 23699 15092 23763 15432
rect 11229 14432 11303 14447
rect 11337 14432 11409 14447
rect 11229 14426 11409 14432
rect 11268 14420 11373 14426
rect 23676 13991 23760 13997
rect 11268 13954 11373 13965
rect 14675 13959 14759 13965
rect 11247 13946 11394 13954
rect 11247 12998 11262 13946
rect 11378 12998 11394 13946
rect 14675 13907 14691 13959
rect 14743 13907 14759 13959
rect 23676 13939 23692 13991
rect 23744 13939 23760 13991
rect 23676 13933 23760 13939
rect 14675 13901 14759 13907
rect 14680 13522 14764 13528
rect 14680 13470 14696 13522
rect 14748 13470 14764 13522
rect 14680 13464 14764 13470
rect 14690 13327 14754 13464
rect 11247 12990 11394 12998
rect 23675 13000 23759 13006
rect 11268 12977 11373 12990
rect 23675 12948 23691 13000
rect 23743 12948 23759 13000
rect 23675 12942 23759 12948
rect 23681 12184 23765 12190
rect 14692 12174 14776 12180
rect 11233 12100 11408 12129
rect 14692 12122 14708 12174
rect 14760 12122 14776 12174
rect 23681 12132 23697 12184
rect 23749 12132 23765 12184
rect 23681 12126 23765 12132
rect 14692 12116 14776 12122
rect 11233 11344 11262 12100
rect 11378 11344 11408 12100
rect 14682 11670 14766 11676
rect 14682 11618 14698 11670
rect 14750 11618 14766 11670
rect 14682 11612 14766 11618
rect 14692 11520 14756 11612
rect 23679 11513 23763 11519
rect 23679 11461 23695 11513
rect 23747 11461 23763 11513
rect 23679 11455 23763 11461
rect 11233 11337 11303 11344
rect 11337 11337 11408 11344
rect 11233 11316 11408 11337
rect 11268 11311 11373 11316
rect 18 10640 197 10668
rect 5662 10402 5714 11030
rect -5855 10401 -678 10402
rect -5855 10349 -5845 10401
rect -5793 10350 -678 10401
rect -626 10350 5714 10402
rect 6484 10472 11218 10536
rect 6484 10438 6572 10472
rect 6606 10438 6644 10472
rect 6678 10438 6716 10472
rect 6750 10438 6788 10472
rect 6822 10438 6860 10472
rect 6894 10438 6932 10472
rect 6966 10438 7004 10472
rect 7038 10438 7076 10472
rect 7110 10438 7148 10472
rect 7182 10438 7220 10472
rect 7254 10438 7292 10472
rect 7326 10438 7364 10472
rect 7398 10438 7436 10472
rect 7470 10438 7508 10472
rect 7542 10438 7580 10472
rect 7614 10438 7652 10472
rect 7686 10438 7724 10472
rect 7758 10438 7796 10472
rect 7830 10438 7868 10472
rect 7902 10438 7940 10472
rect 7974 10438 8012 10472
rect 8046 10438 8084 10472
rect 8118 10438 8156 10472
rect 8190 10438 8228 10472
rect 8262 10438 8300 10472
rect 8334 10438 8372 10472
rect 8406 10438 8444 10472
rect 8478 10438 8516 10472
rect 8550 10438 8588 10472
rect 8622 10438 8660 10472
rect 8694 10438 8732 10472
rect 8766 10438 8804 10472
rect 8838 10438 8876 10472
rect 8910 10438 8948 10472
rect 8982 10438 9020 10472
rect 9054 10438 9092 10472
rect 9126 10438 9164 10472
rect 9198 10438 9236 10472
rect 9270 10438 9308 10472
rect 9342 10438 9380 10472
rect 9414 10438 9452 10472
rect 9486 10438 9524 10472
rect 9558 10438 9596 10472
rect 9630 10438 9668 10472
rect 9702 10438 9740 10472
rect 9774 10438 9812 10472
rect 9846 10438 9884 10472
rect 9918 10438 9956 10472
rect 9990 10438 10028 10472
rect 10062 10438 10100 10472
rect 10134 10438 10172 10472
rect 10206 10438 10244 10472
rect 10278 10438 10316 10472
rect 10350 10438 10388 10472
rect 10422 10438 10460 10472
rect 10494 10438 10532 10472
rect 10566 10438 10604 10472
rect 10638 10438 10676 10472
rect 10710 10438 10748 10472
rect 10782 10438 10820 10472
rect 10854 10438 10892 10472
rect 10926 10438 10964 10472
rect 10998 10438 11036 10472
rect 11070 10438 11218 10472
rect 6484 10357 11218 10438
rect 14681 10377 14765 10383
rect -5793 10349 5714 10350
rect 14681 10325 14697 10377
rect 14749 10325 14765 10377
rect 14681 10319 14765 10325
rect 23681 10374 23765 10380
rect 23681 10322 23697 10374
rect 23749 10322 23765 10374
rect 23681 10316 23765 10322
rect -1769 9917 -1685 9930
rect -1769 9865 -1753 9917
rect -1701 9865 -1685 9917
rect 3748 9911 5267 9945
rect -1769 9853 -1685 9865
rect -1769 9801 -1753 9853
rect -1701 9801 -1685 9853
rect -1769 9789 -1685 9801
rect -1769 9737 -1753 9789
rect -1701 9737 -1685 9789
rect 5233 9756 5267 9911
rect -1769 9725 -1685 9737
rect -1769 9673 -1753 9725
rect -1701 9673 -1685 9725
rect -1769 9661 -1685 9673
rect -1769 9609 -1753 9661
rect -1701 9609 -1685 9661
rect -1769 9597 -1685 9609
rect -6177 9578 -5919 9592
rect -6177 9526 -6138 9578
rect -6086 9526 -6074 9578
rect -6022 9526 -6010 9578
rect -5958 9526 -5919 9578
rect -6177 9513 -5919 9526
rect -5718 9578 -5389 9595
rect -5718 9526 -5708 9578
rect -5656 9526 -5644 9578
rect -5592 9526 -5580 9578
rect -5528 9526 -5516 9578
rect -5464 9526 -5452 9578
rect -5400 9526 -5389 9578
rect -1769 9545 -1753 9597
rect -1701 9545 -1685 9597
rect -1769 9532 -1685 9545
rect 5231 9669 5267 9756
rect -5718 9509 -5389 9526
rect -5855 9400 -5845 9452
rect -5793 9400 -5783 9452
rect -3924 9385 -3914 9437
rect -3862 9385 -3040 9437
rect -1726 9383 -1149 9435
rect -1097 9383 -1087 9435
rect 5231 9418 5265 9669
rect 24534 9418 24618 9424
rect 5213 9417 5286 9418
rect 5213 9365 5223 9417
rect 5275 9365 5286 9417
rect 24534 9366 24550 9418
rect 24602 9366 24618 9418
rect 24534 9360 24618 9366
rect -1779 9119 -1424 9125
rect -1779 9067 -1492 9119
rect -1440 9067 -1424 9119
rect -1779 9061 -1424 9067
rect -1768 8316 -1680 8330
rect -1768 8264 -1750 8316
rect -1698 8264 -1680 8316
rect -1768 8252 -1680 8264
rect -1768 8200 -1750 8252
rect -1698 8200 -1680 8252
rect -1768 8188 -1680 8200
rect -5863 8168 -5779 8174
rect -5863 8116 -5847 8168
rect -5795 8116 -5779 8168
rect -5863 8110 -5779 8116
rect -1768 8136 -1750 8188
rect -1698 8136 -1680 8188
rect -1768 8124 -1680 8136
rect -1768 8072 -1750 8124
rect -1698 8072 -1680 8124
rect -1768 8060 -1680 8072
rect -1768 8008 -1750 8060
rect -1698 8008 -1680 8060
rect -1768 7996 -1680 8008
rect -1768 7944 -1750 7996
rect -1698 7944 -1680 7996
rect -1768 7930 -1680 7944
rect 23198 7844 23271 7845
rect -3425 7783 -3415 7835
rect -3363 7783 -3029 7835
rect -1726 7783 -1149 7835
rect -1097 7783 -1087 7835
rect 23198 7792 23208 7844
rect 23260 7792 23271 7844
rect -6572 7591 -5779 7595
rect -6575 7589 -5779 7591
rect -6575 7585 -5847 7589
rect -6575 7533 -6559 7585
rect -6507 7537 -5847 7585
rect -5795 7537 -5779 7589
rect -6507 7533 -5779 7537
rect -6575 7531 -5779 7533
rect -1796 7580 -1424 7586
rect -6575 7527 -6491 7531
rect -1796 7528 -1492 7580
rect -1440 7528 -1424 7580
rect -1796 7522 -1424 7528
rect -7224 7213 -6741 7243
rect -7224 7033 -7201 7213
rect -6765 7175 -6741 7213
rect -1508 7238 -1424 7258
rect -1508 7186 -1492 7238
rect -1440 7186 -1424 7238
rect -1508 7175 -1424 7186
rect -6765 7174 -1424 7175
rect -6765 7122 -1492 7174
rect -1440 7122 -1424 7174
rect -6765 7110 -1424 7122
rect -6765 7066 -1492 7110
rect -6765 7033 -6741 7066
rect -7224 7003 -6741 7033
rect -1508 7058 -1492 7066
rect -1440 7058 -1424 7110
rect -1508 7046 -1424 7058
rect -1508 6994 -1492 7046
rect -1440 6994 -1424 7046
rect -1508 6974 -1424 6994
rect -25531 6660 -25436 6669
rect -25531 6608 -25510 6660
rect -25458 6608 -25436 6660
rect -25531 6596 -25436 6608
rect -25531 6544 -25510 6596
rect -25458 6544 -25436 6596
rect -25531 6532 -25436 6544
rect -25531 6480 -25510 6532
rect -25458 6480 -25436 6532
rect -25531 6468 -25436 6480
rect -25531 6416 -25510 6468
rect -25458 6416 -25436 6468
rect -25531 6408 -25436 6416
rect -4927 6665 -4826 6695
rect -4927 6613 -4903 6665
rect -4851 6613 -4826 6665
rect -4927 6601 -4826 6613
rect -4927 6549 -4903 6601
rect -4851 6549 -4826 6601
rect -4927 6537 -4826 6549
rect -4927 6485 -4903 6537
rect -4851 6485 -4826 6537
rect -4927 6473 -4826 6485
rect -4927 6421 -4903 6473
rect -4851 6421 -4826 6473
rect -4927 6392 -4826 6421
rect -3114 6445 -1424 6451
rect -3114 6393 -1492 6445
rect -1440 6393 -1424 6445
rect -3114 6387 -1424 6393
rect -31140 6331 -26744 6337
rect -31140 6215 -31124 6331
rect -31008 6215 -26744 6331
rect -25374 6303 -18149 6336
rect -25603 6297 -18149 6303
rect -25603 6245 -18245 6297
rect -18193 6245 -18149 6297
rect -13085 6307 -6261 6313
rect -13085 6255 -13069 6307
rect -13017 6255 -6559 6307
rect -6507 6255 -6261 6307
rect -4806 6258 -3415 6310
rect -3363 6258 -3353 6310
rect -13085 6249 -6261 6255
rect -25603 6239 -18149 6245
rect -31140 6209 -26744 6215
rect -25374 6208 -18149 6239
rect -25532 6173 -25437 6174
rect -25532 6121 -25511 6173
rect -25459 6121 -25437 6173
rect -25532 6109 -25437 6121
rect -25532 6057 -25511 6109
rect -25459 6057 -25437 6109
rect -25532 6045 -25437 6057
rect -25532 5993 -25511 6045
rect -25459 5993 -25437 6045
rect -25532 5981 -25437 5993
rect -25532 5929 -25511 5981
rect -25459 5929 -25437 5981
rect -4917 6146 -4831 6163
rect -3114 6161 -3050 6387
rect -4917 6094 -4900 6146
rect -4848 6094 -4831 6146
rect -4917 6082 -4831 6094
rect -4917 6030 -4900 6082
rect -4848 6030 -4831 6082
rect -4917 6018 -4831 6030
rect -4917 5966 -4900 6018
rect -4848 5966 -4831 6018
rect -4917 5950 -4831 5966
rect -3425 5671 -3415 5723
rect -3363 5671 -2970 5723
rect -1832 5671 -678 5723
rect -626 5671 -616 5723
rect -3203 5558 -3069 5577
rect -3203 5506 -3178 5558
rect -3126 5506 -3069 5558
rect -3203 5494 -3069 5506
rect -3203 5442 -3178 5494
rect -3126 5442 -3069 5494
rect -3203 5430 -3069 5442
rect -3203 5378 -3178 5430
rect -3126 5378 -3069 5430
rect -3203 5366 -3069 5378
rect -3203 5314 -3178 5366
rect -3126 5314 -3069 5366
rect -3203 5296 -3069 5314
rect -1149 5129 899 5130
rect -1159 5077 -1149 5129
rect -1097 5077 899 5129
rect -3437 5041 -3353 5047
rect -3437 4989 -3421 5041
rect -3369 4989 -3353 5041
rect -3437 4983 -3353 4989
rect -3427 4973 -3363 4983
rect 23208 4916 23261 7792
rect 24544 6312 24608 9360
rect 35014 8277 35098 8283
rect 35014 8225 35030 8277
rect 35082 8225 35098 8277
rect 35014 8219 35098 8225
rect 40090 8117 40191 8121
rect 40090 8065 40114 8117
rect 40166 8065 40191 8117
rect 40090 8053 40191 8065
rect 38565 8023 38655 8038
rect 38565 7971 38584 8023
rect 38636 7971 38655 8023
rect 38565 7959 38655 7971
rect 38565 7907 38584 7959
rect 38636 7907 38655 7959
rect 40090 8001 40114 8053
rect 40166 8001 40191 8053
rect 40090 7989 40191 8001
rect 40090 7937 40114 7989
rect 40166 7937 40191 7989
rect 40090 7933 40191 7937
rect 38565 7892 38655 7907
rect 36291 7873 36542 7881
rect 36291 7821 36326 7873
rect 36378 7821 36390 7873
rect 36442 7821 36454 7873
rect 36506 7821 36542 7873
rect 36291 7814 36542 7821
rect 33736 7645 33820 7651
rect 33736 7593 33752 7645
rect 33804 7593 33820 7645
rect 33736 7587 33820 7593
rect 40077 7572 40178 7576
rect 38558 7559 38659 7563
rect 38558 7507 38582 7559
rect 38634 7507 38659 7559
rect 38558 7495 38659 7507
rect 38558 7443 38582 7495
rect 38634 7443 38659 7495
rect 38558 7431 38659 7443
rect 38558 7379 38582 7431
rect 38634 7379 38659 7431
rect 40077 7520 40101 7572
rect 40153 7520 40178 7572
rect 40077 7508 40178 7520
rect 40077 7456 40101 7508
rect 40153 7456 40178 7508
rect 40077 7444 40178 7456
rect 40077 7392 40101 7444
rect 40153 7392 40178 7444
rect 40077 7388 40178 7392
rect 38558 7375 38659 7379
rect 36352 7332 36541 7337
rect 36352 7280 36388 7332
rect 36440 7280 36452 7332
rect 36504 7280 36541 7332
rect 36352 7275 36541 7280
rect 35018 7217 35102 7223
rect 35018 7165 35034 7217
rect 35086 7165 35102 7217
rect 35018 7159 35102 7165
rect 42592 7213 45933 7232
rect 42592 7161 42604 7213
rect 42656 7161 42668 7213
rect 42720 7161 42732 7213
rect 42784 7161 42796 7213
rect 42848 7161 42860 7213
rect 42912 7161 42924 7213
rect 42976 7161 42988 7213
rect 43040 7161 43052 7213
rect 43104 7161 43116 7213
rect 43168 7161 43180 7213
rect 43232 7161 43244 7213
rect 43296 7161 43308 7213
rect 43360 7161 43372 7213
rect 43424 7161 43436 7213
rect 43488 7161 43500 7213
rect 43552 7161 43564 7213
rect 43616 7161 43628 7213
rect 43680 7161 43692 7213
rect 43744 7161 43756 7213
rect 43808 7161 43820 7213
rect 43872 7161 43884 7213
rect 43936 7161 43948 7213
rect 44000 7161 44012 7213
rect 44064 7161 44076 7213
rect 44128 7161 44140 7213
rect 44192 7161 44204 7213
rect 44256 7161 44268 7213
rect 44320 7161 44332 7213
rect 44384 7161 44396 7213
rect 44448 7161 44460 7213
rect 44512 7161 44524 7213
rect 44576 7161 44588 7213
rect 44640 7161 44652 7213
rect 44704 7161 44716 7213
rect 44768 7161 44780 7213
rect 44832 7161 44844 7213
rect 44896 7161 44908 7213
rect 44960 7161 44972 7213
rect 45024 7161 45036 7213
rect 45088 7161 45100 7213
rect 45152 7161 45164 7213
rect 45216 7161 45228 7213
rect 45280 7161 45292 7213
rect 45344 7161 45356 7213
rect 45408 7161 45420 7213
rect 45472 7161 45484 7213
rect 45536 7161 45548 7213
rect 45600 7161 45612 7213
rect 45664 7161 45676 7213
rect 45728 7161 45740 7213
rect 45792 7161 45804 7213
rect 45856 7161 45868 7213
rect 45920 7161 45933 7213
rect 42592 7143 45933 7161
rect 35017 6948 35101 6954
rect 35017 6896 35033 6948
rect 35085 6896 35101 6948
rect 35017 6890 35101 6896
rect 36342 6784 36447 6795
rect 36342 6732 36368 6784
rect 36420 6732 36447 6784
rect 36342 6721 36447 6732
rect 40082 6781 40183 6785
rect 40082 6729 40106 6781
rect 40158 6729 40183 6781
rect 40082 6717 40183 6729
rect 38561 6702 38659 6707
rect 38561 6650 38584 6702
rect 38636 6650 38659 6702
rect 38561 6638 38659 6650
rect 38561 6586 38584 6638
rect 38636 6586 38659 6638
rect 40082 6665 40106 6717
rect 40158 6665 40183 6717
rect 40082 6653 40183 6665
rect 40082 6601 40106 6653
rect 40158 6601 40183 6653
rect 40082 6597 40183 6601
rect 38561 6582 38659 6586
rect 24534 6306 24618 6312
rect 24534 6254 24550 6306
rect 24602 6254 24618 6306
rect 24534 6248 24618 6254
rect 33724 6306 33808 6312
rect 33724 6254 33740 6306
rect 33792 6254 33808 6306
rect 33724 6248 33808 6254
rect 35757 6243 37077 6265
rect 35757 6191 36993 6243
rect 37045 6191 37077 6243
rect 35757 6169 37077 6191
rect 38553 6228 38654 6232
rect 38553 6176 38577 6228
rect 38629 6176 38654 6228
rect 38553 6164 38654 6176
rect 38553 6112 38577 6164
rect 38629 6112 38654 6164
rect 38553 6100 38654 6112
rect 38553 6048 38577 6100
rect 38629 6048 38654 6100
rect 38553 6044 38654 6048
rect 40082 6225 40183 6229
rect 40082 6173 40106 6225
rect 40158 6173 40183 6225
rect 40082 6161 40183 6173
rect 40082 6109 40106 6161
rect 40158 6109 40183 6161
rect 40082 6097 40183 6109
rect 40082 6045 40106 6097
rect 40158 6045 40183 6097
rect 40082 6041 40183 6045
rect 35017 5879 35101 5885
rect 35017 5827 35033 5879
rect 35085 5827 35101 5879
rect 35017 5821 35101 5827
rect 47463 5772 47719 5800
rect 47463 5744 47501 5772
rect 35960 5701 36159 5707
rect 35960 5649 36001 5701
rect 36053 5649 36065 5701
rect 36117 5649 36159 5701
rect 35960 5644 36159 5649
rect 40356 5616 47501 5744
rect 47463 5592 47501 5616
rect 47681 5592 47719 5772
rect 47463 5564 47719 5592
rect 35014 5556 35098 5562
rect 35014 5504 35030 5556
rect 35082 5504 35098 5556
rect 35014 5498 35098 5504
rect 40099 5401 40200 5405
rect 40099 5349 40123 5401
rect 40175 5349 40200 5401
rect 40099 5337 40200 5349
rect 38564 5312 38658 5322
rect 38564 5260 38585 5312
rect 38637 5260 38658 5312
rect 38564 5248 38658 5260
rect 38564 5196 38585 5248
rect 38637 5196 38658 5248
rect 40099 5285 40123 5337
rect 40175 5285 40200 5337
rect 40099 5273 40200 5285
rect 40099 5221 40123 5273
rect 40175 5221 40200 5273
rect 40099 5217 40200 5221
rect 38564 5187 38658 5196
rect 36504 5153 36744 5162
rect 36504 5101 36534 5153
rect 36586 5101 36598 5153
rect 36650 5101 36662 5153
rect 36714 5101 36744 5153
rect 36504 5092 36744 5101
rect 23198 4915 23271 4916
rect 23198 4863 23208 4915
rect 23260 4863 23271 4915
rect 33732 4915 33805 4916
rect 33732 4863 33742 4915
rect 33794 4863 33805 4915
rect 38552 4875 38653 4879
rect 38552 4823 38576 4875
rect 38628 4823 38653 4875
rect 38552 4811 38653 4823
rect 38552 4759 38576 4811
rect 38628 4759 38653 4811
rect 38552 4747 38653 4759
rect 38552 4695 38576 4747
rect 38628 4695 38653 4747
rect 38552 4691 38653 4695
rect 40082 4853 40183 4857
rect 40082 4801 40106 4853
rect 40158 4801 40183 4853
rect 40082 4789 40183 4801
rect 40082 4737 40106 4789
rect 40158 4737 40183 4789
rect 40082 4725 40183 4737
rect 40082 4673 40106 4725
rect 40158 4673 40183 4725
rect 40082 4669 40183 4673
rect 36354 4610 36519 4613
rect 36354 4558 36378 4610
rect 36430 4558 36442 4610
rect 36494 4558 36519 4610
rect 36354 4555 36519 4558
rect 35025 4486 35109 4492
rect 35025 4434 35041 4486
rect 35093 4434 35109 4486
rect 35025 4428 35109 4434
rect -253 3789 867 3790
rect -289 3737 -279 3789
rect -227 3737 867 3789
rect -2121 3298 3361 3416
rect -2121 3180 1661 3298
rect -2121 -6585 -1885 3180
rect 23422 2406 23495 2407
rect 23422 2354 23432 2406
rect 23484 2354 23495 2406
rect 22579 1096 22652 1097
rect 22579 1044 22589 1096
rect 22641 1044 22652 1096
rect 230 292 21384 391
rect 59 207 21384 292
rect 59 183 352 207
rect 312 91 352 183
rect 21076 183 21384 207
rect 21076 91 21117 183
rect 312 67 21117 91
rect 22589 -2017 22642 1044
rect 23432 -640 23485 2354
rect 26001 716 26076 4397
rect 42589 4214 45969 4233
rect 35014 4181 35098 4187
rect 35014 4129 35030 4181
rect 35082 4129 35098 4181
rect 42589 4162 42621 4214
rect 42673 4162 42685 4214
rect 42737 4162 42749 4214
rect 42801 4162 42813 4214
rect 42865 4162 42877 4214
rect 42929 4162 42941 4214
rect 42993 4162 43005 4214
rect 43057 4162 43069 4214
rect 43121 4162 43133 4214
rect 43185 4162 43197 4214
rect 43249 4162 43261 4214
rect 43313 4162 43325 4214
rect 43377 4162 43389 4214
rect 43441 4162 43453 4214
rect 43505 4162 43517 4214
rect 43569 4162 43581 4214
rect 43633 4162 43645 4214
rect 43697 4162 43709 4214
rect 43761 4162 43773 4214
rect 43825 4162 43837 4214
rect 43889 4162 43901 4214
rect 43953 4162 43965 4214
rect 44017 4162 44029 4214
rect 44081 4162 44093 4214
rect 44145 4162 44157 4214
rect 44209 4162 44221 4214
rect 44273 4162 44285 4214
rect 44337 4162 44349 4214
rect 44401 4162 44413 4214
rect 44465 4162 44477 4214
rect 44529 4162 44541 4214
rect 44593 4162 44605 4214
rect 44657 4162 44669 4214
rect 44721 4162 44733 4214
rect 44785 4162 44797 4214
rect 44849 4162 44861 4214
rect 44913 4162 44925 4214
rect 44977 4162 44989 4214
rect 45041 4162 45053 4214
rect 45105 4162 45117 4214
rect 45169 4162 45181 4214
rect 45233 4162 45245 4214
rect 45297 4162 45309 4214
rect 45361 4162 45373 4214
rect 45425 4162 45437 4214
rect 45489 4162 45501 4214
rect 45553 4162 45565 4214
rect 45617 4162 45629 4214
rect 45681 4162 45693 4214
rect 45745 4162 45757 4214
rect 45809 4162 45821 4214
rect 45873 4162 45885 4214
rect 45937 4162 45969 4214
rect 42589 4144 45969 4162
rect 35014 4123 35098 4129
rect 36299 4067 37078 4089
rect 36299 4015 36994 4067
rect 37046 4015 37078 4067
rect 36299 3993 37078 4015
rect 40089 4022 40190 4026
rect 40089 3970 40113 4022
rect 40165 3970 40190 4022
rect 40089 3958 40190 3970
rect 38562 3915 38661 3934
rect 38562 3863 38585 3915
rect 38637 3863 38661 3915
rect 38562 3851 38661 3863
rect 38562 3799 38585 3851
rect 38637 3799 38661 3851
rect 40089 3906 40113 3958
rect 40165 3906 40190 3958
rect 40089 3894 40190 3906
rect 40089 3842 40113 3894
rect 40165 3842 40190 3894
rect 40089 3838 40190 3842
rect 38562 3781 38661 3799
rect 36349 3521 36496 3531
rect 36349 3469 36364 3521
rect 36416 3469 36428 3521
rect 36480 3469 36496 3521
rect 36349 3459 36496 3469
rect 38555 3475 38656 3479
rect 38555 3423 38579 3475
rect 38631 3423 38656 3475
rect 38555 3411 38656 3423
rect 38555 3359 38579 3411
rect 38631 3359 38656 3411
rect 38555 3347 38656 3359
rect 38555 3295 38579 3347
rect 38631 3295 38656 3347
rect 38555 3291 38656 3295
rect 40079 3469 40180 3473
rect 40079 3417 40103 3469
rect 40155 3417 40180 3469
rect 40079 3405 40180 3417
rect 40079 3353 40103 3405
rect 40155 3353 40180 3405
rect 40079 3341 40180 3353
rect 40079 3289 40103 3341
rect 40155 3289 40180 3341
rect 40079 3285 40180 3289
rect 35021 3116 35105 3122
rect 35021 3064 35037 3116
rect 35089 3064 35105 3116
rect 35021 3058 35105 3064
rect 35014 1337 35098 1343
rect 35014 1285 35030 1337
rect 35082 1285 35098 1337
rect 35014 1279 35098 1285
rect 40090 1177 40191 1181
rect 40090 1125 40114 1177
rect 40166 1125 40191 1177
rect 40090 1113 40191 1125
rect 38565 1083 38655 1098
rect 38565 1031 38584 1083
rect 38636 1031 38655 1083
rect 38565 1019 38655 1031
rect 38565 967 38584 1019
rect 38636 967 38655 1019
rect 40090 1061 40114 1113
rect 40166 1061 40191 1113
rect 40090 1049 40191 1061
rect 40090 997 40114 1049
rect 40166 997 40191 1049
rect 40090 993 40191 997
rect 38565 952 38655 967
rect 36291 933 36542 941
rect 36291 881 36326 933
rect 36378 881 36390 933
rect 36442 881 36454 933
rect 36506 881 36542 933
rect 36291 874 36542 881
rect 25991 704 26086 716
rect 25991 652 26012 704
rect 26064 652 26086 704
rect 25991 641 26086 652
rect 33720 711 33815 716
rect 33720 704 33820 711
rect 33720 652 33741 704
rect 33793 652 33820 704
rect 33720 647 33820 652
rect 33720 641 33815 647
rect 40077 632 40178 636
rect 38558 619 38659 623
rect 38558 567 38582 619
rect 38634 567 38659 619
rect 38558 555 38659 567
rect 38558 503 38582 555
rect 38634 503 38659 555
rect 38558 491 38659 503
rect 38558 439 38582 491
rect 38634 439 38659 491
rect 40077 580 40101 632
rect 40153 580 40178 632
rect 40077 568 40178 580
rect 40077 516 40101 568
rect 40153 516 40178 568
rect 40077 504 40178 516
rect 40077 452 40101 504
rect 40153 452 40178 504
rect 40077 448 40178 452
rect 38558 435 38659 439
rect 36352 392 36541 397
rect 36352 340 36388 392
rect 36440 340 36452 392
rect 36504 340 36541 392
rect 36352 335 36541 340
rect 35018 277 35102 283
rect 35018 225 35034 277
rect 35086 225 35102 277
rect 35018 219 35102 225
rect 42589 280 45940 309
rect 42589 228 42606 280
rect 42658 228 42670 280
rect 42722 228 42734 280
rect 42786 228 42798 280
rect 42850 228 42862 280
rect 42914 228 42926 280
rect 42978 228 42990 280
rect 43042 228 43054 280
rect 43106 228 43118 280
rect 43170 228 43182 280
rect 43234 228 43246 280
rect 43298 228 43310 280
rect 43362 228 43374 280
rect 43426 228 43438 280
rect 43490 228 43502 280
rect 43554 228 43566 280
rect 43618 228 43630 280
rect 43682 228 43694 280
rect 43746 228 43758 280
rect 43810 228 43822 280
rect 43874 228 43886 280
rect 43938 228 43950 280
rect 44002 228 44014 280
rect 44066 228 44078 280
rect 44130 228 44142 280
rect 44194 228 44206 280
rect 44258 228 44270 280
rect 44322 228 44334 280
rect 44386 228 44398 280
rect 44450 228 44462 280
rect 44514 228 44526 280
rect 44578 228 44590 280
rect 44642 228 44654 280
rect 44706 228 44718 280
rect 44770 228 44782 280
rect 44834 228 44846 280
rect 44898 228 44910 280
rect 44962 228 44974 280
rect 45026 228 45038 280
rect 45090 228 45102 280
rect 45154 228 45166 280
rect 45218 228 45230 280
rect 45282 228 45294 280
rect 45346 228 45358 280
rect 45410 228 45422 280
rect 45474 228 45486 280
rect 45538 228 45550 280
rect 45602 228 45614 280
rect 45666 228 45678 280
rect 45730 228 45742 280
rect 45794 228 45806 280
rect 45858 228 45870 280
rect 45922 228 45940 280
rect 42589 199 45940 228
rect 35017 8 35101 14
rect 35017 -44 35033 8
rect 35085 -44 35101 8
rect 35017 -50 35101 -44
rect 36342 -156 36447 -145
rect 36342 -208 36368 -156
rect 36420 -208 36447 -156
rect 36342 -219 36447 -208
rect 40082 -159 40183 -155
rect 40082 -211 40106 -159
rect 40158 -211 40183 -159
rect 40082 -223 40183 -211
rect 38561 -238 38659 -233
rect 38561 -290 38584 -238
rect 38636 -290 38659 -238
rect 38561 -302 38659 -290
rect 38561 -354 38584 -302
rect 38636 -354 38659 -302
rect 40082 -275 40106 -223
rect 40158 -275 40183 -223
rect 40082 -287 40183 -275
rect 40082 -339 40106 -287
rect 40158 -339 40183 -287
rect 40082 -343 40183 -339
rect 38561 -358 38659 -354
rect 33724 -635 33808 -628
rect 23422 -641 23495 -640
rect 23422 -693 23432 -641
rect 23484 -693 23495 -641
rect 33724 -687 33741 -635
rect 33793 -687 33808 -635
rect 33724 -692 33808 -687
rect 33731 -693 33804 -692
rect 35757 -697 37077 -675
rect 35757 -749 36993 -697
rect 37045 -749 37077 -697
rect 35757 -771 37077 -749
rect 38553 -712 38654 -708
rect 38553 -764 38577 -712
rect 38629 -764 38654 -712
rect 38553 -776 38654 -764
rect 38553 -828 38577 -776
rect 38629 -828 38654 -776
rect 38553 -840 38654 -828
rect 38553 -892 38577 -840
rect 38629 -892 38654 -840
rect 38553 -896 38654 -892
rect 40082 -715 40183 -711
rect 40082 -767 40106 -715
rect 40158 -767 40183 -715
rect 40082 -779 40183 -767
rect 40082 -831 40106 -779
rect 40158 -831 40183 -779
rect 40082 -843 40183 -831
rect 40082 -895 40106 -843
rect 40158 -895 40183 -843
rect 40082 -899 40183 -895
rect 35017 -1061 35101 -1055
rect 35017 -1113 35033 -1061
rect 35085 -1113 35101 -1061
rect 35017 -1119 35101 -1113
rect 47479 -1168 47735 -1140
rect 47479 -1196 47517 -1168
rect 35960 -1239 36159 -1233
rect 35960 -1291 36001 -1239
rect 36053 -1291 36065 -1239
rect 36117 -1291 36159 -1239
rect 35960 -1296 36159 -1291
rect 40356 -1324 47517 -1196
rect 47479 -1348 47517 -1324
rect 47697 -1348 47735 -1168
rect 47479 -1376 47735 -1348
rect 35014 -1384 35098 -1378
rect 35014 -1436 35030 -1384
rect 35082 -1436 35098 -1384
rect 35014 -1442 35098 -1436
rect 40099 -1539 40200 -1535
rect 40099 -1591 40123 -1539
rect 40175 -1591 40200 -1539
rect 40099 -1603 40200 -1591
rect 38564 -1628 38658 -1618
rect 38564 -1680 38585 -1628
rect 38637 -1680 38658 -1628
rect 38564 -1692 38658 -1680
rect 38564 -1744 38585 -1692
rect 38637 -1744 38658 -1692
rect 40099 -1655 40123 -1603
rect 40175 -1655 40200 -1603
rect 40099 -1667 40200 -1655
rect 40099 -1719 40123 -1667
rect 40175 -1719 40200 -1667
rect 40099 -1723 40200 -1719
rect 38564 -1753 38658 -1744
rect 36504 -1787 36744 -1778
rect 36504 -1839 36534 -1787
rect 36586 -1839 36598 -1787
rect 36650 -1839 36662 -1787
rect 36714 -1839 36744 -1787
rect 36504 -1848 36744 -1839
rect 22579 -2018 22653 -2017
rect 22579 -2070 22590 -2018
rect 22642 -2070 22653 -2018
rect 33736 -2021 33816 -2017
rect 22589 -2073 22642 -2070
rect 33736 -2073 33750 -2021
rect 33802 -2073 33816 -2021
rect 33736 -2077 33816 -2073
rect 38552 -2065 38653 -2061
rect 38552 -2117 38576 -2065
rect 38628 -2117 38653 -2065
rect 38552 -2129 38653 -2117
rect 38552 -2181 38576 -2129
rect 38628 -2181 38653 -2129
rect 38552 -2193 38653 -2181
rect 38552 -2245 38576 -2193
rect 38628 -2245 38653 -2193
rect 38552 -2249 38653 -2245
rect 40082 -2087 40183 -2083
rect 40082 -2139 40106 -2087
rect 40158 -2139 40183 -2087
rect 40082 -2151 40183 -2139
rect 40082 -2203 40106 -2151
rect 40158 -2203 40183 -2151
rect 40082 -2215 40183 -2203
rect 40082 -2267 40106 -2215
rect 40158 -2267 40183 -2215
rect 40082 -2271 40183 -2267
rect 36354 -2330 36519 -2327
rect 36354 -2382 36378 -2330
rect 36430 -2382 36442 -2330
rect 36494 -2382 36519 -2330
rect 36354 -2385 36519 -2382
rect 35025 -2454 35109 -2448
rect 35025 -2506 35041 -2454
rect 35093 -2506 35109 -2454
rect 35025 -2512 35109 -2506
rect 42577 -2726 45943 -2708
rect 35014 -2759 35098 -2753
rect 35014 -2811 35030 -2759
rect 35082 -2811 35098 -2759
rect 42577 -2778 42602 -2726
rect 42654 -2778 42666 -2726
rect 42718 -2778 42730 -2726
rect 42782 -2778 42794 -2726
rect 42846 -2778 42858 -2726
rect 42910 -2778 42922 -2726
rect 42974 -2778 42986 -2726
rect 43038 -2778 43050 -2726
rect 43102 -2778 43114 -2726
rect 43166 -2778 43178 -2726
rect 43230 -2778 43242 -2726
rect 43294 -2778 43306 -2726
rect 43358 -2778 43370 -2726
rect 43422 -2778 43434 -2726
rect 43486 -2778 43498 -2726
rect 43550 -2778 43562 -2726
rect 43614 -2778 43626 -2726
rect 43678 -2778 43690 -2726
rect 43742 -2778 43754 -2726
rect 43806 -2778 43818 -2726
rect 43870 -2778 43882 -2726
rect 43934 -2778 43946 -2726
rect 43998 -2778 44010 -2726
rect 44062 -2778 44074 -2726
rect 44126 -2778 44138 -2726
rect 44190 -2778 44202 -2726
rect 44254 -2778 44266 -2726
rect 44318 -2778 44330 -2726
rect 44382 -2778 44394 -2726
rect 44446 -2778 44458 -2726
rect 44510 -2778 44522 -2726
rect 44574 -2778 44586 -2726
rect 44638 -2778 44650 -2726
rect 44702 -2778 44714 -2726
rect 44766 -2778 44778 -2726
rect 44830 -2778 44842 -2726
rect 44894 -2778 44906 -2726
rect 44958 -2778 44970 -2726
rect 45022 -2778 45034 -2726
rect 45086 -2778 45098 -2726
rect 45150 -2778 45162 -2726
rect 45214 -2778 45226 -2726
rect 45278 -2778 45290 -2726
rect 45342 -2778 45354 -2726
rect 45406 -2778 45418 -2726
rect 45470 -2778 45482 -2726
rect 45534 -2778 45546 -2726
rect 45598 -2778 45610 -2726
rect 45662 -2778 45674 -2726
rect 45726 -2778 45738 -2726
rect 45790 -2778 45802 -2726
rect 45854 -2778 45866 -2726
rect 45918 -2778 45943 -2726
rect 42577 -2796 45943 -2778
rect 35014 -2817 35098 -2811
rect 36299 -2873 37078 -2851
rect 36299 -2925 36994 -2873
rect 37046 -2925 37078 -2873
rect 36299 -2947 37078 -2925
rect 40089 -2918 40190 -2914
rect 40089 -2970 40113 -2918
rect 40165 -2970 40190 -2918
rect 40089 -2982 40190 -2970
rect 38562 -3025 38661 -3006
rect 38562 -3077 38585 -3025
rect 38637 -3077 38661 -3025
rect 38562 -3089 38661 -3077
rect 38562 -3141 38585 -3089
rect 38637 -3141 38661 -3089
rect 40089 -3034 40113 -2982
rect 40165 -3034 40190 -2982
rect 40089 -3046 40190 -3034
rect 40089 -3098 40113 -3046
rect 40165 -3098 40190 -3046
rect 40089 -3102 40190 -3098
rect 38562 -3159 38661 -3141
rect 36349 -3419 36496 -3409
rect 36349 -3471 36364 -3419
rect 36416 -3471 36428 -3419
rect 36480 -3471 36496 -3419
rect 36349 -3481 36496 -3471
rect 38555 -3465 38656 -3461
rect 38555 -3517 38579 -3465
rect 38631 -3517 38656 -3465
rect 38555 -3529 38656 -3517
rect 38555 -3581 38579 -3529
rect 38631 -3581 38656 -3529
rect 38555 -3593 38656 -3581
rect 38555 -3645 38579 -3593
rect 38631 -3645 38656 -3593
rect 38555 -3649 38656 -3645
rect 40079 -3471 40180 -3467
rect 40079 -3523 40103 -3471
rect 40155 -3523 40180 -3471
rect 40079 -3535 40180 -3523
rect 40079 -3587 40103 -3535
rect 40155 -3587 40180 -3535
rect 40079 -3599 40180 -3587
rect 40079 -3651 40103 -3599
rect 40155 -3651 40180 -3599
rect 40079 -3655 40180 -3651
rect 35021 -3824 35105 -3818
rect 35021 -3876 35037 -3824
rect 35089 -3876 35105 -3824
rect 35021 -3882 35105 -3876
rect -2121 -6799 -1993 -6585
rect -3605 -6850 -3493 -6822
rect -3605 -6902 -3575 -6850
rect -3523 -6902 -3493 -6850
rect -3605 -6914 -3493 -6902
rect -3605 -6966 -3575 -6914
rect -3523 -6966 -3493 -6914
rect -3605 -6978 -3493 -6966
rect -3605 -7030 -3575 -6978
rect -3523 -7030 -3493 -6978
rect -3605 -7042 -3493 -7030
rect -3605 -7094 -3575 -7042
rect -3523 -7094 -3493 -7042
rect -3605 -7106 -3493 -7094
rect -3605 -7158 -3575 -7106
rect -3523 -7158 -3493 -7106
rect -3605 -7170 -3493 -7158
rect -3605 -7222 -3575 -7170
rect -3523 -7222 -3493 -7170
rect -3605 -7234 -3493 -7222
rect -3605 -7286 -3575 -7234
rect -3523 -7286 -3493 -7234
rect -3605 -7298 -3493 -7286
rect -3605 -7350 -3575 -7298
rect -3523 -7350 -3493 -7298
rect -3605 -7362 -3493 -7350
rect -3605 -7414 -3575 -7362
rect -3523 -7414 -3493 -7362
rect -3605 -7426 -3493 -7414
rect -3605 -7478 -3575 -7426
rect -3523 -7478 -3493 -7426
rect -3605 -7490 -3493 -7478
rect -3605 -7542 -3575 -7490
rect -3523 -7542 -3493 -7490
rect -3605 -7554 -3493 -7542
rect -3605 -7606 -3575 -7554
rect -3523 -7606 -3493 -7554
rect -3605 -7618 -3493 -7606
rect -3605 -7670 -3575 -7618
rect -3523 -7670 -3493 -7618
rect -3605 -7682 -3493 -7670
rect -3605 -7734 -3575 -7682
rect -3523 -7734 -3493 -7682
rect -3605 -7746 -3493 -7734
rect -3605 -7798 -3575 -7746
rect -3523 -7798 -3493 -7746
rect -3605 -7810 -3493 -7798
rect -3605 -7862 -3575 -7810
rect -3523 -7862 -3493 -7810
rect -3605 -7874 -3493 -7862
rect -3605 -7926 -3575 -7874
rect -3523 -7926 -3493 -7874
rect -3605 -7938 -3493 -7926
rect -3605 -7990 -3575 -7938
rect -3523 -7990 -3493 -7938
rect -3605 -8002 -3493 -7990
rect -3605 -8054 -3575 -8002
rect -3523 -8054 -3493 -8002
rect -3605 -8066 -3493 -8054
rect -3605 -8118 -3575 -8066
rect -3523 -8118 -3493 -8066
rect -3605 -8130 -3493 -8118
rect -3605 -8182 -3575 -8130
rect -3523 -8182 -3493 -8130
rect -3605 -8194 -3493 -8182
rect -3605 -8246 -3575 -8194
rect -3523 -8246 -3493 -8194
rect -3605 -8258 -3493 -8246
rect -3605 -8310 -3575 -8258
rect -3523 -8310 -3493 -8258
rect -3605 -8322 -3493 -8310
rect -3605 -8374 -3575 -8322
rect -3523 -8374 -3493 -8322
rect -3605 -8386 -3493 -8374
rect -3605 -8438 -3575 -8386
rect -3523 -8438 -3493 -8386
rect -3605 -8450 -3493 -8438
rect -3605 -8502 -3575 -8450
rect -3523 -8502 -3493 -8450
rect -3605 -8514 -3493 -8502
rect -3605 -8566 -3575 -8514
rect -3523 -8566 -3493 -8514
rect -3605 -8578 -3493 -8566
rect -3605 -8630 -3575 -8578
rect -3523 -8630 -3493 -8578
rect -3605 -8642 -3493 -8630
rect -3605 -8694 -3575 -8642
rect -3523 -8694 -3493 -8642
rect -3605 -8706 -3493 -8694
rect -3605 -8758 -3575 -8706
rect -3523 -8758 -3493 -8706
rect -3605 -8770 -3493 -8758
rect -3605 -8822 -3575 -8770
rect -3523 -8822 -3493 -8770
rect -3605 -8834 -3493 -8822
rect -3605 -8886 -3575 -8834
rect -3523 -8886 -3493 -8834
rect -3605 -8898 -3493 -8886
rect -3605 -8950 -3575 -8898
rect -3523 -8950 -3493 -8898
rect -3605 -8962 -3493 -8950
rect -3605 -9014 -3575 -8962
rect -3523 -9014 -3493 -8962
rect -3605 -9026 -3493 -9014
rect -3605 -9078 -3575 -9026
rect -3523 -9078 -3493 -9026
rect -3605 -9090 -3493 -9078
rect -3605 -9142 -3575 -9090
rect -3523 -9142 -3493 -9090
rect -3605 -9154 -3493 -9142
rect -3605 -9206 -3575 -9154
rect -3523 -9206 -3493 -9154
rect -3605 -9218 -3493 -9206
rect -3605 -9270 -3575 -9218
rect -3523 -9270 -3493 -9218
rect -3605 -9282 -3493 -9270
rect -3605 -9334 -3575 -9282
rect -3523 -9334 -3493 -9282
rect -3605 -9346 -3493 -9334
rect -3605 -9398 -3575 -9346
rect -3523 -9398 -3493 -9346
rect -3605 -9410 -3493 -9398
rect -3605 -9462 -3575 -9410
rect -3523 -9462 -3493 -9410
rect -3605 -9474 -3493 -9462
rect -3605 -9526 -3575 -9474
rect -3523 -9526 -3493 -9474
rect -3605 -9538 -3493 -9526
rect -3605 -9590 -3575 -9538
rect -3523 -9590 -3493 -9538
rect -3605 -9602 -3493 -9590
rect -3605 -9654 -3575 -9602
rect -3523 -9654 -3493 -9602
rect -3605 -9666 -3493 -9654
rect -3605 -9718 -3575 -9666
rect -3523 -9718 -3493 -9666
rect -3605 -9730 -3493 -9718
rect -3605 -9782 -3575 -9730
rect -3523 -9782 -3493 -9730
rect -3605 -9794 -3493 -9782
rect -3605 -9846 -3575 -9794
rect -3523 -9846 -3493 -9794
rect -3605 -9858 -3493 -9846
rect -3605 -9910 -3575 -9858
rect -3523 -9910 -3493 -9858
rect -3605 -9922 -3493 -9910
rect -3605 -9974 -3575 -9922
rect -3523 -9974 -3493 -9922
rect -3605 -9986 -3493 -9974
rect -3605 -10038 -3575 -9986
rect -3523 -10038 -3493 -9986
rect -3605 -10050 -3493 -10038
rect -3605 -10102 -3575 -10050
rect -3523 -10102 -3493 -10050
rect -3605 -10130 -3493 -10102
rect -2121 -10365 -2003 -6799
rect -610 -6857 -476 -6825
rect -610 -6909 -569 -6857
rect -517 -6909 -476 -6857
rect -610 -6921 -476 -6909
rect -610 -6973 -569 -6921
rect -517 -6973 -476 -6921
rect -610 -6985 -476 -6973
rect -610 -7037 -569 -6985
rect -517 -7037 -476 -6985
rect -610 -7049 -476 -7037
rect -610 -7101 -569 -7049
rect -517 -7101 -476 -7049
rect -610 -7113 -476 -7101
rect -610 -7165 -569 -7113
rect -517 -7165 -476 -7113
rect -610 -7177 -476 -7165
rect -610 -7229 -569 -7177
rect -517 -7229 -476 -7177
rect -610 -7241 -476 -7229
rect -610 -7293 -569 -7241
rect -517 -7293 -476 -7241
rect -610 -7305 -476 -7293
rect -610 -7357 -569 -7305
rect -517 -7357 -476 -7305
rect -610 -7369 -476 -7357
rect -610 -7421 -569 -7369
rect -517 -7421 -476 -7369
rect -610 -7433 -476 -7421
rect -610 -7485 -569 -7433
rect -517 -7485 -476 -7433
rect -610 -7497 -476 -7485
rect -610 -7549 -569 -7497
rect -517 -7549 -476 -7497
rect -610 -7561 -476 -7549
rect -610 -7613 -569 -7561
rect -517 -7613 -476 -7561
rect -610 -7625 -476 -7613
rect -610 -7677 -569 -7625
rect -517 -7677 -476 -7625
rect -610 -7689 -476 -7677
rect -610 -7741 -569 -7689
rect -517 -7741 -476 -7689
rect -610 -7753 -476 -7741
rect -610 -7805 -569 -7753
rect -517 -7805 -476 -7753
rect -610 -7817 -476 -7805
rect -610 -7869 -569 -7817
rect -517 -7869 -476 -7817
rect -610 -7881 -476 -7869
rect -610 -7933 -569 -7881
rect -517 -7933 -476 -7881
rect -610 -7945 -476 -7933
rect -610 -7997 -569 -7945
rect -517 -7997 -476 -7945
rect -610 -8009 -476 -7997
rect -610 -8061 -569 -8009
rect -517 -8061 -476 -8009
rect -610 -8073 -476 -8061
rect -610 -8125 -569 -8073
rect -517 -8125 -476 -8073
rect -610 -8137 -476 -8125
rect -610 -8189 -569 -8137
rect -517 -8189 -476 -8137
rect -610 -8201 -476 -8189
rect -610 -8253 -569 -8201
rect -517 -8253 -476 -8201
rect -610 -8265 -476 -8253
rect -610 -8317 -569 -8265
rect -517 -8317 -476 -8265
rect -610 -8329 -476 -8317
rect -610 -8381 -569 -8329
rect -517 -8381 -476 -8329
rect -610 -8393 -476 -8381
rect -610 -8445 -569 -8393
rect -517 -8445 -476 -8393
rect -610 -8457 -476 -8445
rect -610 -8509 -569 -8457
rect -517 -8509 -476 -8457
rect -610 -8521 -476 -8509
rect -610 -8573 -569 -8521
rect -517 -8573 -476 -8521
rect -610 -8585 -476 -8573
rect -610 -8637 -569 -8585
rect -517 -8637 -476 -8585
rect -610 -8649 -476 -8637
rect -610 -8701 -569 -8649
rect -517 -8701 -476 -8649
rect -610 -8713 -476 -8701
rect -610 -8765 -569 -8713
rect -517 -8765 -476 -8713
rect -610 -8777 -476 -8765
rect -610 -8829 -569 -8777
rect -517 -8829 -476 -8777
rect -610 -8841 -476 -8829
rect -610 -8893 -569 -8841
rect -517 -8893 -476 -8841
rect -610 -8905 -476 -8893
rect -610 -8957 -569 -8905
rect -517 -8957 -476 -8905
rect -610 -8969 -476 -8957
rect -610 -9021 -569 -8969
rect -517 -9021 -476 -8969
rect -610 -9033 -476 -9021
rect -610 -9085 -569 -9033
rect -517 -9085 -476 -9033
rect -610 -9097 -476 -9085
rect -610 -9149 -569 -9097
rect -517 -9149 -476 -9097
rect -610 -9161 -476 -9149
rect -610 -9213 -569 -9161
rect -517 -9213 -476 -9161
rect -610 -9225 -476 -9213
rect -610 -9277 -569 -9225
rect -517 -9277 -476 -9225
rect -610 -9289 -476 -9277
rect -610 -9341 -569 -9289
rect -517 -9341 -476 -9289
rect -610 -9353 -476 -9341
rect -610 -9405 -569 -9353
rect -517 -9405 -476 -9353
rect -610 -9417 -476 -9405
rect -610 -9469 -569 -9417
rect -517 -9469 -476 -9417
rect -610 -9481 -476 -9469
rect -610 -9533 -569 -9481
rect -517 -9533 -476 -9481
rect -610 -9545 -476 -9533
rect -610 -9597 -569 -9545
rect -517 -9597 -476 -9545
rect -610 -9609 -476 -9597
rect -610 -9661 -569 -9609
rect -517 -9661 -476 -9609
rect -610 -9673 -476 -9661
rect -610 -9725 -569 -9673
rect -517 -9725 -476 -9673
rect -610 -9737 -476 -9725
rect -610 -9789 -569 -9737
rect -517 -9789 -476 -9737
rect -610 -9801 -476 -9789
rect -610 -9853 -569 -9801
rect -517 -9853 -476 -9801
rect -610 -9865 -476 -9853
rect -610 -9917 -569 -9865
rect -517 -9917 -476 -9865
rect -610 -9929 -476 -9917
rect -610 -9981 -569 -9929
rect -517 -9981 -476 -9929
rect -610 -9993 -476 -9981
rect -610 -10045 -569 -9993
rect -517 -10045 -476 -9993
rect -610 -10057 -476 -10045
rect -610 -10109 -569 -10057
rect -517 -10109 -476 -10057
rect -610 -10140 -476 -10109
rect -2179 -12082 -1943 -10365
rect -2189 -12110 -1933 -12082
rect -2189 -12290 -2151 -12110
rect -1971 -12290 -1933 -12110
rect -2189 -12318 -1933 -12290
<< via1 >>
rect -15382 77932 -15202 78112
rect -16825 76666 -16773 76718
rect -16825 76602 -16773 76654
rect -16825 76538 -16773 76590
rect -16825 76474 -16773 76526
rect -16825 76410 -16773 76462
rect -16825 76346 -16773 76398
rect -16825 76282 -16773 76334
rect -16825 76218 -16773 76270
rect -16825 76154 -16773 76206
rect -16825 76090 -16773 76142
rect -16825 76026 -16773 76078
rect -16825 75962 -16773 76014
rect -16825 75898 -16773 75950
rect -16825 75834 -16773 75886
rect -16825 75770 -16773 75822
rect -16825 75706 -16773 75758
rect -16825 75642 -16773 75694
rect -16825 75578 -16773 75630
rect -16825 75514 -16773 75566
rect -16825 75450 -16773 75502
rect -16825 75386 -16773 75438
rect -16825 75322 -16773 75374
rect -16825 75258 -16773 75310
rect 12634 77903 12814 78083
rect 24684 77904 24864 78084
rect -13824 76672 -13772 76724
rect -13824 76608 -13772 76660
rect -13824 76544 -13772 76596
rect -13824 76480 -13772 76532
rect -13824 76416 -13772 76468
rect -13824 76352 -13772 76404
rect -13824 76288 -13772 76340
rect -13824 76224 -13772 76276
rect -13824 76160 -13772 76212
rect -13824 76096 -13772 76148
rect -13824 76032 -13772 76084
rect -13824 75968 -13772 76020
rect -13824 75904 -13772 75956
rect -13824 75840 -13772 75892
rect -13824 75776 -13772 75828
rect -13824 75712 -13772 75764
rect -13824 75648 -13772 75700
rect -13824 75584 -13772 75636
rect -13824 75520 -13772 75572
rect -13824 75456 -13772 75508
rect -13824 75392 -13772 75444
rect -13824 75328 -13772 75380
rect -13824 75264 -13772 75316
rect -16825 75194 -16773 75246
rect -16825 75130 -16773 75182
rect -16825 75066 -16773 75118
rect -16825 75002 -16773 75054
rect -16825 74938 -16773 74990
rect -16825 74874 -16773 74926
rect -16825 74810 -16773 74862
rect -13824 75200 -13772 75252
rect -13824 75136 -13772 75188
rect -13824 75072 -13772 75124
rect -13824 75008 -13772 75060
rect -13824 74944 -13772 74996
rect -13824 74880 -13772 74932
rect -13824 74816 -13772 74868
rect -16825 74746 -16773 74798
rect -16825 74682 -16773 74734
rect -16825 74618 -16773 74670
rect -16825 74554 -16773 74606
rect -16825 74490 -16773 74542
rect -16825 74426 -16773 74478
rect -16825 74362 -16773 74414
rect -16825 74298 -16773 74350
rect -16825 74234 -16773 74286
rect -16825 74170 -16773 74222
rect -16825 74106 -16773 74158
rect -16825 74042 -16773 74094
rect -16825 73978 -16773 74030
rect -16825 73914 -16773 73966
rect -16825 73850 -16773 73902
rect -16825 73786 -16773 73838
rect -16825 73722 -16773 73774
rect -16825 73658 -16773 73710
rect -16825 73594 -16773 73646
rect -16825 73530 -16773 73582
rect -16825 73466 -16773 73518
rect -16825 73402 -16773 73454
rect -13824 74752 -13772 74804
rect -13824 74688 -13772 74740
rect -13824 74624 -13772 74676
rect -13824 74560 -13772 74612
rect -13824 74496 -13772 74548
rect -13824 74432 -13772 74484
rect -13824 74368 -13772 74420
rect -13824 74304 -13772 74356
rect -13824 74240 -13772 74292
rect -13824 74176 -13772 74228
rect -13824 74112 -13772 74164
rect -13824 74048 -13772 74100
rect -13824 73984 -13772 74036
rect -13824 73920 -13772 73972
rect -13824 73856 -13772 73908
rect -13824 73792 -13772 73844
rect -13824 73728 -13772 73780
rect -13824 73664 -13772 73716
rect -13824 73600 -13772 73652
rect -13824 73536 -13772 73588
rect -13824 73472 -13772 73524
rect -13824 73408 -13772 73460
rect 11149 76664 11265 76720
rect 11149 76630 11189 76664
rect 11189 76630 11223 76664
rect 11223 76630 11265 76664
rect 11149 76592 11265 76630
rect 11149 76558 11189 76592
rect 11189 76558 11223 76592
rect 11223 76558 11265 76592
rect 11149 76520 11265 76558
rect 11149 76486 11189 76520
rect 11189 76486 11223 76520
rect 11223 76486 11265 76520
rect 11149 76448 11265 76486
rect 11149 76414 11189 76448
rect 11189 76414 11223 76448
rect 11223 76414 11265 76448
rect 11149 76376 11265 76414
rect 11149 76342 11189 76376
rect 11189 76342 11223 76376
rect 11223 76342 11265 76376
rect 11149 76304 11265 76342
rect 11149 76270 11189 76304
rect 11189 76270 11223 76304
rect 11223 76270 11265 76304
rect 11149 76232 11265 76270
rect 11149 76198 11189 76232
rect 11189 76198 11223 76232
rect 11223 76198 11265 76232
rect 11149 76160 11265 76198
rect 11149 76126 11189 76160
rect 11189 76126 11223 76160
rect 11223 76126 11265 76160
rect 11149 76088 11265 76126
rect 11149 76054 11189 76088
rect 11189 76054 11223 76088
rect 11223 76054 11265 76088
rect 11149 76016 11265 76054
rect 11149 75982 11189 76016
rect 11189 75982 11223 76016
rect 11223 75982 11265 76016
rect 11149 75944 11265 75982
rect 11149 75910 11189 75944
rect 11189 75910 11223 75944
rect 11223 75910 11265 75944
rect 11149 75872 11265 75910
rect 11149 75838 11189 75872
rect 11189 75838 11223 75872
rect 11223 75838 11265 75872
rect 11149 75800 11265 75838
rect 11149 75766 11189 75800
rect 11189 75766 11223 75800
rect 11223 75766 11265 75800
rect 11149 75728 11265 75766
rect 11149 75694 11189 75728
rect 11189 75694 11223 75728
rect 11223 75694 11265 75728
rect 11149 75656 11265 75694
rect 11149 75622 11189 75656
rect 11189 75622 11223 75656
rect 11223 75622 11265 75656
rect 11149 75584 11265 75622
rect 11149 75550 11189 75584
rect 11189 75550 11223 75584
rect 11223 75550 11265 75584
rect 11149 75512 11265 75550
rect 11149 75478 11189 75512
rect 11189 75478 11223 75512
rect 11223 75478 11265 75512
rect 11149 75440 11265 75478
rect 11149 75406 11189 75440
rect 11189 75406 11223 75440
rect 11223 75406 11265 75440
rect 11149 75368 11265 75406
rect 11149 75334 11189 75368
rect 11189 75334 11223 75368
rect 11223 75334 11265 75368
rect 11149 75296 11265 75334
rect 11149 75262 11189 75296
rect 11189 75262 11223 75296
rect 11223 75262 11265 75296
rect 11149 75224 11265 75262
rect 11149 75190 11189 75224
rect 11189 75190 11223 75224
rect 11223 75190 11265 75224
rect 11149 75152 11265 75190
rect 11149 75118 11189 75152
rect 11189 75118 11223 75152
rect 11223 75118 11265 75152
rect 11149 75080 11265 75118
rect 11149 75046 11189 75080
rect 11189 75046 11223 75080
rect 11223 75046 11265 75080
rect 11149 75008 11265 75046
rect 11149 74974 11189 75008
rect 11189 74974 11223 75008
rect 11223 74974 11265 75008
rect 11149 74936 11265 74974
rect 11149 74902 11189 74936
rect 11189 74902 11223 74936
rect 11223 74902 11265 74936
rect 11149 74864 11265 74902
rect 11149 74830 11189 74864
rect 11189 74830 11223 74864
rect 11223 74830 11265 74864
rect 11149 74792 11265 74830
rect 11149 74758 11189 74792
rect 11189 74758 11223 74792
rect 11223 74758 11265 74792
rect 11149 74720 11265 74758
rect 11149 74686 11189 74720
rect 11189 74686 11223 74720
rect 11223 74686 11265 74720
rect 11149 74648 11265 74686
rect 11149 74614 11189 74648
rect 11189 74614 11223 74648
rect 11223 74614 11265 74648
rect 11149 74576 11265 74614
rect 11149 74542 11189 74576
rect 11189 74542 11223 74576
rect 11223 74542 11265 74576
rect 11149 74504 11265 74542
rect 11149 74470 11189 74504
rect 11189 74470 11223 74504
rect 11223 74470 11265 74504
rect 11149 74432 11265 74470
rect 11149 74398 11189 74432
rect 11189 74398 11223 74432
rect 11223 74398 11265 74432
rect 11149 74360 11265 74398
rect 11149 74326 11189 74360
rect 11189 74326 11223 74360
rect 11223 74326 11265 74360
rect 11149 74288 11265 74326
rect 11149 74254 11189 74288
rect 11189 74254 11223 74288
rect 11223 74254 11265 74288
rect 11149 74216 11265 74254
rect 11149 74182 11189 74216
rect 11189 74182 11223 74216
rect 11223 74182 11265 74216
rect 11149 74144 11265 74182
rect 11149 74110 11189 74144
rect 11189 74110 11223 74144
rect 11223 74110 11265 74144
rect 11149 74072 11265 74110
rect 11149 74038 11189 74072
rect 11189 74038 11223 74072
rect 11223 74038 11265 74072
rect 11149 74000 11265 74038
rect 11149 73966 11189 74000
rect 11189 73966 11223 74000
rect 11223 73966 11265 74000
rect 11149 73928 11265 73966
rect 11149 73894 11189 73928
rect 11189 73894 11223 73928
rect 11223 73894 11265 73928
rect 11149 73856 11265 73894
rect 11149 73822 11189 73856
rect 11189 73822 11223 73856
rect 11223 73822 11265 73856
rect 11149 73784 11265 73822
rect 11149 73750 11189 73784
rect 11189 73750 11223 73784
rect 11223 73750 11265 73784
rect 11149 73712 11265 73750
rect 11149 73678 11189 73712
rect 11189 73678 11223 73712
rect 11223 73678 11265 73712
rect 11149 73640 11265 73678
rect 11149 73606 11189 73640
rect 11189 73606 11223 73640
rect 11223 73606 11265 73640
rect 11149 73568 11265 73606
rect 11149 73534 11189 73568
rect 11189 73534 11223 73568
rect 11223 73534 11265 73568
rect 11149 73496 11265 73534
rect 11149 73462 11189 73496
rect 11189 73462 11223 73496
rect 11223 73462 11265 73496
rect 11149 73404 11265 73462
rect 14150 73417 14266 76733
rect -16658 71744 -16606 71796
rect -15480 71740 -15428 71792
rect -15263 71747 -15211 71799
rect -14129 71744 -14077 71796
rect -16548 70240 -16496 70292
rect -15434 70226 -15382 70278
rect -15221 70227 -15169 70279
rect -14057 70227 -14005 70279
rect -15416 68442 -15364 68494
rect -15416 68378 -15364 68430
rect -15416 68314 -15364 68366
rect -15953 68189 -15901 68241
rect -15953 68125 -15901 68177
rect -15416 68250 -15364 68302
rect -15416 68186 -15364 68238
rect -14869 68192 -14817 68244
rect -14869 68128 -14817 68180
rect -16571 67555 -16519 67607
rect -15416 67549 -15364 67601
rect -14298 67560 -14246 67612
rect -9881 63344 -9829 63396
rect -9817 63344 -9765 63396
rect -9753 63344 -9701 63396
rect -9689 63344 -9637 63396
rect -9625 63344 -9573 63396
rect -9561 63344 -9509 63396
rect -9497 63344 -9445 63396
rect -8070 63346 -8018 63398
rect -8006 63346 -7954 63398
rect -7942 63346 -7890 63398
rect -7878 63346 -7826 63398
rect -7814 63346 -7762 63398
rect -7750 63346 -7698 63398
rect -7686 63346 -7634 63398
rect -6275 63342 -6223 63394
rect -6211 63342 -6159 63394
rect -6147 63342 -6095 63394
rect -6083 63342 -6031 63394
rect -6019 63342 -5967 63394
rect -5955 63342 -5903 63394
rect -5891 63342 -5839 63394
rect -4476 63340 -4424 63392
rect -4412 63340 -4360 63392
rect -4348 63340 -4296 63392
rect -4284 63340 -4232 63392
rect -4220 63340 -4168 63392
rect -4156 63340 -4104 63392
rect -4092 63340 -4040 63392
rect -6909 62996 -6729 63176
rect -2685 63344 -2633 63396
rect -2621 63344 -2569 63396
rect -2557 63344 -2505 63396
rect -2493 63344 -2441 63396
rect -2429 63344 -2377 63396
rect -2365 63344 -2313 63396
rect -2301 63344 -2249 63396
rect -883 63340 -831 63392
rect -819 63340 -767 63392
rect -755 63340 -703 63392
rect -691 63340 -639 63392
rect -627 63340 -575 63392
rect -563 63340 -511 63392
rect -499 63340 -447 63392
rect 772 63022 1272 63202
rect -8551 54537 -8499 54589
rect -6860 54538 -6808 54590
rect -5155 54537 -5103 54589
rect -3359 54537 -3307 54589
rect -1530 54537 -1478 54589
rect -9673 54345 -9621 54397
rect -9609 54345 -9557 54397
rect -9545 54345 -9493 54397
rect -7878 54344 -7826 54396
rect -7814 54344 -7762 54396
rect -7750 54344 -7698 54396
rect -6078 54346 -6026 54398
rect -6014 54346 -5962 54398
rect -5950 54346 -5898 54398
rect -4280 54345 -4228 54397
rect -4216 54345 -4164 54397
rect -4152 54345 -4100 54397
rect -2482 54346 -2430 54398
rect -2418 54346 -2366 54398
rect -2354 54346 -2302 54398
rect -679 54345 -627 54397
rect -615 54345 -563 54397
rect -551 54345 -499 54397
rect 182 54346 234 54398
rect -14777 53542 -14725 53594
rect -14713 53542 -14661 53594
rect -7544 53542 -7492 53594
rect -6983 53542 -6931 53594
rect -6919 53542 -6867 53594
rect 375 60746 491 60808
rect 375 60712 410 60746
rect 410 60712 444 60746
rect 444 60712 491 60746
rect 375 60674 491 60712
rect 375 60640 410 60674
rect 410 60640 444 60674
rect 444 60640 491 60674
rect 375 60602 491 60640
rect 375 60568 410 60602
rect 410 60568 444 60602
rect 444 60568 491 60602
rect 375 60530 491 60568
rect 375 60496 410 60530
rect 410 60496 444 60530
rect 444 60496 491 60530
rect 375 60458 491 60496
rect 375 60424 410 60458
rect 410 60424 444 60458
rect 444 60424 491 60458
rect 375 60386 491 60424
rect 375 60352 410 60386
rect 410 60352 444 60386
rect 444 60352 491 60386
rect 375 60314 491 60352
rect 375 60280 410 60314
rect 410 60280 444 60314
rect 444 60280 491 60314
rect 375 60242 491 60280
rect 375 60208 410 60242
rect 410 60208 444 60242
rect 444 60208 491 60242
rect 375 60170 491 60208
rect 375 60136 410 60170
rect 410 60136 444 60170
rect 444 60136 491 60170
rect 375 60098 491 60136
rect 375 60064 410 60098
rect 410 60064 444 60098
rect 444 60064 491 60098
rect 375 60026 491 60064
rect 375 59992 410 60026
rect 410 59992 444 60026
rect 444 59992 491 60026
rect 375 59954 491 59992
rect 375 59920 410 59954
rect 410 59920 444 59954
rect 444 59920 491 59954
rect 375 59882 491 59920
rect 375 59848 410 59882
rect 410 59848 444 59882
rect 444 59848 491 59882
rect 375 59810 491 59848
rect 375 59776 410 59810
rect 410 59776 444 59810
rect 444 59776 491 59810
rect 375 59738 491 59776
rect 375 59704 410 59738
rect 410 59704 444 59738
rect 444 59704 491 59738
rect 375 59666 491 59704
rect 375 59632 410 59666
rect 410 59632 444 59666
rect 444 59632 491 59666
rect 375 59594 491 59632
rect 375 59560 410 59594
rect 410 59560 444 59594
rect 444 59560 491 59594
rect 375 59522 491 59560
rect 375 59488 410 59522
rect 410 59488 444 59522
rect 444 59488 491 59522
rect 375 59450 491 59488
rect 375 59416 410 59450
rect 410 59416 444 59450
rect 444 59416 491 59450
rect 375 59378 491 59416
rect 375 59344 410 59378
rect 410 59344 444 59378
rect 444 59344 491 59378
rect 375 59306 491 59344
rect 375 59272 410 59306
rect 410 59272 444 59306
rect 444 59272 491 59306
rect 375 59234 491 59272
rect 375 59200 410 59234
rect 410 59200 444 59234
rect 444 59200 491 59234
rect 375 59162 491 59200
rect 375 59128 410 59162
rect 410 59128 444 59162
rect 444 59128 491 59162
rect 375 59090 491 59128
rect 375 59056 410 59090
rect 410 59056 444 59090
rect 444 59056 491 59090
rect 375 59018 491 59056
rect 375 58984 410 59018
rect 410 58984 444 59018
rect 444 58984 491 59018
rect 375 58946 491 58984
rect 375 58912 410 58946
rect 410 58912 444 58946
rect 444 58912 491 58946
rect 375 58874 491 58912
rect 375 58840 410 58874
rect 410 58840 444 58874
rect 444 58840 491 58874
rect 375 58802 491 58840
rect 375 58768 410 58802
rect 410 58768 444 58802
rect 444 58768 491 58802
rect 375 58730 491 58768
rect 375 58696 410 58730
rect 410 58696 444 58730
rect 444 58696 491 58730
rect 375 58658 491 58696
rect 375 58624 410 58658
rect 410 58624 444 58658
rect 444 58624 491 58658
rect 375 58586 491 58624
rect 375 58552 410 58586
rect 410 58552 444 58586
rect 444 58552 491 58586
rect 375 58514 491 58552
rect 375 58480 410 58514
rect 410 58480 444 58514
rect 444 58480 491 58514
rect 375 58442 491 58480
rect 375 58408 410 58442
rect 410 58408 444 58442
rect 444 58408 491 58442
rect 375 58370 491 58408
rect 375 58336 410 58370
rect 410 58336 444 58370
rect 444 58336 491 58370
rect 375 58298 491 58336
rect 375 58264 410 58298
rect 410 58264 444 58298
rect 444 58264 491 58298
rect 375 58226 491 58264
rect 375 58192 410 58226
rect 410 58192 444 58226
rect 444 58192 491 58226
rect 375 58154 491 58192
rect 375 58120 410 58154
rect 410 58120 444 58154
rect 444 58120 491 58154
rect 375 58082 491 58120
rect 375 58048 410 58082
rect 410 58048 444 58082
rect 444 58048 491 58082
rect 375 58010 491 58048
rect 375 57976 410 58010
rect 410 57976 444 58010
rect 444 57976 491 58010
rect 375 57938 491 57976
rect 375 57904 410 57938
rect 410 57904 444 57938
rect 444 57904 491 57938
rect 375 57866 491 57904
rect 375 57832 410 57866
rect 410 57832 444 57866
rect 444 57832 491 57866
rect 375 57794 491 57832
rect 375 57760 410 57794
rect 410 57760 444 57794
rect 444 57760 491 57794
rect 375 57722 491 57760
rect 375 57688 410 57722
rect 410 57688 444 57722
rect 444 57688 491 57722
rect 375 57650 491 57688
rect 375 57616 410 57650
rect 410 57616 444 57650
rect 444 57616 491 57650
rect 375 57578 491 57616
rect 375 57544 410 57578
rect 410 57544 444 57578
rect 444 57544 491 57578
rect 375 57506 491 57544
rect 375 57472 410 57506
rect 410 57472 444 57506
rect 444 57472 491 57506
rect 375 57434 491 57472
rect 375 57400 410 57434
rect 410 57400 444 57434
rect 444 57400 491 57434
rect 375 57362 491 57400
rect 375 57328 410 57362
rect 410 57328 444 57362
rect 444 57328 491 57362
rect 375 57290 491 57328
rect 375 57256 410 57290
rect 410 57256 444 57290
rect 444 57256 491 57290
rect 375 57218 491 57256
rect 375 57184 410 57218
rect 410 57184 444 57218
rect 444 57184 491 57218
rect 375 57146 491 57184
rect 375 57112 410 57146
rect 410 57112 444 57146
rect 444 57112 491 57146
rect 375 57074 491 57112
rect 375 57040 410 57074
rect 410 57040 444 57074
rect 444 57040 491 57074
rect 375 57002 491 57040
rect 375 56968 410 57002
rect 410 56968 444 57002
rect 444 56968 491 57002
rect 375 56930 491 56968
rect 375 56896 410 56930
rect 410 56896 444 56930
rect 444 56896 491 56930
rect 375 56858 491 56896
rect 375 56824 410 56858
rect 410 56824 444 56858
rect 444 56824 491 56858
rect 375 56786 491 56824
rect 375 56752 410 56786
rect 410 56752 444 56786
rect 444 56752 491 56786
rect 375 56714 491 56752
rect 375 56680 410 56714
rect 410 56680 444 56714
rect 444 56680 491 56714
rect 375 56642 491 56680
rect 375 56608 410 56642
rect 410 56608 444 56642
rect 444 56608 491 56642
rect 375 56570 491 56608
rect 375 56536 410 56570
rect 410 56536 444 56570
rect 444 56536 491 56570
rect 375 56498 491 56536
rect 375 56464 410 56498
rect 410 56464 444 56498
rect 444 56464 491 56498
rect 375 56426 491 56464
rect 375 56392 410 56426
rect 410 56392 444 56426
rect 444 56392 491 56426
rect 375 56354 491 56392
rect 375 56320 410 56354
rect 410 56320 444 56354
rect 444 56320 491 56354
rect 375 56282 491 56320
rect 375 56248 410 56282
rect 410 56248 444 56282
rect 444 56248 491 56282
rect 375 56210 491 56248
rect 375 56176 410 56210
rect 410 56176 444 56210
rect 444 56176 491 56210
rect 375 56138 491 56176
rect 375 56104 410 56138
rect 410 56104 444 56138
rect 444 56104 491 56138
rect 375 56066 491 56104
rect 375 56032 410 56066
rect 410 56032 444 56066
rect 444 56032 491 56066
rect 375 55994 491 56032
rect 375 55960 410 55994
rect 410 55960 444 55994
rect 444 55960 491 55994
rect 375 55922 491 55960
rect 375 55888 410 55922
rect 410 55888 444 55922
rect 444 55888 491 55922
rect 375 55850 491 55888
rect 375 55816 410 55850
rect 410 55816 444 55850
rect 444 55816 491 55850
rect 375 55778 491 55816
rect 375 55744 410 55778
rect 410 55744 444 55778
rect 444 55744 491 55778
rect 375 55706 491 55744
rect 375 55672 410 55706
rect 410 55672 444 55706
rect 444 55672 491 55706
rect 375 55634 491 55672
rect 375 55600 410 55634
rect 410 55600 444 55634
rect 444 55600 491 55634
rect 375 55562 491 55600
rect 375 55528 410 55562
rect 410 55528 444 55562
rect 444 55528 491 55562
rect 375 55490 491 55528
rect 375 55456 410 55490
rect 410 55456 444 55490
rect 444 55456 491 55490
rect 375 55418 491 55456
rect 375 55384 410 55418
rect 410 55384 444 55418
rect 444 55384 491 55418
rect 375 55346 491 55384
rect 375 55312 410 55346
rect 410 55312 444 55346
rect 444 55312 491 55346
rect 375 55274 491 55312
rect 375 55240 410 55274
rect 410 55240 444 55274
rect 444 55240 491 55274
rect 375 55202 491 55240
rect 375 55168 410 55202
rect 410 55168 444 55202
rect 444 55168 491 55202
rect 375 55130 491 55168
rect 375 55096 410 55130
rect 410 55096 444 55130
rect 444 55096 491 55130
rect 375 55058 491 55096
rect 375 55024 410 55058
rect 410 55024 444 55058
rect 444 55024 491 55058
rect 375 54986 491 55024
rect 375 54952 410 54986
rect 410 54952 444 54986
rect 444 54952 491 54986
rect 375 54914 491 54952
rect 375 54880 410 54914
rect 410 54880 444 54914
rect 444 54880 491 54914
rect 375 54842 491 54880
rect 375 54808 410 54842
rect 410 54808 444 54842
rect 444 54808 491 54842
rect 375 54770 491 54808
rect 375 54736 410 54770
rect 410 54736 444 54770
rect 444 54736 491 54770
rect 375 54698 491 54736
rect 375 54664 410 54698
rect 410 54664 444 54698
rect 444 54664 491 54698
rect 375 54626 491 54664
rect 375 54592 410 54626
rect 410 54592 444 54626
rect 444 54592 491 54626
rect 375 54554 491 54592
rect 375 54520 410 54554
rect 410 54520 444 54554
rect 444 54520 491 54554
rect 375 54482 491 54520
rect 375 54448 410 54482
rect 410 54448 444 54482
rect 444 54448 491 54482
rect 375 54410 491 54448
rect 375 54376 410 54410
rect 410 54376 444 54410
rect 444 54376 491 54410
rect 375 54338 491 54376
rect 375 54304 410 54338
rect 410 54304 444 54338
rect 444 54304 491 54338
rect 375 54266 491 54304
rect 375 54232 410 54266
rect 410 54232 444 54266
rect 444 54232 491 54266
rect 375 54194 491 54232
rect 375 54160 410 54194
rect 410 54160 444 54194
rect 444 54160 491 54194
rect 375 54122 491 54160
rect 375 54088 410 54122
rect 410 54088 444 54122
rect 444 54088 491 54122
rect 375 54050 491 54088
rect 375 54016 410 54050
rect 410 54016 444 54050
rect 444 54016 491 54050
rect 375 53978 491 54016
rect 375 53944 410 53978
rect 410 53944 444 53978
rect 444 53944 491 53978
rect 375 53906 491 53944
rect 375 53872 410 53906
rect 410 53872 444 53906
rect 444 53872 491 53906
rect 375 53834 491 53872
rect 375 53800 410 53834
rect 410 53800 444 53834
rect 444 53800 491 53834
rect 375 53762 491 53800
rect 375 53728 410 53762
rect 410 53728 444 53762
rect 444 53728 491 53762
rect 375 53690 491 53728
rect 375 53656 410 53690
rect 410 53656 444 53690
rect 444 53656 491 53690
rect 375 53618 491 53656
rect 375 53584 410 53618
rect 410 53584 444 53618
rect 444 53584 491 53618
rect 375 53546 491 53584
rect 375 53512 410 53546
rect 410 53512 444 53546
rect 444 53512 491 53546
rect 375 53474 491 53512
rect 375 53440 410 53474
rect 410 53440 444 53474
rect 444 53440 491 53474
rect 375 53402 491 53440
rect 375 53368 410 53402
rect 410 53368 444 53402
rect 444 53368 491 53402
rect 375 53330 491 53368
rect 375 53296 410 53330
rect 410 53296 444 53330
rect 444 53296 491 53330
rect 375 53258 491 53296
rect 375 53224 410 53258
rect 410 53224 444 53258
rect 444 53224 491 53258
rect 375 53186 491 53224
rect 375 53152 410 53186
rect 410 53152 444 53186
rect 444 53152 491 53186
rect 375 53140 491 53152
rect -9392 52934 -9340 52986
rect -9328 52934 -9276 52986
rect -8838 51169 -8786 51221
rect -8838 51105 -8786 51157
rect -8838 51041 -8786 51093
rect -9392 50879 -9340 50931
rect -9328 50879 -9276 50931
rect -6983 50877 -6931 50929
rect -6919 50877 -6867 50929
rect -5678 50988 -3898 51064
rect -3359 50988 -2539 51043
rect -1652 50988 -768 51033
rect -5678 50954 -5607 50988
rect -5607 50954 -5573 50988
rect -5573 50954 -5535 50988
rect -5535 50954 -5501 50988
rect -5501 50954 -5463 50988
rect -5463 50954 -5429 50988
rect -5429 50954 -5391 50988
rect -5391 50954 -5357 50988
rect -5357 50954 -5319 50988
rect -5319 50954 -5285 50988
rect -5285 50954 -5247 50988
rect -5247 50954 -5213 50988
rect -5213 50954 -5175 50988
rect -5175 50954 -5141 50988
rect -5141 50954 -5103 50988
rect -5103 50954 -5069 50988
rect -5069 50954 -5031 50988
rect -5031 50954 -4997 50988
rect -4997 50954 -4959 50988
rect -4959 50954 -4925 50988
rect -4925 50954 -4887 50988
rect -4887 50954 -4853 50988
rect -4853 50954 -4815 50988
rect -4815 50954 -4781 50988
rect -4781 50954 -4743 50988
rect -4743 50954 -4709 50988
rect -4709 50954 -4671 50988
rect -4671 50954 -4637 50988
rect -4637 50954 -4599 50988
rect -4599 50954 -4565 50988
rect -4565 50954 -4527 50988
rect -4527 50954 -4493 50988
rect -4493 50954 -4455 50988
rect -4455 50954 -4421 50988
rect -4421 50954 -4383 50988
rect -4383 50954 -4349 50988
rect -4349 50954 -4311 50988
rect -4311 50954 -4277 50988
rect -4277 50954 -4239 50988
rect -4239 50954 -4205 50988
rect -4205 50954 -4167 50988
rect -4167 50954 -4133 50988
rect -4133 50954 -4095 50988
rect -4095 50954 -4061 50988
rect -4061 50954 -4023 50988
rect -4023 50954 -3989 50988
rect -3989 50954 -3951 50988
rect -3951 50954 -3917 50988
rect -3917 50954 -3898 50988
rect -3359 50954 -3341 50988
rect -3341 50954 -3303 50988
rect -3303 50954 -3269 50988
rect -3269 50954 -3231 50988
rect -3231 50954 -3197 50988
rect -3197 50954 -3159 50988
rect -3159 50954 -3125 50988
rect -3125 50954 -3087 50988
rect -3087 50954 -3053 50988
rect -3053 50954 -3015 50988
rect -3015 50954 -2981 50988
rect -2981 50954 -2943 50988
rect -2943 50954 -2909 50988
rect -2909 50954 -2871 50988
rect -2871 50954 -2837 50988
rect -2837 50954 -2799 50988
rect -2799 50954 -2765 50988
rect -2765 50954 -2727 50988
rect -2727 50954 -2693 50988
rect -2693 50954 -2655 50988
rect -2655 50954 -2621 50988
rect -2621 50954 -2583 50988
rect -2583 50954 -2549 50988
rect -2549 50954 -2539 50988
rect -1652 50954 -1647 50988
rect -1647 50954 -1613 50988
rect -1613 50954 -1575 50988
rect -1575 50954 -1541 50988
rect -1541 50954 -1503 50988
rect -1503 50954 -1469 50988
rect -1469 50954 -1431 50988
rect -1431 50954 -1397 50988
rect -1397 50954 -1359 50988
rect -1359 50954 -1325 50988
rect -1325 50954 -1287 50988
rect -1287 50954 -1253 50988
rect -1253 50954 -1215 50988
rect -1215 50954 -1181 50988
rect -1181 50954 -1143 50988
rect -1143 50954 -1109 50988
rect -1109 50954 -1071 50988
rect -1071 50954 -1037 50988
rect -1037 50954 -999 50988
rect -999 50954 -965 50988
rect -965 50954 -927 50988
rect -927 50954 -893 50988
rect -893 50954 -855 50988
rect -855 50954 -821 50988
rect -821 50954 -783 50988
rect -783 50954 -768 50988
rect -5678 50884 -3898 50954
rect -3359 50927 -2539 50954
rect -1652 50917 -768 50954
rect -8853 50718 -8801 50770
rect -8853 50654 -8801 50706
rect -8853 50590 -8801 50642
rect -8853 50526 -8801 50578
rect -8853 50462 -8801 50514
rect -8853 50398 -8801 50450
rect -27052 49662 -27000 49714
rect -26988 49662 -26936 49714
rect -26924 49662 -26872 49714
rect -26860 49662 -26808 49714
rect -26796 49662 -26744 49714
rect -26405 49398 -26353 49407
rect -26341 49398 -26289 49407
rect -26277 49398 -26225 49407
rect -26213 49398 -26161 49407
rect -26405 49364 -26377 49398
rect -26377 49364 -26353 49398
rect -26341 49364 -26305 49398
rect -26305 49364 -26289 49398
rect -26277 49364 -26271 49398
rect -26271 49364 -26233 49398
rect -26233 49364 -26225 49398
rect -26213 49364 -26199 49398
rect -26199 49364 -26161 49398
rect -26405 49355 -26353 49364
rect -26341 49355 -26289 49364
rect -26277 49355 -26225 49364
rect -26213 49355 -26161 49364
rect -26054 49413 -26047 49418
rect -26047 49413 -26013 49418
rect -26013 49413 -26002 49418
rect -26054 49366 -26002 49413
rect -25966 49120 -25914 49172
rect -25902 49120 -25850 49172
rect -25838 49120 -25786 49172
rect -25774 49120 -25722 49172
rect -25710 49120 -25658 49172
rect -5930 47782 -5750 50714
rect -69 50713 111 50761
rect -69 50679 25 50713
rect 25 50679 59 50713
rect 59 50679 111 50713
rect -69 50641 111 50679
rect -69 50607 25 50641
rect 25 50607 59 50641
rect 59 50607 111 50641
rect -69 50569 111 50607
rect -69 50535 25 50569
rect 25 50535 59 50569
rect 59 50535 111 50569
rect -69 50497 111 50535
rect -69 50463 25 50497
rect 25 50463 59 50497
rect 59 50463 111 50497
rect -69 50425 111 50463
rect -69 50391 25 50425
rect 25 50391 59 50425
rect 59 50391 111 50425
rect -69 50353 111 50391
rect -69 50319 25 50353
rect 25 50319 59 50353
rect 59 50319 111 50353
rect -69 50281 111 50319
rect -69 50247 25 50281
rect 25 50247 59 50281
rect 59 50247 111 50281
rect -69 50209 111 50247
rect -69 50175 25 50209
rect 25 50175 59 50209
rect 59 50175 111 50209
rect -69 50137 111 50175
rect -69 50103 25 50137
rect 25 50103 59 50137
rect 59 50103 111 50137
rect -69 50065 111 50103
rect -69 50031 25 50065
rect 25 50031 59 50065
rect 59 50031 111 50065
rect -69 49993 111 50031
rect -69 49959 25 49993
rect 25 49959 59 49993
rect 59 49959 111 49993
rect -69 49921 111 49959
rect -69 49887 25 49921
rect 25 49887 59 49921
rect 59 49887 111 49921
rect -69 49849 111 49887
rect -69 49815 25 49849
rect 25 49815 59 49849
rect 59 49815 111 49849
rect -69 49777 111 49815
rect -69 49743 25 49777
rect 25 49743 59 49777
rect 59 49743 111 49777
rect -69 49705 111 49743
rect -69 49671 25 49705
rect 25 49671 59 49705
rect 59 49671 111 49705
rect -69 49633 111 49671
rect -69 49599 25 49633
rect 25 49599 59 49633
rect 59 49599 111 49633
rect -69 49561 111 49599
rect -69 49527 25 49561
rect 25 49527 59 49561
rect 59 49527 111 49561
rect -69 49489 111 49527
rect -69 49455 25 49489
rect 25 49455 59 49489
rect 59 49455 111 49489
rect -69 49417 111 49455
rect -69 49383 25 49417
rect 25 49383 59 49417
rect 59 49383 111 49417
rect -69 49345 111 49383
rect -69 49311 25 49345
rect 25 49311 59 49345
rect 59 49311 111 49345
rect -69 49273 111 49311
rect -69 49239 25 49273
rect 25 49239 59 49273
rect 59 49239 111 49273
rect -69 49201 111 49239
rect -69 49167 25 49201
rect 25 49167 59 49201
rect 59 49167 111 49201
rect -69 49129 111 49167
rect -69 49095 25 49129
rect 25 49095 59 49129
rect 59 49095 111 49129
rect -69 49057 111 49095
rect -69 49023 25 49057
rect 25 49023 59 49057
rect 59 49023 111 49057
rect -69 48985 111 49023
rect -69 48951 25 48985
rect 25 48951 59 48985
rect 59 48951 111 48985
rect -69 48913 111 48951
rect -69 48879 25 48913
rect 25 48879 59 48913
rect 59 48879 111 48913
rect -69 48841 111 48879
rect -69 48807 25 48841
rect 25 48807 59 48841
rect 59 48807 111 48841
rect -69 48769 111 48807
rect -69 48735 25 48769
rect 25 48735 59 48769
rect 59 48735 111 48769
rect -69 48697 111 48735
rect -69 48663 25 48697
rect 25 48663 59 48697
rect 59 48663 111 48697
rect -69 48625 111 48663
rect -69 48591 25 48625
rect 25 48591 59 48625
rect 59 48591 111 48625
rect -69 48553 111 48591
rect -69 48519 25 48553
rect 25 48519 59 48553
rect 59 48519 111 48553
rect -69 48481 111 48519
rect -69 48447 25 48481
rect 25 48447 59 48481
rect 59 48447 111 48481
rect -69 48409 111 48447
rect -69 48375 25 48409
rect 25 48375 59 48409
rect 59 48375 111 48409
rect -69 48337 111 48375
rect -69 48303 25 48337
rect 25 48303 59 48337
rect 59 48303 111 48337
rect -69 48265 111 48303
rect -69 48231 25 48265
rect 25 48231 59 48265
rect 59 48231 111 48265
rect -69 48193 111 48231
rect -69 48159 25 48193
rect 25 48159 59 48193
rect 59 48159 111 48193
rect -69 48121 111 48159
rect -69 48087 25 48121
rect 25 48087 59 48121
rect 59 48087 111 48121
rect -69 48049 111 48087
rect -69 48015 25 48049
rect 25 48015 59 48049
rect 59 48015 111 48049
rect -69 47977 111 48015
rect -69 47943 25 47977
rect 25 47943 59 47977
rect 59 47943 111 47977
rect -69 47905 111 47943
rect -69 47871 25 47905
rect 25 47871 59 47905
rect 59 47871 111 47905
rect -69 47833 111 47871
rect -69 47799 25 47833
rect 25 47799 59 47833
rect 59 47799 111 47833
rect -69 47765 111 47799
rect 10178 47640 10550 60812
rect -27065 43244 -27013 43296
rect -27065 43180 -27013 43232
rect -27065 43116 -27013 43168
rect -27065 43052 -27013 43104
rect -27065 42988 -27013 43040
rect -13463 43003 -13411 43055
rect -27065 42924 -27013 42976
rect -27065 42860 -27013 42912
rect -27065 42796 -27013 42848
rect -27065 42103 -27013 42155
rect -27065 42039 -27013 42091
rect -27065 41975 -27013 42027
rect -27065 41911 -27013 41963
rect -27065 41847 -27013 41899
rect -27065 41783 -27013 41835
rect -27065 41719 -27013 41771
rect -27065 41655 -27013 41707
rect -27065 41591 -27013 41643
rect -27065 41527 -27013 41579
rect -27065 41463 -27013 41515
rect -27065 41399 -27013 41451
rect -27065 41335 -27013 41387
rect -27065 41271 -27013 41323
rect -27065 41207 -27013 41259
rect -27065 41143 -27013 41195
rect -27065 41079 -27013 41131
rect -27065 41015 -27013 41067
rect -27060 40577 -27008 40629
rect -27060 40513 -27008 40565
rect -27060 40449 -27008 40501
rect -27060 40385 -27008 40437
rect -27060 40321 -27008 40373
rect -27060 40257 -27008 40309
rect -27060 40193 -27008 40245
rect -27060 40129 -27008 40181
rect -27060 40065 -27008 40117
rect -27060 40001 -27008 40053
rect -27060 39937 -27008 39989
rect -27060 39873 -27008 39925
rect -27060 39809 -27008 39861
rect -27060 39745 -27008 39797
rect -27060 39681 -27008 39733
rect -27060 39617 -27008 39669
rect -27060 39553 -27008 39605
rect -27060 39489 -27008 39541
rect -18871 39468 -18819 39520
rect -18871 39404 -18819 39456
rect -18871 39340 -18819 39392
rect -18871 39276 -18819 39328
rect -18871 39212 -18819 39264
rect -31806 39114 -31754 39150
rect -31806 39098 -31795 39114
rect -31795 39098 -31761 39114
rect -31761 39098 -31754 39114
rect -18871 39148 -18819 39200
rect -31806 39080 -31795 39086
rect -31795 39080 -31761 39086
rect -31761 39080 -31754 39086
rect -31806 39042 -31754 39080
rect -31806 39034 -31795 39042
rect -31795 39034 -31761 39042
rect -31761 39034 -31754 39042
rect -31806 39008 -31795 39022
rect -31795 39008 -31761 39022
rect -31761 39008 -31754 39022
rect -31806 38970 -31754 39008
rect -31806 38936 -31795 38958
rect -31795 38936 -31761 38958
rect -31761 38936 -31754 38958
rect -31806 38906 -31754 38936
rect -31806 38864 -31795 38894
rect -31795 38864 -31761 38894
rect -31761 38864 -31754 38894
rect -31806 38842 -31754 38864
rect -31805 38550 -31753 38595
rect -31805 38543 -31795 38550
rect -31795 38543 -31761 38550
rect -31761 38543 -31753 38550
rect -31805 38516 -31795 38531
rect -31795 38516 -31761 38531
rect -31761 38516 -31753 38531
rect -31805 38479 -31753 38516
rect -31805 38444 -31795 38467
rect -31795 38444 -31761 38467
rect -31761 38444 -31753 38467
rect -31805 38415 -31753 38444
rect -31805 38372 -31795 38403
rect -31795 38372 -31761 38403
rect -31761 38372 -31753 38403
rect -31805 38351 -31753 38372
rect -31805 38334 -31753 38339
rect -31805 38300 -31795 38334
rect -31795 38300 -31761 38334
rect -31761 38300 -31753 38334
rect -31805 38287 -31753 38300
rect -31805 38262 -31753 38275
rect -31805 38228 -31795 38262
rect -31795 38228 -31761 38262
rect -31761 38228 -31753 38262
rect -31805 38223 -31753 38228
rect -27066 39066 -27014 39118
rect -27066 39002 -27014 39054
rect -27066 38938 -27014 38990
rect -27066 38874 -27014 38926
rect -27066 38810 -27014 38862
rect -27066 38746 -27014 38798
rect -27066 38682 -27014 38734
rect -27066 38618 -27014 38670
rect -27066 38554 -27014 38606
rect -27066 38490 -27014 38542
rect -27066 38426 -27014 38478
rect -29600 38355 -29548 38407
rect -29536 38355 -29484 38407
rect -29472 38355 -29420 38407
rect -29408 38355 -29356 38407
rect -29344 38355 -29292 38407
rect -29280 38355 -29228 38407
rect -29216 38355 -29164 38407
rect -27066 38362 -27014 38414
rect -27066 38298 -27014 38350
rect -31805 38159 -31753 38211
rect -31024 38198 -30972 38250
rect -30960 38198 -30908 38250
rect -27066 38234 -27014 38286
rect -18871 39084 -18819 39136
rect -18871 39020 -18819 39072
rect -18871 38956 -18819 39008
rect -18871 38892 -18819 38944
rect -18871 38828 -18819 38880
rect -18871 38764 -18819 38816
rect -18871 38700 -18819 38752
rect -18871 38636 -18819 38688
rect -18871 38572 -18819 38624
rect -18871 38508 -18819 38560
rect -18871 38444 -18819 38496
rect -18871 38380 -18819 38432
rect -18871 38316 -18819 38368
rect -18871 38252 -18819 38304
rect -18871 38188 -18819 38240
rect -18871 38124 -18819 38176
rect -18871 38060 -18819 38112
rect -18871 37996 -18819 38048
rect -18871 37932 -18819 37984
rect -18871 37868 -18819 37920
rect -18871 37804 -18819 37856
rect -18871 37740 -18819 37792
rect -18871 37676 -18819 37728
rect -18871 37612 -18819 37664
rect -35490 37360 -35310 37540
rect -18871 37548 -18819 37600
rect -18871 37484 -18819 37536
rect -30193 37417 -30141 37469
rect -30129 37417 -30077 37469
rect -18871 37420 -18819 37472
rect -18871 37356 -18819 37408
rect -29648 37265 -29596 37317
rect -29584 37265 -29532 37317
rect -29520 37265 -29468 37317
rect -29456 37265 -29404 37317
rect -29392 37265 -29340 37317
rect -29328 37265 -29276 37317
rect -29264 37265 -29212 37317
rect -29200 37265 -29148 37317
rect -27063 37299 -27011 37351
rect -27063 37235 -27011 37287
rect -27063 37171 -27011 37223
rect -27063 37107 -27011 37159
rect -27063 37043 -27011 37095
rect -27063 36979 -27011 37031
rect -27063 36915 -27011 36967
rect -27063 36851 -27011 36903
rect -27063 36787 -27011 36839
rect -27063 36723 -27011 36775
rect -27063 36659 -27011 36711
rect -27063 36595 -27011 36647
rect -27063 36531 -27011 36583
rect -27063 36467 -27011 36519
rect -18871 37292 -18819 37344
rect -18871 37228 -18819 37280
rect -18871 37164 -18819 37216
rect -18871 37100 -18819 37152
rect -18871 37036 -18819 37088
rect -18871 36972 -18819 37024
rect -18871 36908 -18819 36960
rect -18871 36844 -18819 36896
rect -18871 36780 -18819 36832
rect -18871 36716 -18819 36768
rect -18871 36652 -18819 36704
rect -18871 36588 -18819 36640
rect -18871 36524 -18819 36576
rect -18871 36460 -18819 36512
rect -18871 36396 -18819 36448
rect -18871 36332 -18819 36384
rect -18871 36268 -18819 36320
rect -18871 36204 -18819 36256
rect -27063 36090 -27011 36142
rect -18871 36140 -18819 36192
rect -27063 36026 -27011 36078
rect -27063 35962 -27011 36014
rect -27063 35898 -27011 35950
rect -27063 35834 -27011 35886
rect -27063 35770 -27011 35822
rect -27063 35706 -27011 35758
rect -27063 35642 -27011 35694
rect -27063 35578 -27011 35630
rect -27063 35514 -27011 35566
rect -27063 35450 -27011 35502
rect -27063 35386 -27011 35438
rect -27063 35322 -27011 35374
rect -27063 35258 -27011 35310
rect -27063 35194 -27011 35246
rect -27063 35130 -27011 35182
rect -27063 35066 -27011 35118
rect -27063 35002 -27011 35054
rect -27066 34612 -27014 34664
rect -27066 34548 -27014 34600
rect -27066 34484 -27014 34536
rect -27066 34420 -27014 34472
rect -27066 34356 -27014 34408
rect -27066 34292 -27014 34344
rect -27066 34228 -27014 34280
rect -27066 34164 -27014 34216
rect -27066 34100 -27014 34152
rect -27066 34036 -27014 34088
rect -27066 33972 -27014 34024
rect -27066 33908 -27014 33960
rect -27066 33844 -27014 33896
rect -27066 33780 -27014 33832
rect -27066 33716 -27014 33768
rect -27066 33652 -27014 33704
rect -27066 33588 -27014 33640
rect -27066 33524 -27014 33576
rect -27071 32830 -27019 32882
rect -27071 32766 -27019 32818
rect -27071 32702 -27019 32754
rect -27071 32638 -27019 32690
rect -27071 32574 -27019 32626
rect -27071 32510 -27019 32562
rect -27071 32446 -27019 32498
rect -27071 32382 -27019 32434
rect -12687 42340 -12635 42392
rect -5913 39820 -5733 46272
rect -9392 39747 -9340 39799
rect -9328 39747 -9276 39799
rect -6983 39747 -6931 39799
rect -6919 39747 -6867 39799
rect -9363 34618 -9311 34670
rect -5662 39773 -170 39846
rect -5662 39739 -5620 39773
rect -5620 39739 -5586 39773
rect -5586 39739 -5548 39773
rect -5548 39739 -5514 39773
rect -5514 39739 -5476 39773
rect -5476 39739 -5442 39773
rect -5442 39739 -5404 39773
rect -5404 39739 -5370 39773
rect -5370 39739 -5332 39773
rect -5332 39739 -5298 39773
rect -5298 39739 -5260 39773
rect -5260 39739 -5226 39773
rect -5226 39739 -5188 39773
rect -5188 39739 -5154 39773
rect -5154 39739 -5116 39773
rect -5116 39739 -5082 39773
rect -5082 39739 -5044 39773
rect -5044 39739 -5010 39773
rect -5010 39739 -4972 39773
rect -4972 39739 -4938 39773
rect -4938 39739 -4900 39773
rect -4900 39739 -4866 39773
rect -4866 39739 -4828 39773
rect -4828 39739 -4794 39773
rect -4794 39739 -4756 39773
rect -4756 39739 -4722 39773
rect -4722 39739 -4684 39773
rect -4684 39739 -4650 39773
rect -4650 39739 -4612 39773
rect -4612 39739 -4578 39773
rect -4578 39739 -4540 39773
rect -4540 39739 -4506 39773
rect -4506 39739 -4468 39773
rect -4468 39739 -4434 39773
rect -4434 39739 -4396 39773
rect -4396 39739 -4362 39773
rect -4362 39739 -4324 39773
rect -4324 39739 -4290 39773
rect -4290 39739 -4252 39773
rect -4252 39739 -4218 39773
rect -4218 39739 -4180 39773
rect -4180 39739 -4146 39773
rect -4146 39739 -4108 39773
rect -4108 39739 -4074 39773
rect -4074 39739 -4036 39773
rect -4036 39739 -4002 39773
rect -4002 39739 -3964 39773
rect -3964 39739 -3930 39773
rect -3930 39739 -3892 39773
rect -3892 39739 -3858 39773
rect -3858 39739 -3820 39773
rect -3820 39739 -3786 39773
rect -3786 39739 -3748 39773
rect -3748 39739 -3714 39773
rect -3714 39739 -3676 39773
rect -3676 39739 -3642 39773
rect -3642 39739 -3604 39773
rect -3604 39739 -3570 39773
rect -3570 39739 -3532 39773
rect -3532 39739 -3498 39773
rect -3498 39739 -3460 39773
rect -3460 39739 -3426 39773
rect -3426 39739 -3388 39773
rect -3388 39739 -3354 39773
rect -3354 39739 -3316 39773
rect -3316 39739 -3282 39773
rect -3282 39739 -3244 39773
rect -3244 39739 -3210 39773
rect -3210 39739 -3172 39773
rect -3172 39739 -3138 39773
rect -3138 39739 -3100 39773
rect -3100 39739 -3066 39773
rect -3066 39739 -3028 39773
rect -3028 39739 -2994 39773
rect -2994 39739 -2956 39773
rect -2956 39739 -2922 39773
rect -2922 39739 -2884 39773
rect -2884 39739 -2850 39773
rect -2850 39739 -2812 39773
rect -2812 39739 -2778 39773
rect -2778 39739 -2740 39773
rect -2740 39739 -2706 39773
rect -2706 39739 -2668 39773
rect -2668 39739 -2634 39773
rect -2634 39739 -2596 39773
rect -2596 39739 -2562 39773
rect -2562 39739 -2524 39773
rect -2524 39739 -2490 39773
rect -2490 39739 -2452 39773
rect -2452 39739 -2418 39773
rect -2418 39739 -2380 39773
rect -2380 39739 -2346 39773
rect -2346 39739 -2308 39773
rect -2308 39739 -2274 39773
rect -2274 39739 -2236 39773
rect -2236 39739 -2202 39773
rect -2202 39739 -2164 39773
rect -2164 39739 -2130 39773
rect -2130 39739 -2092 39773
rect -2092 39739 -2058 39773
rect -2058 39739 -2020 39773
rect -2020 39739 -1986 39773
rect -1986 39739 -1948 39773
rect -1948 39739 -1914 39773
rect -1914 39739 -1876 39773
rect -1876 39739 -1842 39773
rect -1842 39739 -1804 39773
rect -1804 39739 -1770 39773
rect -1770 39739 -1732 39773
rect -1732 39739 -1698 39773
rect -1698 39739 -1660 39773
rect -1660 39739 -1626 39773
rect -1626 39739 -1588 39773
rect -1588 39739 -1554 39773
rect -1554 39739 -1516 39773
rect -1516 39739 -1482 39773
rect -1482 39739 -1444 39773
rect -1444 39739 -1410 39773
rect -1410 39739 -1372 39773
rect -1372 39739 -1338 39773
rect -1338 39739 -1300 39773
rect -1300 39739 -1266 39773
rect -1266 39739 -1228 39773
rect -1228 39739 -1194 39773
rect -1194 39739 -1156 39773
rect -1156 39739 -1122 39773
rect -1122 39739 -1084 39773
rect -1084 39739 -1050 39773
rect -1050 39739 -1012 39773
rect -1012 39739 -978 39773
rect -978 39739 -940 39773
rect -940 39739 -906 39773
rect -906 39739 -868 39773
rect -868 39739 -834 39773
rect -834 39739 -796 39773
rect -796 39739 -762 39773
rect -762 39739 -724 39773
rect -724 39739 -690 39773
rect -690 39739 -652 39773
rect -652 39739 -618 39773
rect -618 39739 -580 39773
rect -580 39739 -546 39773
rect -546 39739 -508 39773
rect -508 39739 -474 39773
rect -474 39739 -436 39773
rect -436 39739 -402 39773
rect -402 39739 -364 39773
rect -364 39739 -330 39773
rect -330 39739 -292 39773
rect -292 39739 -258 39773
rect -258 39739 -220 39773
rect -220 39739 -186 39773
rect -186 39739 -170 39773
rect -5662 39666 -170 39739
rect 361 45785 541 45843
rect 361 45751 410 45785
rect 410 45751 444 45785
rect 444 45751 541 45785
rect 361 45713 541 45751
rect 361 45679 410 45713
rect 410 45679 444 45713
rect 444 45679 541 45713
rect 361 45641 541 45679
rect 361 45607 410 45641
rect 410 45607 444 45641
rect 444 45607 541 45641
rect 361 45569 541 45607
rect 361 45535 410 45569
rect 410 45535 444 45569
rect 444 45535 541 45569
rect 361 45497 541 45535
rect 361 45463 410 45497
rect 410 45463 444 45497
rect 444 45463 541 45497
rect 361 45425 541 45463
rect 361 45391 410 45425
rect 410 45391 444 45425
rect 444 45391 541 45425
rect 361 45353 541 45391
rect 361 45319 410 45353
rect 410 45319 444 45353
rect 444 45319 541 45353
rect 361 45281 541 45319
rect 361 45247 410 45281
rect 410 45247 444 45281
rect 444 45247 541 45281
rect 361 45209 541 45247
rect 361 45175 410 45209
rect 410 45175 444 45209
rect 444 45175 541 45209
rect 361 45137 541 45175
rect 361 45103 410 45137
rect 410 45103 444 45137
rect 444 45103 541 45137
rect 361 45065 541 45103
rect 361 45031 410 45065
rect 410 45031 444 45065
rect 444 45031 541 45065
rect 361 44993 541 45031
rect 361 44959 410 44993
rect 410 44959 444 44993
rect 444 44959 541 44993
rect 361 44921 541 44959
rect 361 44887 410 44921
rect 410 44887 444 44921
rect 444 44887 541 44921
rect 361 44849 541 44887
rect 361 44815 410 44849
rect 410 44815 444 44849
rect 444 44815 541 44849
rect 361 44777 541 44815
rect 361 44743 410 44777
rect 410 44743 444 44777
rect 444 44743 541 44777
rect 361 44705 541 44743
rect 361 44671 410 44705
rect 410 44671 444 44705
rect 444 44671 541 44705
rect 361 44633 541 44671
rect 361 44599 410 44633
rect 410 44599 444 44633
rect 444 44599 541 44633
rect 361 44561 541 44599
rect 361 44527 410 44561
rect 410 44527 444 44561
rect 444 44527 541 44561
rect 361 44489 541 44527
rect 361 44455 410 44489
rect 410 44455 444 44489
rect 444 44455 541 44489
rect 361 44417 541 44455
rect 361 44383 410 44417
rect 410 44383 444 44417
rect 444 44383 541 44417
rect 361 44319 541 44383
rect 374 41326 490 41381
rect 374 41292 410 41326
rect 410 41292 444 41326
rect 444 41292 490 41326
rect 374 41254 490 41292
rect 374 41220 410 41254
rect 410 41220 444 41254
rect 444 41220 490 41254
rect 374 41182 490 41220
rect 374 41148 410 41182
rect 410 41148 444 41182
rect 444 41148 490 41182
rect 374 41110 490 41148
rect 374 41076 410 41110
rect 410 41076 444 41110
rect 444 41076 490 41110
rect 374 41038 490 41076
rect 374 41004 410 41038
rect 410 41004 444 41038
rect 444 41004 490 41038
rect 374 40966 490 41004
rect 374 40932 410 40966
rect 410 40932 444 40966
rect 444 40932 490 40966
rect 374 40894 490 40932
rect 374 40860 410 40894
rect 410 40860 444 40894
rect 444 40860 490 40894
rect 374 40822 490 40860
rect 374 40788 410 40822
rect 410 40788 444 40822
rect 444 40788 490 40822
rect 374 40750 490 40788
rect 374 40716 410 40750
rect 410 40716 444 40750
rect 444 40716 490 40750
rect 374 40678 490 40716
rect 374 40644 410 40678
rect 410 40644 444 40678
rect 444 40644 490 40678
rect 374 40606 490 40644
rect 374 40572 410 40606
rect 410 40572 444 40606
rect 444 40572 490 40606
rect 374 40534 490 40572
rect 374 40500 410 40534
rect 410 40500 444 40534
rect 444 40500 490 40534
rect 374 40462 490 40500
rect 374 40428 410 40462
rect 410 40428 444 40462
rect 444 40428 490 40462
rect 374 40390 490 40428
rect 374 40356 410 40390
rect 410 40356 444 40390
rect 444 40356 490 40390
rect 374 40318 490 40356
rect 374 40284 410 40318
rect 410 40284 444 40318
rect 444 40284 490 40318
rect 374 40246 490 40284
rect 374 40212 410 40246
rect 410 40212 444 40246
rect 444 40212 490 40246
rect 374 40174 490 40212
rect 374 40140 410 40174
rect 410 40140 444 40174
rect 444 40140 490 40174
rect 374 40102 490 40140
rect 374 40068 410 40102
rect 410 40068 444 40102
rect 444 40068 490 40102
rect 374 39857 490 40068
rect 2528 38799 2580 38851
rect 2528 38735 2580 38787
rect 2528 38671 2580 38723
rect 99 38508 151 38560
rect 1236 38508 1288 38560
rect 2632 38510 2684 38562
rect 5367 38510 5419 38562
rect 2538 38342 2590 38394
rect 2538 38278 2590 38330
rect 2538 38214 2590 38266
rect 2538 38150 2590 38202
rect 2538 38086 2590 38138
rect 5367 38097 5419 38149
rect 2538 38022 2590 38074
rect 99 37593 151 37645
rect 3433 37593 3485 37645
rect 2650 37149 2702 37201
rect 2174 37093 2226 37145
rect 2174 37029 2226 37081
rect 2174 36965 2226 37017
rect 2174 36901 2226 36953
rect 99 36758 151 36810
rect 889 36758 941 36810
rect 2175 36593 2227 36645
rect 2175 36529 2227 36581
rect 2175 36465 2227 36517
rect 2175 36401 2227 36453
rect 2175 36337 2227 36389
rect 2175 36273 2227 36325
rect 2954 36033 3006 36085
rect 3018 36033 3070 36085
rect 3082 36033 3134 36085
rect 3146 36033 3198 36085
rect 3210 36033 3262 36085
rect 3274 36033 3326 36085
rect 10211 39867 10519 46127
rect 17437 64686 17489 64738
rect 17437 64622 17489 64674
rect 17437 64558 17489 64610
rect 17437 64494 17489 64546
rect 17437 64430 17489 64482
rect 17437 64366 17489 64418
rect 17437 64302 17489 64354
rect 17437 64238 17489 64290
rect 17437 64174 17489 64226
rect 23965 64686 24017 64738
rect 23965 64622 24017 64674
rect 23965 64558 24017 64610
rect 23965 64494 24017 64546
rect 23965 64430 24017 64482
rect 23965 64366 24017 64418
rect 23965 64302 24017 64354
rect 23965 64238 24017 64290
rect 23965 64174 24017 64226
rect 31581 64686 31633 64738
rect 31581 64622 31633 64674
rect 31581 64558 31633 64610
rect 31581 64494 31633 64546
rect 31581 64430 31633 64482
rect 31581 64366 31633 64418
rect 31581 64302 31633 64354
rect 31581 64238 31633 64290
rect 31581 64174 31633 64226
rect 17982 62683 18034 62735
rect 17982 62619 18034 62671
rect 17982 62555 18034 62607
rect 17982 62491 18034 62543
rect 17982 62427 18034 62479
rect 17982 62363 18034 62415
rect 17982 62299 18034 62351
rect 17982 62235 18034 62287
rect 17982 62171 18034 62223
rect 19070 62683 19122 62735
rect 19070 62619 19122 62671
rect 19070 62555 19122 62607
rect 19070 62491 19122 62543
rect 19070 62427 19122 62479
rect 19070 62363 19122 62415
rect 19070 62299 19122 62351
rect 19070 62235 19122 62287
rect 19070 62171 19122 62223
rect 21246 62683 21298 62735
rect 21246 62619 21298 62671
rect 21246 62555 21298 62607
rect 21246 62491 21298 62543
rect 21246 62427 21298 62479
rect 21246 62363 21298 62415
rect 21246 62299 21298 62351
rect 21246 62235 21298 62287
rect 21246 62171 21298 62223
rect 22334 62683 22386 62735
rect 22334 62619 22386 62671
rect 22334 62555 22386 62607
rect 22334 62491 22386 62543
rect 22334 62427 22386 62479
rect 22334 62363 22386 62415
rect 22334 62299 22386 62351
rect 22334 62235 22386 62287
rect 22334 62171 22386 62223
rect 23422 62683 23474 62735
rect 23422 62619 23474 62671
rect 23422 62555 23474 62607
rect 23422 62491 23474 62543
rect 23422 62427 23474 62479
rect 23422 62363 23474 62415
rect 23422 62299 23474 62351
rect 23422 62235 23474 62287
rect 23422 62171 23474 62223
rect 24510 62683 24562 62735
rect 24510 62619 24562 62671
rect 24510 62555 24562 62607
rect 24510 62491 24562 62543
rect 24510 62427 24562 62479
rect 24510 62363 24562 62415
rect 24510 62299 24562 62351
rect 24510 62235 24562 62287
rect 24510 62171 24562 62223
rect 25598 62683 25650 62735
rect 25598 62619 25650 62671
rect 25598 62555 25650 62607
rect 25598 62491 25650 62543
rect 25598 62427 25650 62479
rect 25598 62363 25650 62415
rect 25598 62299 25650 62351
rect 25598 62235 25650 62287
rect 25598 62171 25650 62223
rect 26686 62683 26738 62735
rect 26686 62619 26738 62671
rect 26686 62555 26738 62607
rect 26686 62491 26738 62543
rect 26686 62427 26738 62479
rect 26686 62363 26738 62415
rect 26686 62299 26738 62351
rect 26686 62235 26738 62287
rect 26686 62171 26738 62223
rect 28862 62683 28914 62735
rect 28862 62619 28914 62671
rect 28862 62555 28914 62607
rect 28862 62491 28914 62543
rect 28862 62427 28914 62479
rect 28862 62363 28914 62415
rect 28862 62299 28914 62351
rect 28862 62235 28914 62287
rect 28862 62171 28914 62223
rect 29950 62683 30002 62735
rect 29950 62619 30002 62671
rect 29950 62555 30002 62607
rect 29950 62491 30002 62543
rect 29950 62427 30002 62479
rect 29950 62363 30002 62415
rect 29950 62299 30002 62351
rect 29950 62235 30002 62287
rect 29950 62171 30002 62223
rect 31038 62683 31090 62735
rect 31038 62619 31090 62671
rect 31038 62555 31090 62607
rect 31038 62491 31090 62543
rect 31038 62427 31090 62479
rect 31038 62363 31090 62415
rect 31038 62299 31090 62351
rect 31038 62235 31090 62287
rect 31038 62171 31090 62223
rect 17437 60686 17489 60738
rect 17437 60622 17489 60674
rect 17437 60558 17489 60610
rect 17437 60494 17489 60546
rect 17437 60430 17489 60482
rect 17437 60366 17489 60418
rect 17437 60302 17489 60354
rect 17437 60238 17489 60290
rect 17437 60174 17489 60226
rect 18525 60686 18577 60738
rect 18525 60622 18577 60674
rect 18525 60558 18577 60610
rect 18525 60494 18577 60546
rect 18525 60430 18577 60482
rect 18525 60366 18577 60418
rect 18525 60302 18577 60354
rect 18525 60238 18577 60290
rect 18525 60174 18577 60226
rect 19613 60686 19665 60738
rect 19613 60622 19665 60674
rect 19613 60558 19665 60610
rect 19613 60494 19665 60546
rect 19613 60430 19665 60482
rect 19613 60366 19665 60418
rect 19613 60302 19665 60354
rect 19613 60238 19665 60290
rect 19613 60174 19665 60226
rect 20701 60686 20753 60738
rect 20701 60622 20753 60674
rect 20701 60558 20753 60610
rect 20701 60494 20753 60546
rect 20701 60430 20753 60482
rect 20701 60366 20753 60418
rect 20701 60302 20753 60354
rect 20701 60238 20753 60290
rect 20701 60174 20753 60226
rect 21789 60686 21841 60738
rect 21789 60622 21841 60674
rect 21789 60558 21841 60610
rect 21789 60494 21841 60546
rect 21789 60430 21841 60482
rect 21789 60366 21841 60418
rect 21789 60302 21841 60354
rect 21789 60238 21841 60290
rect 21789 60174 21841 60226
rect 22877 60686 22929 60738
rect 22877 60622 22929 60674
rect 22877 60558 22929 60610
rect 22877 60494 22929 60546
rect 22877 60430 22929 60482
rect 22877 60366 22929 60418
rect 22877 60302 22929 60354
rect 22877 60238 22929 60290
rect 22877 60174 22929 60226
rect 23965 60686 24017 60738
rect 23965 60622 24017 60674
rect 23965 60558 24017 60610
rect 23965 60494 24017 60546
rect 23965 60430 24017 60482
rect 23965 60366 24017 60418
rect 23965 60302 24017 60354
rect 23965 60238 24017 60290
rect 23965 60174 24017 60226
rect 25053 60686 25105 60738
rect 25053 60622 25105 60674
rect 25053 60558 25105 60610
rect 25053 60494 25105 60546
rect 25053 60430 25105 60482
rect 25053 60366 25105 60418
rect 25053 60302 25105 60354
rect 25053 60238 25105 60290
rect 25053 60174 25105 60226
rect 26141 60686 26193 60738
rect 26141 60622 26193 60674
rect 26141 60558 26193 60610
rect 26141 60494 26193 60546
rect 26141 60430 26193 60482
rect 26141 60366 26193 60418
rect 26141 60302 26193 60354
rect 26141 60238 26193 60290
rect 26141 60174 26193 60226
rect 27229 60686 27281 60738
rect 27229 60622 27281 60674
rect 27229 60558 27281 60610
rect 27229 60494 27281 60546
rect 27229 60430 27281 60482
rect 27229 60366 27281 60418
rect 27229 60302 27281 60354
rect 27229 60238 27281 60290
rect 27229 60174 27281 60226
rect 28317 60686 28369 60738
rect 28317 60622 28369 60674
rect 28317 60558 28369 60610
rect 28317 60494 28369 60546
rect 28317 60430 28369 60482
rect 28317 60366 28369 60418
rect 28317 60302 28369 60354
rect 28317 60238 28369 60290
rect 28317 60174 28369 60226
rect 29405 60686 29457 60738
rect 29405 60622 29457 60674
rect 29405 60558 29457 60610
rect 29405 60494 29457 60546
rect 29405 60430 29457 60482
rect 29405 60366 29457 60418
rect 29405 60302 29457 60354
rect 29405 60238 29457 60290
rect 29405 60174 29457 60226
rect 30493 60686 30545 60738
rect 30493 60622 30545 60674
rect 30493 60558 30545 60610
rect 30493 60494 30545 60546
rect 30493 60430 30545 60482
rect 30493 60366 30545 60418
rect 30493 60302 30545 60354
rect 30493 60238 30545 60290
rect 30493 60174 30545 60226
rect 31581 60686 31633 60738
rect 31581 60622 31633 60674
rect 31581 60558 31633 60610
rect 31581 60494 31633 60546
rect 31581 60430 31633 60482
rect 31581 60366 31633 60418
rect 31581 60302 31633 60354
rect 31581 60238 31633 60290
rect 31581 60174 31633 60226
rect 17982 58683 18034 58735
rect 17982 58619 18034 58671
rect 17982 58555 18034 58607
rect 17982 58491 18034 58543
rect 17982 58427 18034 58479
rect 17982 58363 18034 58415
rect 17982 58299 18034 58351
rect 17982 58235 18034 58287
rect 17982 58171 18034 58223
rect 19070 58683 19122 58735
rect 19070 58619 19122 58671
rect 19070 58555 19122 58607
rect 19070 58491 19122 58543
rect 19070 58427 19122 58479
rect 19070 58363 19122 58415
rect 19070 58299 19122 58351
rect 19070 58235 19122 58287
rect 19070 58171 19122 58223
rect 20158 58683 20210 58735
rect 20158 58619 20210 58671
rect 20158 58555 20210 58607
rect 20158 58491 20210 58543
rect 20158 58427 20210 58479
rect 20158 58363 20210 58415
rect 20158 58299 20210 58351
rect 20158 58235 20210 58287
rect 20158 58171 20210 58223
rect 21246 58683 21298 58735
rect 21246 58619 21298 58671
rect 21246 58555 21298 58607
rect 21246 58491 21298 58543
rect 21246 58427 21298 58479
rect 21246 58363 21298 58415
rect 21246 58299 21298 58351
rect 21246 58235 21298 58287
rect 21246 58171 21298 58223
rect 22334 58683 22386 58735
rect 22334 58619 22386 58671
rect 22334 58555 22386 58607
rect 22334 58491 22386 58543
rect 22334 58427 22386 58479
rect 22334 58363 22386 58415
rect 22334 58299 22386 58351
rect 22334 58235 22386 58287
rect 22334 58171 22386 58223
rect 23422 58683 23474 58735
rect 23422 58619 23474 58671
rect 23422 58555 23474 58607
rect 23422 58491 23474 58543
rect 23422 58427 23474 58479
rect 23422 58363 23474 58415
rect 23422 58299 23474 58351
rect 23422 58235 23474 58287
rect 23422 58171 23474 58223
rect 24510 58683 24562 58735
rect 24510 58619 24562 58671
rect 24510 58555 24562 58607
rect 24510 58491 24562 58543
rect 24510 58427 24562 58479
rect 24510 58363 24562 58415
rect 24510 58299 24562 58351
rect 24510 58235 24562 58287
rect 24510 58171 24562 58223
rect 25598 58683 25650 58735
rect 25598 58619 25650 58671
rect 25598 58555 25650 58607
rect 25598 58491 25650 58543
rect 25598 58427 25650 58479
rect 25598 58363 25650 58415
rect 25598 58299 25650 58351
rect 25598 58235 25650 58287
rect 25598 58171 25650 58223
rect 26686 58683 26738 58735
rect 26686 58619 26738 58671
rect 26686 58555 26738 58607
rect 26686 58491 26738 58543
rect 26686 58427 26738 58479
rect 26686 58363 26738 58415
rect 26686 58299 26738 58351
rect 26686 58235 26738 58287
rect 26686 58171 26738 58223
rect 27774 58683 27826 58735
rect 27774 58619 27826 58671
rect 27774 58555 27826 58607
rect 27774 58491 27826 58543
rect 27774 58427 27826 58479
rect 27774 58363 27826 58415
rect 27774 58299 27826 58351
rect 27774 58235 27826 58287
rect 27774 58171 27826 58223
rect 28862 58683 28914 58735
rect 28862 58619 28914 58671
rect 28862 58555 28914 58607
rect 28862 58491 28914 58543
rect 28862 58427 28914 58479
rect 28862 58363 28914 58415
rect 28862 58299 28914 58351
rect 28862 58235 28914 58287
rect 28862 58171 28914 58223
rect 29950 58683 30002 58735
rect 29950 58619 30002 58671
rect 29950 58555 30002 58607
rect 29950 58491 30002 58543
rect 29950 58427 30002 58479
rect 29950 58363 30002 58415
rect 29950 58299 30002 58351
rect 29950 58235 30002 58287
rect 29950 58171 30002 58223
rect 31038 58683 31090 58735
rect 31038 58619 31090 58671
rect 31038 58555 31090 58607
rect 31038 58491 31090 58543
rect 31038 58427 31090 58479
rect 31038 58363 31090 58415
rect 31038 58299 31090 58351
rect 31038 58235 31090 58287
rect 31038 58171 31090 58223
rect 17437 56686 17489 56738
rect 17437 56622 17489 56674
rect 17437 56558 17489 56610
rect 17437 56494 17489 56546
rect 17437 56430 17489 56482
rect 17437 56366 17489 56418
rect 17437 56302 17489 56354
rect 17437 56238 17489 56290
rect 17437 56174 17489 56226
rect 18525 56686 18577 56738
rect 18525 56622 18577 56674
rect 18525 56558 18577 56610
rect 18525 56494 18577 56546
rect 18525 56430 18577 56482
rect 18525 56366 18577 56418
rect 18525 56302 18577 56354
rect 18525 56238 18577 56290
rect 18525 56174 18577 56226
rect 19613 56686 19665 56738
rect 19613 56622 19665 56674
rect 19613 56558 19665 56610
rect 19613 56494 19665 56546
rect 19613 56430 19665 56482
rect 19613 56366 19665 56418
rect 19613 56302 19665 56354
rect 19613 56238 19665 56290
rect 19613 56174 19665 56226
rect 20701 56686 20753 56738
rect 20701 56622 20753 56674
rect 20701 56558 20753 56610
rect 20701 56494 20753 56546
rect 20701 56430 20753 56482
rect 20701 56366 20753 56418
rect 20701 56302 20753 56354
rect 20701 56238 20753 56290
rect 20701 56174 20753 56226
rect 21789 56686 21841 56738
rect 21789 56622 21841 56674
rect 21789 56558 21841 56610
rect 21789 56494 21841 56546
rect 21789 56430 21841 56482
rect 21789 56366 21841 56418
rect 21789 56302 21841 56354
rect 21789 56238 21841 56290
rect 21789 56174 21841 56226
rect 22877 56686 22929 56738
rect 22877 56622 22929 56674
rect 22877 56558 22929 56610
rect 22877 56494 22929 56546
rect 22877 56430 22929 56482
rect 22877 56366 22929 56418
rect 22877 56302 22929 56354
rect 22877 56238 22929 56290
rect 22877 56174 22929 56226
rect 23965 56686 24017 56738
rect 23965 56622 24017 56674
rect 23965 56558 24017 56610
rect 23965 56494 24017 56546
rect 23965 56430 24017 56482
rect 23965 56366 24017 56418
rect 23965 56302 24017 56354
rect 23965 56238 24017 56290
rect 23965 56174 24017 56226
rect 25053 56686 25105 56738
rect 25053 56622 25105 56674
rect 25053 56558 25105 56610
rect 25053 56494 25105 56546
rect 25053 56430 25105 56482
rect 25053 56366 25105 56418
rect 25053 56302 25105 56354
rect 25053 56238 25105 56290
rect 25053 56174 25105 56226
rect 26141 56686 26193 56738
rect 26141 56622 26193 56674
rect 26141 56558 26193 56610
rect 26141 56494 26193 56546
rect 26141 56430 26193 56482
rect 26141 56366 26193 56418
rect 26141 56302 26193 56354
rect 26141 56238 26193 56290
rect 26141 56174 26193 56226
rect 27229 56686 27281 56738
rect 27229 56622 27281 56674
rect 27229 56558 27281 56610
rect 27229 56494 27281 56546
rect 27229 56430 27281 56482
rect 27229 56366 27281 56418
rect 27229 56302 27281 56354
rect 27229 56238 27281 56290
rect 27229 56174 27281 56226
rect 28317 56686 28369 56738
rect 28317 56622 28369 56674
rect 28317 56558 28369 56610
rect 28317 56494 28369 56546
rect 28317 56430 28369 56482
rect 28317 56366 28369 56418
rect 28317 56302 28369 56354
rect 28317 56238 28369 56290
rect 28317 56174 28369 56226
rect 29405 56686 29457 56738
rect 29405 56622 29457 56674
rect 29405 56558 29457 56610
rect 29405 56494 29457 56546
rect 29405 56430 29457 56482
rect 29405 56366 29457 56418
rect 29405 56302 29457 56354
rect 29405 56238 29457 56290
rect 29405 56174 29457 56226
rect 30493 56686 30545 56738
rect 30493 56622 30545 56674
rect 30493 56558 30545 56610
rect 30493 56494 30545 56546
rect 30493 56430 30545 56482
rect 30493 56366 30545 56418
rect 30493 56302 30545 56354
rect 30493 56238 30545 56290
rect 30493 56174 30545 56226
rect 31581 56686 31633 56738
rect 31581 56622 31633 56674
rect 31581 56558 31633 56610
rect 31581 56494 31633 56546
rect 31581 56430 31633 56482
rect 31581 56366 31633 56418
rect 31581 56302 31633 56354
rect 31581 56238 31633 56290
rect 31581 56174 31633 56226
rect 17982 54683 18034 54735
rect 17982 54619 18034 54671
rect 17982 54555 18034 54607
rect 17982 54491 18034 54543
rect 17982 54427 18034 54479
rect 17982 54363 18034 54415
rect 17982 54299 18034 54351
rect 17982 54235 18034 54287
rect 17982 54171 18034 54223
rect 19070 54683 19122 54735
rect 19070 54619 19122 54671
rect 19070 54555 19122 54607
rect 19070 54491 19122 54543
rect 19070 54427 19122 54479
rect 19070 54363 19122 54415
rect 19070 54299 19122 54351
rect 19070 54235 19122 54287
rect 19070 54171 19122 54223
rect 20158 54683 20210 54735
rect 20158 54619 20210 54671
rect 20158 54555 20210 54607
rect 20158 54491 20210 54543
rect 20158 54427 20210 54479
rect 20158 54363 20210 54415
rect 20158 54299 20210 54351
rect 20158 54235 20210 54287
rect 20158 54171 20210 54223
rect 21246 54683 21298 54735
rect 21246 54619 21298 54671
rect 21246 54555 21298 54607
rect 21246 54491 21298 54543
rect 21246 54427 21298 54479
rect 21246 54363 21298 54415
rect 21246 54299 21298 54351
rect 21246 54235 21298 54287
rect 21246 54171 21298 54223
rect 22334 54683 22386 54735
rect 22334 54619 22386 54671
rect 22334 54555 22386 54607
rect 22334 54491 22386 54543
rect 22334 54427 22386 54479
rect 22334 54363 22386 54415
rect 22334 54299 22386 54351
rect 22334 54235 22386 54287
rect 22334 54171 22386 54223
rect 23422 54683 23474 54735
rect 23422 54619 23474 54671
rect 23422 54555 23474 54607
rect 23422 54491 23474 54543
rect 23422 54427 23474 54479
rect 23422 54363 23474 54415
rect 23422 54299 23474 54351
rect 23422 54235 23474 54287
rect 23422 54171 23474 54223
rect 24510 54683 24562 54735
rect 24510 54619 24562 54671
rect 24510 54555 24562 54607
rect 24510 54491 24562 54543
rect 24510 54427 24562 54479
rect 24510 54363 24562 54415
rect 24510 54299 24562 54351
rect 24510 54235 24562 54287
rect 24510 54171 24562 54223
rect 25598 54683 25650 54735
rect 25598 54619 25650 54671
rect 25598 54555 25650 54607
rect 25598 54491 25650 54543
rect 25598 54427 25650 54479
rect 25598 54363 25650 54415
rect 25598 54299 25650 54351
rect 25598 54235 25650 54287
rect 25598 54171 25650 54223
rect 26686 54683 26738 54735
rect 26686 54619 26738 54671
rect 26686 54555 26738 54607
rect 26686 54491 26738 54543
rect 26686 54427 26738 54479
rect 26686 54363 26738 54415
rect 26686 54299 26738 54351
rect 26686 54235 26738 54287
rect 26686 54171 26738 54223
rect 27774 54683 27826 54735
rect 27774 54619 27826 54671
rect 27774 54555 27826 54607
rect 27774 54491 27826 54543
rect 27774 54427 27826 54479
rect 27774 54363 27826 54415
rect 27774 54299 27826 54351
rect 27774 54235 27826 54287
rect 27774 54171 27826 54223
rect 28862 54683 28914 54735
rect 28862 54619 28914 54671
rect 28862 54555 28914 54607
rect 28862 54491 28914 54543
rect 28862 54427 28914 54479
rect 28862 54363 28914 54415
rect 28862 54299 28914 54351
rect 28862 54235 28914 54287
rect 28862 54171 28914 54223
rect 29950 54683 30002 54735
rect 29950 54619 30002 54671
rect 29950 54555 30002 54607
rect 29950 54491 30002 54543
rect 29950 54427 30002 54479
rect 29950 54363 30002 54415
rect 29950 54299 30002 54351
rect 29950 54235 30002 54287
rect 29950 54171 30002 54223
rect 31038 54683 31090 54735
rect 31038 54619 31090 54671
rect 31038 54555 31090 54607
rect 31038 54491 31090 54543
rect 31038 54427 31090 54479
rect 31038 54363 31090 54415
rect 31038 54299 31090 54351
rect 31038 54235 31090 54287
rect 31038 54171 31090 54223
rect 17437 52686 17489 52738
rect 17437 52622 17489 52674
rect 17437 52558 17489 52610
rect 17437 52494 17489 52546
rect 17437 52430 17489 52482
rect 17437 52366 17489 52418
rect 17437 52302 17489 52354
rect 17437 52238 17489 52290
rect 17437 52174 17489 52226
rect 18525 52686 18577 52738
rect 18525 52622 18577 52674
rect 18525 52558 18577 52610
rect 18525 52494 18577 52546
rect 18525 52430 18577 52482
rect 18525 52366 18577 52418
rect 18525 52302 18577 52354
rect 18525 52238 18577 52290
rect 18525 52174 18577 52226
rect 19613 52686 19665 52738
rect 19613 52622 19665 52674
rect 19613 52558 19665 52610
rect 19613 52494 19665 52546
rect 19613 52430 19665 52482
rect 19613 52366 19665 52418
rect 19613 52302 19665 52354
rect 19613 52238 19665 52290
rect 19613 52174 19665 52226
rect 20701 52686 20753 52738
rect 20701 52622 20753 52674
rect 20701 52558 20753 52610
rect 20701 52494 20753 52546
rect 20701 52430 20753 52482
rect 20701 52366 20753 52418
rect 20701 52302 20753 52354
rect 20701 52238 20753 52290
rect 20701 52174 20753 52226
rect 21789 52686 21841 52738
rect 21789 52622 21841 52674
rect 21789 52558 21841 52610
rect 21789 52494 21841 52546
rect 21789 52430 21841 52482
rect 21789 52366 21841 52418
rect 21789 52302 21841 52354
rect 21789 52238 21841 52290
rect 21789 52174 21841 52226
rect 22877 52686 22929 52738
rect 22877 52622 22929 52674
rect 22877 52558 22929 52610
rect 22877 52494 22929 52546
rect 22877 52430 22929 52482
rect 22877 52366 22929 52418
rect 22877 52302 22929 52354
rect 22877 52238 22929 52290
rect 22877 52174 22929 52226
rect 23965 52686 24017 52738
rect 23965 52622 24017 52674
rect 23965 52558 24017 52610
rect 23965 52494 24017 52546
rect 23965 52430 24017 52482
rect 23965 52366 24017 52418
rect 23965 52302 24017 52354
rect 23965 52238 24017 52290
rect 23965 52174 24017 52226
rect 25053 52686 25105 52738
rect 25053 52622 25105 52674
rect 25053 52558 25105 52610
rect 25053 52494 25105 52546
rect 25053 52430 25105 52482
rect 25053 52366 25105 52418
rect 25053 52302 25105 52354
rect 25053 52238 25105 52290
rect 25053 52174 25105 52226
rect 26141 52686 26193 52738
rect 26141 52622 26193 52674
rect 26141 52558 26193 52610
rect 26141 52494 26193 52546
rect 26141 52430 26193 52482
rect 26141 52366 26193 52418
rect 26141 52302 26193 52354
rect 26141 52238 26193 52290
rect 26141 52174 26193 52226
rect 27229 52686 27281 52738
rect 27229 52622 27281 52674
rect 27229 52558 27281 52610
rect 27229 52494 27281 52546
rect 27229 52430 27281 52482
rect 27229 52366 27281 52418
rect 27229 52302 27281 52354
rect 27229 52238 27281 52290
rect 27229 52174 27281 52226
rect 28317 52686 28369 52738
rect 28317 52622 28369 52674
rect 28317 52558 28369 52610
rect 28317 52494 28369 52546
rect 28317 52430 28369 52482
rect 28317 52366 28369 52418
rect 28317 52302 28369 52354
rect 28317 52238 28369 52290
rect 28317 52174 28369 52226
rect 29405 52686 29457 52738
rect 29405 52622 29457 52674
rect 29405 52558 29457 52610
rect 29405 52494 29457 52546
rect 29405 52430 29457 52482
rect 29405 52366 29457 52418
rect 29405 52302 29457 52354
rect 29405 52238 29457 52290
rect 29405 52174 29457 52226
rect 30493 52686 30545 52738
rect 30493 52622 30545 52674
rect 30493 52558 30545 52610
rect 30493 52494 30545 52546
rect 30493 52430 30545 52482
rect 30493 52366 30545 52418
rect 30493 52302 30545 52354
rect 30493 52238 30545 52290
rect 30493 52174 30545 52226
rect 31581 52686 31633 52738
rect 31581 52622 31633 52674
rect 31581 52558 31633 52610
rect 31581 52494 31633 52546
rect 31581 52430 31633 52482
rect 31581 52366 31633 52418
rect 31581 52302 31633 52354
rect 31581 52238 31633 52290
rect 31581 52174 31633 52226
rect 17982 50683 18034 50735
rect 17982 50619 18034 50671
rect 17982 50555 18034 50607
rect 17982 50491 18034 50543
rect 17982 50427 18034 50479
rect 17982 50363 18034 50415
rect 17982 50299 18034 50351
rect 17982 50235 18034 50287
rect 17982 50171 18034 50223
rect 20158 50683 20210 50735
rect 20158 50619 20210 50671
rect 20158 50555 20210 50607
rect 20158 50491 20210 50543
rect 20158 50427 20210 50479
rect 20158 50363 20210 50415
rect 20158 50299 20210 50351
rect 20158 50235 20210 50287
rect 20158 50171 20210 50223
rect 21246 50683 21298 50735
rect 21246 50619 21298 50671
rect 21246 50555 21298 50607
rect 21246 50491 21298 50543
rect 21246 50427 21298 50479
rect 21246 50363 21298 50415
rect 21246 50299 21298 50351
rect 21246 50235 21298 50287
rect 21246 50171 21298 50223
rect 23422 50683 23474 50735
rect 23422 50619 23474 50671
rect 23422 50555 23474 50607
rect 23422 50491 23474 50543
rect 23422 50427 23474 50479
rect 23422 50363 23474 50415
rect 23422 50299 23474 50351
rect 23422 50235 23474 50287
rect 23422 50171 23474 50223
rect 24510 50683 24562 50735
rect 24510 50619 24562 50671
rect 24510 50555 24562 50607
rect 24510 50491 24562 50543
rect 24510 50427 24562 50479
rect 24510 50363 24562 50415
rect 24510 50299 24562 50351
rect 24510 50235 24562 50287
rect 24510 50171 24562 50223
rect 25598 50683 25650 50735
rect 25598 50619 25650 50671
rect 25598 50555 25650 50607
rect 25598 50491 25650 50543
rect 25598 50427 25650 50479
rect 25598 50363 25650 50415
rect 25598 50299 25650 50351
rect 25598 50235 25650 50287
rect 25598 50171 25650 50223
rect 27774 50683 27826 50735
rect 27774 50619 27826 50671
rect 27774 50555 27826 50607
rect 27774 50491 27826 50543
rect 27774 50427 27826 50479
rect 27774 50363 27826 50415
rect 27774 50299 27826 50351
rect 27774 50235 27826 50287
rect 27774 50171 27826 50223
rect 28862 50683 28914 50735
rect 28862 50619 28914 50671
rect 28862 50555 28914 50607
rect 28862 50491 28914 50543
rect 28862 50427 28914 50479
rect 28862 50363 28914 50415
rect 28862 50299 28914 50351
rect 28862 50235 28914 50287
rect 28862 50171 28914 50223
rect 31038 50683 31090 50735
rect 31038 50619 31090 50671
rect 31038 50555 31090 50607
rect 31038 50491 31090 50543
rect 31038 50427 31090 50479
rect 31038 50363 31090 50415
rect 31038 50299 31090 50351
rect 31038 50235 31090 50287
rect 31038 50171 31090 50223
rect 17437 48686 17489 48738
rect 17437 48622 17489 48674
rect 17437 48558 17489 48610
rect 17437 48494 17489 48546
rect 17437 48430 17489 48482
rect 17437 48366 17489 48418
rect 17437 48302 17489 48354
rect 17437 48238 17489 48290
rect 17437 48174 17489 48226
rect 18525 48686 18577 48738
rect 18525 48622 18577 48674
rect 18525 48558 18577 48610
rect 18525 48494 18577 48546
rect 18525 48430 18577 48482
rect 18525 48366 18577 48418
rect 18525 48302 18577 48354
rect 18525 48238 18577 48290
rect 18525 48174 18577 48226
rect 19613 48686 19665 48738
rect 19613 48622 19665 48674
rect 19613 48558 19665 48610
rect 19613 48494 19665 48546
rect 19613 48430 19665 48482
rect 19613 48366 19665 48418
rect 19613 48302 19665 48354
rect 19613 48238 19665 48290
rect 19613 48174 19665 48226
rect 20701 48686 20753 48738
rect 20701 48622 20753 48674
rect 20701 48558 20753 48610
rect 20701 48494 20753 48546
rect 20701 48430 20753 48482
rect 20701 48366 20753 48418
rect 20701 48302 20753 48354
rect 20701 48238 20753 48290
rect 20701 48174 20753 48226
rect 21789 48686 21841 48738
rect 21789 48622 21841 48674
rect 21789 48558 21841 48610
rect 21789 48494 21841 48546
rect 21789 48430 21841 48482
rect 21789 48366 21841 48418
rect 21789 48302 21841 48354
rect 21789 48238 21841 48290
rect 21789 48174 21841 48226
rect 22877 48686 22929 48738
rect 22877 48622 22929 48674
rect 22877 48558 22929 48610
rect 22877 48494 22929 48546
rect 22877 48430 22929 48482
rect 22877 48366 22929 48418
rect 22877 48302 22929 48354
rect 22877 48238 22929 48290
rect 22877 48174 22929 48226
rect 23965 48686 24017 48738
rect 23965 48622 24017 48674
rect 23965 48558 24017 48610
rect 23965 48494 24017 48546
rect 23965 48430 24017 48482
rect 23965 48366 24017 48418
rect 23965 48302 24017 48354
rect 23965 48238 24017 48290
rect 23965 48174 24017 48226
rect 29405 48686 29457 48738
rect 29405 48622 29457 48674
rect 29405 48558 29457 48610
rect 29405 48494 29457 48546
rect 29405 48430 29457 48482
rect 29405 48366 29457 48418
rect 29405 48302 29457 48354
rect 29405 48238 29457 48290
rect 29405 48174 29457 48226
rect 30493 48686 30545 48738
rect 30493 48622 30545 48674
rect 30493 48558 30545 48610
rect 30493 48494 30545 48546
rect 30493 48430 30545 48482
rect 30493 48366 30545 48418
rect 30493 48302 30545 48354
rect 30493 48238 30545 48290
rect 30493 48174 30545 48226
rect 31581 48686 31633 48738
rect 31581 48622 31633 48674
rect 31581 48558 31633 48610
rect 31581 48494 31633 48546
rect 31581 48430 31633 48482
rect 31581 48366 31633 48418
rect 31581 48302 31633 48354
rect 31581 48238 31633 48290
rect 31581 48174 31633 48226
rect 17982 46683 18034 46735
rect 17982 46619 18034 46671
rect 17982 46555 18034 46607
rect 17982 46491 18034 46543
rect 17982 46427 18034 46479
rect 17982 46363 18034 46415
rect 17982 46299 18034 46351
rect 17982 46235 18034 46287
rect 17982 46171 18034 46223
rect 19070 46683 19122 46735
rect 19070 46619 19122 46671
rect 19070 46555 19122 46607
rect 19070 46491 19122 46543
rect 19070 46427 19122 46479
rect 19070 46363 19122 46415
rect 19070 46299 19122 46351
rect 19070 46235 19122 46287
rect 19070 46171 19122 46223
rect 20158 46683 20210 46735
rect 20158 46619 20210 46671
rect 20158 46555 20210 46607
rect 20158 46491 20210 46543
rect 20158 46427 20210 46479
rect 20158 46363 20210 46415
rect 20158 46299 20210 46351
rect 20158 46235 20210 46287
rect 20158 46171 20210 46223
rect 21246 46683 21298 46735
rect 21246 46619 21298 46671
rect 21246 46555 21298 46607
rect 21246 46491 21298 46543
rect 21246 46427 21298 46479
rect 21246 46363 21298 46415
rect 21246 46299 21298 46351
rect 21246 46235 21298 46287
rect 21246 46171 21298 46223
rect 22334 46683 22386 46735
rect 22334 46619 22386 46671
rect 22334 46555 22386 46607
rect 22334 46491 22386 46543
rect 22334 46427 22386 46479
rect 22334 46363 22386 46415
rect 22334 46299 22386 46351
rect 22334 46235 22386 46287
rect 22334 46171 22386 46223
rect 24510 46683 24562 46735
rect 24510 46619 24562 46671
rect 24510 46555 24562 46607
rect 24510 46491 24562 46543
rect 24510 46427 24562 46479
rect 24510 46363 24562 46415
rect 24510 46299 24562 46351
rect 24510 46235 24562 46287
rect 24510 46171 24562 46223
rect 25598 46683 25650 46735
rect 25598 46619 25650 46671
rect 25598 46555 25650 46607
rect 25598 46491 25650 46543
rect 25598 46427 25650 46479
rect 25598 46363 25650 46415
rect 25598 46299 25650 46351
rect 25598 46235 25650 46287
rect 25598 46171 25650 46223
rect 26686 46683 26738 46735
rect 26686 46619 26738 46671
rect 26686 46555 26738 46607
rect 26686 46491 26738 46543
rect 26686 46427 26738 46479
rect 26686 46363 26738 46415
rect 26686 46299 26738 46351
rect 26686 46235 26738 46287
rect 26686 46171 26738 46223
rect 27774 46683 27826 46735
rect 27774 46619 27826 46671
rect 27774 46555 27826 46607
rect 27774 46491 27826 46543
rect 27774 46427 27826 46479
rect 27774 46363 27826 46415
rect 27774 46299 27826 46351
rect 27774 46235 27826 46287
rect 27774 46171 27826 46223
rect 28862 46683 28914 46735
rect 28862 46619 28914 46671
rect 28862 46555 28914 46607
rect 28862 46491 28914 46543
rect 28862 46427 28914 46479
rect 28862 46363 28914 46415
rect 28862 46299 28914 46351
rect 28862 46235 28914 46287
rect 28862 46171 28914 46223
rect 29950 46683 30002 46735
rect 29950 46619 30002 46671
rect 29950 46555 30002 46607
rect 29950 46491 30002 46543
rect 29950 46427 30002 46479
rect 29950 46363 30002 46415
rect 29950 46299 30002 46351
rect 29950 46235 30002 46287
rect 29950 46171 30002 46223
rect 31038 46683 31090 46735
rect 31038 46619 31090 46671
rect 31038 46555 31090 46607
rect 31038 46491 31090 46543
rect 31038 46427 31090 46479
rect 31038 46363 31090 46415
rect 31038 46299 31090 46351
rect 31038 46235 31090 46287
rect 31038 46171 31090 46223
rect 18251 45690 18303 45742
rect 18797 45690 18849 45742
rect 19343 45681 19395 45733
rect 19888 45680 19940 45732
rect 21519 45668 21571 45720
rect 22062 45665 22114 45717
rect 22604 45664 22656 45716
rect 23151 45669 23203 45721
rect 25869 45680 25921 45732
rect 26412 45684 26464 45736
rect 26954 45678 27006 45730
rect 27511 45669 27563 45721
rect 29135 45680 29187 45732
rect 29679 45673 29731 45725
rect 30229 45677 30281 45729
rect 30762 45677 30814 45729
rect 44780 45014 44832 45066
rect 44844 45014 44896 45066
rect 44908 45014 44960 45066
rect 44972 45014 45024 45066
rect 45036 45014 45088 45066
rect 45100 45014 45152 45066
rect 45164 45014 45216 45066
rect 45228 45014 45280 45066
rect 39563 44833 39615 44885
rect 40595 44816 40647 44830
rect 40595 44782 40603 44816
rect 40603 44782 40637 44816
rect 40637 44782 40647 44816
rect 40595 44778 40647 44782
rect 40995 44810 41047 44819
rect 40995 44776 41005 44810
rect 41005 44776 41039 44810
rect 41039 44776 41047 44810
rect 40995 44767 41047 44776
rect 41152 44816 41204 44823
rect 41152 44782 41161 44816
rect 41161 44782 41195 44816
rect 41195 44782 41204 44816
rect 41152 44771 41204 44782
rect 40894 44751 40946 44762
rect 40894 44717 40905 44751
rect 40905 44717 40939 44751
rect 40939 44717 40946 44751
rect 40894 44710 40946 44717
rect 39563 44643 39615 44695
rect 46322 44731 46502 44911
rect 41541 44468 41593 44520
rect 41605 44468 41657 44520
rect 41669 44468 41721 44520
rect 41733 44468 41785 44520
rect 41797 44468 41849 44520
rect 44779 43863 44831 43915
rect 44843 43863 44895 43915
rect 44907 43863 44959 43915
rect 44971 43863 45023 43915
rect 45035 43863 45087 43915
rect 45099 43863 45151 43915
rect 45163 43863 45215 43915
rect 45227 43863 45279 43915
rect 39563 43683 39615 43735
rect 40595 43666 40647 43680
rect 40595 43632 40603 43666
rect 40603 43632 40637 43666
rect 40637 43632 40647 43666
rect 40595 43628 40647 43632
rect 40995 43660 41047 43669
rect 40995 43626 41005 43660
rect 41005 43626 41039 43660
rect 41039 43626 41047 43660
rect 40995 43617 41047 43626
rect 41152 43666 41204 43673
rect 41152 43632 41161 43666
rect 41161 43632 41195 43666
rect 41195 43632 41204 43666
rect 41152 43621 41204 43632
rect 40894 43601 40946 43612
rect 40894 43567 40905 43601
rect 40905 43567 40939 43601
rect 40939 43567 40946 43601
rect 40894 43560 40946 43567
rect 39563 43493 39615 43545
rect 46310 43580 46490 43760
rect 41539 43318 41591 43370
rect 41603 43318 41655 43370
rect 41667 43318 41719 43370
rect 41731 43318 41783 43370
rect 41795 43318 41847 43370
rect 44769 41321 44821 41373
rect 44833 41321 44885 41373
rect 44897 41321 44949 41373
rect 44961 41321 45013 41373
rect 45025 41321 45077 41373
rect 45089 41321 45141 41373
rect 45153 41321 45205 41373
rect 45217 41321 45269 41373
rect 39563 41143 39615 41195
rect 40595 41126 40647 41140
rect 40595 41092 40603 41126
rect 40603 41092 40637 41126
rect 40637 41092 40647 41126
rect 40595 41088 40647 41092
rect 40995 41120 41047 41129
rect 40995 41086 41005 41120
rect 41005 41086 41039 41120
rect 41039 41086 41047 41120
rect 40995 41077 41047 41086
rect 41152 41126 41204 41133
rect 41152 41092 41161 41126
rect 41161 41092 41195 41126
rect 41195 41092 41204 41126
rect 41152 41081 41204 41092
rect 40894 41061 40946 41072
rect 40894 41027 40905 41061
rect 40905 41027 40939 41061
rect 40939 41027 40946 41061
rect 40894 41020 40946 41027
rect 39563 40953 39615 41005
rect 46168 41048 46348 41228
rect 41457 40777 41509 40829
rect 41521 40777 41573 40829
rect 41585 40777 41637 40829
rect 41649 40777 41701 40829
rect 41713 40777 41765 40829
rect 44769 40051 44821 40103
rect 44833 40051 44885 40103
rect 44897 40051 44949 40103
rect 44961 40051 45013 40103
rect 45025 40051 45077 40103
rect 45089 40051 45141 40103
rect 45153 40051 45205 40103
rect 45217 40051 45269 40103
rect 39563 39873 39615 39925
rect 40595 39856 40647 39870
rect 40595 39822 40603 39856
rect 40603 39822 40637 39856
rect 40637 39822 40647 39856
rect 40595 39818 40647 39822
rect 40995 39850 41047 39859
rect 40995 39816 41005 39850
rect 41005 39816 41039 39850
rect 41039 39816 41047 39850
rect 40995 39807 41047 39816
rect 41152 39856 41204 39863
rect 41152 39822 41161 39856
rect 41161 39822 41195 39856
rect 41195 39822 41204 39856
rect 41152 39811 41204 39822
rect 40894 39791 40946 39802
rect 40894 39757 40905 39791
rect 40905 39757 40939 39791
rect 40939 39757 40946 39791
rect 40894 39750 40946 39757
rect 39563 39683 39615 39735
rect 46139 39758 46319 39938
rect 41455 39508 41507 39560
rect 41519 39508 41571 39560
rect 41583 39508 41635 39560
rect 41647 39508 41699 39560
rect 41711 39508 41763 39560
rect 7110 39002 7290 39182
rect 12570 39002 12750 39182
rect 7242 38097 7294 38149
rect 5435 37149 5487 37201
rect 6707 37149 6759 37201
rect 3606 36036 3658 36088
rect 3670 36036 3722 36088
rect 3734 36036 3786 36088
rect 5081 36035 5133 36087
rect 5145 36035 5197 36087
rect 5209 36035 5261 36087
rect 5273 36035 5325 36087
rect 9434 37593 9486 37645
rect 5597 36036 5649 36088
rect 5661 36036 5713 36088
rect 5725 36036 5777 36088
rect 6956 36028 7008 36080
rect 7020 36028 7072 36080
rect 7084 36028 7136 36080
rect 7410 36035 7462 36087
rect 7474 36035 7526 36087
rect 7538 36035 7590 36087
rect 7602 36035 7654 36087
rect 8948 36034 9000 36086
rect 9012 36034 9064 36086
rect 9076 36034 9128 36086
rect 9140 36034 9192 36086
rect 9204 36034 9256 36086
rect 9268 36034 9320 36086
rect 9598 36031 9650 36083
rect 9662 36031 9714 36083
rect 9726 36031 9778 36083
rect 5436 34962 5488 35014
rect 7248 34960 7300 35012
rect 3745 33798 3797 33850
rect -6942 33121 -6890 33173
rect -6983 31753 -6931 31805
rect -6919 31753 -6867 31805
rect 5436 34367 5488 34419
rect 7248 34367 7300 34419
rect 5436 33503 5488 33555
rect 7434 33511 7486 33563
rect 9745 33798 9797 33850
rect 4360 30374 4412 30426
rect 8334 30379 8386 30431
rect -9391 30247 -9339 30299
rect -9327 30247 -9275 30299
rect -12687 29694 -12635 29746
rect -30193 29165 -30077 29281
rect -18517 29165 -18401 29281
rect -13463 29271 -13411 29323
rect 1957 28750 2009 28802
rect 2021 28750 2073 28802
rect 7966 28788 8018 28840
rect -6080 28550 -6028 28602
rect -6016 28550 -5964 28602
rect 3405 28537 3457 28589
rect -15689 28037 -15637 28089
rect -15689 27973 -15637 28025
rect -13983 28014 -13931 28066
rect -31024 27807 -30908 27923
rect -19377 27807 -19261 27923
rect -15689 27909 -15637 27961
rect -15689 27845 -15637 27897
rect -15689 27781 -15637 27833
rect -15689 27717 -15637 27769
rect -15689 27653 -15637 27705
rect -12379 28007 -12327 28059
rect -12379 27943 -12327 27995
rect -12379 27879 -12327 27931
rect -12379 27815 -12327 27867
rect -12379 27751 -12327 27803
rect -12379 27687 -12327 27739
rect -18320 27517 -18268 27569
rect -17629 27522 -17513 27638
rect -14906 27519 -14854 27571
rect -12372 27350 -12320 27402
rect -12372 27286 -12320 27338
rect -14404 27207 -14352 27259
rect -12372 27222 -12320 27274
rect -18320 27040 -18268 27092
rect -18875 26702 -18823 26754
rect -38181 26536 -38129 26588
rect -38117 26536 -38065 26588
rect -38053 26536 -38001 26588
rect -37989 26536 -37937 26588
rect -37925 26536 -37873 26588
rect -37861 26536 -37809 26588
rect -37797 26536 -37745 26588
rect -37733 26536 -37681 26588
rect -37669 26536 -37617 26588
rect -37605 26536 -37553 26588
rect -37541 26536 -37489 26588
rect -37477 26536 -37425 26588
rect -37413 26536 -37361 26588
rect -37349 26536 -37297 26588
rect -37285 26536 -37233 26588
rect -37221 26536 -37169 26588
rect -37157 26536 -37105 26588
rect -37093 26536 -37041 26588
rect -37029 26536 -36977 26588
rect -36965 26536 -36913 26588
rect -36901 26536 -36849 26588
rect -36837 26536 -36785 26588
rect -36773 26536 -36721 26588
rect -36709 26536 -36657 26588
rect -36645 26536 -36593 26588
rect -36581 26536 -36529 26588
rect -36517 26536 -36465 26588
rect -36453 26536 -36401 26588
rect -36389 26536 -36337 26588
rect -36325 26536 -36273 26588
rect -36261 26536 -36209 26588
rect -36197 26536 -36145 26588
rect -36133 26536 -36081 26588
rect -36069 26536 -36017 26588
rect -36005 26536 -35953 26588
rect -35941 26536 -35889 26588
rect -35877 26536 -35825 26588
rect -35813 26536 -35761 26588
rect -35749 26536 -35697 26588
rect -35685 26536 -35633 26588
rect -35621 26536 -35569 26588
rect -35557 26536 -35505 26588
rect -35493 26536 -35441 26588
rect -35429 26536 -35377 26588
rect -35365 26536 -35313 26588
rect -35301 26536 -35249 26588
rect -35237 26536 -35185 26588
rect -35173 26536 -35121 26588
rect -35109 26536 -35057 26588
rect -35045 26536 -34993 26588
rect -34981 26536 -34929 26588
rect -34917 26536 -34865 26588
rect -18876 25919 -18824 25971
rect -25435 25398 -25383 25450
rect -25435 25334 -25383 25386
rect -25435 25270 -25383 25322
rect -25435 25206 -25383 25258
rect -40565 24963 -40385 25143
rect -32985 24990 -32869 25106
rect -25435 24867 -25383 24919
rect -25435 24803 -25383 24855
rect -25435 24739 -25383 24791
rect -38175 23528 -38123 23580
rect -38111 23528 -38059 23580
rect -38047 23528 -37995 23580
rect -37983 23528 -37931 23580
rect -37919 23528 -37867 23580
rect -37855 23528 -37803 23580
rect -37791 23528 -37739 23580
rect -37727 23528 -37675 23580
rect -37663 23528 -37611 23580
rect -37599 23528 -37547 23580
rect -37535 23528 -37483 23580
rect -37471 23528 -37419 23580
rect -37407 23528 -37355 23580
rect -37343 23528 -37291 23580
rect -37279 23528 -37227 23580
rect -37215 23528 -37163 23580
rect -37151 23528 -37099 23580
rect -37087 23528 -37035 23580
rect -37023 23528 -36971 23580
rect -36959 23528 -36907 23580
rect -36895 23528 -36843 23580
rect -36831 23528 -36779 23580
rect -36767 23528 -36715 23580
rect -36703 23528 -36651 23580
rect -36639 23528 -36587 23580
rect -36575 23528 -36523 23580
rect -36511 23528 -36459 23580
rect -36447 23528 -36395 23580
rect -36383 23528 -36331 23580
rect -36319 23528 -36267 23580
rect -36255 23528 -36203 23580
rect -36191 23528 -36139 23580
rect -36127 23528 -36075 23580
rect -36063 23528 -36011 23580
rect -35999 23528 -35947 23580
rect -35935 23528 -35883 23580
rect -35871 23528 -35819 23580
rect -35807 23528 -35755 23580
rect -35743 23528 -35691 23580
rect -35679 23528 -35627 23580
rect -35615 23528 -35563 23580
rect -35551 23528 -35499 23580
rect -35487 23528 -35435 23580
rect -35423 23528 -35371 23580
rect -35359 23528 -35307 23580
rect -35295 23528 -35243 23580
rect -35231 23528 -35179 23580
rect -35167 23528 -35115 23580
rect -35103 23528 -35051 23580
rect -35039 23528 -34987 23580
rect -34975 23528 -34923 23580
rect -34911 23528 -34859 23580
rect -14906 27031 -14854 27083
rect -17250 26702 -17198 26754
rect -10010 26530 -9958 26582
rect -9946 26530 -9894 26582
rect -13983 26414 -13931 26466
rect -17629 26293 -17513 26409
rect -12375 26405 -12323 26457
rect -12375 26341 -12323 26393
rect -15707 26200 -15655 26252
rect -15707 26136 -15655 26188
rect -15707 26072 -15655 26124
rect -12375 26277 -12323 26329
rect -12375 26213 -12323 26265
rect -12375 26149 -12323 26201
rect -12375 26085 -12323 26137
rect -14906 25915 -14854 25967
rect -12379 25751 -12327 25803
rect 1958 25762 2010 25814
rect 2022 25762 2074 25814
rect -12379 25687 -12327 25739
rect -14404 25607 -14352 25659
rect -12379 25623 -12327 25675
rect -15706 25366 -15654 25418
rect -15706 25302 -15654 25354
rect -15706 25238 -15654 25290
rect -15706 25174 -15654 25226
rect -15706 25110 -15654 25162
rect -15706 25046 -15654 25098
rect -3495 25356 -3443 25408
rect -3431 25356 -3379 25408
rect -17629 24880 -17513 24996
rect -13983 24814 -13931 24866
rect -12387 24655 -12335 24707
rect -12387 24591 -12335 24643
rect -12387 24527 -12335 24579
rect -12387 24463 -12335 24515
rect -18320 24399 -18268 24451
rect -14908 24389 -14856 24441
rect -12383 24159 -12331 24211
rect -18875 24060 -18823 24112
rect -17257 24060 -17205 24112
rect -12383 24095 -12331 24147
rect -14404 24007 -14352 24059
rect -12383 24031 -12331 24083
rect 9405 28534 9457 28586
rect 7966 25762 8018 25814
rect 5723 24524 5775 24576
rect 5723 24460 5775 24512
rect 5723 24396 5775 24448
rect 5723 24332 5775 24384
rect 5723 24268 5775 24320
rect 5723 24204 5775 24256
rect 3405 24043 3457 24095
rect -17629 23651 -17513 23767
rect -15718 23559 -15666 23611
rect -15718 23495 -15666 23547
rect -15718 23431 -15666 23483
rect 5649 24039 5701 24091
rect 7023 24043 7075 24095
rect 9405 24043 9457 24095
rect 42865 24093 42917 24145
rect 42929 24093 42981 24145
rect 42993 24093 43045 24145
rect 43057 24093 43109 24145
rect 43121 24093 43173 24145
rect 43185 24093 43237 24145
rect 43249 24093 43301 24145
rect 43313 24093 43365 24145
rect 43377 24093 43429 24145
rect 43441 24093 43493 24145
rect 43505 24093 43557 24145
rect 43569 24093 43621 24145
rect 43633 24093 43685 24145
rect 43697 24093 43749 24145
rect 43761 24093 43813 24145
rect 43825 24093 43877 24145
rect 43889 24093 43941 24145
rect 43953 24093 44005 24145
rect 44017 24093 44069 24145
rect 44081 24093 44133 24145
rect 44145 24093 44197 24145
rect 44209 24093 44261 24145
rect 44273 24093 44325 24145
rect 44337 24093 44389 24145
rect 44401 24093 44453 24145
rect 44465 24093 44517 24145
rect 44529 24093 44581 24145
rect 44593 24093 44645 24145
rect 44657 24093 44709 24145
rect 44721 24093 44773 24145
rect 44785 24093 44837 24145
rect 44849 24093 44901 24145
rect 44913 24093 44965 24145
rect 44977 24093 45029 24145
rect 45041 24093 45093 24145
rect 45105 24093 45157 24145
rect 45169 24093 45221 24145
rect 45233 24093 45285 24145
rect 45297 24093 45349 24145
rect 45361 24093 45413 24145
rect 45425 24093 45477 24145
rect 45489 24093 45541 24145
rect 45553 24093 45605 24145
rect 45617 24093 45669 24145
rect 45681 24093 45733 24145
rect 45745 24093 45797 24145
rect 45809 24093 45861 24145
rect 45873 24093 45925 24145
rect 45937 24093 45989 24145
rect 46001 24093 46053 24145
rect 46065 24093 46117 24145
rect 46129 24093 46181 24145
rect 35158 23808 35210 23860
rect 39357 23641 39409 23693
rect 37829 23557 37881 23609
rect 37829 23493 37881 23545
rect 39357 23577 39409 23629
rect 39357 23513 39409 23565
rect -13983 23214 -13931 23266
rect -12380 23201 -12328 23253
rect -12380 23137 -12328 23189
rect -12380 23073 -12328 23125
rect 8807 23275 8859 23327
rect 8871 23275 8923 23327
rect -12380 23009 -12328 23061
rect 2556 23005 2608 23057
rect 10208 23005 10260 23057
rect -12380 22945 -12328 22997
rect -12380 22881 -12328 22933
rect -14908 22719 -14856 22771
rect -11595 22718 -11543 22770
rect -11531 22718 -11479 22770
rect -12383 22549 -12331 22601
rect -12383 22485 -12331 22537
rect -14404 22407 -14352 22459
rect -12383 22421 -12331 22473
rect -6080 21613 -6028 21665
rect -6016 21613 -5964 21665
rect -3495 20751 -3443 20803
rect -3431 20751 -3379 20803
rect -38141 19000 -38089 19052
rect -38077 19000 -38025 19052
rect -38013 19000 -37961 19052
rect -37949 19000 -37897 19052
rect -37885 19000 -37833 19052
rect -37821 19000 -37769 19052
rect -37757 19000 -37705 19052
rect -37693 19000 -37641 19052
rect -37629 19000 -37577 19052
rect -37565 19000 -37513 19052
rect -37501 19000 -37449 19052
rect -37437 19000 -37385 19052
rect -37373 19000 -37321 19052
rect -37309 19000 -37257 19052
rect -37245 19000 -37193 19052
rect -37181 19000 -37129 19052
rect -37117 19000 -37065 19052
rect -37053 19000 -37001 19052
rect -36989 19000 -36937 19052
rect -36925 19000 -36873 19052
rect -36861 19000 -36809 19052
rect -36797 19000 -36745 19052
rect -36733 19000 -36681 19052
rect -36669 19000 -36617 19052
rect -36605 19000 -36553 19052
rect -36541 19000 -36489 19052
rect -36477 19000 -36425 19052
rect -36413 19000 -36361 19052
rect -36349 19000 -36297 19052
rect -36285 19000 -36233 19052
rect -36221 19000 -36169 19052
rect -36157 19000 -36105 19052
rect -36093 19000 -36041 19052
rect -36029 19000 -35977 19052
rect -35965 19000 -35913 19052
rect -35901 19000 -35849 19052
rect -35837 19000 -35785 19052
rect -35773 19000 -35721 19052
rect -35709 19000 -35657 19052
rect -35645 19000 -35593 19052
rect -35581 19000 -35529 19052
rect -35517 19000 -35465 19052
rect -35453 19000 -35401 19052
rect -35389 19000 -35337 19052
rect -35325 19000 -35273 19052
rect -35261 19000 -35209 19052
rect -35197 19000 -35145 19052
rect -35133 19000 -35081 19052
rect -35069 19000 -35017 19052
rect -35005 19000 -34953 19052
rect -34941 19000 -34889 19052
rect -25446 17844 -25394 17896
rect -25446 17780 -25394 17832
rect -25446 17716 -25394 17768
rect -25446 17652 -25394 17704
rect -40568 17422 -40388 17602
rect -438 20051 -386 20103
rect -438 19987 -386 20039
rect 1690 19352 1742 19404
rect 1690 19288 1742 19340
rect -31124 17460 -31008 17576
rect 239 17714 291 17766
rect -815 17467 -763 17519
rect -25440 17324 -25388 17376
rect -25440 17260 -25388 17312
rect -25440 17196 -25388 17248
rect 4397 21985 4449 22037
rect 8228 21985 8280 22037
rect 4397 20893 4449 20945
rect 8228 20893 8280 20945
rect 5400 20051 5452 20103
rect 5400 19987 5452 20039
rect 9400 20051 9452 20103
rect 9400 19987 9452 20039
rect 3401 19288 3453 19340
rect 3067 19048 3119 19100
rect 4871 19042 5179 19158
rect 7400 19352 7452 19404
rect 7400 19288 7452 19340
rect 7091 19048 7143 19100
rect -439 17163 -387 17215
rect -439 17099 -387 17151
rect 1690 17163 1742 17215
rect 1690 17099 1742 17151
rect 4301 17231 4353 17283
rect 8987 19048 9039 19100
rect 37836 23140 37888 23192
rect 37836 23076 37888 23128
rect 37836 23012 37888 23064
rect 37836 22948 37888 23000
rect 39352 23146 39404 23198
rect 39352 23082 39404 23134
rect 39352 23018 39404 23070
rect 39352 22954 39404 23006
rect 35100 22610 35280 22790
rect 35768 22673 35820 22725
rect 35832 22673 35884 22725
rect 35896 22673 35948 22725
rect 35960 22673 36012 22725
rect 39357 22315 39409 22367
rect 37835 22221 37887 22273
rect 37835 22157 37887 22209
rect 39357 22251 39409 22303
rect 39357 22187 39409 22239
rect 47584 22526 47764 22706
rect 37830 21760 37882 21812
rect 37830 21696 37882 21748
rect 37830 21632 37882 21684
rect 39358 21780 39410 21832
rect 39358 21716 39410 21768
rect 39358 21652 39410 21704
rect 39358 21588 39410 21640
rect 35158 21527 35210 21579
rect 42863 21097 42915 21149
rect 42927 21097 42979 21149
rect 42991 21097 43043 21149
rect 43055 21097 43107 21149
rect 43119 21097 43171 21149
rect 43183 21097 43235 21149
rect 43247 21097 43299 21149
rect 43311 21097 43363 21149
rect 43375 21097 43427 21149
rect 43439 21097 43491 21149
rect 43503 21097 43555 21149
rect 43567 21097 43619 21149
rect 43631 21097 43683 21149
rect 43695 21097 43747 21149
rect 43759 21097 43811 21149
rect 43823 21097 43875 21149
rect 43887 21097 43939 21149
rect 43951 21097 44003 21149
rect 44015 21097 44067 21149
rect 44079 21097 44131 21149
rect 44143 21097 44195 21149
rect 44207 21097 44259 21149
rect 44271 21097 44323 21149
rect 44335 21097 44387 21149
rect 44399 21097 44451 21149
rect 44463 21097 44515 21149
rect 44527 21097 44579 21149
rect 44591 21097 44643 21149
rect 44655 21097 44707 21149
rect 44719 21097 44771 21149
rect 44783 21097 44835 21149
rect 44847 21097 44899 21149
rect 44911 21097 44963 21149
rect 44975 21097 45027 21149
rect 45039 21097 45091 21149
rect 45103 21097 45155 21149
rect 45167 21097 45219 21149
rect 45231 21097 45283 21149
rect 45295 21097 45347 21149
rect 45359 21097 45411 21149
rect 45423 21097 45475 21149
rect 45487 21097 45539 21149
rect 45551 21097 45603 21149
rect 45615 21097 45667 21149
rect 45679 21097 45731 21149
rect 45743 21097 45795 21149
rect 45807 21097 45859 21149
rect 45871 21097 45923 21149
rect 45935 21097 45987 21149
rect 45999 21097 46051 21149
rect 46063 21097 46115 21149
rect 46127 21097 46179 21149
rect 14694 20969 14746 21021
rect 23676 20158 23728 20210
rect 12379 19989 12495 20105
rect 11301 19290 11417 19406
rect 23695 19324 23747 19376
rect 10238 19000 10290 19052
rect 8286 18660 8338 18712
rect 13580 18630 13632 18682
rect 23664 18370 23716 18422
rect 23695 17494 23747 17546
rect 7399 17301 7451 17353
rect 6233 17231 6285 17283
rect 7399 17237 7451 17289
rect 9402 17301 9454 17353
rect 9402 17237 9454 17289
rect 13891 17301 13943 17353
rect 13891 17237 13943 17289
rect 14696 17025 14748 17077
rect 3399 16808 3451 16860
rect 3399 16744 3451 16796
rect 5399 16808 5451 16860
rect 5399 16744 5451 16796
rect 13283 16808 13335 16860
rect 13283 16744 13335 16796
rect -3920 16230 -3868 16282
rect 261 16252 11129 16432
rect -38171 16005 -38119 16057
rect -38107 16005 -38055 16057
rect -38043 16005 -37991 16057
rect -37979 16005 -37927 16057
rect -37915 16005 -37863 16057
rect -37851 16005 -37799 16057
rect -37787 16005 -37735 16057
rect -37723 16005 -37671 16057
rect -37659 16005 -37607 16057
rect -37595 16005 -37543 16057
rect -37531 16005 -37479 16057
rect -37467 16005 -37415 16057
rect -37403 16005 -37351 16057
rect -37339 16005 -37287 16057
rect -37275 16005 -37223 16057
rect -37211 16005 -37159 16057
rect -37147 16005 -37095 16057
rect -37083 16005 -37031 16057
rect -37019 16005 -36967 16057
rect -36955 16005 -36903 16057
rect -36891 16005 -36839 16057
rect -36827 16005 -36775 16057
rect -36763 16005 -36711 16057
rect -36699 16005 -36647 16057
rect -36635 16005 -36583 16057
rect -36571 16005 -36519 16057
rect -36507 16005 -36455 16057
rect -36443 16005 -36391 16057
rect -36379 16005 -36327 16057
rect -36315 16005 -36263 16057
rect -36251 16005 -36199 16057
rect -36187 16005 -36135 16057
rect -36123 16005 -36071 16057
rect -36059 16005 -36007 16057
rect -35995 16005 -35943 16057
rect -35931 16005 -35879 16057
rect -35867 16005 -35815 16057
rect -35803 16005 -35751 16057
rect -35739 16005 -35687 16057
rect -35675 16005 -35623 16057
rect -35611 16005 -35559 16057
rect -35547 16005 -35495 16057
rect -35483 16005 -35431 16057
rect -35419 16005 -35367 16057
rect -35355 16005 -35303 16057
rect -35291 16005 -35239 16057
rect -35227 16005 -35175 16057
rect -35163 16005 -35111 16057
rect -35099 16005 -35047 16057
rect -35035 16005 -34983 16057
rect -34971 16005 -34919 16057
rect -34907 16005 -34855 16057
rect -5780 15650 -5728 15702
rect -3914 15083 -3862 15135
rect -678 15084 -626 15136
rect -3129 14928 -3077 14980
rect -3129 14864 -3077 14916
rect -3129 14800 -3077 14852
rect -3129 14736 -3077 14788
rect -25507 14371 -25455 14423
rect -25507 14307 -25455 14359
rect -25507 14243 -25455 14295
rect -4893 14379 -4841 14431
rect -4893 14315 -4841 14367
rect -4893 14251 -4841 14303
rect -25507 14179 -25455 14231
rect -32985 13980 -32869 14096
rect -13058 14083 -13006 14135
rect -6538 14083 -6486 14135
rect -3914 14087 -3862 14139
rect -18217 14015 -18165 14067
rect -25508 13845 -25456 13897
rect -25508 13781 -25456 13833
rect -25508 13717 -25456 13769
rect -4901 13922 -4849 13974
rect -4901 13858 -4849 13910
rect -4901 13794 -4849 13846
rect -4901 13730 -4849 13782
rect -1793 13063 -1741 13115
rect -1793 12999 -1741 13051
rect -1793 12935 -1741 12987
rect -6538 12834 -6486 12886
rect -5845 12834 -5793 12886
rect -1793 12871 -1741 12923
rect -1793 12807 -1741 12859
rect -1793 12743 -1741 12795
rect -3914 12583 -3862 12635
rect -279 12585 -227 12637
rect -1492 12351 -1440 12403
rect -5845 12161 -5793 12213
rect -1752 11468 -1700 11520
rect -1752 11404 -1700 11456
rect -1752 11340 -1700 11392
rect -1752 11276 -1700 11328
rect -1752 11212 -1700 11264
rect -1752 11148 -1700 11200
rect -3415 10982 -3363 11034
rect -279 10983 -227 11035
rect -5845 10891 -5793 10943
rect -6140 10769 -6088 10821
rect -6076 10769 -6024 10821
rect -6012 10769 -5960 10821
rect -5676 10768 -5624 10820
rect -5612 10768 -5560 10820
rect -5548 10768 -5496 10820
rect -5484 10768 -5432 10820
rect -1492 10725 -1440 10777
rect 49 16117 165 16160
rect 49 16083 88 16117
rect 88 16083 122 16117
rect 122 16083 165 16117
rect 49 16045 165 16083
rect 49 16011 88 16045
rect 88 16011 122 16045
rect 122 16011 165 16045
rect 49 15973 165 16011
rect 49 15939 88 15973
rect 88 15939 122 15973
rect 122 15939 165 15973
rect 49 15901 165 15939
rect 49 15867 88 15901
rect 88 15867 122 15901
rect 122 15867 165 15901
rect 49 15829 165 15867
rect 49 15795 88 15829
rect 88 15795 122 15829
rect 122 15795 165 15829
rect 49 15757 165 15795
rect 49 15723 88 15757
rect 88 15723 122 15757
rect 122 15723 165 15757
rect 49 15685 165 15723
rect 49 15651 88 15685
rect 88 15651 122 15685
rect 122 15651 165 15685
rect 49 15613 165 15651
rect 49 15579 88 15613
rect 88 15579 122 15613
rect 122 15579 165 15613
rect 49 15541 165 15579
rect 49 15507 88 15541
rect 88 15507 122 15541
rect 122 15507 165 15541
rect 49 15469 165 15507
rect 49 15435 88 15469
rect 88 15435 122 15469
rect 122 15435 165 15469
rect 49 15397 165 15435
rect 49 15363 88 15397
rect 88 15363 122 15397
rect 122 15363 165 15397
rect 49 15325 165 15363
rect 49 15291 88 15325
rect 88 15291 122 15325
rect 122 15291 165 15325
rect 49 15253 165 15291
rect 49 15219 88 15253
rect 88 15219 122 15253
rect 122 15219 165 15253
rect 49 15181 165 15219
rect 49 15147 88 15181
rect 88 15147 122 15181
rect 122 15147 165 15181
rect 49 15109 165 15147
rect 49 15075 88 15109
rect 88 15075 122 15109
rect 122 15075 165 15109
rect 49 15037 165 15075
rect 49 15003 88 15037
rect 88 15003 122 15037
rect 122 15003 165 15037
rect 49 14965 165 15003
rect 49 14931 88 14965
rect 88 14931 122 14965
rect 122 14931 165 14965
rect 49 14893 165 14931
rect 49 14859 88 14893
rect 88 14859 122 14893
rect 122 14859 165 14893
rect 49 14821 165 14859
rect 49 14787 88 14821
rect 88 14787 122 14821
rect 122 14787 165 14821
rect 49 14749 165 14787
rect 49 14715 88 14749
rect 88 14715 122 14749
rect 122 14715 165 14749
rect 49 14677 165 14715
rect 49 14643 88 14677
rect 88 14643 122 14677
rect 122 14643 165 14677
rect 49 14605 165 14643
rect 49 14571 88 14605
rect 88 14571 122 14605
rect 122 14571 165 14605
rect 49 14533 165 14571
rect 49 14499 88 14533
rect 88 14499 122 14533
rect 122 14499 165 14533
rect 49 14461 165 14499
rect 49 14427 88 14461
rect 88 14427 122 14461
rect 122 14427 165 14461
rect 49 14389 165 14427
rect 49 14355 88 14389
rect 88 14355 122 14389
rect 122 14355 165 14389
rect 49 14317 165 14355
rect 49 14283 88 14317
rect 88 14283 122 14317
rect 122 14283 165 14317
rect 49 14245 165 14283
rect 49 14211 88 14245
rect 88 14211 122 14245
rect 122 14211 165 14245
rect 49 14173 165 14211
rect 49 14139 88 14173
rect 88 14139 122 14173
rect 122 14139 165 14173
rect 49 14101 165 14139
rect 49 14067 88 14101
rect 88 14067 122 14101
rect 122 14067 165 14101
rect 49 14029 165 14067
rect 49 13995 88 14029
rect 88 13995 122 14029
rect 122 13995 165 14029
rect 49 13957 165 13995
rect 49 13923 88 13957
rect 88 13923 122 13957
rect 122 13923 165 13957
rect 49 13885 165 13923
rect 49 13851 88 13885
rect 88 13851 122 13885
rect 122 13851 165 13885
rect 49 13813 165 13851
rect 49 13779 88 13813
rect 88 13779 122 13813
rect 122 13779 165 13813
rect 49 13741 165 13779
rect 49 13707 88 13741
rect 88 13707 122 13741
rect 122 13707 165 13741
rect 49 13669 165 13707
rect 49 13635 88 13669
rect 88 13635 122 13669
rect 122 13635 165 13669
rect 49 13597 165 13635
rect 49 13563 88 13597
rect 88 13563 122 13597
rect 122 13563 165 13597
rect 49 13525 165 13563
rect 49 13491 88 13525
rect 88 13491 122 13525
rect 122 13491 165 13525
rect 49 13453 165 13491
rect 49 13419 88 13453
rect 88 13419 122 13453
rect 122 13419 165 13453
rect 49 13381 165 13419
rect 49 13347 88 13381
rect 88 13347 122 13381
rect 122 13347 165 13381
rect 49 13309 165 13347
rect 49 13275 88 13309
rect 88 13275 122 13309
rect 122 13275 165 13309
rect 49 13237 165 13275
rect 49 13203 88 13237
rect 88 13203 122 13237
rect 122 13203 165 13237
rect 49 13165 165 13203
rect 49 13131 88 13165
rect 88 13131 122 13165
rect 122 13131 165 13165
rect 49 13093 165 13131
rect 49 13059 88 13093
rect 88 13059 122 13093
rect 122 13059 165 13093
rect 49 13021 165 13059
rect 49 12987 88 13021
rect 88 12987 122 13021
rect 122 12987 165 13021
rect 49 12949 165 12987
rect 49 12915 88 12949
rect 88 12915 122 12949
rect 122 12915 165 12949
rect 49 12877 165 12915
rect 49 12843 88 12877
rect 88 12843 122 12877
rect 122 12843 165 12877
rect 49 12805 165 12843
rect 49 12771 88 12805
rect 88 12771 122 12805
rect 122 12771 165 12805
rect 49 12733 165 12771
rect 49 12699 88 12733
rect 88 12699 122 12733
rect 122 12699 165 12733
rect 49 12661 165 12699
rect 49 12627 88 12661
rect 88 12627 122 12661
rect 122 12627 165 12661
rect 49 12589 165 12627
rect 49 12555 88 12589
rect 88 12555 122 12589
rect 122 12555 165 12589
rect 49 12517 165 12555
rect 49 12483 88 12517
rect 88 12483 122 12517
rect 122 12483 165 12517
rect 49 12445 165 12483
rect 49 12411 88 12445
rect 88 12411 122 12445
rect 122 12411 165 12445
rect 49 12373 165 12411
rect 49 12339 88 12373
rect 88 12339 122 12373
rect 122 12339 165 12373
rect 49 12301 165 12339
rect 49 12267 88 12301
rect 88 12267 122 12301
rect 122 12267 165 12301
rect 49 12229 165 12267
rect 49 12195 88 12229
rect 88 12195 122 12229
rect 122 12195 165 12229
rect 49 12157 165 12195
rect 49 12123 88 12157
rect 88 12123 122 12157
rect 122 12123 165 12157
rect 49 12085 165 12123
rect 49 12051 88 12085
rect 88 12051 122 12085
rect 122 12051 165 12085
rect 49 12013 165 12051
rect 49 11979 88 12013
rect 88 11979 122 12013
rect 122 11979 165 12013
rect 49 11941 165 11979
rect 49 11907 88 11941
rect 88 11907 122 11941
rect 122 11907 165 11941
rect 49 11869 165 11907
rect 49 11835 88 11869
rect 88 11835 122 11869
rect 122 11835 165 11869
rect 49 11797 165 11835
rect 49 11763 88 11797
rect 88 11763 122 11797
rect 122 11763 165 11797
rect 49 11725 165 11763
rect 49 11691 88 11725
rect 88 11691 122 11725
rect 122 11691 165 11725
rect 49 11653 165 11691
rect 49 11619 88 11653
rect 88 11619 122 11653
rect 122 11619 165 11653
rect 49 11581 165 11619
rect 49 11547 88 11581
rect 88 11547 122 11581
rect 122 11547 165 11581
rect 49 11509 165 11547
rect 49 11475 88 11509
rect 88 11475 122 11509
rect 122 11475 165 11509
rect 49 11437 165 11475
rect 49 11403 88 11437
rect 88 11403 122 11437
rect 122 11403 165 11437
rect 49 11365 165 11403
rect 49 11331 88 11365
rect 88 11331 122 11365
rect 122 11331 165 11365
rect 49 11293 165 11331
rect 49 11259 88 11293
rect 88 11259 122 11293
rect 122 11259 165 11293
rect 49 11221 165 11259
rect 49 11187 88 11221
rect 88 11187 122 11221
rect 122 11187 165 11221
rect 49 11149 165 11187
rect 49 11115 88 11149
rect 88 11115 122 11149
rect 122 11115 165 11149
rect 49 11077 165 11115
rect 49 11043 88 11077
rect 88 11043 122 11077
rect 122 11043 165 11077
rect 49 11005 165 11043
rect 49 10971 88 11005
rect 88 10971 122 11005
rect 122 10971 165 11005
rect 49 10933 165 10971
rect 49 10899 88 10933
rect 88 10899 122 10933
rect 122 10899 165 10933
rect 49 10861 165 10899
rect 49 10827 88 10861
rect 88 10827 122 10861
rect 122 10827 165 10861
rect 49 10789 165 10827
rect 49 10755 88 10789
rect 88 10755 122 10789
rect 122 10755 165 10789
rect 49 10717 165 10755
rect 49 10683 88 10717
rect 88 10683 122 10717
rect 122 10683 165 10717
rect 49 10668 165 10683
rect 11261 16122 11377 16163
rect 11261 16088 11303 16122
rect 11303 16088 11337 16122
rect 11337 16088 11377 16122
rect 11261 16050 11377 16088
rect 11261 16016 11303 16050
rect 11303 16016 11337 16050
rect 11337 16016 11377 16050
rect 11261 15978 11377 16016
rect 11261 15944 11303 15978
rect 11303 15944 11337 15978
rect 11337 15944 11377 15978
rect 11261 15906 11377 15944
rect 11261 15872 11303 15906
rect 11303 15872 11337 15906
rect 11337 15872 11377 15906
rect 11261 15834 11377 15872
rect 11261 15800 11303 15834
rect 11303 15800 11337 15834
rect 11337 15800 11377 15834
rect 11261 15762 11377 15800
rect 11261 15728 11303 15762
rect 11303 15728 11337 15762
rect 11337 15728 11377 15762
rect 11261 15690 11377 15728
rect 11261 15656 11303 15690
rect 11303 15656 11337 15690
rect 11337 15656 11377 15690
rect 11261 15618 11377 15656
rect 11261 15584 11303 15618
rect 11303 15584 11337 15618
rect 11337 15584 11377 15618
rect 11261 15546 11377 15584
rect 11261 15512 11303 15546
rect 11303 15512 11337 15546
rect 11337 15512 11377 15546
rect 11261 15474 11377 15512
rect 11261 15440 11303 15474
rect 11303 15440 11337 15474
rect 11337 15440 11377 15474
rect 11261 15402 11377 15440
rect 11261 15368 11303 15402
rect 11303 15368 11337 15402
rect 11337 15368 11377 15402
rect 11261 15330 11377 15368
rect 11261 15296 11303 15330
rect 11303 15296 11337 15330
rect 11337 15296 11377 15330
rect 11261 15258 11377 15296
rect 11261 15224 11303 15258
rect 11303 15224 11337 15258
rect 11337 15224 11377 15258
rect 11261 15186 11377 15224
rect 11261 15152 11303 15186
rect 11303 15152 11337 15186
rect 11337 15152 11377 15186
rect 11261 15114 11377 15152
rect 11261 15080 11303 15114
rect 11303 15080 11337 15114
rect 11337 15080 11377 15114
rect 11261 15042 11377 15080
rect 11261 15008 11303 15042
rect 11303 15008 11337 15042
rect 11337 15008 11377 15042
rect 11261 14970 11377 15008
rect 11261 14936 11303 14970
rect 11303 14936 11337 14970
rect 11337 14936 11377 14970
rect 11261 14898 11377 14936
rect 11261 14864 11303 14898
rect 11303 14864 11337 14898
rect 11337 14864 11377 14898
rect 11261 14826 11377 14864
rect 11261 14792 11303 14826
rect 11303 14792 11337 14826
rect 11337 14792 11377 14826
rect 11261 14754 11377 14792
rect 11261 14720 11303 14754
rect 11303 14720 11337 14754
rect 11337 14720 11377 14754
rect 11261 14682 11377 14720
rect 11261 14648 11303 14682
rect 11303 14648 11337 14682
rect 11337 14648 11377 14682
rect 11261 14610 11377 14648
rect 11261 14576 11303 14610
rect 11303 14576 11337 14610
rect 11337 14576 11377 14610
rect 11261 14538 11377 14576
rect 11261 14504 11303 14538
rect 11303 14504 11337 14538
rect 11337 14504 11377 14538
rect 11261 14466 11377 14504
rect 11261 14447 11303 14466
rect 11303 14447 11337 14466
rect 11337 14447 11377 14466
rect 23692 15730 23744 15782
rect 20934 15438 20986 15490
rect 14696 15170 14748 15222
rect 11262 13920 11378 13946
rect 11262 13886 11303 13920
rect 11303 13886 11337 13920
rect 11337 13886 11378 13920
rect 11262 13848 11378 13886
rect 11262 13814 11303 13848
rect 11303 13814 11337 13848
rect 11337 13814 11378 13848
rect 11262 13776 11378 13814
rect 11262 13742 11303 13776
rect 11303 13742 11337 13776
rect 11337 13742 11378 13776
rect 11262 13704 11378 13742
rect 11262 13670 11303 13704
rect 11303 13670 11337 13704
rect 11337 13670 11378 13704
rect 11262 13632 11378 13670
rect 11262 13598 11303 13632
rect 11303 13598 11337 13632
rect 11337 13598 11378 13632
rect 11262 13560 11378 13598
rect 11262 13526 11303 13560
rect 11303 13526 11337 13560
rect 11337 13526 11378 13560
rect 11262 13488 11378 13526
rect 11262 13454 11303 13488
rect 11303 13454 11337 13488
rect 11337 13454 11378 13488
rect 11262 13416 11378 13454
rect 11262 13382 11303 13416
rect 11303 13382 11337 13416
rect 11337 13382 11378 13416
rect 11262 13344 11378 13382
rect 11262 13310 11303 13344
rect 11303 13310 11337 13344
rect 11337 13310 11378 13344
rect 11262 13272 11378 13310
rect 11262 13238 11303 13272
rect 11303 13238 11337 13272
rect 11337 13238 11378 13272
rect 11262 13200 11378 13238
rect 11262 13166 11303 13200
rect 11303 13166 11337 13200
rect 11337 13166 11378 13200
rect 11262 13128 11378 13166
rect 11262 13094 11303 13128
rect 11303 13094 11337 13128
rect 11337 13094 11378 13128
rect 11262 13056 11378 13094
rect 11262 13022 11303 13056
rect 11303 13022 11337 13056
rect 11337 13022 11378 13056
rect 11262 12998 11378 13022
rect 14691 13907 14743 13959
rect 23692 13939 23744 13991
rect 14696 13470 14748 13522
rect 23691 12948 23743 13000
rect 14708 12122 14760 12174
rect 23697 12132 23749 12184
rect 11262 12091 11378 12100
rect 11262 12057 11303 12091
rect 11303 12057 11337 12091
rect 11337 12057 11378 12091
rect 11262 12019 11378 12057
rect 11262 11985 11303 12019
rect 11303 11985 11337 12019
rect 11337 11985 11378 12019
rect 11262 11947 11378 11985
rect 11262 11913 11303 11947
rect 11303 11913 11337 11947
rect 11337 11913 11378 11947
rect 11262 11875 11378 11913
rect 11262 11841 11303 11875
rect 11303 11841 11337 11875
rect 11337 11841 11378 11875
rect 11262 11803 11378 11841
rect 11262 11769 11303 11803
rect 11303 11769 11337 11803
rect 11337 11769 11378 11803
rect 11262 11731 11378 11769
rect 11262 11697 11303 11731
rect 11303 11697 11337 11731
rect 11337 11697 11378 11731
rect 11262 11659 11378 11697
rect 11262 11625 11303 11659
rect 11303 11625 11337 11659
rect 11337 11625 11378 11659
rect 11262 11587 11378 11625
rect 11262 11553 11303 11587
rect 11303 11553 11337 11587
rect 11337 11553 11378 11587
rect 11262 11515 11378 11553
rect 11262 11481 11303 11515
rect 11303 11481 11337 11515
rect 11337 11481 11378 11515
rect 11262 11443 11378 11481
rect 11262 11409 11303 11443
rect 11303 11409 11337 11443
rect 11337 11409 11378 11443
rect 11262 11371 11378 11409
rect 11262 11344 11303 11371
rect 11303 11344 11337 11371
rect 11337 11344 11378 11371
rect 14698 11618 14750 11670
rect 23695 11461 23747 11513
rect -5845 10349 -5793 10401
rect -678 10350 -626 10402
rect 14697 10325 14749 10377
rect 23697 10322 23749 10374
rect -1753 9865 -1701 9917
rect -1753 9801 -1701 9853
rect -1753 9737 -1701 9789
rect -1753 9673 -1701 9725
rect -1753 9609 -1701 9661
rect -6138 9526 -6086 9578
rect -6074 9526 -6022 9578
rect -6010 9526 -5958 9578
rect -5708 9526 -5656 9578
rect -5644 9526 -5592 9578
rect -5580 9526 -5528 9578
rect -5516 9526 -5464 9578
rect -5452 9526 -5400 9578
rect -1753 9545 -1701 9597
rect -5845 9400 -5793 9452
rect -3914 9385 -3862 9437
rect -1149 9383 -1097 9435
rect 5223 9365 5275 9417
rect 24550 9366 24602 9418
rect -1492 9067 -1440 9119
rect -1750 8264 -1698 8316
rect -1750 8200 -1698 8252
rect -5847 8116 -5795 8168
rect -1750 8136 -1698 8188
rect -1750 8072 -1698 8124
rect -1750 8008 -1698 8060
rect -1750 7944 -1698 7996
rect -3415 7783 -3363 7835
rect -1149 7783 -1097 7835
rect 23208 7792 23260 7844
rect -6559 7533 -6507 7585
rect -5847 7537 -5795 7589
rect -1492 7528 -1440 7580
rect -7201 7033 -6765 7213
rect -1492 7186 -1440 7238
rect -1492 7122 -1440 7174
rect -1492 7058 -1440 7110
rect -1492 6994 -1440 7046
rect -25510 6608 -25458 6660
rect -25510 6544 -25458 6596
rect -25510 6480 -25458 6532
rect -25510 6416 -25458 6468
rect -4903 6613 -4851 6665
rect -4903 6549 -4851 6601
rect -4903 6485 -4851 6537
rect -4903 6421 -4851 6473
rect -1492 6393 -1440 6445
rect -31124 6215 -31008 6331
rect -18245 6245 -18193 6297
rect -13069 6255 -13017 6307
rect -6559 6255 -6507 6307
rect -3415 6258 -3363 6310
rect -25511 6121 -25459 6173
rect -25511 6057 -25459 6109
rect -25511 5993 -25459 6045
rect -25511 5929 -25459 5981
rect -4900 6094 -4848 6146
rect -4900 6030 -4848 6082
rect -4900 5966 -4848 6018
rect -3415 5671 -3363 5723
rect -678 5671 -626 5723
rect -3178 5506 -3126 5558
rect -3178 5442 -3126 5494
rect -3178 5378 -3126 5430
rect -3178 5314 -3126 5366
rect -1149 5077 -1097 5129
rect -3421 4989 -3369 5041
rect 35030 8225 35082 8277
rect 40114 8065 40166 8117
rect 38584 7971 38636 8023
rect 38584 7907 38636 7959
rect 40114 8001 40166 8053
rect 40114 7937 40166 7989
rect 36326 7821 36378 7873
rect 36390 7821 36442 7873
rect 36454 7821 36506 7873
rect 33752 7593 33804 7645
rect 38582 7507 38634 7559
rect 38582 7443 38634 7495
rect 38582 7379 38634 7431
rect 40101 7520 40153 7572
rect 40101 7456 40153 7508
rect 40101 7392 40153 7444
rect 36388 7280 36440 7332
rect 36452 7280 36504 7332
rect 35034 7165 35086 7217
rect 42604 7161 42656 7213
rect 42668 7161 42720 7213
rect 42732 7161 42784 7213
rect 42796 7161 42848 7213
rect 42860 7161 42912 7213
rect 42924 7161 42976 7213
rect 42988 7161 43040 7213
rect 43052 7161 43104 7213
rect 43116 7161 43168 7213
rect 43180 7161 43232 7213
rect 43244 7161 43296 7213
rect 43308 7161 43360 7213
rect 43372 7161 43424 7213
rect 43436 7161 43488 7213
rect 43500 7161 43552 7213
rect 43564 7161 43616 7213
rect 43628 7161 43680 7213
rect 43692 7161 43744 7213
rect 43756 7161 43808 7213
rect 43820 7161 43872 7213
rect 43884 7161 43936 7213
rect 43948 7161 44000 7213
rect 44012 7161 44064 7213
rect 44076 7161 44128 7213
rect 44140 7161 44192 7213
rect 44204 7161 44256 7213
rect 44268 7161 44320 7213
rect 44332 7161 44384 7213
rect 44396 7161 44448 7213
rect 44460 7161 44512 7213
rect 44524 7161 44576 7213
rect 44588 7161 44640 7213
rect 44652 7161 44704 7213
rect 44716 7161 44768 7213
rect 44780 7161 44832 7213
rect 44844 7161 44896 7213
rect 44908 7161 44960 7213
rect 44972 7161 45024 7213
rect 45036 7161 45088 7213
rect 45100 7161 45152 7213
rect 45164 7161 45216 7213
rect 45228 7161 45280 7213
rect 45292 7161 45344 7213
rect 45356 7161 45408 7213
rect 45420 7161 45472 7213
rect 45484 7161 45536 7213
rect 45548 7161 45600 7213
rect 45612 7161 45664 7213
rect 45676 7161 45728 7213
rect 45740 7161 45792 7213
rect 45804 7161 45856 7213
rect 45868 7161 45920 7213
rect 35033 6896 35085 6948
rect 36368 6732 36420 6784
rect 40106 6729 40158 6781
rect 38584 6650 38636 6702
rect 38584 6586 38636 6638
rect 40106 6665 40158 6717
rect 40106 6601 40158 6653
rect 24550 6254 24602 6306
rect 33740 6254 33792 6306
rect 36993 6191 37045 6243
rect 38577 6176 38629 6228
rect 38577 6112 38629 6164
rect 38577 6048 38629 6100
rect 40106 6173 40158 6225
rect 40106 6109 40158 6161
rect 40106 6045 40158 6097
rect 35033 5827 35085 5879
rect 36001 5649 36053 5701
rect 36065 5649 36117 5701
rect 47501 5592 47681 5772
rect 35030 5504 35082 5556
rect 40123 5349 40175 5401
rect 38585 5260 38637 5312
rect 38585 5196 38637 5248
rect 40123 5285 40175 5337
rect 40123 5221 40175 5273
rect 36534 5101 36586 5153
rect 36598 5101 36650 5153
rect 36662 5101 36714 5153
rect 23208 4863 23260 4915
rect 33742 4863 33794 4915
rect 38576 4823 38628 4875
rect 38576 4759 38628 4811
rect 38576 4695 38628 4747
rect 40106 4801 40158 4853
rect 40106 4737 40158 4789
rect 40106 4673 40158 4725
rect 36378 4558 36430 4610
rect 36442 4558 36494 4610
rect 35041 4434 35093 4486
rect -279 3737 -227 3789
rect 23432 2354 23484 2406
rect 22589 1044 22641 1096
rect 352 91 21076 207
rect 35030 4129 35082 4181
rect 42621 4162 42673 4214
rect 42685 4162 42737 4214
rect 42749 4162 42801 4214
rect 42813 4162 42865 4214
rect 42877 4162 42929 4214
rect 42941 4162 42993 4214
rect 43005 4162 43057 4214
rect 43069 4162 43121 4214
rect 43133 4162 43185 4214
rect 43197 4162 43249 4214
rect 43261 4162 43313 4214
rect 43325 4162 43377 4214
rect 43389 4162 43441 4214
rect 43453 4162 43505 4214
rect 43517 4162 43569 4214
rect 43581 4162 43633 4214
rect 43645 4162 43697 4214
rect 43709 4162 43761 4214
rect 43773 4162 43825 4214
rect 43837 4162 43889 4214
rect 43901 4162 43953 4214
rect 43965 4162 44017 4214
rect 44029 4162 44081 4214
rect 44093 4162 44145 4214
rect 44157 4162 44209 4214
rect 44221 4162 44273 4214
rect 44285 4162 44337 4214
rect 44349 4162 44401 4214
rect 44413 4162 44465 4214
rect 44477 4162 44529 4214
rect 44541 4162 44593 4214
rect 44605 4162 44657 4214
rect 44669 4162 44721 4214
rect 44733 4162 44785 4214
rect 44797 4162 44849 4214
rect 44861 4162 44913 4214
rect 44925 4162 44977 4214
rect 44989 4162 45041 4214
rect 45053 4162 45105 4214
rect 45117 4162 45169 4214
rect 45181 4162 45233 4214
rect 45245 4162 45297 4214
rect 45309 4162 45361 4214
rect 45373 4162 45425 4214
rect 45437 4162 45489 4214
rect 45501 4162 45553 4214
rect 45565 4162 45617 4214
rect 45629 4162 45681 4214
rect 45693 4162 45745 4214
rect 45757 4162 45809 4214
rect 45821 4162 45873 4214
rect 45885 4162 45937 4214
rect 36994 4015 37046 4067
rect 40113 3970 40165 4022
rect 38585 3863 38637 3915
rect 38585 3799 38637 3851
rect 40113 3906 40165 3958
rect 40113 3842 40165 3894
rect 36364 3469 36416 3521
rect 36428 3469 36480 3521
rect 38579 3423 38631 3475
rect 38579 3359 38631 3411
rect 38579 3295 38631 3347
rect 40103 3417 40155 3469
rect 40103 3353 40155 3405
rect 40103 3289 40155 3341
rect 35037 3064 35089 3116
rect 35030 1285 35082 1337
rect 40114 1125 40166 1177
rect 38584 1031 38636 1083
rect 38584 967 38636 1019
rect 40114 1061 40166 1113
rect 40114 997 40166 1049
rect 36326 881 36378 933
rect 36390 881 36442 933
rect 36454 881 36506 933
rect 26012 652 26064 704
rect 33741 652 33793 704
rect 38582 567 38634 619
rect 38582 503 38634 555
rect 38582 439 38634 491
rect 40101 580 40153 632
rect 40101 516 40153 568
rect 40101 452 40153 504
rect 36388 340 36440 392
rect 36452 340 36504 392
rect 35034 225 35086 277
rect 42606 228 42658 280
rect 42670 228 42722 280
rect 42734 228 42786 280
rect 42798 228 42850 280
rect 42862 228 42914 280
rect 42926 228 42978 280
rect 42990 228 43042 280
rect 43054 228 43106 280
rect 43118 228 43170 280
rect 43182 228 43234 280
rect 43246 228 43298 280
rect 43310 228 43362 280
rect 43374 228 43426 280
rect 43438 228 43490 280
rect 43502 228 43554 280
rect 43566 228 43618 280
rect 43630 228 43682 280
rect 43694 228 43746 280
rect 43758 228 43810 280
rect 43822 228 43874 280
rect 43886 228 43938 280
rect 43950 228 44002 280
rect 44014 228 44066 280
rect 44078 228 44130 280
rect 44142 228 44194 280
rect 44206 228 44258 280
rect 44270 228 44322 280
rect 44334 228 44386 280
rect 44398 228 44450 280
rect 44462 228 44514 280
rect 44526 228 44578 280
rect 44590 228 44642 280
rect 44654 228 44706 280
rect 44718 228 44770 280
rect 44782 228 44834 280
rect 44846 228 44898 280
rect 44910 228 44962 280
rect 44974 228 45026 280
rect 45038 228 45090 280
rect 45102 228 45154 280
rect 45166 228 45218 280
rect 45230 228 45282 280
rect 45294 228 45346 280
rect 45358 228 45410 280
rect 45422 228 45474 280
rect 45486 228 45538 280
rect 45550 228 45602 280
rect 45614 228 45666 280
rect 45678 228 45730 280
rect 45742 228 45794 280
rect 45806 228 45858 280
rect 45870 228 45922 280
rect 35033 -44 35085 8
rect 36368 -208 36420 -156
rect 40106 -211 40158 -159
rect 38584 -290 38636 -238
rect 38584 -354 38636 -302
rect 40106 -275 40158 -223
rect 40106 -339 40158 -287
rect 23432 -693 23484 -641
rect 33741 -687 33793 -635
rect 36993 -749 37045 -697
rect 38577 -764 38629 -712
rect 38577 -828 38629 -776
rect 38577 -892 38629 -840
rect 40106 -767 40158 -715
rect 40106 -831 40158 -779
rect 40106 -895 40158 -843
rect 35033 -1113 35085 -1061
rect 36001 -1291 36053 -1239
rect 36065 -1291 36117 -1239
rect 47517 -1348 47697 -1168
rect 35030 -1436 35082 -1384
rect 40123 -1591 40175 -1539
rect 38585 -1680 38637 -1628
rect 38585 -1744 38637 -1692
rect 40123 -1655 40175 -1603
rect 40123 -1719 40175 -1667
rect 36534 -1839 36586 -1787
rect 36598 -1839 36650 -1787
rect 36662 -1839 36714 -1787
rect 22590 -2070 22642 -2018
rect 33750 -2073 33802 -2021
rect 38576 -2117 38628 -2065
rect 38576 -2181 38628 -2129
rect 38576 -2245 38628 -2193
rect 40106 -2139 40158 -2087
rect 40106 -2203 40158 -2151
rect 40106 -2267 40158 -2215
rect 36378 -2382 36430 -2330
rect 36442 -2382 36494 -2330
rect 35041 -2506 35093 -2454
rect 35030 -2811 35082 -2759
rect 42602 -2778 42654 -2726
rect 42666 -2778 42718 -2726
rect 42730 -2778 42782 -2726
rect 42794 -2778 42846 -2726
rect 42858 -2778 42910 -2726
rect 42922 -2778 42974 -2726
rect 42986 -2778 43038 -2726
rect 43050 -2778 43102 -2726
rect 43114 -2778 43166 -2726
rect 43178 -2778 43230 -2726
rect 43242 -2778 43294 -2726
rect 43306 -2778 43358 -2726
rect 43370 -2778 43422 -2726
rect 43434 -2778 43486 -2726
rect 43498 -2778 43550 -2726
rect 43562 -2778 43614 -2726
rect 43626 -2778 43678 -2726
rect 43690 -2778 43742 -2726
rect 43754 -2778 43806 -2726
rect 43818 -2778 43870 -2726
rect 43882 -2778 43934 -2726
rect 43946 -2778 43998 -2726
rect 44010 -2778 44062 -2726
rect 44074 -2778 44126 -2726
rect 44138 -2778 44190 -2726
rect 44202 -2778 44254 -2726
rect 44266 -2778 44318 -2726
rect 44330 -2778 44382 -2726
rect 44394 -2778 44446 -2726
rect 44458 -2778 44510 -2726
rect 44522 -2778 44574 -2726
rect 44586 -2778 44638 -2726
rect 44650 -2778 44702 -2726
rect 44714 -2778 44766 -2726
rect 44778 -2778 44830 -2726
rect 44842 -2778 44894 -2726
rect 44906 -2778 44958 -2726
rect 44970 -2778 45022 -2726
rect 45034 -2778 45086 -2726
rect 45098 -2778 45150 -2726
rect 45162 -2778 45214 -2726
rect 45226 -2778 45278 -2726
rect 45290 -2778 45342 -2726
rect 45354 -2778 45406 -2726
rect 45418 -2778 45470 -2726
rect 45482 -2778 45534 -2726
rect 45546 -2778 45598 -2726
rect 45610 -2778 45662 -2726
rect 45674 -2778 45726 -2726
rect 45738 -2778 45790 -2726
rect 45802 -2778 45854 -2726
rect 45866 -2778 45918 -2726
rect 36994 -2925 37046 -2873
rect 40113 -2970 40165 -2918
rect 38585 -3077 38637 -3025
rect 38585 -3141 38637 -3089
rect 40113 -3034 40165 -2982
rect 40113 -3098 40165 -3046
rect 36364 -3471 36416 -3419
rect 36428 -3471 36480 -3419
rect 38579 -3517 38631 -3465
rect 38579 -3581 38631 -3529
rect 38579 -3645 38631 -3593
rect 40103 -3523 40155 -3471
rect 40103 -3587 40155 -3535
rect 40103 -3651 40155 -3599
rect 35037 -3876 35089 -3824
rect -3575 -6902 -3523 -6850
rect -3575 -6966 -3523 -6914
rect -3575 -7030 -3523 -6978
rect -3575 -7094 -3523 -7042
rect -3575 -7158 -3523 -7106
rect -3575 -7222 -3523 -7170
rect -3575 -7286 -3523 -7234
rect -3575 -7350 -3523 -7298
rect -3575 -7414 -3523 -7362
rect -3575 -7478 -3523 -7426
rect -3575 -7542 -3523 -7490
rect -3575 -7606 -3523 -7554
rect -3575 -7670 -3523 -7618
rect -3575 -7734 -3523 -7682
rect -3575 -7798 -3523 -7746
rect -3575 -7862 -3523 -7810
rect -3575 -7926 -3523 -7874
rect -3575 -7990 -3523 -7938
rect -3575 -8054 -3523 -8002
rect -3575 -8118 -3523 -8066
rect -3575 -8182 -3523 -8130
rect -3575 -8246 -3523 -8194
rect -3575 -8310 -3523 -8258
rect -3575 -8374 -3523 -8322
rect -3575 -8438 -3523 -8386
rect -3575 -8502 -3523 -8450
rect -3575 -8566 -3523 -8514
rect -3575 -8630 -3523 -8578
rect -3575 -8694 -3523 -8642
rect -3575 -8758 -3523 -8706
rect -3575 -8822 -3523 -8770
rect -3575 -8886 -3523 -8834
rect -3575 -8950 -3523 -8898
rect -3575 -9014 -3523 -8962
rect -3575 -9078 -3523 -9026
rect -3575 -9142 -3523 -9090
rect -3575 -9206 -3523 -9154
rect -3575 -9270 -3523 -9218
rect -3575 -9334 -3523 -9282
rect -3575 -9398 -3523 -9346
rect -3575 -9462 -3523 -9410
rect -3575 -9526 -3523 -9474
rect -3575 -9590 -3523 -9538
rect -3575 -9654 -3523 -9602
rect -3575 -9718 -3523 -9666
rect -3575 -9782 -3523 -9730
rect -3575 -9846 -3523 -9794
rect -3575 -9910 -3523 -9858
rect -3575 -9974 -3523 -9922
rect -3575 -10038 -3523 -9986
rect -3575 -10102 -3523 -10050
rect -569 -6909 -517 -6857
rect -569 -6973 -517 -6921
rect -569 -7037 -517 -6985
rect -569 -7101 -517 -7049
rect -569 -7165 -517 -7113
rect -569 -7229 -517 -7177
rect -569 -7293 -517 -7241
rect -569 -7357 -517 -7305
rect -569 -7421 -517 -7369
rect -569 -7485 -517 -7433
rect -569 -7549 -517 -7497
rect -569 -7613 -517 -7561
rect -569 -7677 -517 -7625
rect -569 -7741 -517 -7689
rect -569 -7805 -517 -7753
rect -569 -7869 -517 -7817
rect -569 -7933 -517 -7881
rect -569 -7997 -517 -7945
rect -569 -8061 -517 -8009
rect -569 -8125 -517 -8073
rect -569 -8189 -517 -8137
rect -569 -8253 -517 -8201
rect -569 -8317 -517 -8265
rect -569 -8381 -517 -8329
rect -569 -8445 -517 -8393
rect -569 -8509 -517 -8457
rect -569 -8573 -517 -8521
rect -569 -8637 -517 -8585
rect -569 -8701 -517 -8649
rect -569 -8765 -517 -8713
rect -569 -8829 -517 -8777
rect -569 -8893 -517 -8841
rect -569 -8957 -517 -8905
rect -569 -9021 -517 -8969
rect -569 -9085 -517 -9033
rect -569 -9149 -517 -9097
rect -569 -9213 -517 -9161
rect -569 -9277 -517 -9225
rect -569 -9341 -517 -9289
rect -569 -9405 -517 -9353
rect -569 -9469 -517 -9417
rect -569 -9533 -517 -9481
rect -569 -9597 -517 -9545
rect -569 -9661 -517 -9609
rect -569 -9725 -517 -9673
rect -569 -9789 -517 -9737
rect -569 -9853 -517 -9801
rect -569 -9917 -517 -9865
rect -569 -9981 -517 -9929
rect -569 -10045 -517 -9993
rect -569 -10109 -517 -10057
rect -2151 -12290 -1971 -12110
<< metal2 >>
rect -15410 78130 -15174 78150
rect -15410 77914 -15400 78130
rect -15184 77914 -15174 78130
rect -15410 77894 -15174 77914
rect 12606 78101 12842 78121
rect 12606 77885 12616 78101
rect 12832 77885 12842 78101
rect 12606 77865 12842 77885
rect 24656 78102 24892 78122
rect 24656 77886 24666 78102
rect 24882 77886 24892 78102
rect 24656 77866 24892 77886
rect 14144 76743 14272 76755
rect -16849 76718 -16748 76733
rect -16849 76688 -16825 76718
rect -16773 76688 -16748 76718
rect -16849 76632 -16827 76688
rect -16771 76632 -16748 76688
rect -16849 76608 -16825 76632
rect -16773 76608 -16748 76632
rect -16849 76552 -16827 76608
rect -16771 76552 -16748 76608
rect -16849 76538 -16825 76552
rect -16773 76538 -16748 76552
rect -16849 76528 -16748 76538
rect -16849 76472 -16827 76528
rect -16771 76472 -16748 76528
rect -16849 76462 -16748 76472
rect -16849 76448 -16825 76462
rect -16773 76448 -16748 76462
rect -16849 76392 -16827 76448
rect -16771 76392 -16748 76448
rect -16849 76368 -16825 76392
rect -16773 76368 -16748 76392
rect -16849 76312 -16827 76368
rect -16771 76312 -16748 76368
rect -16849 76288 -16825 76312
rect -16773 76288 -16748 76312
rect -16849 76232 -16827 76288
rect -16771 76232 -16748 76288
rect -16849 76218 -16825 76232
rect -16773 76218 -16748 76232
rect -16849 76208 -16748 76218
rect -16849 76152 -16827 76208
rect -16771 76152 -16748 76208
rect -16849 76142 -16748 76152
rect -16849 76128 -16825 76142
rect -16773 76128 -16748 76142
rect -16849 76072 -16827 76128
rect -16771 76072 -16748 76128
rect -16849 76048 -16825 76072
rect -16773 76048 -16748 76072
rect -16849 75992 -16827 76048
rect -16771 75992 -16748 76048
rect -16849 75968 -16825 75992
rect -16773 75968 -16748 75992
rect -16849 75912 -16827 75968
rect -16771 75912 -16748 75968
rect -16849 75898 -16825 75912
rect -16773 75898 -16748 75912
rect -16849 75888 -16748 75898
rect -16849 75832 -16827 75888
rect -16771 75832 -16748 75888
rect -16849 75822 -16748 75832
rect -16849 75808 -16825 75822
rect -16773 75808 -16748 75822
rect -16849 75752 -16827 75808
rect -16771 75752 -16748 75808
rect -16849 75728 -16825 75752
rect -16773 75728 -16748 75752
rect -16849 75672 -16827 75728
rect -16771 75672 -16748 75728
rect -16849 75648 -16825 75672
rect -16773 75648 -16748 75672
rect -16849 75592 -16827 75648
rect -16771 75592 -16748 75648
rect -16849 75578 -16825 75592
rect -16773 75578 -16748 75592
rect -16849 75568 -16748 75578
rect -16849 75512 -16827 75568
rect -16771 75512 -16748 75568
rect -16849 75502 -16748 75512
rect -16849 75488 -16825 75502
rect -16773 75488 -16748 75502
rect -16849 75432 -16827 75488
rect -16771 75432 -16748 75488
rect -16849 75408 -16825 75432
rect -16773 75408 -16748 75432
rect -16849 75352 -16827 75408
rect -16771 75352 -16748 75408
rect -16849 75328 -16825 75352
rect -16773 75328 -16748 75352
rect -16849 75272 -16827 75328
rect -16771 75272 -16748 75328
rect -16849 75258 -16825 75272
rect -16773 75258 -16748 75272
rect -16849 75248 -16748 75258
rect -16849 75192 -16827 75248
rect -16771 75192 -16748 75248
rect -16849 75182 -16748 75192
rect -16849 75168 -16825 75182
rect -16773 75168 -16748 75182
rect -16849 75112 -16827 75168
rect -16771 75112 -16748 75168
rect -16849 75088 -16825 75112
rect -16773 75088 -16748 75112
rect -16849 75032 -16827 75088
rect -16771 75032 -16748 75088
rect -16849 75008 -16825 75032
rect -16773 75008 -16748 75032
rect -16849 74952 -16827 75008
rect -16771 74952 -16748 75008
rect -16849 74938 -16825 74952
rect -16773 74938 -16748 74952
rect -16849 74928 -16748 74938
rect -16849 74872 -16827 74928
rect -16771 74872 -16748 74928
rect -16849 74862 -16748 74872
rect -16849 74848 -16825 74862
rect -16773 74848 -16748 74862
rect -16849 74792 -16827 74848
rect -16771 74792 -16748 74848
rect -16849 74768 -16825 74792
rect -16773 74768 -16748 74792
rect -16849 74712 -16827 74768
rect -16771 74712 -16748 74768
rect -16849 74688 -16825 74712
rect -16773 74688 -16748 74712
rect -16849 74632 -16827 74688
rect -16771 74632 -16748 74688
rect -16849 74618 -16825 74632
rect -16773 74618 -16748 74632
rect -16849 74608 -16748 74618
rect -16849 74552 -16827 74608
rect -16771 74552 -16748 74608
rect -16849 74542 -16748 74552
rect -16849 74528 -16825 74542
rect -16773 74528 -16748 74542
rect -16849 74472 -16827 74528
rect -16771 74472 -16748 74528
rect -16849 74448 -16825 74472
rect -16773 74448 -16748 74472
rect -16849 74392 -16827 74448
rect -16771 74392 -16748 74448
rect -16849 74368 -16825 74392
rect -16773 74368 -16748 74392
rect -16849 74312 -16827 74368
rect -16771 74312 -16748 74368
rect -16849 74298 -16825 74312
rect -16773 74298 -16748 74312
rect -16849 74288 -16748 74298
rect -16849 74232 -16827 74288
rect -16771 74232 -16748 74288
rect -16849 74222 -16748 74232
rect -16849 74208 -16825 74222
rect -16773 74208 -16748 74222
rect -16849 74152 -16827 74208
rect -16771 74152 -16748 74208
rect -16849 74128 -16825 74152
rect -16773 74128 -16748 74152
rect -16849 74072 -16827 74128
rect -16771 74072 -16748 74128
rect -16849 74048 -16825 74072
rect -16773 74048 -16748 74072
rect -16849 73992 -16827 74048
rect -16771 73992 -16748 74048
rect -16849 73978 -16825 73992
rect -16773 73978 -16748 73992
rect -16849 73968 -16748 73978
rect -16849 73912 -16827 73968
rect -16771 73912 -16748 73968
rect -16849 73902 -16748 73912
rect -16849 73888 -16825 73902
rect -16773 73888 -16748 73902
rect -16849 73832 -16827 73888
rect -16771 73832 -16748 73888
rect -16849 73808 -16825 73832
rect -16773 73808 -16748 73832
rect -16849 73752 -16827 73808
rect -16771 73752 -16748 73808
rect -16849 73728 -16825 73752
rect -16773 73728 -16748 73752
rect -16849 73672 -16827 73728
rect -16771 73672 -16748 73728
rect -16849 73658 -16825 73672
rect -16773 73658 -16748 73672
rect -16849 73648 -16748 73658
rect -16849 73592 -16827 73648
rect -16771 73592 -16748 73648
rect -16849 73582 -16748 73592
rect -16849 73568 -16825 73582
rect -16773 73568 -16748 73582
rect -16849 73512 -16827 73568
rect -16771 73512 -16748 73568
rect -16849 73488 -16825 73512
rect -16773 73488 -16748 73512
rect -16849 73432 -16827 73488
rect -16771 73432 -16748 73488
rect -16849 73402 -16825 73432
rect -16773 73402 -16748 73432
rect -16849 73388 -16748 73402
rect -13848 76724 -13747 76739
rect -13848 76694 -13824 76724
rect -13772 76694 -13747 76724
rect -13848 76638 -13826 76694
rect -13770 76638 -13747 76694
rect -13848 76614 -13824 76638
rect -13772 76614 -13747 76638
rect -13848 76558 -13826 76614
rect -13770 76558 -13747 76614
rect -13848 76544 -13824 76558
rect -13772 76544 -13747 76558
rect -13848 76534 -13747 76544
rect -13848 76478 -13826 76534
rect -13770 76478 -13747 76534
rect -13848 76468 -13747 76478
rect -13848 76454 -13824 76468
rect -13772 76454 -13747 76468
rect -13848 76398 -13826 76454
rect -13770 76398 -13747 76454
rect -13848 76374 -13824 76398
rect -13772 76374 -13747 76398
rect -13848 76318 -13826 76374
rect -13770 76318 -13747 76374
rect -13848 76294 -13824 76318
rect -13772 76294 -13747 76318
rect -13848 76238 -13826 76294
rect -13770 76238 -13747 76294
rect -13848 76224 -13824 76238
rect -13772 76224 -13747 76238
rect -13848 76214 -13747 76224
rect -13848 76158 -13826 76214
rect -13770 76158 -13747 76214
rect -13848 76148 -13747 76158
rect -13848 76134 -13824 76148
rect -13772 76134 -13747 76148
rect -13848 76078 -13826 76134
rect -13770 76078 -13747 76134
rect -13848 76054 -13824 76078
rect -13772 76054 -13747 76078
rect -13848 75998 -13826 76054
rect -13770 75998 -13747 76054
rect -13848 75974 -13824 75998
rect -13772 75974 -13747 75998
rect -13848 75918 -13826 75974
rect -13770 75918 -13747 75974
rect -13848 75904 -13824 75918
rect -13772 75904 -13747 75918
rect -13848 75894 -13747 75904
rect -13848 75838 -13826 75894
rect -13770 75838 -13747 75894
rect -13848 75828 -13747 75838
rect -13848 75814 -13824 75828
rect -13772 75814 -13747 75828
rect -13848 75758 -13826 75814
rect -13770 75758 -13747 75814
rect -13848 75734 -13824 75758
rect -13772 75734 -13747 75758
rect -13848 75678 -13826 75734
rect -13770 75678 -13747 75734
rect -13848 75654 -13824 75678
rect -13772 75654 -13747 75678
rect -13848 75598 -13826 75654
rect -13770 75598 -13747 75654
rect -13848 75584 -13824 75598
rect -13772 75584 -13747 75598
rect -13848 75574 -13747 75584
rect -13848 75518 -13826 75574
rect -13770 75518 -13747 75574
rect -13848 75508 -13747 75518
rect -13848 75494 -13824 75508
rect -13772 75494 -13747 75508
rect -13848 75438 -13826 75494
rect -13770 75438 -13747 75494
rect -13848 75414 -13824 75438
rect -13772 75414 -13747 75438
rect -13848 75358 -13826 75414
rect -13770 75358 -13747 75414
rect -13848 75334 -13824 75358
rect -13772 75334 -13747 75358
rect -13848 75278 -13826 75334
rect -13770 75278 -13747 75334
rect -13848 75264 -13824 75278
rect -13772 75264 -13747 75278
rect -13848 75254 -13747 75264
rect -13848 75198 -13826 75254
rect -13770 75198 -13747 75254
rect -13848 75188 -13747 75198
rect -13848 75174 -13824 75188
rect -13772 75174 -13747 75188
rect -13848 75118 -13826 75174
rect -13770 75118 -13747 75174
rect -13848 75094 -13824 75118
rect -13772 75094 -13747 75118
rect -13848 75038 -13826 75094
rect -13770 75038 -13747 75094
rect -13848 75014 -13824 75038
rect -13772 75014 -13747 75038
rect -13848 74958 -13826 75014
rect -13770 74958 -13747 75014
rect -13848 74944 -13824 74958
rect -13772 74944 -13747 74958
rect -13848 74934 -13747 74944
rect -13848 74878 -13826 74934
rect -13770 74878 -13747 74934
rect -13848 74868 -13747 74878
rect -13848 74854 -13824 74868
rect -13772 74854 -13747 74868
rect -13848 74798 -13826 74854
rect -13770 74798 -13747 74854
rect -13848 74774 -13824 74798
rect -13772 74774 -13747 74798
rect -13848 74718 -13826 74774
rect -13770 74718 -13747 74774
rect -13848 74694 -13824 74718
rect -13772 74694 -13747 74718
rect -13848 74638 -13826 74694
rect -13770 74638 -13747 74694
rect -13848 74624 -13824 74638
rect -13772 74624 -13747 74638
rect -13848 74614 -13747 74624
rect -13848 74558 -13826 74614
rect -13770 74558 -13747 74614
rect -13848 74548 -13747 74558
rect -13848 74534 -13824 74548
rect -13772 74534 -13747 74548
rect -13848 74478 -13826 74534
rect -13770 74478 -13747 74534
rect -13848 74454 -13824 74478
rect -13772 74454 -13747 74478
rect -13848 74398 -13826 74454
rect -13770 74398 -13747 74454
rect -13848 74374 -13824 74398
rect -13772 74374 -13747 74398
rect -13848 74318 -13826 74374
rect -13770 74318 -13747 74374
rect -13848 74304 -13824 74318
rect -13772 74304 -13747 74318
rect -13848 74294 -13747 74304
rect -13848 74238 -13826 74294
rect -13770 74238 -13747 74294
rect -13848 74228 -13747 74238
rect -13848 74214 -13824 74228
rect -13772 74214 -13747 74228
rect -13848 74158 -13826 74214
rect -13770 74158 -13747 74214
rect -13848 74134 -13824 74158
rect -13772 74134 -13747 74158
rect -13848 74078 -13826 74134
rect -13770 74078 -13747 74134
rect -13848 74054 -13824 74078
rect -13772 74054 -13747 74078
rect -13848 73998 -13826 74054
rect -13770 73998 -13747 74054
rect -13848 73984 -13824 73998
rect -13772 73984 -13747 73998
rect -13848 73974 -13747 73984
rect -13848 73918 -13826 73974
rect -13770 73918 -13747 73974
rect -13848 73908 -13747 73918
rect -13848 73894 -13824 73908
rect -13772 73894 -13747 73908
rect -13848 73838 -13826 73894
rect -13770 73838 -13747 73894
rect -13848 73814 -13824 73838
rect -13772 73814 -13747 73838
rect -13848 73758 -13826 73814
rect -13770 73758 -13747 73814
rect -13848 73734 -13824 73758
rect -13772 73734 -13747 73758
rect -13848 73678 -13826 73734
rect -13770 73678 -13747 73734
rect -13848 73664 -13824 73678
rect -13772 73664 -13747 73678
rect -13848 73654 -13747 73664
rect -13848 73598 -13826 73654
rect -13770 73598 -13747 73654
rect -13848 73588 -13747 73598
rect -13848 73574 -13824 73588
rect -13772 73574 -13747 73588
rect -13848 73518 -13826 73574
rect -13770 73518 -13747 73574
rect -13848 73494 -13824 73518
rect -13772 73494 -13747 73518
rect -13848 73438 -13826 73494
rect -13770 73438 -13747 73494
rect -13848 73408 -13824 73438
rect -13772 73408 -13747 73438
rect -13848 73394 -13747 73408
rect 11143 76730 11271 76742
rect 11143 76720 11179 76730
rect 11235 76720 11271 76730
rect 11143 73404 11149 76720
rect 11265 73404 11271 76720
rect 11143 73394 11179 73404
rect 11235 73394 11271 73404
rect 14144 76733 14180 76743
rect 14236 76733 14272 76743
rect 14144 73417 14150 76733
rect 14266 73417 14272 76733
rect 14144 73407 14180 73417
rect 14236 73407 14272 73417
rect 14144 73395 14272 73407
rect 11143 73382 11271 73394
rect -16664 71798 -16600 71812
rect -16664 71742 -16660 71798
rect -16604 71742 -16600 71798
rect -16664 71728 -16600 71742
rect -15486 71794 -15422 71808
rect -15486 71738 -15482 71794
rect -15426 71738 -15422 71794
rect -15486 71724 -15422 71738
rect -15269 71801 -15205 71815
rect -15269 71745 -15265 71801
rect -15209 71745 -15205 71801
rect -15269 71731 -15205 71745
rect -14135 71798 -14071 71812
rect -14135 71742 -14131 71798
rect -14075 71742 -14071 71798
rect -14135 71728 -14071 71742
rect -16554 70294 -16490 70308
rect -16554 70238 -16550 70294
rect -16494 70238 -16490 70294
rect -16554 70224 -16490 70238
rect -15440 70280 -15376 70294
rect -15440 70224 -15436 70280
rect -15380 70224 -15376 70280
rect -15440 70210 -15376 70224
rect -15227 70281 -15163 70295
rect -15227 70225 -15223 70281
rect -15167 70225 -15163 70281
rect -15227 70211 -15163 70225
rect -14063 70281 -13999 70295
rect -14063 70225 -14059 70281
rect -14003 70225 -13999 70281
rect -14063 70211 -13999 70225
rect -16708 68699 -16644 68713
rect -16708 68643 -16704 68699
rect -16648 68643 -16644 68699
rect -16708 68629 -16644 68643
rect -16699 68335 -16647 68629
rect -15422 68494 -15358 68525
rect -15422 68488 -15416 68494
rect -15364 68488 -15358 68494
rect -15422 68432 -15418 68488
rect -15362 68432 -15358 68488
rect -15422 68430 -15358 68432
rect -15422 68408 -15416 68430
rect -15364 68408 -15358 68430
rect -15422 68352 -15418 68408
rect -15362 68352 -15358 68408
rect -15422 68328 -15416 68352
rect -15364 68328 -15358 68352
rect -15422 68272 -15418 68328
rect -15362 68272 -15358 68328
rect -15963 68251 -15890 68271
rect -15963 68195 -15955 68251
rect -15899 68195 -15890 68251
rect -15963 68189 -15953 68195
rect -15901 68189 -15890 68195
rect -15963 68177 -15890 68189
rect -15963 68171 -15953 68177
rect -15901 68171 -15890 68177
rect -15963 68115 -15955 68171
rect -15899 68115 -15890 68171
rect -15422 68250 -15416 68272
rect -15364 68250 -15358 68272
rect -15422 68248 -15358 68250
rect -15422 68192 -15418 68248
rect -15362 68192 -15358 68248
rect -15422 68186 -15416 68192
rect -15364 68186 -15358 68192
rect -15422 68156 -15358 68186
rect -14879 68254 -14806 68274
rect -14879 68198 -14871 68254
rect -14815 68198 -14806 68254
rect -14879 68192 -14869 68198
rect -14817 68192 -14806 68198
rect -14879 68180 -14806 68192
rect -14879 68174 -14869 68180
rect -14817 68174 -14806 68180
rect -15963 68095 -15890 68115
rect -14879 68118 -14871 68174
rect -14815 68118 -14806 68174
rect -14879 68098 -14806 68118
rect -14192 68083 -14140 68387
rect -14199 68069 -14135 68083
rect -14199 68013 -14195 68069
rect -14139 68013 -14135 68069
rect -14199 67999 -14135 68013
rect -14192 67996 -14140 67999
rect -16577 67609 -16513 67623
rect -16577 67553 -16573 67609
rect -16517 67553 -16513 67609
rect -16577 67539 -16513 67553
rect -15422 67603 -15358 67617
rect -15422 67547 -15418 67603
rect -15362 67547 -15358 67603
rect -15422 67533 -15358 67547
rect -14304 67614 -14240 67628
rect -14304 67558 -14300 67614
rect -14244 67558 -14240 67614
rect -14304 67544 -14240 67558
rect 17430 64738 17496 64753
rect 17430 64724 17437 64738
rect 17489 64724 17496 64738
rect 17430 64668 17435 64724
rect 17491 64668 17496 64724
rect 17430 64644 17437 64668
rect 17489 64644 17496 64668
rect 17430 64588 17435 64644
rect 17491 64588 17496 64644
rect 17430 64564 17437 64588
rect 17489 64564 17496 64588
rect 17430 64508 17435 64564
rect 17491 64508 17496 64564
rect 17430 64494 17437 64508
rect 17489 64494 17496 64508
rect 17430 64484 17496 64494
rect 17430 64428 17435 64484
rect 17491 64428 17496 64484
rect 17430 64418 17496 64428
rect 17430 64404 17437 64418
rect 17489 64404 17496 64418
rect 17430 64348 17435 64404
rect 17491 64348 17496 64404
rect 17430 64324 17437 64348
rect 17489 64324 17496 64348
rect 17430 64268 17435 64324
rect 17491 64268 17496 64324
rect 17430 64244 17437 64268
rect 17489 64244 17496 64268
rect 17430 64188 17435 64244
rect 17491 64188 17496 64244
rect 17430 64174 17437 64188
rect 17489 64174 17496 64188
rect 17430 64159 17496 64174
rect 23958 64738 24024 64753
rect 23958 64724 23965 64738
rect 24017 64724 24024 64738
rect 23958 64668 23963 64724
rect 24019 64668 24024 64724
rect 23958 64644 23965 64668
rect 24017 64644 24024 64668
rect 23958 64588 23963 64644
rect 24019 64588 24024 64644
rect 23958 64564 23965 64588
rect 24017 64564 24024 64588
rect 23958 64508 23963 64564
rect 24019 64508 24024 64564
rect 23958 64494 23965 64508
rect 24017 64494 24024 64508
rect 23958 64484 24024 64494
rect 23958 64428 23963 64484
rect 24019 64428 24024 64484
rect 23958 64418 24024 64428
rect 23958 64404 23965 64418
rect 24017 64404 24024 64418
rect 23958 64348 23963 64404
rect 24019 64348 24024 64404
rect 23958 64324 23965 64348
rect 24017 64324 24024 64348
rect 23958 64268 23963 64324
rect 24019 64268 24024 64324
rect 23958 64244 23965 64268
rect 24017 64244 24024 64268
rect 23958 64188 23963 64244
rect 24019 64188 24024 64244
rect 23958 64174 23965 64188
rect 24017 64174 24024 64188
rect 23958 64159 24024 64174
rect 31574 64738 31640 64753
rect 31574 64724 31581 64738
rect 31633 64724 31640 64738
rect 31574 64668 31579 64724
rect 31635 64668 31640 64724
rect 31574 64644 31581 64668
rect 31633 64644 31640 64668
rect 31574 64588 31579 64644
rect 31635 64588 31640 64644
rect 31574 64564 31581 64588
rect 31633 64564 31640 64588
rect 31574 64508 31579 64564
rect 31635 64508 31640 64564
rect 31574 64494 31581 64508
rect 31633 64494 31640 64508
rect 31574 64484 31640 64494
rect 31574 64428 31579 64484
rect 31635 64428 31640 64484
rect 31574 64418 31640 64428
rect 31574 64404 31581 64418
rect 31633 64404 31640 64418
rect 31574 64348 31579 64404
rect 31635 64348 31640 64404
rect 31574 64324 31581 64348
rect 31633 64324 31640 64348
rect 31574 64268 31579 64324
rect 31635 64268 31640 64324
rect 31574 64244 31581 64268
rect 31633 64244 31640 64268
rect 31574 64188 31579 64244
rect 31635 64188 31640 64244
rect 31574 64174 31581 64188
rect 31633 64174 31640 64188
rect 31574 64159 31640 64174
rect -9884 63398 -9442 63412
rect -9884 63396 -9851 63398
rect -9795 63396 -9771 63398
rect -9715 63396 -9691 63398
rect -9635 63396 -9611 63398
rect -9555 63396 -9531 63398
rect -9475 63396 -9442 63398
rect -9884 63344 -9881 63396
rect -9701 63344 -9691 63396
rect -9635 63344 -9625 63396
rect -9445 63344 -9442 63396
rect -9884 63342 -9851 63344
rect -9795 63342 -9771 63344
rect -9715 63342 -9691 63344
rect -9635 63342 -9611 63344
rect -9555 63342 -9531 63344
rect -9475 63342 -9442 63344
rect -9884 63328 -9442 63342
rect -8073 63400 -7631 63414
rect -8073 63398 -8040 63400
rect -7984 63398 -7960 63400
rect -7904 63398 -7880 63400
rect -7824 63398 -7800 63400
rect -7744 63398 -7720 63400
rect -7664 63398 -7631 63400
rect -8073 63346 -8070 63398
rect -7890 63346 -7880 63398
rect -7824 63346 -7814 63398
rect -7634 63346 -7631 63398
rect -8073 63344 -8040 63346
rect -7984 63344 -7960 63346
rect -7904 63344 -7880 63346
rect -7824 63344 -7800 63346
rect -7744 63344 -7720 63346
rect -7664 63344 -7631 63346
rect -8073 63330 -7631 63344
rect -6278 63396 -5836 63410
rect -6278 63394 -6245 63396
rect -6189 63394 -6165 63396
rect -6109 63394 -6085 63396
rect -6029 63394 -6005 63396
rect -5949 63394 -5925 63396
rect -5869 63394 -5836 63396
rect -6278 63342 -6275 63394
rect -6095 63342 -6085 63394
rect -6029 63342 -6019 63394
rect -5839 63342 -5836 63394
rect -6278 63340 -6245 63342
rect -6189 63340 -6165 63342
rect -6109 63340 -6085 63342
rect -6029 63340 -6005 63342
rect -5949 63340 -5925 63342
rect -5869 63340 -5836 63342
rect -6278 63326 -5836 63340
rect -4479 63394 -4037 63408
rect -4479 63392 -4446 63394
rect -4390 63392 -4366 63394
rect -4310 63392 -4286 63394
rect -4230 63392 -4206 63394
rect -4150 63392 -4126 63394
rect -4070 63392 -4037 63394
rect -4479 63340 -4476 63392
rect -4296 63340 -4286 63392
rect -4230 63340 -4220 63392
rect -4040 63340 -4037 63392
rect -4479 63338 -4446 63340
rect -4390 63338 -4366 63340
rect -4310 63338 -4286 63340
rect -4230 63338 -4206 63340
rect -4150 63338 -4126 63340
rect -4070 63338 -4037 63340
rect -4479 63324 -4037 63338
rect -2688 63398 -2246 63412
rect -2688 63396 -2655 63398
rect -2599 63396 -2575 63398
rect -2519 63396 -2495 63398
rect -2439 63396 -2415 63398
rect -2359 63396 -2335 63398
rect -2279 63396 -2246 63398
rect -2688 63344 -2685 63396
rect -2505 63344 -2495 63396
rect -2439 63344 -2429 63396
rect -2249 63344 -2246 63396
rect -2688 63342 -2655 63344
rect -2599 63342 -2575 63344
rect -2519 63342 -2495 63344
rect -2439 63342 -2415 63344
rect -2359 63342 -2335 63344
rect -2279 63342 -2246 63344
rect -2688 63328 -2246 63342
rect -886 63394 -444 63408
rect -886 63392 -853 63394
rect -797 63392 -773 63394
rect -717 63392 -693 63394
rect -637 63392 -613 63394
rect -557 63392 -533 63394
rect -477 63392 -444 63394
rect -886 63340 -883 63392
rect -703 63340 -693 63392
rect -637 63340 -627 63392
rect -447 63340 -444 63392
rect -886 63338 -853 63340
rect -797 63338 -773 63340
rect -717 63338 -693 63340
rect -637 63338 -613 63340
rect -557 63338 -533 63340
rect -477 63338 -444 63340
rect -886 63324 -444 63338
rect 757 63220 1287 63242
rect -6939 63194 -6699 63216
rect -6939 62978 -6927 63194
rect -6711 62978 -6699 63194
rect 757 63202 794 63220
rect 1250 63202 1287 63220
rect 757 63022 772 63202
rect 1272 63022 1287 63202
rect 757 63004 794 63022
rect 1250 63004 1287 63022
rect 757 62982 1287 63004
rect -6939 62956 -6699 62978
rect 17975 62735 18041 62750
rect 17975 62721 17982 62735
rect 18034 62721 18041 62735
rect 17975 62665 17980 62721
rect 18036 62665 18041 62721
rect 17975 62641 17982 62665
rect 18034 62641 18041 62665
rect 17975 62585 17980 62641
rect 18036 62585 18041 62641
rect 17975 62561 17982 62585
rect 18034 62561 18041 62585
rect 17975 62505 17980 62561
rect 18036 62505 18041 62561
rect 17975 62491 17982 62505
rect 18034 62491 18041 62505
rect 17975 62481 18041 62491
rect 17975 62425 17980 62481
rect 18036 62425 18041 62481
rect 17975 62415 18041 62425
rect 17975 62401 17982 62415
rect 18034 62401 18041 62415
rect 17975 62345 17980 62401
rect 18036 62345 18041 62401
rect 17975 62321 17982 62345
rect 18034 62321 18041 62345
rect 17975 62265 17980 62321
rect 18036 62265 18041 62321
rect 17975 62241 17982 62265
rect 18034 62241 18041 62265
rect 17975 62185 17980 62241
rect 18036 62185 18041 62241
rect 17975 62171 17982 62185
rect 18034 62171 18041 62185
rect 17975 62156 18041 62171
rect 19063 62735 19129 62750
rect 19063 62721 19070 62735
rect 19122 62721 19129 62735
rect 19063 62665 19068 62721
rect 19124 62665 19129 62721
rect 19063 62641 19070 62665
rect 19122 62641 19129 62665
rect 19063 62585 19068 62641
rect 19124 62585 19129 62641
rect 19063 62561 19070 62585
rect 19122 62561 19129 62585
rect 19063 62505 19068 62561
rect 19124 62505 19129 62561
rect 19063 62491 19070 62505
rect 19122 62491 19129 62505
rect 19063 62481 19129 62491
rect 19063 62425 19068 62481
rect 19124 62425 19129 62481
rect 19063 62415 19129 62425
rect 19063 62401 19070 62415
rect 19122 62401 19129 62415
rect 19063 62345 19068 62401
rect 19124 62345 19129 62401
rect 19063 62321 19070 62345
rect 19122 62321 19129 62345
rect 19063 62265 19068 62321
rect 19124 62265 19129 62321
rect 19063 62241 19070 62265
rect 19122 62241 19129 62265
rect 19063 62185 19068 62241
rect 19124 62185 19129 62241
rect 19063 62171 19070 62185
rect 19122 62171 19129 62185
rect 19063 62156 19129 62171
rect 21239 62735 21305 62750
rect 21239 62721 21246 62735
rect 21298 62721 21305 62735
rect 21239 62665 21244 62721
rect 21300 62665 21305 62721
rect 21239 62641 21246 62665
rect 21298 62641 21305 62665
rect 21239 62585 21244 62641
rect 21300 62585 21305 62641
rect 21239 62561 21246 62585
rect 21298 62561 21305 62585
rect 21239 62505 21244 62561
rect 21300 62505 21305 62561
rect 21239 62491 21246 62505
rect 21298 62491 21305 62505
rect 21239 62481 21305 62491
rect 21239 62425 21244 62481
rect 21300 62425 21305 62481
rect 21239 62415 21305 62425
rect 21239 62401 21246 62415
rect 21298 62401 21305 62415
rect 21239 62345 21244 62401
rect 21300 62345 21305 62401
rect 21239 62321 21246 62345
rect 21298 62321 21305 62345
rect 21239 62265 21244 62321
rect 21300 62265 21305 62321
rect 21239 62241 21246 62265
rect 21298 62241 21305 62265
rect 21239 62185 21244 62241
rect 21300 62185 21305 62241
rect 21239 62171 21246 62185
rect 21298 62171 21305 62185
rect 21239 62156 21305 62171
rect 22327 62735 22393 62750
rect 22327 62721 22334 62735
rect 22386 62721 22393 62735
rect 22327 62665 22332 62721
rect 22388 62665 22393 62721
rect 22327 62641 22334 62665
rect 22386 62641 22393 62665
rect 22327 62585 22332 62641
rect 22388 62585 22393 62641
rect 22327 62561 22334 62585
rect 22386 62561 22393 62585
rect 22327 62505 22332 62561
rect 22388 62505 22393 62561
rect 22327 62491 22334 62505
rect 22386 62491 22393 62505
rect 22327 62481 22393 62491
rect 22327 62425 22332 62481
rect 22388 62425 22393 62481
rect 22327 62415 22393 62425
rect 22327 62401 22334 62415
rect 22386 62401 22393 62415
rect 22327 62345 22332 62401
rect 22388 62345 22393 62401
rect 22327 62321 22334 62345
rect 22386 62321 22393 62345
rect 22327 62265 22332 62321
rect 22388 62265 22393 62321
rect 22327 62241 22334 62265
rect 22386 62241 22393 62265
rect 22327 62185 22332 62241
rect 22388 62185 22393 62241
rect 22327 62171 22334 62185
rect 22386 62171 22393 62185
rect 22327 62156 22393 62171
rect 23415 62735 23481 62750
rect 23415 62721 23422 62735
rect 23474 62721 23481 62735
rect 23415 62665 23420 62721
rect 23476 62665 23481 62721
rect 23415 62641 23422 62665
rect 23474 62641 23481 62665
rect 23415 62585 23420 62641
rect 23476 62585 23481 62641
rect 23415 62561 23422 62585
rect 23474 62561 23481 62585
rect 23415 62505 23420 62561
rect 23476 62505 23481 62561
rect 23415 62491 23422 62505
rect 23474 62491 23481 62505
rect 23415 62481 23481 62491
rect 23415 62425 23420 62481
rect 23476 62425 23481 62481
rect 23415 62415 23481 62425
rect 23415 62401 23422 62415
rect 23474 62401 23481 62415
rect 23415 62345 23420 62401
rect 23476 62345 23481 62401
rect 23415 62321 23422 62345
rect 23474 62321 23481 62345
rect 23415 62265 23420 62321
rect 23476 62265 23481 62321
rect 23415 62241 23422 62265
rect 23474 62241 23481 62265
rect 23415 62185 23420 62241
rect 23476 62185 23481 62241
rect 23415 62171 23422 62185
rect 23474 62171 23481 62185
rect 23415 62156 23481 62171
rect 24503 62735 24569 62750
rect 24503 62721 24510 62735
rect 24562 62721 24569 62735
rect 24503 62665 24508 62721
rect 24564 62665 24569 62721
rect 24503 62641 24510 62665
rect 24562 62641 24569 62665
rect 24503 62585 24508 62641
rect 24564 62585 24569 62641
rect 24503 62561 24510 62585
rect 24562 62561 24569 62585
rect 24503 62505 24508 62561
rect 24564 62505 24569 62561
rect 24503 62491 24510 62505
rect 24562 62491 24569 62505
rect 24503 62481 24569 62491
rect 24503 62425 24508 62481
rect 24564 62425 24569 62481
rect 24503 62415 24569 62425
rect 24503 62401 24510 62415
rect 24562 62401 24569 62415
rect 24503 62345 24508 62401
rect 24564 62345 24569 62401
rect 24503 62321 24510 62345
rect 24562 62321 24569 62345
rect 24503 62265 24508 62321
rect 24564 62265 24569 62321
rect 24503 62241 24510 62265
rect 24562 62241 24569 62265
rect 24503 62185 24508 62241
rect 24564 62185 24569 62241
rect 24503 62171 24510 62185
rect 24562 62171 24569 62185
rect 24503 62156 24569 62171
rect 25591 62735 25657 62750
rect 25591 62721 25598 62735
rect 25650 62721 25657 62735
rect 25591 62665 25596 62721
rect 25652 62665 25657 62721
rect 25591 62641 25598 62665
rect 25650 62641 25657 62665
rect 25591 62585 25596 62641
rect 25652 62585 25657 62641
rect 25591 62561 25598 62585
rect 25650 62561 25657 62585
rect 25591 62505 25596 62561
rect 25652 62505 25657 62561
rect 25591 62491 25598 62505
rect 25650 62491 25657 62505
rect 25591 62481 25657 62491
rect 25591 62425 25596 62481
rect 25652 62425 25657 62481
rect 25591 62415 25657 62425
rect 25591 62401 25598 62415
rect 25650 62401 25657 62415
rect 25591 62345 25596 62401
rect 25652 62345 25657 62401
rect 25591 62321 25598 62345
rect 25650 62321 25657 62345
rect 25591 62265 25596 62321
rect 25652 62265 25657 62321
rect 25591 62241 25598 62265
rect 25650 62241 25657 62265
rect 25591 62185 25596 62241
rect 25652 62185 25657 62241
rect 25591 62171 25598 62185
rect 25650 62171 25657 62185
rect 25591 62156 25657 62171
rect 26679 62735 26745 62750
rect 26679 62721 26686 62735
rect 26738 62721 26745 62735
rect 26679 62665 26684 62721
rect 26740 62665 26745 62721
rect 26679 62641 26686 62665
rect 26738 62641 26745 62665
rect 26679 62585 26684 62641
rect 26740 62585 26745 62641
rect 26679 62561 26686 62585
rect 26738 62561 26745 62585
rect 26679 62505 26684 62561
rect 26740 62505 26745 62561
rect 26679 62491 26686 62505
rect 26738 62491 26745 62505
rect 26679 62481 26745 62491
rect 26679 62425 26684 62481
rect 26740 62425 26745 62481
rect 26679 62415 26745 62425
rect 26679 62401 26686 62415
rect 26738 62401 26745 62415
rect 26679 62345 26684 62401
rect 26740 62345 26745 62401
rect 26679 62321 26686 62345
rect 26738 62321 26745 62345
rect 26679 62265 26684 62321
rect 26740 62265 26745 62321
rect 26679 62241 26686 62265
rect 26738 62241 26745 62265
rect 26679 62185 26684 62241
rect 26740 62185 26745 62241
rect 26679 62171 26686 62185
rect 26738 62171 26745 62185
rect 26679 62156 26745 62171
rect 28855 62735 28921 62750
rect 28855 62721 28862 62735
rect 28914 62721 28921 62735
rect 28855 62665 28860 62721
rect 28916 62665 28921 62721
rect 28855 62641 28862 62665
rect 28914 62641 28921 62665
rect 28855 62585 28860 62641
rect 28916 62585 28921 62641
rect 28855 62561 28862 62585
rect 28914 62561 28921 62585
rect 28855 62505 28860 62561
rect 28916 62505 28921 62561
rect 28855 62491 28862 62505
rect 28914 62491 28921 62505
rect 28855 62481 28921 62491
rect 28855 62425 28860 62481
rect 28916 62425 28921 62481
rect 28855 62415 28921 62425
rect 28855 62401 28862 62415
rect 28914 62401 28921 62415
rect 28855 62345 28860 62401
rect 28916 62345 28921 62401
rect 28855 62321 28862 62345
rect 28914 62321 28921 62345
rect 28855 62265 28860 62321
rect 28916 62265 28921 62321
rect 28855 62241 28862 62265
rect 28914 62241 28921 62265
rect 28855 62185 28860 62241
rect 28916 62185 28921 62241
rect 28855 62171 28862 62185
rect 28914 62171 28921 62185
rect 28855 62156 28921 62171
rect 29943 62735 30009 62750
rect 29943 62721 29950 62735
rect 30002 62721 30009 62735
rect 29943 62665 29948 62721
rect 30004 62665 30009 62721
rect 29943 62641 29950 62665
rect 30002 62641 30009 62665
rect 29943 62585 29948 62641
rect 30004 62585 30009 62641
rect 29943 62561 29950 62585
rect 30002 62561 30009 62585
rect 29943 62505 29948 62561
rect 30004 62505 30009 62561
rect 29943 62491 29950 62505
rect 30002 62491 30009 62505
rect 29943 62481 30009 62491
rect 29943 62425 29948 62481
rect 30004 62425 30009 62481
rect 29943 62415 30009 62425
rect 29943 62401 29950 62415
rect 30002 62401 30009 62415
rect 29943 62345 29948 62401
rect 30004 62345 30009 62401
rect 29943 62321 29950 62345
rect 30002 62321 30009 62345
rect 29943 62265 29948 62321
rect 30004 62265 30009 62321
rect 29943 62241 29950 62265
rect 30002 62241 30009 62265
rect 29943 62185 29948 62241
rect 30004 62185 30009 62241
rect 29943 62171 29950 62185
rect 30002 62171 30009 62185
rect 29943 62156 30009 62171
rect 31031 62735 31097 62750
rect 31031 62721 31038 62735
rect 31090 62721 31097 62735
rect 31031 62665 31036 62721
rect 31092 62665 31097 62721
rect 31031 62641 31038 62665
rect 31090 62641 31097 62665
rect 31031 62585 31036 62641
rect 31092 62585 31097 62641
rect 31031 62561 31038 62585
rect 31090 62561 31097 62585
rect 31031 62505 31036 62561
rect 31092 62505 31097 62561
rect 31031 62491 31038 62505
rect 31090 62491 31097 62505
rect 31031 62481 31097 62491
rect 31031 62425 31036 62481
rect 31092 62425 31097 62481
rect 31031 62415 31097 62425
rect 31031 62401 31038 62415
rect 31090 62401 31097 62415
rect 31031 62345 31036 62401
rect 31092 62345 31097 62401
rect 31031 62321 31038 62345
rect 31090 62321 31097 62345
rect 31031 62265 31036 62321
rect 31092 62265 31097 62321
rect 31031 62241 31038 62265
rect 31090 62241 31097 62265
rect 31031 62185 31036 62241
rect 31092 62185 31097 62241
rect 31031 62171 31038 62185
rect 31090 62171 31097 62185
rect 31031 62156 31097 62171
rect 347 60808 519 60837
rect 347 60802 375 60808
rect 491 60802 519 60808
rect -8557 54591 -8493 54605
rect -8557 54535 -8553 54591
rect -8497 54535 -8493 54591
rect -8557 54521 -8493 54535
rect -6866 54592 -6802 54606
rect -6866 54536 -6862 54592
rect -6806 54536 -6802 54592
rect -6866 54522 -6802 54536
rect -5161 54591 -5097 54605
rect -5161 54535 -5157 54591
rect -5101 54535 -5097 54591
rect -5161 54521 -5097 54535
rect -3365 54591 -3301 54605
rect -3365 54535 -3361 54591
rect -3305 54535 -3301 54591
rect -3365 54521 -3301 54535
rect -1536 54591 -1472 54605
rect -1536 54535 -1532 54591
rect -1476 54535 -1472 54591
rect -1536 54521 -1472 54535
rect -9704 54399 -9462 54413
rect -9704 54343 -9691 54399
rect -9635 54397 -9611 54399
rect -9555 54397 -9531 54399
rect -9621 54345 -9611 54397
rect -9555 54345 -9545 54397
rect -9635 54343 -9611 54345
rect -9555 54343 -9531 54345
rect -9475 54343 -9462 54399
rect -9704 54329 -9462 54343
rect -7909 54398 -7667 54412
rect -7909 54342 -7896 54398
rect -7840 54396 -7816 54398
rect -7760 54396 -7736 54398
rect -7826 54344 -7816 54396
rect -7760 54344 -7750 54396
rect -7840 54342 -7816 54344
rect -7760 54342 -7736 54344
rect -7680 54342 -7667 54398
rect -7909 54328 -7667 54342
rect -6109 54400 -5867 54414
rect -6109 54344 -6096 54400
rect -6040 54398 -6016 54400
rect -5960 54398 -5936 54400
rect -6026 54346 -6016 54398
rect -5960 54346 -5950 54398
rect -6040 54344 -6016 54346
rect -5960 54344 -5936 54346
rect -5880 54344 -5867 54400
rect -6109 54330 -5867 54344
rect -4311 54399 -4069 54413
rect -4311 54343 -4298 54399
rect -4242 54397 -4218 54399
rect -4162 54397 -4138 54399
rect -4228 54345 -4218 54397
rect -4162 54345 -4152 54397
rect -4242 54343 -4218 54345
rect -4162 54343 -4138 54345
rect -4082 54343 -4069 54399
rect -4311 54329 -4069 54343
rect -2513 54400 -2271 54414
rect -2513 54344 -2500 54400
rect -2444 54398 -2420 54400
rect -2364 54398 -2340 54400
rect -2430 54346 -2420 54398
rect -2364 54346 -2354 54398
rect -2444 54344 -2420 54346
rect -2364 54344 -2340 54346
rect -2284 54344 -2271 54400
rect -2513 54330 -2271 54344
rect -710 54399 -468 54413
rect -710 54343 -697 54399
rect -641 54397 -617 54399
rect -561 54397 -537 54399
rect -627 54345 -617 54397
rect -561 54345 -551 54397
rect -641 54343 -617 54345
rect -561 54343 -537 54345
rect -481 54343 -468 54399
rect -710 54329 -468 54343
rect 176 54400 240 54414
rect 176 54344 180 54400
rect 236 54344 240 54400
rect 176 54330 240 54344
rect -14783 53600 -14655 53610
rect -7550 53600 -7486 53610
rect -14783 53594 -7486 53600
rect -14783 53542 -14777 53594
rect -14725 53542 -14713 53594
rect -14661 53542 -7544 53594
rect -7492 53542 -7486 53594
rect -14783 53536 -7486 53542
rect -14783 53526 -14655 53536
rect -7550 53526 -7486 53536
rect -6989 53594 -6861 53610
rect -6989 53542 -6983 53594
rect -6931 53542 -6919 53594
rect -6867 53542 -6861 53594
rect -9398 52986 -9270 53002
rect -9398 52934 -9392 52986
rect -9340 52934 -9328 52986
rect -9276 52934 -9270 52986
rect -9398 50931 -9270 52934
rect -8854 51239 -8770 51259
rect -8854 51183 -8840 51239
rect -8784 51183 -8770 51239
rect -8854 51169 -8838 51183
rect -8786 51169 -8770 51183
rect -7722 51243 -7658 51257
rect -7722 51187 -7718 51243
rect -7662 51187 -7658 51243
rect -7722 51173 -7658 51187
rect -8854 51159 -8770 51169
rect -8854 51103 -8840 51159
rect -8784 51103 -8770 51159
rect -8854 51093 -8770 51103
rect -8854 51079 -8838 51093
rect -8786 51079 -8770 51093
rect -8854 51023 -8840 51079
rect -8784 51023 -8770 51079
rect -8854 51004 -8770 51023
rect -9398 50879 -9392 50931
rect -9340 50879 -9328 50931
rect -9276 50879 -9270 50931
rect -27070 49716 -26726 49730
rect -27070 49714 -27046 49716
rect -26990 49714 -26966 49716
rect -26910 49714 -26886 49716
rect -26830 49714 -26806 49716
rect -26750 49714 -26726 49716
rect -27070 49662 -27052 49714
rect -26990 49662 -26988 49714
rect -26808 49662 -26806 49714
rect -26744 49662 -26726 49714
rect -27070 49660 -27046 49662
rect -26990 49660 -26966 49662
rect -26910 49660 -26886 49662
rect -26830 49660 -26806 49662
rect -26750 49660 -26726 49662
rect -27070 49646 -26726 49660
rect -26408 49409 -26157 49423
rect -26408 49407 -26391 49409
rect -26335 49407 -26311 49409
rect -26255 49407 -26231 49409
rect -26175 49407 -26157 49409
rect -26408 49355 -26405 49407
rect -26161 49355 -26157 49407
rect -26408 49353 -26391 49355
rect -26335 49353 -26311 49355
rect -26255 49353 -26231 49355
rect -26175 49353 -26157 49355
rect -26408 49339 -26157 49353
rect -26060 49420 -25996 49434
rect -26060 49364 -26056 49420
rect -26000 49364 -25996 49420
rect -26060 49350 -25996 49364
rect -25984 49174 -25640 49188
rect -25984 49172 -25960 49174
rect -25904 49172 -25880 49174
rect -25824 49172 -25800 49174
rect -25744 49172 -25720 49174
rect -25664 49172 -25640 49174
rect -25984 49120 -25966 49172
rect -25904 49120 -25902 49172
rect -25722 49120 -25720 49172
rect -25658 49120 -25640 49172
rect -25984 49118 -25960 49120
rect -25904 49118 -25880 49120
rect -25824 49118 -25800 49120
rect -25744 49118 -25720 49120
rect -25664 49118 -25640 49120
rect -25984 49104 -25640 49118
rect -27087 43296 -26990 43323
rect -27087 43274 -27065 43296
rect -27013 43274 -26990 43296
rect -27087 43218 -27067 43274
rect -27011 43218 -26990 43274
rect -27087 43194 -27065 43218
rect -27013 43194 -26990 43218
rect -27087 43138 -27067 43194
rect -27011 43138 -26990 43194
rect -27087 43116 -27065 43138
rect -27013 43116 -26990 43138
rect -27087 43114 -26990 43116
rect -27087 43058 -27067 43114
rect -27011 43058 -26990 43114
rect -27087 43052 -27065 43058
rect -27013 43052 -26990 43058
rect -27087 43040 -26990 43052
rect -27087 43034 -27065 43040
rect -27013 43034 -26990 43040
rect -27087 42978 -27067 43034
rect -27011 42978 -26990 43034
rect -13469 43057 -13405 43071
rect -13469 43001 -13465 43057
rect -13409 43001 -13405 43057
rect -13469 42987 -13405 43001
rect -27087 42976 -26990 42978
rect -27087 42954 -27065 42976
rect -27013 42954 -26990 42976
rect -27087 42898 -27067 42954
rect -27011 42898 -26990 42954
rect -27087 42874 -27065 42898
rect -27013 42874 -26990 42898
rect -27087 42818 -27067 42874
rect -27011 42818 -26990 42874
rect -27087 42796 -27065 42818
rect -27013 42796 -26990 42818
rect -27087 42769 -26990 42796
rect -12693 42394 -12629 42408
rect -12693 42338 -12689 42394
rect -12633 42338 -12629 42394
rect -12693 42324 -12629 42338
rect -27082 42155 -26995 42179
rect -27082 42133 -27065 42155
rect -27013 42133 -26995 42155
rect -27082 42077 -27067 42133
rect -27011 42077 -26995 42133
rect -21475 42159 -21411 42173
rect -21475 42103 -21471 42159
rect -21415 42103 -21411 42159
rect -21475 42089 -21411 42103
rect -27082 42053 -27065 42077
rect -27013 42053 -26995 42077
rect -27082 41997 -27067 42053
rect -27011 41997 -26995 42053
rect -27082 41975 -27065 41997
rect -27013 41975 -26995 41997
rect -27082 41973 -26995 41975
rect -27082 41917 -27067 41973
rect -27011 41917 -26995 41973
rect -27082 41911 -27065 41917
rect -27013 41911 -26995 41917
rect -27082 41899 -26995 41911
rect -27082 41893 -27065 41899
rect -27013 41893 -26995 41899
rect -27082 41837 -27067 41893
rect -27011 41837 -26995 41893
rect -27082 41835 -26995 41837
rect -27082 41813 -27065 41835
rect -27013 41813 -26995 41835
rect -27082 41757 -27067 41813
rect -27011 41757 -26995 41813
rect -27082 41733 -27065 41757
rect -27013 41733 -26995 41757
rect -27082 41677 -27067 41733
rect -27011 41677 -26995 41733
rect -27082 41655 -27065 41677
rect -27013 41655 -26995 41677
rect -27082 41653 -26995 41655
rect -27082 41597 -27067 41653
rect -27011 41597 -26995 41653
rect -27082 41591 -27065 41597
rect -27013 41591 -26995 41597
rect -27082 41579 -26995 41591
rect -27082 41573 -27065 41579
rect -27013 41573 -26995 41579
rect -27082 41517 -27067 41573
rect -27011 41517 -26995 41573
rect -27082 41515 -26995 41517
rect -27082 41493 -27065 41515
rect -27013 41493 -26995 41515
rect -27082 41437 -27067 41493
rect -27011 41437 -26995 41493
rect -27082 41413 -27065 41437
rect -27013 41413 -26995 41437
rect -27082 41357 -27067 41413
rect -27011 41357 -26995 41413
rect -27082 41335 -27065 41357
rect -27013 41335 -26995 41357
rect -27082 41333 -26995 41335
rect -27082 41277 -27067 41333
rect -27011 41277 -26995 41333
rect -27082 41271 -27065 41277
rect -27013 41271 -26995 41277
rect -27082 41259 -26995 41271
rect -27082 41253 -27065 41259
rect -27013 41253 -26995 41259
rect -27082 41197 -27067 41253
rect -27011 41197 -26995 41253
rect -27082 41195 -26995 41197
rect -27082 41173 -27065 41195
rect -27013 41173 -26995 41195
rect -27082 41117 -27067 41173
rect -27011 41117 -26995 41173
rect -27082 41093 -27065 41117
rect -27013 41093 -26995 41117
rect -27082 41037 -27067 41093
rect -27011 41037 -26995 41093
rect -27082 41015 -27065 41037
rect -27013 41015 -26995 41037
rect -27082 40992 -26995 41015
rect -27077 40629 -26990 40653
rect -27077 40607 -27060 40629
rect -27008 40607 -26990 40629
rect -27077 40551 -27062 40607
rect -27006 40551 -26990 40607
rect -27077 40527 -27060 40551
rect -27008 40527 -26990 40551
rect -27077 40471 -27062 40527
rect -27006 40471 -26990 40527
rect -27077 40449 -27060 40471
rect -27008 40449 -26990 40471
rect -27077 40447 -26990 40449
rect -27077 40391 -27062 40447
rect -27006 40391 -26990 40447
rect -27077 40385 -27060 40391
rect -27008 40385 -26990 40391
rect -27077 40373 -26990 40385
rect -27077 40367 -27060 40373
rect -27008 40367 -26990 40373
rect -27077 40311 -27062 40367
rect -27006 40311 -26990 40367
rect -27077 40309 -26990 40311
rect -27077 40287 -27060 40309
rect -27008 40287 -26990 40309
rect -27077 40231 -27062 40287
rect -27006 40231 -26990 40287
rect -27077 40207 -27060 40231
rect -27008 40207 -26990 40231
rect -27077 40151 -27062 40207
rect -27006 40151 -26990 40207
rect -27077 40129 -27060 40151
rect -27008 40129 -26990 40151
rect -27077 40127 -26990 40129
rect -27077 40071 -27062 40127
rect -27006 40071 -26990 40127
rect -27077 40065 -27060 40071
rect -27008 40065 -26990 40071
rect -27077 40053 -26990 40065
rect -27077 40047 -27060 40053
rect -27008 40047 -26990 40053
rect -27077 39991 -27062 40047
rect -27006 39991 -26990 40047
rect -27077 39989 -26990 39991
rect -27077 39967 -27060 39989
rect -27008 39967 -26990 39989
rect -27077 39911 -27062 39967
rect -27006 39911 -26990 39967
rect -27077 39887 -27060 39911
rect -27008 39887 -26990 39911
rect -27077 39831 -27062 39887
rect -27006 39831 -26990 39887
rect -27077 39809 -27060 39831
rect -27008 39809 -26990 39831
rect -27077 39807 -26990 39809
rect -27077 39751 -27062 39807
rect -27006 39751 -26990 39807
rect -27077 39745 -27060 39751
rect -27008 39745 -26990 39751
rect -27077 39733 -26990 39745
rect -27077 39727 -27060 39733
rect -27008 39727 -26990 39733
rect -9398 39799 -9270 50879
rect -6989 50929 -6861 53542
rect 347 53146 365 60802
rect 501 53146 519 60802
rect 347 53140 375 53146
rect 491 53140 519 53146
rect 347 53111 519 53140
rect 10177 60814 10551 60846
rect 10177 60812 10216 60814
rect 10512 60812 10551 60814
rect -6989 50877 -6983 50929
rect -6931 50877 -6919 50929
rect -6867 50877 -6861 50929
rect -8874 50772 -8780 50801
rect -8874 50716 -8855 50772
rect -8799 50716 -8780 50772
rect -8874 50706 -8780 50716
rect -8874 50692 -8853 50706
rect -8801 50692 -8780 50706
rect -8874 50636 -8855 50692
rect -8799 50636 -8780 50692
rect -8874 50612 -8853 50636
rect -8801 50612 -8780 50636
rect -8874 50556 -8855 50612
rect -8799 50556 -8780 50612
rect -8874 50532 -8853 50556
rect -8801 50532 -8780 50556
rect -8874 50476 -8855 50532
rect -8799 50476 -8780 50532
rect -8874 50462 -8853 50476
rect -8801 50462 -8780 50476
rect -8874 50452 -8780 50462
rect -8874 50396 -8855 50452
rect -8799 50396 -8780 50452
rect -8874 50368 -8780 50396
rect -8480 50437 -8416 50451
rect -8480 50381 -8476 50437
rect -8420 50381 -8416 50437
rect -8480 50367 -8416 50381
rect -9398 39747 -9392 39799
rect -9340 39747 -9328 39799
rect -9276 39747 -9270 39799
rect -9398 39728 -9270 39747
rect -6989 39799 -6861 50877
rect -5688 51064 -3888 51076
rect -5688 50884 -5678 51064
rect -3898 50884 -3888 51064
rect -3362 51053 -2536 51084
rect -3362 51043 -3337 51053
rect -2561 51043 -2536 51053
rect -3362 50927 -3359 51043
rect -2539 50927 -2536 51043
rect -3362 50917 -3337 50927
rect -2561 50917 -2536 50927
rect -3362 50886 -2536 50917
rect -1655 51043 -765 51074
rect -1655 51033 -1638 51043
rect -782 51033 -765 51043
rect -1655 50917 -1652 51033
rect -768 50917 -765 51033
rect -1655 50907 -1638 50917
rect -782 50907 -765 50917
rect -5688 50873 -3888 50884
rect -1655 50876 -765 50907
rect -78 50771 121 50784
rect -78 50761 -47 50771
rect 89 50761 121 50771
rect -5932 50716 -5748 50730
rect -5932 50714 -5908 50716
rect -5772 50714 -5748 50716
rect -5932 47782 -5930 50714
rect -5750 47782 -5748 50714
rect -5932 47780 -5908 47782
rect -5772 47780 -5748 47782
rect -5932 47766 -5748 47780
rect -78 47765 -69 50761
rect 111 47765 121 50761
rect -78 47755 -47 47765
rect 89 47755 121 47765
rect -78 47742 121 47755
rect 10177 47640 10178 60812
rect 10550 47640 10551 60812
rect 17430 60738 17496 60753
rect 17430 60724 17437 60738
rect 17489 60724 17496 60738
rect 17430 60668 17435 60724
rect 17491 60668 17496 60724
rect 17430 60644 17437 60668
rect 17489 60644 17496 60668
rect 17430 60588 17435 60644
rect 17491 60588 17496 60644
rect 17430 60564 17437 60588
rect 17489 60564 17496 60588
rect 17430 60508 17435 60564
rect 17491 60508 17496 60564
rect 17430 60494 17437 60508
rect 17489 60494 17496 60508
rect 17430 60484 17496 60494
rect 17430 60428 17435 60484
rect 17491 60428 17496 60484
rect 17430 60418 17496 60428
rect 17430 60404 17437 60418
rect 17489 60404 17496 60418
rect 17430 60348 17435 60404
rect 17491 60348 17496 60404
rect 17430 60324 17437 60348
rect 17489 60324 17496 60348
rect 17430 60268 17435 60324
rect 17491 60268 17496 60324
rect 17430 60244 17437 60268
rect 17489 60244 17496 60268
rect 17430 60188 17435 60244
rect 17491 60188 17496 60244
rect 17430 60174 17437 60188
rect 17489 60174 17496 60188
rect 17430 60159 17496 60174
rect 18518 60738 18584 60753
rect 18518 60724 18525 60738
rect 18577 60724 18584 60738
rect 18518 60668 18523 60724
rect 18579 60668 18584 60724
rect 18518 60644 18525 60668
rect 18577 60644 18584 60668
rect 18518 60588 18523 60644
rect 18579 60588 18584 60644
rect 18518 60564 18525 60588
rect 18577 60564 18584 60588
rect 18518 60508 18523 60564
rect 18579 60508 18584 60564
rect 18518 60494 18525 60508
rect 18577 60494 18584 60508
rect 18518 60484 18584 60494
rect 18518 60428 18523 60484
rect 18579 60428 18584 60484
rect 18518 60418 18584 60428
rect 18518 60404 18525 60418
rect 18577 60404 18584 60418
rect 18518 60348 18523 60404
rect 18579 60348 18584 60404
rect 18518 60324 18525 60348
rect 18577 60324 18584 60348
rect 18518 60268 18523 60324
rect 18579 60268 18584 60324
rect 18518 60244 18525 60268
rect 18577 60244 18584 60268
rect 18518 60188 18523 60244
rect 18579 60188 18584 60244
rect 18518 60174 18525 60188
rect 18577 60174 18584 60188
rect 18518 60159 18584 60174
rect 19606 60738 19672 60753
rect 19606 60724 19613 60738
rect 19665 60724 19672 60738
rect 19606 60668 19611 60724
rect 19667 60668 19672 60724
rect 19606 60644 19613 60668
rect 19665 60644 19672 60668
rect 19606 60588 19611 60644
rect 19667 60588 19672 60644
rect 19606 60564 19613 60588
rect 19665 60564 19672 60588
rect 19606 60508 19611 60564
rect 19667 60508 19672 60564
rect 19606 60494 19613 60508
rect 19665 60494 19672 60508
rect 19606 60484 19672 60494
rect 19606 60428 19611 60484
rect 19667 60428 19672 60484
rect 19606 60418 19672 60428
rect 19606 60404 19613 60418
rect 19665 60404 19672 60418
rect 19606 60348 19611 60404
rect 19667 60348 19672 60404
rect 19606 60324 19613 60348
rect 19665 60324 19672 60348
rect 19606 60268 19611 60324
rect 19667 60268 19672 60324
rect 19606 60244 19613 60268
rect 19665 60244 19672 60268
rect 19606 60188 19611 60244
rect 19667 60188 19672 60244
rect 19606 60174 19613 60188
rect 19665 60174 19672 60188
rect 19606 60159 19672 60174
rect 20694 60738 20760 60753
rect 20694 60724 20701 60738
rect 20753 60724 20760 60738
rect 20694 60668 20699 60724
rect 20755 60668 20760 60724
rect 20694 60644 20701 60668
rect 20753 60644 20760 60668
rect 20694 60588 20699 60644
rect 20755 60588 20760 60644
rect 20694 60564 20701 60588
rect 20753 60564 20760 60588
rect 20694 60508 20699 60564
rect 20755 60508 20760 60564
rect 20694 60494 20701 60508
rect 20753 60494 20760 60508
rect 20694 60484 20760 60494
rect 20694 60428 20699 60484
rect 20755 60428 20760 60484
rect 20694 60418 20760 60428
rect 20694 60404 20701 60418
rect 20753 60404 20760 60418
rect 20694 60348 20699 60404
rect 20755 60348 20760 60404
rect 20694 60324 20701 60348
rect 20753 60324 20760 60348
rect 20694 60268 20699 60324
rect 20755 60268 20760 60324
rect 20694 60244 20701 60268
rect 20753 60244 20760 60268
rect 20694 60188 20699 60244
rect 20755 60188 20760 60244
rect 20694 60174 20701 60188
rect 20753 60174 20760 60188
rect 20694 60159 20760 60174
rect 21782 60738 21848 60753
rect 21782 60724 21789 60738
rect 21841 60724 21848 60738
rect 21782 60668 21787 60724
rect 21843 60668 21848 60724
rect 21782 60644 21789 60668
rect 21841 60644 21848 60668
rect 21782 60588 21787 60644
rect 21843 60588 21848 60644
rect 21782 60564 21789 60588
rect 21841 60564 21848 60588
rect 21782 60508 21787 60564
rect 21843 60508 21848 60564
rect 21782 60494 21789 60508
rect 21841 60494 21848 60508
rect 21782 60484 21848 60494
rect 21782 60428 21787 60484
rect 21843 60428 21848 60484
rect 21782 60418 21848 60428
rect 21782 60404 21789 60418
rect 21841 60404 21848 60418
rect 21782 60348 21787 60404
rect 21843 60348 21848 60404
rect 21782 60324 21789 60348
rect 21841 60324 21848 60348
rect 21782 60268 21787 60324
rect 21843 60268 21848 60324
rect 21782 60244 21789 60268
rect 21841 60244 21848 60268
rect 21782 60188 21787 60244
rect 21843 60188 21848 60244
rect 21782 60174 21789 60188
rect 21841 60174 21848 60188
rect 21782 60159 21848 60174
rect 22870 60738 22936 60753
rect 22870 60724 22877 60738
rect 22929 60724 22936 60738
rect 22870 60668 22875 60724
rect 22931 60668 22936 60724
rect 22870 60644 22877 60668
rect 22929 60644 22936 60668
rect 22870 60588 22875 60644
rect 22931 60588 22936 60644
rect 22870 60564 22877 60588
rect 22929 60564 22936 60588
rect 22870 60508 22875 60564
rect 22931 60508 22936 60564
rect 22870 60494 22877 60508
rect 22929 60494 22936 60508
rect 22870 60484 22936 60494
rect 22870 60428 22875 60484
rect 22931 60428 22936 60484
rect 22870 60418 22936 60428
rect 22870 60404 22877 60418
rect 22929 60404 22936 60418
rect 22870 60348 22875 60404
rect 22931 60348 22936 60404
rect 22870 60324 22877 60348
rect 22929 60324 22936 60348
rect 22870 60268 22875 60324
rect 22931 60268 22936 60324
rect 22870 60244 22877 60268
rect 22929 60244 22936 60268
rect 22870 60188 22875 60244
rect 22931 60188 22936 60244
rect 22870 60174 22877 60188
rect 22929 60174 22936 60188
rect 22870 60159 22936 60174
rect 23958 60738 24024 60753
rect 23958 60724 23965 60738
rect 24017 60724 24024 60738
rect 23958 60668 23963 60724
rect 24019 60668 24024 60724
rect 23958 60644 23965 60668
rect 24017 60644 24024 60668
rect 23958 60588 23963 60644
rect 24019 60588 24024 60644
rect 23958 60564 23965 60588
rect 24017 60564 24024 60588
rect 23958 60508 23963 60564
rect 24019 60508 24024 60564
rect 23958 60494 23965 60508
rect 24017 60494 24024 60508
rect 23958 60484 24024 60494
rect 23958 60428 23963 60484
rect 24019 60428 24024 60484
rect 23958 60418 24024 60428
rect 23958 60404 23965 60418
rect 24017 60404 24024 60418
rect 23958 60348 23963 60404
rect 24019 60348 24024 60404
rect 23958 60324 23965 60348
rect 24017 60324 24024 60348
rect 23958 60268 23963 60324
rect 24019 60268 24024 60324
rect 23958 60244 23965 60268
rect 24017 60244 24024 60268
rect 23958 60188 23963 60244
rect 24019 60188 24024 60244
rect 23958 60174 23965 60188
rect 24017 60174 24024 60188
rect 23958 60159 24024 60174
rect 25046 60738 25112 60753
rect 25046 60724 25053 60738
rect 25105 60724 25112 60738
rect 25046 60668 25051 60724
rect 25107 60668 25112 60724
rect 25046 60644 25053 60668
rect 25105 60644 25112 60668
rect 25046 60588 25051 60644
rect 25107 60588 25112 60644
rect 25046 60564 25053 60588
rect 25105 60564 25112 60588
rect 25046 60508 25051 60564
rect 25107 60508 25112 60564
rect 25046 60494 25053 60508
rect 25105 60494 25112 60508
rect 25046 60484 25112 60494
rect 25046 60428 25051 60484
rect 25107 60428 25112 60484
rect 25046 60418 25112 60428
rect 25046 60404 25053 60418
rect 25105 60404 25112 60418
rect 25046 60348 25051 60404
rect 25107 60348 25112 60404
rect 25046 60324 25053 60348
rect 25105 60324 25112 60348
rect 25046 60268 25051 60324
rect 25107 60268 25112 60324
rect 25046 60244 25053 60268
rect 25105 60244 25112 60268
rect 25046 60188 25051 60244
rect 25107 60188 25112 60244
rect 25046 60174 25053 60188
rect 25105 60174 25112 60188
rect 25046 60159 25112 60174
rect 26134 60738 26200 60753
rect 26134 60724 26141 60738
rect 26193 60724 26200 60738
rect 26134 60668 26139 60724
rect 26195 60668 26200 60724
rect 26134 60644 26141 60668
rect 26193 60644 26200 60668
rect 26134 60588 26139 60644
rect 26195 60588 26200 60644
rect 26134 60564 26141 60588
rect 26193 60564 26200 60588
rect 26134 60508 26139 60564
rect 26195 60508 26200 60564
rect 26134 60494 26141 60508
rect 26193 60494 26200 60508
rect 26134 60484 26200 60494
rect 26134 60428 26139 60484
rect 26195 60428 26200 60484
rect 26134 60418 26200 60428
rect 26134 60404 26141 60418
rect 26193 60404 26200 60418
rect 26134 60348 26139 60404
rect 26195 60348 26200 60404
rect 26134 60324 26141 60348
rect 26193 60324 26200 60348
rect 26134 60268 26139 60324
rect 26195 60268 26200 60324
rect 26134 60244 26141 60268
rect 26193 60244 26200 60268
rect 26134 60188 26139 60244
rect 26195 60188 26200 60244
rect 26134 60174 26141 60188
rect 26193 60174 26200 60188
rect 26134 60159 26200 60174
rect 27222 60738 27288 60753
rect 27222 60724 27229 60738
rect 27281 60724 27288 60738
rect 27222 60668 27227 60724
rect 27283 60668 27288 60724
rect 27222 60644 27229 60668
rect 27281 60644 27288 60668
rect 27222 60588 27227 60644
rect 27283 60588 27288 60644
rect 27222 60564 27229 60588
rect 27281 60564 27288 60588
rect 27222 60508 27227 60564
rect 27283 60508 27288 60564
rect 27222 60494 27229 60508
rect 27281 60494 27288 60508
rect 27222 60484 27288 60494
rect 27222 60428 27227 60484
rect 27283 60428 27288 60484
rect 27222 60418 27288 60428
rect 27222 60404 27229 60418
rect 27281 60404 27288 60418
rect 27222 60348 27227 60404
rect 27283 60348 27288 60404
rect 27222 60324 27229 60348
rect 27281 60324 27288 60348
rect 27222 60268 27227 60324
rect 27283 60268 27288 60324
rect 27222 60244 27229 60268
rect 27281 60244 27288 60268
rect 27222 60188 27227 60244
rect 27283 60188 27288 60244
rect 27222 60174 27229 60188
rect 27281 60174 27288 60188
rect 27222 60159 27288 60174
rect 28310 60738 28376 60753
rect 28310 60724 28317 60738
rect 28369 60724 28376 60738
rect 28310 60668 28315 60724
rect 28371 60668 28376 60724
rect 28310 60644 28317 60668
rect 28369 60644 28376 60668
rect 28310 60588 28315 60644
rect 28371 60588 28376 60644
rect 28310 60564 28317 60588
rect 28369 60564 28376 60588
rect 28310 60508 28315 60564
rect 28371 60508 28376 60564
rect 28310 60494 28317 60508
rect 28369 60494 28376 60508
rect 28310 60484 28376 60494
rect 28310 60428 28315 60484
rect 28371 60428 28376 60484
rect 28310 60418 28376 60428
rect 28310 60404 28317 60418
rect 28369 60404 28376 60418
rect 28310 60348 28315 60404
rect 28371 60348 28376 60404
rect 28310 60324 28317 60348
rect 28369 60324 28376 60348
rect 28310 60268 28315 60324
rect 28371 60268 28376 60324
rect 28310 60244 28317 60268
rect 28369 60244 28376 60268
rect 28310 60188 28315 60244
rect 28371 60188 28376 60244
rect 28310 60174 28317 60188
rect 28369 60174 28376 60188
rect 28310 60159 28376 60174
rect 29398 60738 29464 60753
rect 29398 60724 29405 60738
rect 29457 60724 29464 60738
rect 29398 60668 29403 60724
rect 29459 60668 29464 60724
rect 29398 60644 29405 60668
rect 29457 60644 29464 60668
rect 29398 60588 29403 60644
rect 29459 60588 29464 60644
rect 29398 60564 29405 60588
rect 29457 60564 29464 60588
rect 29398 60508 29403 60564
rect 29459 60508 29464 60564
rect 29398 60494 29405 60508
rect 29457 60494 29464 60508
rect 29398 60484 29464 60494
rect 29398 60428 29403 60484
rect 29459 60428 29464 60484
rect 29398 60418 29464 60428
rect 29398 60404 29405 60418
rect 29457 60404 29464 60418
rect 29398 60348 29403 60404
rect 29459 60348 29464 60404
rect 29398 60324 29405 60348
rect 29457 60324 29464 60348
rect 29398 60268 29403 60324
rect 29459 60268 29464 60324
rect 29398 60244 29405 60268
rect 29457 60244 29464 60268
rect 29398 60188 29403 60244
rect 29459 60188 29464 60244
rect 29398 60174 29405 60188
rect 29457 60174 29464 60188
rect 29398 60159 29464 60174
rect 30486 60738 30552 60753
rect 30486 60724 30493 60738
rect 30545 60724 30552 60738
rect 30486 60668 30491 60724
rect 30547 60668 30552 60724
rect 30486 60644 30493 60668
rect 30545 60644 30552 60668
rect 30486 60588 30491 60644
rect 30547 60588 30552 60644
rect 30486 60564 30493 60588
rect 30545 60564 30552 60588
rect 30486 60508 30491 60564
rect 30547 60508 30552 60564
rect 30486 60494 30493 60508
rect 30545 60494 30552 60508
rect 30486 60484 30552 60494
rect 30486 60428 30491 60484
rect 30547 60428 30552 60484
rect 30486 60418 30552 60428
rect 30486 60404 30493 60418
rect 30545 60404 30552 60418
rect 30486 60348 30491 60404
rect 30547 60348 30552 60404
rect 30486 60324 30493 60348
rect 30545 60324 30552 60348
rect 30486 60268 30491 60324
rect 30547 60268 30552 60324
rect 30486 60244 30493 60268
rect 30545 60244 30552 60268
rect 30486 60188 30491 60244
rect 30547 60188 30552 60244
rect 30486 60174 30493 60188
rect 30545 60174 30552 60188
rect 30486 60159 30552 60174
rect 31574 60738 31640 60753
rect 31574 60724 31581 60738
rect 31633 60724 31640 60738
rect 31574 60668 31579 60724
rect 31635 60668 31640 60724
rect 31574 60644 31581 60668
rect 31633 60644 31640 60668
rect 31574 60588 31579 60644
rect 31635 60588 31640 60644
rect 31574 60564 31581 60588
rect 31633 60564 31640 60588
rect 31574 60508 31579 60564
rect 31635 60508 31640 60564
rect 31574 60494 31581 60508
rect 31633 60494 31640 60508
rect 31574 60484 31640 60494
rect 31574 60428 31579 60484
rect 31635 60428 31640 60484
rect 31574 60418 31640 60428
rect 31574 60404 31581 60418
rect 31633 60404 31640 60418
rect 31574 60348 31579 60404
rect 31635 60348 31640 60404
rect 31574 60324 31581 60348
rect 31633 60324 31640 60348
rect 31574 60268 31579 60324
rect 31635 60268 31640 60324
rect 31574 60244 31581 60268
rect 31633 60244 31640 60268
rect 31574 60188 31579 60244
rect 31635 60188 31640 60244
rect 31574 60174 31581 60188
rect 31633 60174 31640 60188
rect 31574 60159 31640 60174
rect 17975 58735 18041 58750
rect 17975 58721 17982 58735
rect 18034 58721 18041 58735
rect 17975 58665 17980 58721
rect 18036 58665 18041 58721
rect 17975 58641 17982 58665
rect 18034 58641 18041 58665
rect 17975 58585 17980 58641
rect 18036 58585 18041 58641
rect 17975 58561 17982 58585
rect 18034 58561 18041 58585
rect 17975 58505 17980 58561
rect 18036 58505 18041 58561
rect 17975 58491 17982 58505
rect 18034 58491 18041 58505
rect 17975 58481 18041 58491
rect 17975 58425 17980 58481
rect 18036 58425 18041 58481
rect 17975 58415 18041 58425
rect 17975 58401 17982 58415
rect 18034 58401 18041 58415
rect 17975 58345 17980 58401
rect 18036 58345 18041 58401
rect 17975 58321 17982 58345
rect 18034 58321 18041 58345
rect 17975 58265 17980 58321
rect 18036 58265 18041 58321
rect 17975 58241 17982 58265
rect 18034 58241 18041 58265
rect 17975 58185 17980 58241
rect 18036 58185 18041 58241
rect 17975 58171 17982 58185
rect 18034 58171 18041 58185
rect 17975 58156 18041 58171
rect 19063 58735 19129 58750
rect 19063 58721 19070 58735
rect 19122 58721 19129 58735
rect 19063 58665 19068 58721
rect 19124 58665 19129 58721
rect 19063 58641 19070 58665
rect 19122 58641 19129 58665
rect 19063 58585 19068 58641
rect 19124 58585 19129 58641
rect 19063 58561 19070 58585
rect 19122 58561 19129 58585
rect 19063 58505 19068 58561
rect 19124 58505 19129 58561
rect 19063 58491 19070 58505
rect 19122 58491 19129 58505
rect 19063 58481 19129 58491
rect 19063 58425 19068 58481
rect 19124 58425 19129 58481
rect 19063 58415 19129 58425
rect 19063 58401 19070 58415
rect 19122 58401 19129 58415
rect 19063 58345 19068 58401
rect 19124 58345 19129 58401
rect 19063 58321 19070 58345
rect 19122 58321 19129 58345
rect 19063 58265 19068 58321
rect 19124 58265 19129 58321
rect 19063 58241 19070 58265
rect 19122 58241 19129 58265
rect 19063 58185 19068 58241
rect 19124 58185 19129 58241
rect 19063 58171 19070 58185
rect 19122 58171 19129 58185
rect 19063 58156 19129 58171
rect 20151 58735 20217 58750
rect 20151 58721 20158 58735
rect 20210 58721 20217 58735
rect 20151 58665 20156 58721
rect 20212 58665 20217 58721
rect 20151 58641 20158 58665
rect 20210 58641 20217 58665
rect 20151 58585 20156 58641
rect 20212 58585 20217 58641
rect 20151 58561 20158 58585
rect 20210 58561 20217 58585
rect 20151 58505 20156 58561
rect 20212 58505 20217 58561
rect 20151 58491 20158 58505
rect 20210 58491 20217 58505
rect 20151 58481 20217 58491
rect 20151 58425 20156 58481
rect 20212 58425 20217 58481
rect 20151 58415 20217 58425
rect 20151 58401 20158 58415
rect 20210 58401 20217 58415
rect 20151 58345 20156 58401
rect 20212 58345 20217 58401
rect 20151 58321 20158 58345
rect 20210 58321 20217 58345
rect 20151 58265 20156 58321
rect 20212 58265 20217 58321
rect 20151 58241 20158 58265
rect 20210 58241 20217 58265
rect 20151 58185 20156 58241
rect 20212 58185 20217 58241
rect 20151 58171 20158 58185
rect 20210 58171 20217 58185
rect 20151 58156 20217 58171
rect 21239 58735 21305 58750
rect 21239 58721 21246 58735
rect 21298 58721 21305 58735
rect 21239 58665 21244 58721
rect 21300 58665 21305 58721
rect 21239 58641 21246 58665
rect 21298 58641 21305 58665
rect 21239 58585 21244 58641
rect 21300 58585 21305 58641
rect 21239 58561 21246 58585
rect 21298 58561 21305 58585
rect 21239 58505 21244 58561
rect 21300 58505 21305 58561
rect 21239 58491 21246 58505
rect 21298 58491 21305 58505
rect 21239 58481 21305 58491
rect 21239 58425 21244 58481
rect 21300 58425 21305 58481
rect 21239 58415 21305 58425
rect 21239 58401 21246 58415
rect 21298 58401 21305 58415
rect 21239 58345 21244 58401
rect 21300 58345 21305 58401
rect 21239 58321 21246 58345
rect 21298 58321 21305 58345
rect 21239 58265 21244 58321
rect 21300 58265 21305 58321
rect 21239 58241 21246 58265
rect 21298 58241 21305 58265
rect 21239 58185 21244 58241
rect 21300 58185 21305 58241
rect 21239 58171 21246 58185
rect 21298 58171 21305 58185
rect 21239 58156 21305 58171
rect 22327 58735 22393 58750
rect 22327 58721 22334 58735
rect 22386 58721 22393 58735
rect 22327 58665 22332 58721
rect 22388 58665 22393 58721
rect 22327 58641 22334 58665
rect 22386 58641 22393 58665
rect 22327 58585 22332 58641
rect 22388 58585 22393 58641
rect 22327 58561 22334 58585
rect 22386 58561 22393 58585
rect 22327 58505 22332 58561
rect 22388 58505 22393 58561
rect 22327 58491 22334 58505
rect 22386 58491 22393 58505
rect 22327 58481 22393 58491
rect 22327 58425 22332 58481
rect 22388 58425 22393 58481
rect 22327 58415 22393 58425
rect 22327 58401 22334 58415
rect 22386 58401 22393 58415
rect 22327 58345 22332 58401
rect 22388 58345 22393 58401
rect 22327 58321 22334 58345
rect 22386 58321 22393 58345
rect 22327 58265 22332 58321
rect 22388 58265 22393 58321
rect 22327 58241 22334 58265
rect 22386 58241 22393 58265
rect 22327 58185 22332 58241
rect 22388 58185 22393 58241
rect 22327 58171 22334 58185
rect 22386 58171 22393 58185
rect 22327 58156 22393 58171
rect 23415 58735 23481 58750
rect 23415 58721 23422 58735
rect 23474 58721 23481 58735
rect 23415 58665 23420 58721
rect 23476 58665 23481 58721
rect 23415 58641 23422 58665
rect 23474 58641 23481 58665
rect 23415 58585 23420 58641
rect 23476 58585 23481 58641
rect 23415 58561 23422 58585
rect 23474 58561 23481 58585
rect 23415 58505 23420 58561
rect 23476 58505 23481 58561
rect 23415 58491 23422 58505
rect 23474 58491 23481 58505
rect 23415 58481 23481 58491
rect 23415 58425 23420 58481
rect 23476 58425 23481 58481
rect 23415 58415 23481 58425
rect 23415 58401 23422 58415
rect 23474 58401 23481 58415
rect 23415 58345 23420 58401
rect 23476 58345 23481 58401
rect 23415 58321 23422 58345
rect 23474 58321 23481 58345
rect 23415 58265 23420 58321
rect 23476 58265 23481 58321
rect 23415 58241 23422 58265
rect 23474 58241 23481 58265
rect 23415 58185 23420 58241
rect 23476 58185 23481 58241
rect 23415 58171 23422 58185
rect 23474 58171 23481 58185
rect 23415 58156 23481 58171
rect 24503 58735 24569 58750
rect 24503 58721 24510 58735
rect 24562 58721 24569 58735
rect 24503 58665 24508 58721
rect 24564 58665 24569 58721
rect 24503 58641 24510 58665
rect 24562 58641 24569 58665
rect 24503 58585 24508 58641
rect 24564 58585 24569 58641
rect 24503 58561 24510 58585
rect 24562 58561 24569 58585
rect 24503 58505 24508 58561
rect 24564 58505 24569 58561
rect 24503 58491 24510 58505
rect 24562 58491 24569 58505
rect 24503 58481 24569 58491
rect 24503 58425 24508 58481
rect 24564 58425 24569 58481
rect 24503 58415 24569 58425
rect 24503 58401 24510 58415
rect 24562 58401 24569 58415
rect 24503 58345 24508 58401
rect 24564 58345 24569 58401
rect 24503 58321 24510 58345
rect 24562 58321 24569 58345
rect 24503 58265 24508 58321
rect 24564 58265 24569 58321
rect 24503 58241 24510 58265
rect 24562 58241 24569 58265
rect 24503 58185 24508 58241
rect 24564 58185 24569 58241
rect 24503 58171 24510 58185
rect 24562 58171 24569 58185
rect 24503 58156 24569 58171
rect 25591 58735 25657 58750
rect 25591 58721 25598 58735
rect 25650 58721 25657 58735
rect 25591 58665 25596 58721
rect 25652 58665 25657 58721
rect 25591 58641 25598 58665
rect 25650 58641 25657 58665
rect 25591 58585 25596 58641
rect 25652 58585 25657 58641
rect 25591 58561 25598 58585
rect 25650 58561 25657 58585
rect 25591 58505 25596 58561
rect 25652 58505 25657 58561
rect 25591 58491 25598 58505
rect 25650 58491 25657 58505
rect 25591 58481 25657 58491
rect 25591 58425 25596 58481
rect 25652 58425 25657 58481
rect 25591 58415 25657 58425
rect 25591 58401 25598 58415
rect 25650 58401 25657 58415
rect 25591 58345 25596 58401
rect 25652 58345 25657 58401
rect 25591 58321 25598 58345
rect 25650 58321 25657 58345
rect 25591 58265 25596 58321
rect 25652 58265 25657 58321
rect 25591 58241 25598 58265
rect 25650 58241 25657 58265
rect 25591 58185 25596 58241
rect 25652 58185 25657 58241
rect 25591 58171 25598 58185
rect 25650 58171 25657 58185
rect 25591 58156 25657 58171
rect 26679 58735 26745 58750
rect 26679 58721 26686 58735
rect 26738 58721 26745 58735
rect 26679 58665 26684 58721
rect 26740 58665 26745 58721
rect 26679 58641 26686 58665
rect 26738 58641 26745 58665
rect 26679 58585 26684 58641
rect 26740 58585 26745 58641
rect 26679 58561 26686 58585
rect 26738 58561 26745 58585
rect 26679 58505 26684 58561
rect 26740 58505 26745 58561
rect 26679 58491 26686 58505
rect 26738 58491 26745 58505
rect 26679 58481 26745 58491
rect 26679 58425 26684 58481
rect 26740 58425 26745 58481
rect 26679 58415 26745 58425
rect 26679 58401 26686 58415
rect 26738 58401 26745 58415
rect 26679 58345 26684 58401
rect 26740 58345 26745 58401
rect 26679 58321 26686 58345
rect 26738 58321 26745 58345
rect 26679 58265 26684 58321
rect 26740 58265 26745 58321
rect 26679 58241 26686 58265
rect 26738 58241 26745 58265
rect 26679 58185 26684 58241
rect 26740 58185 26745 58241
rect 26679 58171 26686 58185
rect 26738 58171 26745 58185
rect 26679 58156 26745 58171
rect 27767 58735 27833 58750
rect 27767 58721 27774 58735
rect 27826 58721 27833 58735
rect 27767 58665 27772 58721
rect 27828 58665 27833 58721
rect 27767 58641 27774 58665
rect 27826 58641 27833 58665
rect 27767 58585 27772 58641
rect 27828 58585 27833 58641
rect 27767 58561 27774 58585
rect 27826 58561 27833 58585
rect 27767 58505 27772 58561
rect 27828 58505 27833 58561
rect 27767 58491 27774 58505
rect 27826 58491 27833 58505
rect 27767 58481 27833 58491
rect 27767 58425 27772 58481
rect 27828 58425 27833 58481
rect 27767 58415 27833 58425
rect 27767 58401 27774 58415
rect 27826 58401 27833 58415
rect 27767 58345 27772 58401
rect 27828 58345 27833 58401
rect 27767 58321 27774 58345
rect 27826 58321 27833 58345
rect 27767 58265 27772 58321
rect 27828 58265 27833 58321
rect 27767 58241 27774 58265
rect 27826 58241 27833 58265
rect 27767 58185 27772 58241
rect 27828 58185 27833 58241
rect 27767 58171 27774 58185
rect 27826 58171 27833 58185
rect 27767 58156 27833 58171
rect 28855 58735 28921 58750
rect 28855 58721 28862 58735
rect 28914 58721 28921 58735
rect 28855 58665 28860 58721
rect 28916 58665 28921 58721
rect 28855 58641 28862 58665
rect 28914 58641 28921 58665
rect 28855 58585 28860 58641
rect 28916 58585 28921 58641
rect 28855 58561 28862 58585
rect 28914 58561 28921 58585
rect 28855 58505 28860 58561
rect 28916 58505 28921 58561
rect 28855 58491 28862 58505
rect 28914 58491 28921 58505
rect 28855 58481 28921 58491
rect 28855 58425 28860 58481
rect 28916 58425 28921 58481
rect 28855 58415 28921 58425
rect 28855 58401 28862 58415
rect 28914 58401 28921 58415
rect 28855 58345 28860 58401
rect 28916 58345 28921 58401
rect 28855 58321 28862 58345
rect 28914 58321 28921 58345
rect 28855 58265 28860 58321
rect 28916 58265 28921 58321
rect 28855 58241 28862 58265
rect 28914 58241 28921 58265
rect 28855 58185 28860 58241
rect 28916 58185 28921 58241
rect 28855 58171 28862 58185
rect 28914 58171 28921 58185
rect 28855 58156 28921 58171
rect 29943 58735 30009 58750
rect 29943 58721 29950 58735
rect 30002 58721 30009 58735
rect 29943 58665 29948 58721
rect 30004 58665 30009 58721
rect 29943 58641 29950 58665
rect 30002 58641 30009 58665
rect 29943 58585 29948 58641
rect 30004 58585 30009 58641
rect 29943 58561 29950 58585
rect 30002 58561 30009 58585
rect 29943 58505 29948 58561
rect 30004 58505 30009 58561
rect 29943 58491 29950 58505
rect 30002 58491 30009 58505
rect 29943 58481 30009 58491
rect 29943 58425 29948 58481
rect 30004 58425 30009 58481
rect 29943 58415 30009 58425
rect 29943 58401 29950 58415
rect 30002 58401 30009 58415
rect 29943 58345 29948 58401
rect 30004 58345 30009 58401
rect 29943 58321 29950 58345
rect 30002 58321 30009 58345
rect 29943 58265 29948 58321
rect 30004 58265 30009 58321
rect 29943 58241 29950 58265
rect 30002 58241 30009 58265
rect 29943 58185 29948 58241
rect 30004 58185 30009 58241
rect 29943 58171 29950 58185
rect 30002 58171 30009 58185
rect 29943 58156 30009 58171
rect 31031 58735 31097 58750
rect 31031 58721 31038 58735
rect 31090 58721 31097 58735
rect 31031 58665 31036 58721
rect 31092 58665 31097 58721
rect 31031 58641 31038 58665
rect 31090 58641 31097 58665
rect 31031 58585 31036 58641
rect 31092 58585 31097 58641
rect 31031 58561 31038 58585
rect 31090 58561 31097 58585
rect 31031 58505 31036 58561
rect 31092 58505 31097 58561
rect 31031 58491 31038 58505
rect 31090 58491 31097 58505
rect 31031 58481 31097 58491
rect 31031 58425 31036 58481
rect 31092 58425 31097 58481
rect 31031 58415 31097 58425
rect 31031 58401 31038 58415
rect 31090 58401 31097 58415
rect 31031 58345 31036 58401
rect 31092 58345 31097 58401
rect 31031 58321 31038 58345
rect 31090 58321 31097 58345
rect 31031 58265 31036 58321
rect 31092 58265 31097 58321
rect 31031 58241 31038 58265
rect 31090 58241 31097 58265
rect 31031 58185 31036 58241
rect 31092 58185 31097 58241
rect 31031 58171 31038 58185
rect 31090 58171 31097 58185
rect 31031 58156 31097 58171
rect 17430 56738 17496 56753
rect 17430 56724 17437 56738
rect 17489 56724 17496 56738
rect 17430 56668 17435 56724
rect 17491 56668 17496 56724
rect 17430 56644 17437 56668
rect 17489 56644 17496 56668
rect 17430 56588 17435 56644
rect 17491 56588 17496 56644
rect 17430 56564 17437 56588
rect 17489 56564 17496 56588
rect 17430 56508 17435 56564
rect 17491 56508 17496 56564
rect 17430 56494 17437 56508
rect 17489 56494 17496 56508
rect 17430 56484 17496 56494
rect 17430 56428 17435 56484
rect 17491 56428 17496 56484
rect 17430 56418 17496 56428
rect 17430 56404 17437 56418
rect 17489 56404 17496 56418
rect 17430 56348 17435 56404
rect 17491 56348 17496 56404
rect 17430 56324 17437 56348
rect 17489 56324 17496 56348
rect 17430 56268 17435 56324
rect 17491 56268 17496 56324
rect 17430 56244 17437 56268
rect 17489 56244 17496 56268
rect 17430 56188 17435 56244
rect 17491 56188 17496 56244
rect 17430 56174 17437 56188
rect 17489 56174 17496 56188
rect 17430 56159 17496 56174
rect 18518 56738 18584 56753
rect 18518 56724 18525 56738
rect 18577 56724 18584 56738
rect 18518 56668 18523 56724
rect 18579 56668 18584 56724
rect 18518 56644 18525 56668
rect 18577 56644 18584 56668
rect 18518 56588 18523 56644
rect 18579 56588 18584 56644
rect 18518 56564 18525 56588
rect 18577 56564 18584 56588
rect 18518 56508 18523 56564
rect 18579 56508 18584 56564
rect 18518 56494 18525 56508
rect 18577 56494 18584 56508
rect 18518 56484 18584 56494
rect 18518 56428 18523 56484
rect 18579 56428 18584 56484
rect 18518 56418 18584 56428
rect 18518 56404 18525 56418
rect 18577 56404 18584 56418
rect 18518 56348 18523 56404
rect 18579 56348 18584 56404
rect 18518 56324 18525 56348
rect 18577 56324 18584 56348
rect 18518 56268 18523 56324
rect 18579 56268 18584 56324
rect 18518 56244 18525 56268
rect 18577 56244 18584 56268
rect 18518 56188 18523 56244
rect 18579 56188 18584 56244
rect 18518 56174 18525 56188
rect 18577 56174 18584 56188
rect 18518 56159 18584 56174
rect 19606 56738 19672 56753
rect 19606 56724 19613 56738
rect 19665 56724 19672 56738
rect 19606 56668 19611 56724
rect 19667 56668 19672 56724
rect 19606 56644 19613 56668
rect 19665 56644 19672 56668
rect 19606 56588 19611 56644
rect 19667 56588 19672 56644
rect 19606 56564 19613 56588
rect 19665 56564 19672 56588
rect 19606 56508 19611 56564
rect 19667 56508 19672 56564
rect 19606 56494 19613 56508
rect 19665 56494 19672 56508
rect 19606 56484 19672 56494
rect 19606 56428 19611 56484
rect 19667 56428 19672 56484
rect 19606 56418 19672 56428
rect 19606 56404 19613 56418
rect 19665 56404 19672 56418
rect 19606 56348 19611 56404
rect 19667 56348 19672 56404
rect 19606 56324 19613 56348
rect 19665 56324 19672 56348
rect 19606 56268 19611 56324
rect 19667 56268 19672 56324
rect 19606 56244 19613 56268
rect 19665 56244 19672 56268
rect 19606 56188 19611 56244
rect 19667 56188 19672 56244
rect 19606 56174 19613 56188
rect 19665 56174 19672 56188
rect 19606 56159 19672 56174
rect 20694 56738 20760 56753
rect 20694 56724 20701 56738
rect 20753 56724 20760 56738
rect 20694 56668 20699 56724
rect 20755 56668 20760 56724
rect 20694 56644 20701 56668
rect 20753 56644 20760 56668
rect 20694 56588 20699 56644
rect 20755 56588 20760 56644
rect 20694 56564 20701 56588
rect 20753 56564 20760 56588
rect 20694 56508 20699 56564
rect 20755 56508 20760 56564
rect 20694 56494 20701 56508
rect 20753 56494 20760 56508
rect 20694 56484 20760 56494
rect 20694 56428 20699 56484
rect 20755 56428 20760 56484
rect 20694 56418 20760 56428
rect 20694 56404 20701 56418
rect 20753 56404 20760 56418
rect 20694 56348 20699 56404
rect 20755 56348 20760 56404
rect 20694 56324 20701 56348
rect 20753 56324 20760 56348
rect 20694 56268 20699 56324
rect 20755 56268 20760 56324
rect 20694 56244 20701 56268
rect 20753 56244 20760 56268
rect 20694 56188 20699 56244
rect 20755 56188 20760 56244
rect 20694 56174 20701 56188
rect 20753 56174 20760 56188
rect 20694 56159 20760 56174
rect 21782 56738 21848 56753
rect 21782 56724 21789 56738
rect 21841 56724 21848 56738
rect 21782 56668 21787 56724
rect 21843 56668 21848 56724
rect 21782 56644 21789 56668
rect 21841 56644 21848 56668
rect 21782 56588 21787 56644
rect 21843 56588 21848 56644
rect 21782 56564 21789 56588
rect 21841 56564 21848 56588
rect 21782 56508 21787 56564
rect 21843 56508 21848 56564
rect 21782 56494 21789 56508
rect 21841 56494 21848 56508
rect 21782 56484 21848 56494
rect 21782 56428 21787 56484
rect 21843 56428 21848 56484
rect 21782 56418 21848 56428
rect 21782 56404 21789 56418
rect 21841 56404 21848 56418
rect 21782 56348 21787 56404
rect 21843 56348 21848 56404
rect 21782 56324 21789 56348
rect 21841 56324 21848 56348
rect 21782 56268 21787 56324
rect 21843 56268 21848 56324
rect 21782 56244 21789 56268
rect 21841 56244 21848 56268
rect 21782 56188 21787 56244
rect 21843 56188 21848 56244
rect 21782 56174 21789 56188
rect 21841 56174 21848 56188
rect 21782 56159 21848 56174
rect 22870 56738 22936 56753
rect 22870 56724 22877 56738
rect 22929 56724 22936 56738
rect 22870 56668 22875 56724
rect 22931 56668 22936 56724
rect 22870 56644 22877 56668
rect 22929 56644 22936 56668
rect 22870 56588 22875 56644
rect 22931 56588 22936 56644
rect 22870 56564 22877 56588
rect 22929 56564 22936 56588
rect 22870 56508 22875 56564
rect 22931 56508 22936 56564
rect 22870 56494 22877 56508
rect 22929 56494 22936 56508
rect 22870 56484 22936 56494
rect 22870 56428 22875 56484
rect 22931 56428 22936 56484
rect 22870 56418 22936 56428
rect 22870 56404 22877 56418
rect 22929 56404 22936 56418
rect 22870 56348 22875 56404
rect 22931 56348 22936 56404
rect 22870 56324 22877 56348
rect 22929 56324 22936 56348
rect 22870 56268 22875 56324
rect 22931 56268 22936 56324
rect 22870 56244 22877 56268
rect 22929 56244 22936 56268
rect 22870 56188 22875 56244
rect 22931 56188 22936 56244
rect 22870 56174 22877 56188
rect 22929 56174 22936 56188
rect 22870 56159 22936 56174
rect 23958 56738 24024 56753
rect 23958 56724 23965 56738
rect 24017 56724 24024 56738
rect 23958 56668 23963 56724
rect 24019 56668 24024 56724
rect 23958 56644 23965 56668
rect 24017 56644 24024 56668
rect 23958 56588 23963 56644
rect 24019 56588 24024 56644
rect 23958 56564 23965 56588
rect 24017 56564 24024 56588
rect 23958 56508 23963 56564
rect 24019 56508 24024 56564
rect 23958 56494 23965 56508
rect 24017 56494 24024 56508
rect 23958 56484 24024 56494
rect 23958 56428 23963 56484
rect 24019 56428 24024 56484
rect 23958 56418 24024 56428
rect 23958 56404 23965 56418
rect 24017 56404 24024 56418
rect 23958 56348 23963 56404
rect 24019 56348 24024 56404
rect 23958 56324 23965 56348
rect 24017 56324 24024 56348
rect 23958 56268 23963 56324
rect 24019 56268 24024 56324
rect 23958 56244 23965 56268
rect 24017 56244 24024 56268
rect 23958 56188 23963 56244
rect 24019 56188 24024 56244
rect 23958 56174 23965 56188
rect 24017 56174 24024 56188
rect 23958 56159 24024 56174
rect 25046 56738 25112 56753
rect 25046 56724 25053 56738
rect 25105 56724 25112 56738
rect 25046 56668 25051 56724
rect 25107 56668 25112 56724
rect 25046 56644 25053 56668
rect 25105 56644 25112 56668
rect 25046 56588 25051 56644
rect 25107 56588 25112 56644
rect 25046 56564 25053 56588
rect 25105 56564 25112 56588
rect 25046 56508 25051 56564
rect 25107 56508 25112 56564
rect 25046 56494 25053 56508
rect 25105 56494 25112 56508
rect 25046 56484 25112 56494
rect 25046 56428 25051 56484
rect 25107 56428 25112 56484
rect 25046 56418 25112 56428
rect 25046 56404 25053 56418
rect 25105 56404 25112 56418
rect 25046 56348 25051 56404
rect 25107 56348 25112 56404
rect 25046 56324 25053 56348
rect 25105 56324 25112 56348
rect 25046 56268 25051 56324
rect 25107 56268 25112 56324
rect 25046 56244 25053 56268
rect 25105 56244 25112 56268
rect 25046 56188 25051 56244
rect 25107 56188 25112 56244
rect 25046 56174 25053 56188
rect 25105 56174 25112 56188
rect 25046 56159 25112 56174
rect 26134 56738 26200 56753
rect 26134 56724 26141 56738
rect 26193 56724 26200 56738
rect 26134 56668 26139 56724
rect 26195 56668 26200 56724
rect 26134 56644 26141 56668
rect 26193 56644 26200 56668
rect 26134 56588 26139 56644
rect 26195 56588 26200 56644
rect 26134 56564 26141 56588
rect 26193 56564 26200 56588
rect 26134 56508 26139 56564
rect 26195 56508 26200 56564
rect 26134 56494 26141 56508
rect 26193 56494 26200 56508
rect 26134 56484 26200 56494
rect 26134 56428 26139 56484
rect 26195 56428 26200 56484
rect 26134 56418 26200 56428
rect 26134 56404 26141 56418
rect 26193 56404 26200 56418
rect 26134 56348 26139 56404
rect 26195 56348 26200 56404
rect 26134 56324 26141 56348
rect 26193 56324 26200 56348
rect 26134 56268 26139 56324
rect 26195 56268 26200 56324
rect 26134 56244 26141 56268
rect 26193 56244 26200 56268
rect 26134 56188 26139 56244
rect 26195 56188 26200 56244
rect 26134 56174 26141 56188
rect 26193 56174 26200 56188
rect 26134 56159 26200 56174
rect 27222 56738 27288 56753
rect 27222 56724 27229 56738
rect 27281 56724 27288 56738
rect 27222 56668 27227 56724
rect 27283 56668 27288 56724
rect 27222 56644 27229 56668
rect 27281 56644 27288 56668
rect 27222 56588 27227 56644
rect 27283 56588 27288 56644
rect 27222 56564 27229 56588
rect 27281 56564 27288 56588
rect 27222 56508 27227 56564
rect 27283 56508 27288 56564
rect 27222 56494 27229 56508
rect 27281 56494 27288 56508
rect 27222 56484 27288 56494
rect 27222 56428 27227 56484
rect 27283 56428 27288 56484
rect 27222 56418 27288 56428
rect 27222 56404 27229 56418
rect 27281 56404 27288 56418
rect 27222 56348 27227 56404
rect 27283 56348 27288 56404
rect 27222 56324 27229 56348
rect 27281 56324 27288 56348
rect 27222 56268 27227 56324
rect 27283 56268 27288 56324
rect 27222 56244 27229 56268
rect 27281 56244 27288 56268
rect 27222 56188 27227 56244
rect 27283 56188 27288 56244
rect 27222 56174 27229 56188
rect 27281 56174 27288 56188
rect 27222 56159 27288 56174
rect 28310 56738 28376 56753
rect 28310 56724 28317 56738
rect 28369 56724 28376 56738
rect 28310 56668 28315 56724
rect 28371 56668 28376 56724
rect 28310 56644 28317 56668
rect 28369 56644 28376 56668
rect 28310 56588 28315 56644
rect 28371 56588 28376 56644
rect 28310 56564 28317 56588
rect 28369 56564 28376 56588
rect 28310 56508 28315 56564
rect 28371 56508 28376 56564
rect 28310 56494 28317 56508
rect 28369 56494 28376 56508
rect 28310 56484 28376 56494
rect 28310 56428 28315 56484
rect 28371 56428 28376 56484
rect 28310 56418 28376 56428
rect 28310 56404 28317 56418
rect 28369 56404 28376 56418
rect 28310 56348 28315 56404
rect 28371 56348 28376 56404
rect 28310 56324 28317 56348
rect 28369 56324 28376 56348
rect 28310 56268 28315 56324
rect 28371 56268 28376 56324
rect 28310 56244 28317 56268
rect 28369 56244 28376 56268
rect 28310 56188 28315 56244
rect 28371 56188 28376 56244
rect 28310 56174 28317 56188
rect 28369 56174 28376 56188
rect 28310 56159 28376 56174
rect 29398 56738 29464 56753
rect 29398 56724 29405 56738
rect 29457 56724 29464 56738
rect 29398 56668 29403 56724
rect 29459 56668 29464 56724
rect 29398 56644 29405 56668
rect 29457 56644 29464 56668
rect 29398 56588 29403 56644
rect 29459 56588 29464 56644
rect 29398 56564 29405 56588
rect 29457 56564 29464 56588
rect 29398 56508 29403 56564
rect 29459 56508 29464 56564
rect 29398 56494 29405 56508
rect 29457 56494 29464 56508
rect 29398 56484 29464 56494
rect 29398 56428 29403 56484
rect 29459 56428 29464 56484
rect 29398 56418 29464 56428
rect 29398 56404 29405 56418
rect 29457 56404 29464 56418
rect 29398 56348 29403 56404
rect 29459 56348 29464 56404
rect 29398 56324 29405 56348
rect 29457 56324 29464 56348
rect 29398 56268 29403 56324
rect 29459 56268 29464 56324
rect 29398 56244 29405 56268
rect 29457 56244 29464 56268
rect 29398 56188 29403 56244
rect 29459 56188 29464 56244
rect 29398 56174 29405 56188
rect 29457 56174 29464 56188
rect 29398 56159 29464 56174
rect 30486 56738 30552 56753
rect 30486 56724 30493 56738
rect 30545 56724 30552 56738
rect 30486 56668 30491 56724
rect 30547 56668 30552 56724
rect 30486 56644 30493 56668
rect 30545 56644 30552 56668
rect 30486 56588 30491 56644
rect 30547 56588 30552 56644
rect 30486 56564 30493 56588
rect 30545 56564 30552 56588
rect 30486 56508 30491 56564
rect 30547 56508 30552 56564
rect 30486 56494 30493 56508
rect 30545 56494 30552 56508
rect 30486 56484 30552 56494
rect 30486 56428 30491 56484
rect 30547 56428 30552 56484
rect 30486 56418 30552 56428
rect 30486 56404 30493 56418
rect 30545 56404 30552 56418
rect 30486 56348 30491 56404
rect 30547 56348 30552 56404
rect 30486 56324 30493 56348
rect 30545 56324 30552 56348
rect 30486 56268 30491 56324
rect 30547 56268 30552 56324
rect 30486 56244 30493 56268
rect 30545 56244 30552 56268
rect 30486 56188 30491 56244
rect 30547 56188 30552 56244
rect 30486 56174 30493 56188
rect 30545 56174 30552 56188
rect 30486 56159 30552 56174
rect 31574 56738 31640 56753
rect 31574 56724 31581 56738
rect 31633 56724 31640 56738
rect 31574 56668 31579 56724
rect 31635 56668 31640 56724
rect 31574 56644 31581 56668
rect 31633 56644 31640 56668
rect 31574 56588 31579 56644
rect 31635 56588 31640 56644
rect 31574 56564 31581 56588
rect 31633 56564 31640 56588
rect 31574 56508 31579 56564
rect 31635 56508 31640 56564
rect 31574 56494 31581 56508
rect 31633 56494 31640 56508
rect 31574 56484 31640 56494
rect 31574 56428 31579 56484
rect 31635 56428 31640 56484
rect 31574 56418 31640 56428
rect 31574 56404 31581 56418
rect 31633 56404 31640 56418
rect 31574 56348 31579 56404
rect 31635 56348 31640 56404
rect 31574 56324 31581 56348
rect 31633 56324 31640 56348
rect 31574 56268 31579 56324
rect 31635 56268 31640 56324
rect 31574 56244 31581 56268
rect 31633 56244 31640 56268
rect 31574 56188 31579 56244
rect 31635 56188 31640 56244
rect 31574 56174 31581 56188
rect 31633 56174 31640 56188
rect 31574 56159 31640 56174
rect 17975 54735 18041 54750
rect 17975 54721 17982 54735
rect 18034 54721 18041 54735
rect 17975 54665 17980 54721
rect 18036 54665 18041 54721
rect 17975 54641 17982 54665
rect 18034 54641 18041 54665
rect 17975 54585 17980 54641
rect 18036 54585 18041 54641
rect 17975 54561 17982 54585
rect 18034 54561 18041 54585
rect 17975 54505 17980 54561
rect 18036 54505 18041 54561
rect 17975 54491 17982 54505
rect 18034 54491 18041 54505
rect 17975 54481 18041 54491
rect 17975 54425 17980 54481
rect 18036 54425 18041 54481
rect 17975 54415 18041 54425
rect 17975 54401 17982 54415
rect 18034 54401 18041 54415
rect 17975 54345 17980 54401
rect 18036 54345 18041 54401
rect 17975 54321 17982 54345
rect 18034 54321 18041 54345
rect 17975 54265 17980 54321
rect 18036 54265 18041 54321
rect 17975 54241 17982 54265
rect 18034 54241 18041 54265
rect 17975 54185 17980 54241
rect 18036 54185 18041 54241
rect 17975 54171 17982 54185
rect 18034 54171 18041 54185
rect 17975 54156 18041 54171
rect 19063 54735 19129 54750
rect 19063 54721 19070 54735
rect 19122 54721 19129 54735
rect 19063 54665 19068 54721
rect 19124 54665 19129 54721
rect 19063 54641 19070 54665
rect 19122 54641 19129 54665
rect 19063 54585 19068 54641
rect 19124 54585 19129 54641
rect 19063 54561 19070 54585
rect 19122 54561 19129 54585
rect 19063 54505 19068 54561
rect 19124 54505 19129 54561
rect 19063 54491 19070 54505
rect 19122 54491 19129 54505
rect 19063 54481 19129 54491
rect 19063 54425 19068 54481
rect 19124 54425 19129 54481
rect 19063 54415 19129 54425
rect 19063 54401 19070 54415
rect 19122 54401 19129 54415
rect 19063 54345 19068 54401
rect 19124 54345 19129 54401
rect 19063 54321 19070 54345
rect 19122 54321 19129 54345
rect 19063 54265 19068 54321
rect 19124 54265 19129 54321
rect 19063 54241 19070 54265
rect 19122 54241 19129 54265
rect 19063 54185 19068 54241
rect 19124 54185 19129 54241
rect 19063 54171 19070 54185
rect 19122 54171 19129 54185
rect 19063 54156 19129 54171
rect 20151 54735 20217 54750
rect 20151 54721 20158 54735
rect 20210 54721 20217 54735
rect 20151 54665 20156 54721
rect 20212 54665 20217 54721
rect 20151 54641 20158 54665
rect 20210 54641 20217 54665
rect 20151 54585 20156 54641
rect 20212 54585 20217 54641
rect 20151 54561 20158 54585
rect 20210 54561 20217 54585
rect 20151 54505 20156 54561
rect 20212 54505 20217 54561
rect 20151 54491 20158 54505
rect 20210 54491 20217 54505
rect 20151 54481 20217 54491
rect 20151 54425 20156 54481
rect 20212 54425 20217 54481
rect 20151 54415 20217 54425
rect 20151 54401 20158 54415
rect 20210 54401 20217 54415
rect 20151 54345 20156 54401
rect 20212 54345 20217 54401
rect 20151 54321 20158 54345
rect 20210 54321 20217 54345
rect 20151 54265 20156 54321
rect 20212 54265 20217 54321
rect 20151 54241 20158 54265
rect 20210 54241 20217 54265
rect 20151 54185 20156 54241
rect 20212 54185 20217 54241
rect 20151 54171 20158 54185
rect 20210 54171 20217 54185
rect 20151 54156 20217 54171
rect 21239 54735 21305 54750
rect 21239 54721 21246 54735
rect 21298 54721 21305 54735
rect 21239 54665 21244 54721
rect 21300 54665 21305 54721
rect 21239 54641 21246 54665
rect 21298 54641 21305 54665
rect 21239 54585 21244 54641
rect 21300 54585 21305 54641
rect 21239 54561 21246 54585
rect 21298 54561 21305 54585
rect 21239 54505 21244 54561
rect 21300 54505 21305 54561
rect 21239 54491 21246 54505
rect 21298 54491 21305 54505
rect 21239 54481 21305 54491
rect 21239 54425 21244 54481
rect 21300 54425 21305 54481
rect 21239 54415 21305 54425
rect 21239 54401 21246 54415
rect 21298 54401 21305 54415
rect 21239 54345 21244 54401
rect 21300 54345 21305 54401
rect 21239 54321 21246 54345
rect 21298 54321 21305 54345
rect 21239 54265 21244 54321
rect 21300 54265 21305 54321
rect 21239 54241 21246 54265
rect 21298 54241 21305 54265
rect 21239 54185 21244 54241
rect 21300 54185 21305 54241
rect 21239 54171 21246 54185
rect 21298 54171 21305 54185
rect 21239 54156 21305 54171
rect 22327 54735 22393 54750
rect 22327 54721 22334 54735
rect 22386 54721 22393 54735
rect 22327 54665 22332 54721
rect 22388 54665 22393 54721
rect 22327 54641 22334 54665
rect 22386 54641 22393 54665
rect 22327 54585 22332 54641
rect 22388 54585 22393 54641
rect 22327 54561 22334 54585
rect 22386 54561 22393 54585
rect 22327 54505 22332 54561
rect 22388 54505 22393 54561
rect 22327 54491 22334 54505
rect 22386 54491 22393 54505
rect 22327 54481 22393 54491
rect 22327 54425 22332 54481
rect 22388 54425 22393 54481
rect 22327 54415 22393 54425
rect 22327 54401 22334 54415
rect 22386 54401 22393 54415
rect 22327 54345 22332 54401
rect 22388 54345 22393 54401
rect 22327 54321 22334 54345
rect 22386 54321 22393 54345
rect 22327 54265 22332 54321
rect 22388 54265 22393 54321
rect 22327 54241 22334 54265
rect 22386 54241 22393 54265
rect 22327 54185 22332 54241
rect 22388 54185 22393 54241
rect 22327 54171 22334 54185
rect 22386 54171 22393 54185
rect 22327 54156 22393 54171
rect 23415 54735 23481 54750
rect 23415 54721 23422 54735
rect 23474 54721 23481 54735
rect 23415 54665 23420 54721
rect 23476 54665 23481 54721
rect 23415 54641 23422 54665
rect 23474 54641 23481 54665
rect 23415 54585 23420 54641
rect 23476 54585 23481 54641
rect 23415 54561 23422 54585
rect 23474 54561 23481 54585
rect 23415 54505 23420 54561
rect 23476 54505 23481 54561
rect 23415 54491 23422 54505
rect 23474 54491 23481 54505
rect 23415 54481 23481 54491
rect 23415 54425 23420 54481
rect 23476 54425 23481 54481
rect 23415 54415 23481 54425
rect 23415 54401 23422 54415
rect 23474 54401 23481 54415
rect 23415 54345 23420 54401
rect 23476 54345 23481 54401
rect 23415 54321 23422 54345
rect 23474 54321 23481 54345
rect 23415 54265 23420 54321
rect 23476 54265 23481 54321
rect 23415 54241 23422 54265
rect 23474 54241 23481 54265
rect 23415 54185 23420 54241
rect 23476 54185 23481 54241
rect 23415 54171 23422 54185
rect 23474 54171 23481 54185
rect 23415 54156 23481 54171
rect 24503 54735 24569 54750
rect 24503 54721 24510 54735
rect 24562 54721 24569 54735
rect 24503 54665 24508 54721
rect 24564 54665 24569 54721
rect 24503 54641 24510 54665
rect 24562 54641 24569 54665
rect 24503 54585 24508 54641
rect 24564 54585 24569 54641
rect 24503 54561 24510 54585
rect 24562 54561 24569 54585
rect 24503 54505 24508 54561
rect 24564 54505 24569 54561
rect 24503 54491 24510 54505
rect 24562 54491 24569 54505
rect 24503 54481 24569 54491
rect 24503 54425 24508 54481
rect 24564 54425 24569 54481
rect 24503 54415 24569 54425
rect 24503 54401 24510 54415
rect 24562 54401 24569 54415
rect 24503 54345 24508 54401
rect 24564 54345 24569 54401
rect 24503 54321 24510 54345
rect 24562 54321 24569 54345
rect 24503 54265 24508 54321
rect 24564 54265 24569 54321
rect 24503 54241 24510 54265
rect 24562 54241 24569 54265
rect 24503 54185 24508 54241
rect 24564 54185 24569 54241
rect 24503 54171 24510 54185
rect 24562 54171 24569 54185
rect 24503 54156 24569 54171
rect 25591 54735 25657 54750
rect 25591 54721 25598 54735
rect 25650 54721 25657 54735
rect 25591 54665 25596 54721
rect 25652 54665 25657 54721
rect 25591 54641 25598 54665
rect 25650 54641 25657 54665
rect 25591 54585 25596 54641
rect 25652 54585 25657 54641
rect 25591 54561 25598 54585
rect 25650 54561 25657 54585
rect 25591 54505 25596 54561
rect 25652 54505 25657 54561
rect 25591 54491 25598 54505
rect 25650 54491 25657 54505
rect 25591 54481 25657 54491
rect 25591 54425 25596 54481
rect 25652 54425 25657 54481
rect 25591 54415 25657 54425
rect 25591 54401 25598 54415
rect 25650 54401 25657 54415
rect 25591 54345 25596 54401
rect 25652 54345 25657 54401
rect 25591 54321 25598 54345
rect 25650 54321 25657 54345
rect 25591 54265 25596 54321
rect 25652 54265 25657 54321
rect 25591 54241 25598 54265
rect 25650 54241 25657 54265
rect 25591 54185 25596 54241
rect 25652 54185 25657 54241
rect 25591 54171 25598 54185
rect 25650 54171 25657 54185
rect 25591 54156 25657 54171
rect 26679 54735 26745 54750
rect 26679 54721 26686 54735
rect 26738 54721 26745 54735
rect 26679 54665 26684 54721
rect 26740 54665 26745 54721
rect 26679 54641 26686 54665
rect 26738 54641 26745 54665
rect 26679 54585 26684 54641
rect 26740 54585 26745 54641
rect 26679 54561 26686 54585
rect 26738 54561 26745 54585
rect 26679 54505 26684 54561
rect 26740 54505 26745 54561
rect 26679 54491 26686 54505
rect 26738 54491 26745 54505
rect 26679 54481 26745 54491
rect 26679 54425 26684 54481
rect 26740 54425 26745 54481
rect 26679 54415 26745 54425
rect 26679 54401 26686 54415
rect 26738 54401 26745 54415
rect 26679 54345 26684 54401
rect 26740 54345 26745 54401
rect 26679 54321 26686 54345
rect 26738 54321 26745 54345
rect 26679 54265 26684 54321
rect 26740 54265 26745 54321
rect 26679 54241 26686 54265
rect 26738 54241 26745 54265
rect 26679 54185 26684 54241
rect 26740 54185 26745 54241
rect 26679 54171 26686 54185
rect 26738 54171 26745 54185
rect 26679 54156 26745 54171
rect 27767 54735 27833 54750
rect 27767 54721 27774 54735
rect 27826 54721 27833 54735
rect 27767 54665 27772 54721
rect 27828 54665 27833 54721
rect 27767 54641 27774 54665
rect 27826 54641 27833 54665
rect 27767 54585 27772 54641
rect 27828 54585 27833 54641
rect 27767 54561 27774 54585
rect 27826 54561 27833 54585
rect 27767 54505 27772 54561
rect 27828 54505 27833 54561
rect 27767 54491 27774 54505
rect 27826 54491 27833 54505
rect 27767 54481 27833 54491
rect 27767 54425 27772 54481
rect 27828 54425 27833 54481
rect 27767 54415 27833 54425
rect 27767 54401 27774 54415
rect 27826 54401 27833 54415
rect 27767 54345 27772 54401
rect 27828 54345 27833 54401
rect 27767 54321 27774 54345
rect 27826 54321 27833 54345
rect 27767 54265 27772 54321
rect 27828 54265 27833 54321
rect 27767 54241 27774 54265
rect 27826 54241 27833 54265
rect 27767 54185 27772 54241
rect 27828 54185 27833 54241
rect 27767 54171 27774 54185
rect 27826 54171 27833 54185
rect 27767 54156 27833 54171
rect 28855 54735 28921 54750
rect 28855 54721 28862 54735
rect 28914 54721 28921 54735
rect 28855 54665 28860 54721
rect 28916 54665 28921 54721
rect 28855 54641 28862 54665
rect 28914 54641 28921 54665
rect 28855 54585 28860 54641
rect 28916 54585 28921 54641
rect 28855 54561 28862 54585
rect 28914 54561 28921 54585
rect 28855 54505 28860 54561
rect 28916 54505 28921 54561
rect 28855 54491 28862 54505
rect 28914 54491 28921 54505
rect 28855 54481 28921 54491
rect 28855 54425 28860 54481
rect 28916 54425 28921 54481
rect 28855 54415 28921 54425
rect 28855 54401 28862 54415
rect 28914 54401 28921 54415
rect 28855 54345 28860 54401
rect 28916 54345 28921 54401
rect 28855 54321 28862 54345
rect 28914 54321 28921 54345
rect 28855 54265 28860 54321
rect 28916 54265 28921 54321
rect 28855 54241 28862 54265
rect 28914 54241 28921 54265
rect 28855 54185 28860 54241
rect 28916 54185 28921 54241
rect 28855 54171 28862 54185
rect 28914 54171 28921 54185
rect 28855 54156 28921 54171
rect 29943 54735 30009 54750
rect 29943 54721 29950 54735
rect 30002 54721 30009 54735
rect 29943 54665 29948 54721
rect 30004 54665 30009 54721
rect 29943 54641 29950 54665
rect 30002 54641 30009 54665
rect 29943 54585 29948 54641
rect 30004 54585 30009 54641
rect 29943 54561 29950 54585
rect 30002 54561 30009 54585
rect 29943 54505 29948 54561
rect 30004 54505 30009 54561
rect 29943 54491 29950 54505
rect 30002 54491 30009 54505
rect 29943 54481 30009 54491
rect 29943 54425 29948 54481
rect 30004 54425 30009 54481
rect 29943 54415 30009 54425
rect 29943 54401 29950 54415
rect 30002 54401 30009 54415
rect 29943 54345 29948 54401
rect 30004 54345 30009 54401
rect 29943 54321 29950 54345
rect 30002 54321 30009 54345
rect 29943 54265 29948 54321
rect 30004 54265 30009 54321
rect 29943 54241 29950 54265
rect 30002 54241 30009 54265
rect 29943 54185 29948 54241
rect 30004 54185 30009 54241
rect 29943 54171 29950 54185
rect 30002 54171 30009 54185
rect 29943 54156 30009 54171
rect 31031 54735 31097 54750
rect 31031 54721 31038 54735
rect 31090 54721 31097 54735
rect 31031 54665 31036 54721
rect 31092 54665 31097 54721
rect 31031 54641 31038 54665
rect 31090 54641 31097 54665
rect 31031 54585 31036 54641
rect 31092 54585 31097 54641
rect 31031 54561 31038 54585
rect 31090 54561 31097 54585
rect 31031 54505 31036 54561
rect 31092 54505 31097 54561
rect 31031 54491 31038 54505
rect 31090 54491 31097 54505
rect 31031 54481 31097 54491
rect 31031 54425 31036 54481
rect 31092 54425 31097 54481
rect 31031 54415 31097 54425
rect 31031 54401 31038 54415
rect 31090 54401 31097 54415
rect 31031 54345 31036 54401
rect 31092 54345 31097 54401
rect 31031 54321 31038 54345
rect 31090 54321 31097 54345
rect 31031 54265 31036 54321
rect 31092 54265 31097 54321
rect 31031 54241 31038 54265
rect 31090 54241 31097 54265
rect 31031 54185 31036 54241
rect 31092 54185 31097 54241
rect 31031 54171 31038 54185
rect 31090 54171 31097 54185
rect 31031 54156 31097 54171
rect 17430 52738 17496 52753
rect 17430 52724 17437 52738
rect 17489 52724 17496 52738
rect 17430 52668 17435 52724
rect 17491 52668 17496 52724
rect 17430 52644 17437 52668
rect 17489 52644 17496 52668
rect 17430 52588 17435 52644
rect 17491 52588 17496 52644
rect 17430 52564 17437 52588
rect 17489 52564 17496 52588
rect 17430 52508 17435 52564
rect 17491 52508 17496 52564
rect 17430 52494 17437 52508
rect 17489 52494 17496 52508
rect 17430 52484 17496 52494
rect 17430 52428 17435 52484
rect 17491 52428 17496 52484
rect 17430 52418 17496 52428
rect 17430 52404 17437 52418
rect 17489 52404 17496 52418
rect 17430 52348 17435 52404
rect 17491 52348 17496 52404
rect 17430 52324 17437 52348
rect 17489 52324 17496 52348
rect 17430 52268 17435 52324
rect 17491 52268 17496 52324
rect 17430 52244 17437 52268
rect 17489 52244 17496 52268
rect 17430 52188 17435 52244
rect 17491 52188 17496 52244
rect 17430 52174 17437 52188
rect 17489 52174 17496 52188
rect 17430 52159 17496 52174
rect 18518 52738 18584 52753
rect 18518 52724 18525 52738
rect 18577 52724 18584 52738
rect 18518 52668 18523 52724
rect 18579 52668 18584 52724
rect 18518 52644 18525 52668
rect 18577 52644 18584 52668
rect 18518 52588 18523 52644
rect 18579 52588 18584 52644
rect 18518 52564 18525 52588
rect 18577 52564 18584 52588
rect 18518 52508 18523 52564
rect 18579 52508 18584 52564
rect 18518 52494 18525 52508
rect 18577 52494 18584 52508
rect 18518 52484 18584 52494
rect 18518 52428 18523 52484
rect 18579 52428 18584 52484
rect 18518 52418 18584 52428
rect 18518 52404 18525 52418
rect 18577 52404 18584 52418
rect 18518 52348 18523 52404
rect 18579 52348 18584 52404
rect 18518 52324 18525 52348
rect 18577 52324 18584 52348
rect 18518 52268 18523 52324
rect 18579 52268 18584 52324
rect 18518 52244 18525 52268
rect 18577 52244 18584 52268
rect 18518 52188 18523 52244
rect 18579 52188 18584 52244
rect 18518 52174 18525 52188
rect 18577 52174 18584 52188
rect 18518 52159 18584 52174
rect 19606 52738 19672 52753
rect 19606 52724 19613 52738
rect 19665 52724 19672 52738
rect 19606 52668 19611 52724
rect 19667 52668 19672 52724
rect 19606 52644 19613 52668
rect 19665 52644 19672 52668
rect 19606 52588 19611 52644
rect 19667 52588 19672 52644
rect 19606 52564 19613 52588
rect 19665 52564 19672 52588
rect 19606 52508 19611 52564
rect 19667 52508 19672 52564
rect 19606 52494 19613 52508
rect 19665 52494 19672 52508
rect 19606 52484 19672 52494
rect 19606 52428 19611 52484
rect 19667 52428 19672 52484
rect 19606 52418 19672 52428
rect 19606 52404 19613 52418
rect 19665 52404 19672 52418
rect 19606 52348 19611 52404
rect 19667 52348 19672 52404
rect 19606 52324 19613 52348
rect 19665 52324 19672 52348
rect 19606 52268 19611 52324
rect 19667 52268 19672 52324
rect 19606 52244 19613 52268
rect 19665 52244 19672 52268
rect 19606 52188 19611 52244
rect 19667 52188 19672 52244
rect 19606 52174 19613 52188
rect 19665 52174 19672 52188
rect 19606 52159 19672 52174
rect 20694 52738 20760 52753
rect 20694 52724 20701 52738
rect 20753 52724 20760 52738
rect 20694 52668 20699 52724
rect 20755 52668 20760 52724
rect 20694 52644 20701 52668
rect 20753 52644 20760 52668
rect 20694 52588 20699 52644
rect 20755 52588 20760 52644
rect 20694 52564 20701 52588
rect 20753 52564 20760 52588
rect 20694 52508 20699 52564
rect 20755 52508 20760 52564
rect 20694 52494 20701 52508
rect 20753 52494 20760 52508
rect 20694 52484 20760 52494
rect 20694 52428 20699 52484
rect 20755 52428 20760 52484
rect 20694 52418 20760 52428
rect 20694 52404 20701 52418
rect 20753 52404 20760 52418
rect 20694 52348 20699 52404
rect 20755 52348 20760 52404
rect 20694 52324 20701 52348
rect 20753 52324 20760 52348
rect 20694 52268 20699 52324
rect 20755 52268 20760 52324
rect 20694 52244 20701 52268
rect 20753 52244 20760 52268
rect 20694 52188 20699 52244
rect 20755 52188 20760 52244
rect 20694 52174 20701 52188
rect 20753 52174 20760 52188
rect 20694 52159 20760 52174
rect 21782 52738 21848 52753
rect 21782 52724 21789 52738
rect 21841 52724 21848 52738
rect 21782 52668 21787 52724
rect 21843 52668 21848 52724
rect 21782 52644 21789 52668
rect 21841 52644 21848 52668
rect 21782 52588 21787 52644
rect 21843 52588 21848 52644
rect 21782 52564 21789 52588
rect 21841 52564 21848 52588
rect 21782 52508 21787 52564
rect 21843 52508 21848 52564
rect 21782 52494 21789 52508
rect 21841 52494 21848 52508
rect 21782 52484 21848 52494
rect 21782 52428 21787 52484
rect 21843 52428 21848 52484
rect 21782 52418 21848 52428
rect 21782 52404 21789 52418
rect 21841 52404 21848 52418
rect 21782 52348 21787 52404
rect 21843 52348 21848 52404
rect 21782 52324 21789 52348
rect 21841 52324 21848 52348
rect 21782 52268 21787 52324
rect 21843 52268 21848 52324
rect 21782 52244 21789 52268
rect 21841 52244 21848 52268
rect 21782 52188 21787 52244
rect 21843 52188 21848 52244
rect 21782 52174 21789 52188
rect 21841 52174 21848 52188
rect 21782 52159 21848 52174
rect 22870 52738 22936 52753
rect 22870 52724 22877 52738
rect 22929 52724 22936 52738
rect 22870 52668 22875 52724
rect 22931 52668 22936 52724
rect 22870 52644 22877 52668
rect 22929 52644 22936 52668
rect 22870 52588 22875 52644
rect 22931 52588 22936 52644
rect 22870 52564 22877 52588
rect 22929 52564 22936 52588
rect 22870 52508 22875 52564
rect 22931 52508 22936 52564
rect 22870 52494 22877 52508
rect 22929 52494 22936 52508
rect 22870 52484 22936 52494
rect 22870 52428 22875 52484
rect 22931 52428 22936 52484
rect 22870 52418 22936 52428
rect 22870 52404 22877 52418
rect 22929 52404 22936 52418
rect 22870 52348 22875 52404
rect 22931 52348 22936 52404
rect 22870 52324 22877 52348
rect 22929 52324 22936 52348
rect 22870 52268 22875 52324
rect 22931 52268 22936 52324
rect 22870 52244 22877 52268
rect 22929 52244 22936 52268
rect 22870 52188 22875 52244
rect 22931 52188 22936 52244
rect 22870 52174 22877 52188
rect 22929 52174 22936 52188
rect 22870 52159 22936 52174
rect 23958 52738 24024 52753
rect 23958 52724 23965 52738
rect 24017 52724 24024 52738
rect 23958 52668 23963 52724
rect 24019 52668 24024 52724
rect 23958 52644 23965 52668
rect 24017 52644 24024 52668
rect 23958 52588 23963 52644
rect 24019 52588 24024 52644
rect 23958 52564 23965 52588
rect 24017 52564 24024 52588
rect 23958 52508 23963 52564
rect 24019 52508 24024 52564
rect 23958 52494 23965 52508
rect 24017 52494 24024 52508
rect 23958 52484 24024 52494
rect 23958 52428 23963 52484
rect 24019 52428 24024 52484
rect 23958 52418 24024 52428
rect 23958 52404 23965 52418
rect 24017 52404 24024 52418
rect 23958 52348 23963 52404
rect 24019 52348 24024 52404
rect 23958 52324 23965 52348
rect 24017 52324 24024 52348
rect 23958 52268 23963 52324
rect 24019 52268 24024 52324
rect 23958 52244 23965 52268
rect 24017 52244 24024 52268
rect 23958 52188 23963 52244
rect 24019 52188 24024 52244
rect 23958 52174 23965 52188
rect 24017 52174 24024 52188
rect 23958 52159 24024 52174
rect 25046 52738 25112 52753
rect 25046 52724 25053 52738
rect 25105 52724 25112 52738
rect 25046 52668 25051 52724
rect 25107 52668 25112 52724
rect 25046 52644 25053 52668
rect 25105 52644 25112 52668
rect 25046 52588 25051 52644
rect 25107 52588 25112 52644
rect 25046 52564 25053 52588
rect 25105 52564 25112 52588
rect 25046 52508 25051 52564
rect 25107 52508 25112 52564
rect 25046 52494 25053 52508
rect 25105 52494 25112 52508
rect 25046 52484 25112 52494
rect 25046 52428 25051 52484
rect 25107 52428 25112 52484
rect 25046 52418 25112 52428
rect 25046 52404 25053 52418
rect 25105 52404 25112 52418
rect 25046 52348 25051 52404
rect 25107 52348 25112 52404
rect 25046 52324 25053 52348
rect 25105 52324 25112 52348
rect 25046 52268 25051 52324
rect 25107 52268 25112 52324
rect 25046 52244 25053 52268
rect 25105 52244 25112 52268
rect 25046 52188 25051 52244
rect 25107 52188 25112 52244
rect 25046 52174 25053 52188
rect 25105 52174 25112 52188
rect 25046 52159 25112 52174
rect 26134 52738 26200 52753
rect 26134 52724 26141 52738
rect 26193 52724 26200 52738
rect 26134 52668 26139 52724
rect 26195 52668 26200 52724
rect 26134 52644 26141 52668
rect 26193 52644 26200 52668
rect 26134 52588 26139 52644
rect 26195 52588 26200 52644
rect 26134 52564 26141 52588
rect 26193 52564 26200 52588
rect 26134 52508 26139 52564
rect 26195 52508 26200 52564
rect 26134 52494 26141 52508
rect 26193 52494 26200 52508
rect 26134 52484 26200 52494
rect 26134 52428 26139 52484
rect 26195 52428 26200 52484
rect 26134 52418 26200 52428
rect 26134 52404 26141 52418
rect 26193 52404 26200 52418
rect 26134 52348 26139 52404
rect 26195 52348 26200 52404
rect 26134 52324 26141 52348
rect 26193 52324 26200 52348
rect 26134 52268 26139 52324
rect 26195 52268 26200 52324
rect 26134 52244 26141 52268
rect 26193 52244 26200 52268
rect 26134 52188 26139 52244
rect 26195 52188 26200 52244
rect 26134 52174 26141 52188
rect 26193 52174 26200 52188
rect 26134 52159 26200 52174
rect 27222 52738 27288 52753
rect 27222 52724 27229 52738
rect 27281 52724 27288 52738
rect 27222 52668 27227 52724
rect 27283 52668 27288 52724
rect 27222 52644 27229 52668
rect 27281 52644 27288 52668
rect 27222 52588 27227 52644
rect 27283 52588 27288 52644
rect 27222 52564 27229 52588
rect 27281 52564 27288 52588
rect 27222 52508 27227 52564
rect 27283 52508 27288 52564
rect 27222 52494 27229 52508
rect 27281 52494 27288 52508
rect 27222 52484 27288 52494
rect 27222 52428 27227 52484
rect 27283 52428 27288 52484
rect 27222 52418 27288 52428
rect 27222 52404 27229 52418
rect 27281 52404 27288 52418
rect 27222 52348 27227 52404
rect 27283 52348 27288 52404
rect 27222 52324 27229 52348
rect 27281 52324 27288 52348
rect 27222 52268 27227 52324
rect 27283 52268 27288 52324
rect 27222 52244 27229 52268
rect 27281 52244 27288 52268
rect 27222 52188 27227 52244
rect 27283 52188 27288 52244
rect 27222 52174 27229 52188
rect 27281 52174 27288 52188
rect 27222 52159 27288 52174
rect 28310 52738 28376 52753
rect 28310 52724 28317 52738
rect 28369 52724 28376 52738
rect 28310 52668 28315 52724
rect 28371 52668 28376 52724
rect 28310 52644 28317 52668
rect 28369 52644 28376 52668
rect 28310 52588 28315 52644
rect 28371 52588 28376 52644
rect 28310 52564 28317 52588
rect 28369 52564 28376 52588
rect 28310 52508 28315 52564
rect 28371 52508 28376 52564
rect 28310 52494 28317 52508
rect 28369 52494 28376 52508
rect 28310 52484 28376 52494
rect 28310 52428 28315 52484
rect 28371 52428 28376 52484
rect 28310 52418 28376 52428
rect 28310 52404 28317 52418
rect 28369 52404 28376 52418
rect 28310 52348 28315 52404
rect 28371 52348 28376 52404
rect 28310 52324 28317 52348
rect 28369 52324 28376 52348
rect 28310 52268 28315 52324
rect 28371 52268 28376 52324
rect 28310 52244 28317 52268
rect 28369 52244 28376 52268
rect 28310 52188 28315 52244
rect 28371 52188 28376 52244
rect 28310 52174 28317 52188
rect 28369 52174 28376 52188
rect 28310 52159 28376 52174
rect 29398 52738 29464 52753
rect 29398 52724 29405 52738
rect 29457 52724 29464 52738
rect 29398 52668 29403 52724
rect 29459 52668 29464 52724
rect 29398 52644 29405 52668
rect 29457 52644 29464 52668
rect 29398 52588 29403 52644
rect 29459 52588 29464 52644
rect 29398 52564 29405 52588
rect 29457 52564 29464 52588
rect 29398 52508 29403 52564
rect 29459 52508 29464 52564
rect 29398 52494 29405 52508
rect 29457 52494 29464 52508
rect 29398 52484 29464 52494
rect 29398 52428 29403 52484
rect 29459 52428 29464 52484
rect 29398 52418 29464 52428
rect 29398 52404 29405 52418
rect 29457 52404 29464 52418
rect 29398 52348 29403 52404
rect 29459 52348 29464 52404
rect 29398 52324 29405 52348
rect 29457 52324 29464 52348
rect 29398 52268 29403 52324
rect 29459 52268 29464 52324
rect 29398 52244 29405 52268
rect 29457 52244 29464 52268
rect 29398 52188 29403 52244
rect 29459 52188 29464 52244
rect 29398 52174 29405 52188
rect 29457 52174 29464 52188
rect 29398 52159 29464 52174
rect 30486 52738 30552 52753
rect 30486 52724 30493 52738
rect 30545 52724 30552 52738
rect 30486 52668 30491 52724
rect 30547 52668 30552 52724
rect 30486 52644 30493 52668
rect 30545 52644 30552 52668
rect 30486 52588 30491 52644
rect 30547 52588 30552 52644
rect 30486 52564 30493 52588
rect 30545 52564 30552 52588
rect 30486 52508 30491 52564
rect 30547 52508 30552 52564
rect 30486 52494 30493 52508
rect 30545 52494 30552 52508
rect 30486 52484 30552 52494
rect 30486 52428 30491 52484
rect 30547 52428 30552 52484
rect 30486 52418 30552 52428
rect 30486 52404 30493 52418
rect 30545 52404 30552 52418
rect 30486 52348 30491 52404
rect 30547 52348 30552 52404
rect 30486 52324 30493 52348
rect 30545 52324 30552 52348
rect 30486 52268 30491 52324
rect 30547 52268 30552 52324
rect 30486 52244 30493 52268
rect 30545 52244 30552 52268
rect 30486 52188 30491 52244
rect 30547 52188 30552 52244
rect 30486 52174 30493 52188
rect 30545 52174 30552 52188
rect 30486 52159 30552 52174
rect 31574 52738 31640 52753
rect 31574 52724 31581 52738
rect 31633 52724 31640 52738
rect 31574 52668 31579 52724
rect 31635 52668 31640 52724
rect 31574 52644 31581 52668
rect 31633 52644 31640 52668
rect 31574 52588 31579 52644
rect 31635 52588 31640 52644
rect 31574 52564 31581 52588
rect 31633 52564 31640 52588
rect 31574 52508 31579 52564
rect 31635 52508 31640 52564
rect 31574 52494 31581 52508
rect 31633 52494 31640 52508
rect 31574 52484 31640 52494
rect 31574 52428 31579 52484
rect 31635 52428 31640 52484
rect 31574 52418 31640 52428
rect 31574 52404 31581 52418
rect 31633 52404 31640 52418
rect 31574 52348 31579 52404
rect 31635 52348 31640 52404
rect 31574 52324 31581 52348
rect 31633 52324 31640 52348
rect 31574 52268 31579 52324
rect 31635 52268 31640 52324
rect 31574 52244 31581 52268
rect 31633 52244 31640 52268
rect 31574 52188 31579 52244
rect 31635 52188 31640 52244
rect 31574 52174 31581 52188
rect 31633 52174 31640 52188
rect 31574 52159 31640 52174
rect 17975 50735 18041 50750
rect 17975 50721 17982 50735
rect 18034 50721 18041 50735
rect 17975 50665 17980 50721
rect 18036 50665 18041 50721
rect 17975 50641 17982 50665
rect 18034 50641 18041 50665
rect 17975 50585 17980 50641
rect 18036 50585 18041 50641
rect 17975 50561 17982 50585
rect 18034 50561 18041 50585
rect 17975 50505 17980 50561
rect 18036 50505 18041 50561
rect 17975 50491 17982 50505
rect 18034 50491 18041 50505
rect 17975 50481 18041 50491
rect 17975 50425 17980 50481
rect 18036 50425 18041 50481
rect 17975 50415 18041 50425
rect 17975 50401 17982 50415
rect 18034 50401 18041 50415
rect 17975 50345 17980 50401
rect 18036 50345 18041 50401
rect 17975 50321 17982 50345
rect 18034 50321 18041 50345
rect 17975 50265 17980 50321
rect 18036 50265 18041 50321
rect 17975 50241 17982 50265
rect 18034 50241 18041 50265
rect 17975 50185 17980 50241
rect 18036 50185 18041 50241
rect 17975 50171 17982 50185
rect 18034 50171 18041 50185
rect 17975 50156 18041 50171
rect 20151 50735 20217 50750
rect 20151 50721 20158 50735
rect 20210 50721 20217 50735
rect 20151 50665 20156 50721
rect 20212 50665 20217 50721
rect 20151 50641 20158 50665
rect 20210 50641 20217 50665
rect 20151 50585 20156 50641
rect 20212 50585 20217 50641
rect 20151 50561 20158 50585
rect 20210 50561 20217 50585
rect 20151 50505 20156 50561
rect 20212 50505 20217 50561
rect 20151 50491 20158 50505
rect 20210 50491 20217 50505
rect 20151 50481 20217 50491
rect 20151 50425 20156 50481
rect 20212 50425 20217 50481
rect 20151 50415 20217 50425
rect 20151 50401 20158 50415
rect 20210 50401 20217 50415
rect 20151 50345 20156 50401
rect 20212 50345 20217 50401
rect 20151 50321 20158 50345
rect 20210 50321 20217 50345
rect 20151 50265 20156 50321
rect 20212 50265 20217 50321
rect 20151 50241 20158 50265
rect 20210 50241 20217 50265
rect 20151 50185 20156 50241
rect 20212 50185 20217 50241
rect 20151 50171 20158 50185
rect 20210 50171 20217 50185
rect 20151 50156 20217 50171
rect 21239 50735 21305 50750
rect 21239 50721 21246 50735
rect 21298 50721 21305 50735
rect 21239 50665 21244 50721
rect 21300 50665 21305 50721
rect 21239 50641 21246 50665
rect 21298 50641 21305 50665
rect 21239 50585 21244 50641
rect 21300 50585 21305 50641
rect 21239 50561 21246 50585
rect 21298 50561 21305 50585
rect 21239 50505 21244 50561
rect 21300 50505 21305 50561
rect 21239 50491 21246 50505
rect 21298 50491 21305 50505
rect 21239 50481 21305 50491
rect 21239 50425 21244 50481
rect 21300 50425 21305 50481
rect 21239 50415 21305 50425
rect 21239 50401 21246 50415
rect 21298 50401 21305 50415
rect 21239 50345 21244 50401
rect 21300 50345 21305 50401
rect 21239 50321 21246 50345
rect 21298 50321 21305 50345
rect 21239 50265 21244 50321
rect 21300 50265 21305 50321
rect 21239 50241 21246 50265
rect 21298 50241 21305 50265
rect 21239 50185 21244 50241
rect 21300 50185 21305 50241
rect 21239 50171 21246 50185
rect 21298 50171 21305 50185
rect 21239 50156 21305 50171
rect 23415 50735 23481 50750
rect 23415 50721 23422 50735
rect 23474 50721 23481 50735
rect 23415 50665 23420 50721
rect 23476 50665 23481 50721
rect 23415 50641 23422 50665
rect 23474 50641 23481 50665
rect 23415 50585 23420 50641
rect 23476 50585 23481 50641
rect 23415 50561 23422 50585
rect 23474 50561 23481 50585
rect 23415 50505 23420 50561
rect 23476 50505 23481 50561
rect 23415 50491 23422 50505
rect 23474 50491 23481 50505
rect 23415 50481 23481 50491
rect 23415 50425 23420 50481
rect 23476 50425 23481 50481
rect 23415 50415 23481 50425
rect 23415 50401 23422 50415
rect 23474 50401 23481 50415
rect 23415 50345 23420 50401
rect 23476 50345 23481 50401
rect 23415 50321 23422 50345
rect 23474 50321 23481 50345
rect 23415 50265 23420 50321
rect 23476 50265 23481 50321
rect 23415 50241 23422 50265
rect 23474 50241 23481 50265
rect 23415 50185 23420 50241
rect 23476 50185 23481 50241
rect 23415 50171 23422 50185
rect 23474 50171 23481 50185
rect 23415 50156 23481 50171
rect 24503 50735 24569 50750
rect 24503 50721 24510 50735
rect 24562 50721 24569 50735
rect 24503 50665 24508 50721
rect 24564 50665 24569 50721
rect 24503 50641 24510 50665
rect 24562 50641 24569 50665
rect 24503 50585 24508 50641
rect 24564 50585 24569 50641
rect 24503 50561 24510 50585
rect 24562 50561 24569 50585
rect 24503 50505 24508 50561
rect 24564 50505 24569 50561
rect 24503 50491 24510 50505
rect 24562 50491 24569 50505
rect 24503 50481 24569 50491
rect 24503 50425 24508 50481
rect 24564 50425 24569 50481
rect 24503 50415 24569 50425
rect 24503 50401 24510 50415
rect 24562 50401 24569 50415
rect 24503 50345 24508 50401
rect 24564 50345 24569 50401
rect 24503 50321 24510 50345
rect 24562 50321 24569 50345
rect 24503 50265 24508 50321
rect 24564 50265 24569 50321
rect 24503 50241 24510 50265
rect 24562 50241 24569 50265
rect 24503 50185 24508 50241
rect 24564 50185 24569 50241
rect 24503 50171 24510 50185
rect 24562 50171 24569 50185
rect 24503 50156 24569 50171
rect 25591 50735 25657 50750
rect 25591 50721 25598 50735
rect 25650 50721 25657 50735
rect 25591 50665 25596 50721
rect 25652 50665 25657 50721
rect 25591 50641 25598 50665
rect 25650 50641 25657 50665
rect 25591 50585 25596 50641
rect 25652 50585 25657 50641
rect 25591 50561 25598 50585
rect 25650 50561 25657 50585
rect 25591 50505 25596 50561
rect 25652 50505 25657 50561
rect 25591 50491 25598 50505
rect 25650 50491 25657 50505
rect 25591 50481 25657 50491
rect 25591 50425 25596 50481
rect 25652 50425 25657 50481
rect 25591 50415 25657 50425
rect 25591 50401 25598 50415
rect 25650 50401 25657 50415
rect 25591 50345 25596 50401
rect 25652 50345 25657 50401
rect 25591 50321 25598 50345
rect 25650 50321 25657 50345
rect 25591 50265 25596 50321
rect 25652 50265 25657 50321
rect 25591 50241 25598 50265
rect 25650 50241 25657 50265
rect 25591 50185 25596 50241
rect 25652 50185 25657 50241
rect 25591 50171 25598 50185
rect 25650 50171 25657 50185
rect 25591 50156 25657 50171
rect 27767 50735 27833 50750
rect 27767 50721 27774 50735
rect 27826 50721 27833 50735
rect 27767 50665 27772 50721
rect 27828 50665 27833 50721
rect 27767 50641 27774 50665
rect 27826 50641 27833 50665
rect 27767 50585 27772 50641
rect 27828 50585 27833 50641
rect 27767 50561 27774 50585
rect 27826 50561 27833 50585
rect 27767 50505 27772 50561
rect 27828 50505 27833 50561
rect 27767 50491 27774 50505
rect 27826 50491 27833 50505
rect 27767 50481 27833 50491
rect 27767 50425 27772 50481
rect 27828 50425 27833 50481
rect 27767 50415 27833 50425
rect 27767 50401 27774 50415
rect 27826 50401 27833 50415
rect 27767 50345 27772 50401
rect 27828 50345 27833 50401
rect 27767 50321 27774 50345
rect 27826 50321 27833 50345
rect 27767 50265 27772 50321
rect 27828 50265 27833 50321
rect 27767 50241 27774 50265
rect 27826 50241 27833 50265
rect 27767 50185 27772 50241
rect 27828 50185 27833 50241
rect 27767 50171 27774 50185
rect 27826 50171 27833 50185
rect 27767 50156 27833 50171
rect 28855 50735 28921 50750
rect 28855 50721 28862 50735
rect 28914 50721 28921 50735
rect 28855 50665 28860 50721
rect 28916 50665 28921 50721
rect 28855 50641 28862 50665
rect 28914 50641 28921 50665
rect 28855 50585 28860 50641
rect 28916 50585 28921 50641
rect 28855 50561 28862 50585
rect 28914 50561 28921 50585
rect 28855 50505 28860 50561
rect 28916 50505 28921 50561
rect 28855 50491 28862 50505
rect 28914 50491 28921 50505
rect 28855 50481 28921 50491
rect 28855 50425 28860 50481
rect 28916 50425 28921 50481
rect 28855 50415 28921 50425
rect 28855 50401 28862 50415
rect 28914 50401 28921 50415
rect 28855 50345 28860 50401
rect 28916 50345 28921 50401
rect 28855 50321 28862 50345
rect 28914 50321 28921 50345
rect 28855 50265 28860 50321
rect 28916 50265 28921 50321
rect 28855 50241 28862 50265
rect 28914 50241 28921 50265
rect 28855 50185 28860 50241
rect 28916 50185 28921 50241
rect 28855 50171 28862 50185
rect 28914 50171 28921 50185
rect 28855 50156 28921 50171
rect 31031 50735 31097 50750
rect 31031 50721 31038 50735
rect 31090 50721 31097 50735
rect 31031 50665 31036 50721
rect 31092 50665 31097 50721
rect 31031 50641 31038 50665
rect 31090 50641 31097 50665
rect 31031 50585 31036 50641
rect 31092 50585 31097 50641
rect 31031 50561 31038 50585
rect 31090 50561 31097 50585
rect 31031 50505 31036 50561
rect 31092 50505 31097 50561
rect 31031 50491 31038 50505
rect 31090 50491 31097 50505
rect 31031 50481 31097 50491
rect 31031 50425 31036 50481
rect 31092 50425 31097 50481
rect 31031 50415 31097 50425
rect 31031 50401 31038 50415
rect 31090 50401 31097 50415
rect 31031 50345 31036 50401
rect 31092 50345 31097 50401
rect 31031 50321 31038 50345
rect 31090 50321 31097 50345
rect 31031 50265 31036 50321
rect 31092 50265 31097 50321
rect 31031 50241 31038 50265
rect 31090 50241 31097 50265
rect 31031 50185 31036 50241
rect 31092 50185 31097 50241
rect 31031 50171 31038 50185
rect 31090 50171 31097 50185
rect 31031 50156 31097 50171
rect 17430 48738 17496 48753
rect 17430 48724 17437 48738
rect 17489 48724 17496 48738
rect 17430 48668 17435 48724
rect 17491 48668 17496 48724
rect 17430 48644 17437 48668
rect 17489 48644 17496 48668
rect 17430 48588 17435 48644
rect 17491 48588 17496 48644
rect 17430 48564 17437 48588
rect 17489 48564 17496 48588
rect 17430 48508 17435 48564
rect 17491 48508 17496 48564
rect 17430 48494 17437 48508
rect 17489 48494 17496 48508
rect 17430 48484 17496 48494
rect 17430 48428 17435 48484
rect 17491 48428 17496 48484
rect 17430 48418 17496 48428
rect 17430 48404 17437 48418
rect 17489 48404 17496 48418
rect 17430 48348 17435 48404
rect 17491 48348 17496 48404
rect 17430 48324 17437 48348
rect 17489 48324 17496 48348
rect 17430 48268 17435 48324
rect 17491 48268 17496 48324
rect 17430 48244 17437 48268
rect 17489 48244 17496 48268
rect 17430 48188 17435 48244
rect 17491 48188 17496 48244
rect 17430 48174 17437 48188
rect 17489 48174 17496 48188
rect 17430 48159 17496 48174
rect 18518 48738 18584 48753
rect 18518 48724 18525 48738
rect 18577 48724 18584 48738
rect 18518 48668 18523 48724
rect 18579 48668 18584 48724
rect 18518 48644 18525 48668
rect 18577 48644 18584 48668
rect 18518 48588 18523 48644
rect 18579 48588 18584 48644
rect 18518 48564 18525 48588
rect 18577 48564 18584 48588
rect 18518 48508 18523 48564
rect 18579 48508 18584 48564
rect 18518 48494 18525 48508
rect 18577 48494 18584 48508
rect 18518 48484 18584 48494
rect 18518 48428 18523 48484
rect 18579 48428 18584 48484
rect 18518 48418 18584 48428
rect 18518 48404 18525 48418
rect 18577 48404 18584 48418
rect 18518 48348 18523 48404
rect 18579 48348 18584 48404
rect 18518 48324 18525 48348
rect 18577 48324 18584 48348
rect 18518 48268 18523 48324
rect 18579 48268 18584 48324
rect 18518 48244 18525 48268
rect 18577 48244 18584 48268
rect 18518 48188 18523 48244
rect 18579 48188 18584 48244
rect 18518 48174 18525 48188
rect 18577 48174 18584 48188
rect 18518 48159 18584 48174
rect 19606 48738 19672 48753
rect 19606 48724 19613 48738
rect 19665 48724 19672 48738
rect 19606 48668 19611 48724
rect 19667 48668 19672 48724
rect 19606 48644 19613 48668
rect 19665 48644 19672 48668
rect 19606 48588 19611 48644
rect 19667 48588 19672 48644
rect 19606 48564 19613 48588
rect 19665 48564 19672 48588
rect 19606 48508 19611 48564
rect 19667 48508 19672 48564
rect 19606 48494 19613 48508
rect 19665 48494 19672 48508
rect 19606 48484 19672 48494
rect 19606 48428 19611 48484
rect 19667 48428 19672 48484
rect 19606 48418 19672 48428
rect 19606 48404 19613 48418
rect 19665 48404 19672 48418
rect 19606 48348 19611 48404
rect 19667 48348 19672 48404
rect 19606 48324 19613 48348
rect 19665 48324 19672 48348
rect 19606 48268 19611 48324
rect 19667 48268 19672 48324
rect 19606 48244 19613 48268
rect 19665 48244 19672 48268
rect 19606 48188 19611 48244
rect 19667 48188 19672 48244
rect 19606 48174 19613 48188
rect 19665 48174 19672 48188
rect 19606 48159 19672 48174
rect 20694 48738 20760 48753
rect 20694 48724 20701 48738
rect 20753 48724 20760 48738
rect 20694 48668 20699 48724
rect 20755 48668 20760 48724
rect 20694 48644 20701 48668
rect 20753 48644 20760 48668
rect 20694 48588 20699 48644
rect 20755 48588 20760 48644
rect 20694 48564 20701 48588
rect 20753 48564 20760 48588
rect 20694 48508 20699 48564
rect 20755 48508 20760 48564
rect 20694 48494 20701 48508
rect 20753 48494 20760 48508
rect 20694 48484 20760 48494
rect 20694 48428 20699 48484
rect 20755 48428 20760 48484
rect 20694 48418 20760 48428
rect 20694 48404 20701 48418
rect 20753 48404 20760 48418
rect 20694 48348 20699 48404
rect 20755 48348 20760 48404
rect 20694 48324 20701 48348
rect 20753 48324 20760 48348
rect 20694 48268 20699 48324
rect 20755 48268 20760 48324
rect 20694 48244 20701 48268
rect 20753 48244 20760 48268
rect 20694 48188 20699 48244
rect 20755 48188 20760 48244
rect 20694 48174 20701 48188
rect 20753 48174 20760 48188
rect 20694 48159 20760 48174
rect 21782 48738 21848 48753
rect 21782 48724 21789 48738
rect 21841 48724 21848 48738
rect 21782 48668 21787 48724
rect 21843 48668 21848 48724
rect 21782 48644 21789 48668
rect 21841 48644 21848 48668
rect 21782 48588 21787 48644
rect 21843 48588 21848 48644
rect 21782 48564 21789 48588
rect 21841 48564 21848 48588
rect 21782 48508 21787 48564
rect 21843 48508 21848 48564
rect 21782 48494 21789 48508
rect 21841 48494 21848 48508
rect 21782 48484 21848 48494
rect 21782 48428 21787 48484
rect 21843 48428 21848 48484
rect 21782 48418 21848 48428
rect 21782 48404 21789 48418
rect 21841 48404 21848 48418
rect 21782 48348 21787 48404
rect 21843 48348 21848 48404
rect 21782 48324 21789 48348
rect 21841 48324 21848 48348
rect 21782 48268 21787 48324
rect 21843 48268 21848 48324
rect 21782 48244 21789 48268
rect 21841 48244 21848 48268
rect 21782 48188 21787 48244
rect 21843 48188 21848 48244
rect 21782 48174 21789 48188
rect 21841 48174 21848 48188
rect 21782 48159 21848 48174
rect 22870 48738 22936 48753
rect 22870 48724 22877 48738
rect 22929 48724 22936 48738
rect 22870 48668 22875 48724
rect 22931 48668 22936 48724
rect 22870 48644 22877 48668
rect 22929 48644 22936 48668
rect 22870 48588 22875 48644
rect 22931 48588 22936 48644
rect 22870 48564 22877 48588
rect 22929 48564 22936 48588
rect 22870 48508 22875 48564
rect 22931 48508 22936 48564
rect 22870 48494 22877 48508
rect 22929 48494 22936 48508
rect 22870 48484 22936 48494
rect 22870 48428 22875 48484
rect 22931 48428 22936 48484
rect 22870 48418 22936 48428
rect 22870 48404 22877 48418
rect 22929 48404 22936 48418
rect 22870 48348 22875 48404
rect 22931 48348 22936 48404
rect 22870 48324 22877 48348
rect 22929 48324 22936 48348
rect 22870 48268 22875 48324
rect 22931 48268 22936 48324
rect 22870 48244 22877 48268
rect 22929 48244 22936 48268
rect 22870 48188 22875 48244
rect 22931 48188 22936 48244
rect 22870 48174 22877 48188
rect 22929 48174 22936 48188
rect 22870 48159 22936 48174
rect 23958 48738 24024 48753
rect 23958 48724 23965 48738
rect 24017 48724 24024 48738
rect 23958 48668 23963 48724
rect 24019 48668 24024 48724
rect 23958 48644 23965 48668
rect 24017 48644 24024 48668
rect 23958 48588 23963 48644
rect 24019 48588 24024 48644
rect 23958 48564 23965 48588
rect 24017 48564 24024 48588
rect 23958 48508 23963 48564
rect 24019 48508 24024 48564
rect 23958 48494 23965 48508
rect 24017 48494 24024 48508
rect 23958 48484 24024 48494
rect 23958 48428 23963 48484
rect 24019 48428 24024 48484
rect 23958 48418 24024 48428
rect 23958 48404 23965 48418
rect 24017 48404 24024 48418
rect 23958 48348 23963 48404
rect 24019 48348 24024 48404
rect 23958 48324 23965 48348
rect 24017 48324 24024 48348
rect 23958 48268 23963 48324
rect 24019 48268 24024 48324
rect 23958 48244 23965 48268
rect 24017 48244 24024 48268
rect 23958 48188 23963 48244
rect 24019 48188 24024 48244
rect 23958 48174 23965 48188
rect 24017 48174 24024 48188
rect 23958 48159 24024 48174
rect 29398 48738 29464 48753
rect 29398 48724 29405 48738
rect 29457 48724 29464 48738
rect 29398 48668 29403 48724
rect 29459 48668 29464 48724
rect 29398 48644 29405 48668
rect 29457 48644 29464 48668
rect 29398 48588 29403 48644
rect 29459 48588 29464 48644
rect 29398 48564 29405 48588
rect 29457 48564 29464 48588
rect 29398 48508 29403 48564
rect 29459 48508 29464 48564
rect 29398 48494 29405 48508
rect 29457 48494 29464 48508
rect 29398 48484 29464 48494
rect 29398 48428 29403 48484
rect 29459 48428 29464 48484
rect 29398 48418 29464 48428
rect 29398 48404 29405 48418
rect 29457 48404 29464 48418
rect 29398 48348 29403 48404
rect 29459 48348 29464 48404
rect 29398 48324 29405 48348
rect 29457 48324 29464 48348
rect 29398 48268 29403 48324
rect 29459 48268 29464 48324
rect 29398 48244 29405 48268
rect 29457 48244 29464 48268
rect 29398 48188 29403 48244
rect 29459 48188 29464 48244
rect 29398 48174 29405 48188
rect 29457 48174 29464 48188
rect 29398 48159 29464 48174
rect 30486 48738 30552 48753
rect 30486 48724 30493 48738
rect 30545 48724 30552 48738
rect 30486 48668 30491 48724
rect 30547 48668 30552 48724
rect 30486 48644 30493 48668
rect 30545 48644 30552 48668
rect 30486 48588 30491 48644
rect 30547 48588 30552 48644
rect 30486 48564 30493 48588
rect 30545 48564 30552 48588
rect 30486 48508 30491 48564
rect 30547 48508 30552 48564
rect 30486 48494 30493 48508
rect 30545 48494 30552 48508
rect 30486 48484 30552 48494
rect 30486 48428 30491 48484
rect 30547 48428 30552 48484
rect 30486 48418 30552 48428
rect 30486 48404 30493 48418
rect 30545 48404 30552 48418
rect 30486 48348 30491 48404
rect 30547 48348 30552 48404
rect 30486 48324 30493 48348
rect 30545 48324 30552 48348
rect 30486 48268 30491 48324
rect 30547 48268 30552 48324
rect 30486 48244 30493 48268
rect 30545 48244 30552 48268
rect 30486 48188 30491 48244
rect 30547 48188 30552 48244
rect 30486 48174 30493 48188
rect 30545 48174 30552 48188
rect 30486 48159 30552 48174
rect 31574 48738 31640 48753
rect 31574 48724 31581 48738
rect 31633 48724 31640 48738
rect 31574 48668 31579 48724
rect 31635 48668 31640 48724
rect 31574 48644 31581 48668
rect 31633 48644 31640 48668
rect 31574 48588 31579 48644
rect 31635 48588 31640 48644
rect 31574 48564 31581 48588
rect 31633 48564 31640 48588
rect 31574 48508 31579 48564
rect 31635 48508 31640 48564
rect 31574 48494 31581 48508
rect 31633 48494 31640 48508
rect 31574 48484 31640 48494
rect 31574 48428 31579 48484
rect 31635 48428 31640 48484
rect 31574 48418 31640 48428
rect 31574 48404 31581 48418
rect 31633 48404 31640 48418
rect 31574 48348 31579 48404
rect 31635 48348 31640 48404
rect 31574 48324 31581 48348
rect 31633 48324 31640 48348
rect 31574 48268 31579 48324
rect 31635 48268 31640 48324
rect 31574 48244 31581 48268
rect 31633 48244 31640 48268
rect 31574 48188 31579 48244
rect 31635 48188 31640 48244
rect 31574 48174 31581 48188
rect 31633 48174 31640 48188
rect 31574 48159 31640 48174
rect 10177 47638 10216 47640
rect 10512 47638 10551 47640
rect 10177 47607 10551 47638
rect 17975 46735 18041 46750
rect 17975 46721 17982 46735
rect 18034 46721 18041 46735
rect 17975 46665 17980 46721
rect 18036 46665 18041 46721
rect 17975 46641 17982 46665
rect 18034 46641 18041 46665
rect 17975 46585 17980 46641
rect 18036 46585 18041 46641
rect 17975 46561 17982 46585
rect 18034 46561 18041 46585
rect 17975 46505 17980 46561
rect 18036 46505 18041 46561
rect 17975 46491 17982 46505
rect 18034 46491 18041 46505
rect 17975 46481 18041 46491
rect 17975 46425 17980 46481
rect 18036 46425 18041 46481
rect 17975 46415 18041 46425
rect 17975 46401 17982 46415
rect 18034 46401 18041 46415
rect 17975 46345 17980 46401
rect 18036 46345 18041 46401
rect 17975 46321 17982 46345
rect 18034 46321 18041 46345
rect -5924 46272 -5722 46284
rect -5924 39820 -5913 46272
rect -5733 39820 -5722 46272
rect 17975 46265 17980 46321
rect 18036 46265 18041 46321
rect 17975 46241 17982 46265
rect 18034 46241 18041 46265
rect 17975 46185 17980 46241
rect 18036 46185 18041 46241
rect 17975 46171 17982 46185
rect 18034 46171 18041 46185
rect 17975 46156 18041 46171
rect 19063 46735 19129 46750
rect 19063 46721 19070 46735
rect 19122 46721 19129 46735
rect 19063 46665 19068 46721
rect 19124 46665 19129 46721
rect 19063 46641 19070 46665
rect 19122 46641 19129 46665
rect 19063 46585 19068 46641
rect 19124 46585 19129 46641
rect 19063 46561 19070 46585
rect 19122 46561 19129 46585
rect 19063 46505 19068 46561
rect 19124 46505 19129 46561
rect 19063 46491 19070 46505
rect 19122 46491 19129 46505
rect 19063 46481 19129 46491
rect 19063 46425 19068 46481
rect 19124 46425 19129 46481
rect 19063 46415 19129 46425
rect 19063 46401 19070 46415
rect 19122 46401 19129 46415
rect 19063 46345 19068 46401
rect 19124 46345 19129 46401
rect 19063 46321 19070 46345
rect 19122 46321 19129 46345
rect 19063 46265 19068 46321
rect 19124 46265 19129 46321
rect 19063 46241 19070 46265
rect 19122 46241 19129 46265
rect 19063 46185 19068 46241
rect 19124 46185 19129 46241
rect 19063 46171 19070 46185
rect 19122 46171 19129 46185
rect 19063 46156 19129 46171
rect 20151 46735 20217 46750
rect 20151 46721 20158 46735
rect 20210 46721 20217 46735
rect 20151 46665 20156 46721
rect 20212 46665 20217 46721
rect 20151 46641 20158 46665
rect 20210 46641 20217 46665
rect 20151 46585 20156 46641
rect 20212 46585 20217 46641
rect 20151 46561 20158 46585
rect 20210 46561 20217 46585
rect 20151 46505 20156 46561
rect 20212 46505 20217 46561
rect 20151 46491 20158 46505
rect 20210 46491 20217 46505
rect 20151 46481 20217 46491
rect 20151 46425 20156 46481
rect 20212 46425 20217 46481
rect 20151 46415 20217 46425
rect 20151 46401 20158 46415
rect 20210 46401 20217 46415
rect 20151 46345 20156 46401
rect 20212 46345 20217 46401
rect 20151 46321 20158 46345
rect 20210 46321 20217 46345
rect 20151 46265 20156 46321
rect 20212 46265 20217 46321
rect 20151 46241 20158 46265
rect 20210 46241 20217 46265
rect 20151 46185 20156 46241
rect 20212 46185 20217 46241
rect 20151 46171 20158 46185
rect 20210 46171 20217 46185
rect 20151 46156 20217 46171
rect 21239 46735 21305 46750
rect 21239 46721 21246 46735
rect 21298 46721 21305 46735
rect 21239 46665 21244 46721
rect 21300 46665 21305 46721
rect 21239 46641 21246 46665
rect 21298 46641 21305 46665
rect 21239 46585 21244 46641
rect 21300 46585 21305 46641
rect 21239 46561 21246 46585
rect 21298 46561 21305 46585
rect 21239 46505 21244 46561
rect 21300 46505 21305 46561
rect 21239 46491 21246 46505
rect 21298 46491 21305 46505
rect 21239 46481 21305 46491
rect 21239 46425 21244 46481
rect 21300 46425 21305 46481
rect 21239 46415 21305 46425
rect 21239 46401 21246 46415
rect 21298 46401 21305 46415
rect 21239 46345 21244 46401
rect 21300 46345 21305 46401
rect 21239 46321 21246 46345
rect 21298 46321 21305 46345
rect 21239 46265 21244 46321
rect 21300 46265 21305 46321
rect 21239 46241 21246 46265
rect 21298 46241 21305 46265
rect 21239 46185 21244 46241
rect 21300 46185 21305 46241
rect 21239 46171 21246 46185
rect 21298 46171 21305 46185
rect 21239 46156 21305 46171
rect 22327 46735 22393 46750
rect 22327 46721 22334 46735
rect 22386 46721 22393 46735
rect 22327 46665 22332 46721
rect 22388 46665 22393 46721
rect 22327 46641 22334 46665
rect 22386 46641 22393 46665
rect 22327 46585 22332 46641
rect 22388 46585 22393 46641
rect 22327 46561 22334 46585
rect 22386 46561 22393 46585
rect 22327 46505 22332 46561
rect 22388 46505 22393 46561
rect 22327 46491 22334 46505
rect 22386 46491 22393 46505
rect 22327 46481 22393 46491
rect 22327 46425 22332 46481
rect 22388 46425 22393 46481
rect 22327 46415 22393 46425
rect 22327 46401 22334 46415
rect 22386 46401 22393 46415
rect 22327 46345 22332 46401
rect 22388 46345 22393 46401
rect 22327 46321 22334 46345
rect 22386 46321 22393 46345
rect 22327 46265 22332 46321
rect 22388 46265 22393 46321
rect 22327 46241 22334 46265
rect 22386 46241 22393 46265
rect 22327 46185 22332 46241
rect 22388 46185 22393 46241
rect 22327 46171 22334 46185
rect 22386 46171 22393 46185
rect 22327 46156 22393 46171
rect 24503 46735 24569 46750
rect 24503 46721 24510 46735
rect 24562 46721 24569 46735
rect 24503 46665 24508 46721
rect 24564 46665 24569 46721
rect 24503 46641 24510 46665
rect 24562 46641 24569 46665
rect 24503 46585 24508 46641
rect 24564 46585 24569 46641
rect 24503 46561 24510 46585
rect 24562 46561 24569 46585
rect 24503 46505 24508 46561
rect 24564 46505 24569 46561
rect 24503 46491 24510 46505
rect 24562 46491 24569 46505
rect 24503 46481 24569 46491
rect 24503 46425 24508 46481
rect 24564 46425 24569 46481
rect 24503 46415 24569 46425
rect 24503 46401 24510 46415
rect 24562 46401 24569 46415
rect 24503 46345 24508 46401
rect 24564 46345 24569 46401
rect 24503 46321 24510 46345
rect 24562 46321 24569 46345
rect 24503 46265 24508 46321
rect 24564 46265 24569 46321
rect 24503 46241 24510 46265
rect 24562 46241 24569 46265
rect 24503 46185 24508 46241
rect 24564 46185 24569 46241
rect 24503 46171 24510 46185
rect 24562 46171 24569 46185
rect 24503 46156 24569 46171
rect 25591 46735 25657 46750
rect 25591 46721 25598 46735
rect 25650 46721 25657 46735
rect 25591 46665 25596 46721
rect 25652 46665 25657 46721
rect 25591 46641 25598 46665
rect 25650 46641 25657 46665
rect 25591 46585 25596 46641
rect 25652 46585 25657 46641
rect 25591 46561 25598 46585
rect 25650 46561 25657 46585
rect 25591 46505 25596 46561
rect 25652 46505 25657 46561
rect 25591 46491 25598 46505
rect 25650 46491 25657 46505
rect 25591 46481 25657 46491
rect 25591 46425 25596 46481
rect 25652 46425 25657 46481
rect 25591 46415 25657 46425
rect 25591 46401 25598 46415
rect 25650 46401 25657 46415
rect 25591 46345 25596 46401
rect 25652 46345 25657 46401
rect 25591 46321 25598 46345
rect 25650 46321 25657 46345
rect 25591 46265 25596 46321
rect 25652 46265 25657 46321
rect 25591 46241 25598 46265
rect 25650 46241 25657 46265
rect 25591 46185 25596 46241
rect 25652 46185 25657 46241
rect 25591 46171 25598 46185
rect 25650 46171 25657 46185
rect 25591 46156 25657 46171
rect 26679 46735 26745 46750
rect 26679 46721 26686 46735
rect 26738 46721 26745 46735
rect 26679 46665 26684 46721
rect 26740 46665 26745 46721
rect 26679 46641 26686 46665
rect 26738 46641 26745 46665
rect 26679 46585 26684 46641
rect 26740 46585 26745 46641
rect 26679 46561 26686 46585
rect 26738 46561 26745 46585
rect 26679 46505 26684 46561
rect 26740 46505 26745 46561
rect 26679 46491 26686 46505
rect 26738 46491 26745 46505
rect 26679 46481 26745 46491
rect 26679 46425 26684 46481
rect 26740 46425 26745 46481
rect 26679 46415 26745 46425
rect 26679 46401 26686 46415
rect 26738 46401 26745 46415
rect 26679 46345 26684 46401
rect 26740 46345 26745 46401
rect 26679 46321 26686 46345
rect 26738 46321 26745 46345
rect 26679 46265 26684 46321
rect 26740 46265 26745 46321
rect 26679 46241 26686 46265
rect 26738 46241 26745 46265
rect 26679 46185 26684 46241
rect 26740 46185 26745 46241
rect 26679 46171 26686 46185
rect 26738 46171 26745 46185
rect 26679 46156 26745 46171
rect 27767 46735 27833 46750
rect 27767 46721 27774 46735
rect 27826 46721 27833 46735
rect 27767 46665 27772 46721
rect 27828 46665 27833 46721
rect 27767 46641 27774 46665
rect 27826 46641 27833 46665
rect 27767 46585 27772 46641
rect 27828 46585 27833 46641
rect 27767 46561 27774 46585
rect 27826 46561 27833 46585
rect 27767 46505 27772 46561
rect 27828 46505 27833 46561
rect 27767 46491 27774 46505
rect 27826 46491 27833 46505
rect 27767 46481 27833 46491
rect 27767 46425 27772 46481
rect 27828 46425 27833 46481
rect 27767 46415 27833 46425
rect 27767 46401 27774 46415
rect 27826 46401 27833 46415
rect 27767 46345 27772 46401
rect 27828 46345 27833 46401
rect 27767 46321 27774 46345
rect 27826 46321 27833 46345
rect 27767 46265 27772 46321
rect 27828 46265 27833 46321
rect 27767 46241 27774 46265
rect 27826 46241 27833 46265
rect 27767 46185 27772 46241
rect 27828 46185 27833 46241
rect 27767 46171 27774 46185
rect 27826 46171 27833 46185
rect 27767 46156 27833 46171
rect 28855 46735 28921 46750
rect 28855 46721 28862 46735
rect 28914 46721 28921 46735
rect 28855 46665 28860 46721
rect 28916 46665 28921 46721
rect 28855 46641 28862 46665
rect 28914 46641 28921 46665
rect 28855 46585 28860 46641
rect 28916 46585 28921 46641
rect 28855 46561 28862 46585
rect 28914 46561 28921 46585
rect 28855 46505 28860 46561
rect 28916 46505 28921 46561
rect 28855 46491 28862 46505
rect 28914 46491 28921 46505
rect 28855 46481 28921 46491
rect 28855 46425 28860 46481
rect 28916 46425 28921 46481
rect 28855 46415 28921 46425
rect 28855 46401 28862 46415
rect 28914 46401 28921 46415
rect 28855 46345 28860 46401
rect 28916 46345 28921 46401
rect 28855 46321 28862 46345
rect 28914 46321 28921 46345
rect 28855 46265 28860 46321
rect 28916 46265 28921 46321
rect 28855 46241 28862 46265
rect 28914 46241 28921 46265
rect 28855 46185 28860 46241
rect 28916 46185 28921 46241
rect 28855 46171 28862 46185
rect 28914 46171 28921 46185
rect 28855 46156 28921 46171
rect 29943 46735 30009 46750
rect 29943 46721 29950 46735
rect 30002 46721 30009 46735
rect 29943 46665 29948 46721
rect 30004 46665 30009 46721
rect 29943 46641 29950 46665
rect 30002 46641 30009 46665
rect 29943 46585 29948 46641
rect 30004 46585 30009 46641
rect 29943 46561 29950 46585
rect 30002 46561 30009 46585
rect 29943 46505 29948 46561
rect 30004 46505 30009 46561
rect 29943 46491 29950 46505
rect 30002 46491 30009 46505
rect 29943 46481 30009 46491
rect 29943 46425 29948 46481
rect 30004 46425 30009 46481
rect 29943 46415 30009 46425
rect 29943 46401 29950 46415
rect 30002 46401 30009 46415
rect 29943 46345 29948 46401
rect 30004 46345 30009 46401
rect 29943 46321 29950 46345
rect 30002 46321 30009 46345
rect 29943 46265 29948 46321
rect 30004 46265 30009 46321
rect 29943 46241 29950 46265
rect 30002 46241 30009 46265
rect 29943 46185 29948 46241
rect 30004 46185 30009 46241
rect 29943 46171 29950 46185
rect 30002 46171 30009 46185
rect 29943 46156 30009 46171
rect 31031 46735 31097 46750
rect 31031 46721 31038 46735
rect 31090 46721 31097 46735
rect 31031 46665 31036 46721
rect 31092 46665 31097 46721
rect 31031 46641 31038 46665
rect 31090 46641 31097 46665
rect 31031 46585 31036 46641
rect 31092 46585 31097 46641
rect 31031 46561 31038 46585
rect 31090 46561 31097 46585
rect 31031 46505 31036 46561
rect 31092 46505 31097 46561
rect 31031 46491 31038 46505
rect 31090 46491 31097 46505
rect 31031 46481 31097 46491
rect 31031 46425 31036 46481
rect 31092 46425 31097 46481
rect 31031 46415 31097 46425
rect 31031 46401 31038 46415
rect 31090 46401 31097 46415
rect 31031 46345 31036 46401
rect 31092 46345 31097 46401
rect 31031 46321 31038 46345
rect 31090 46321 31097 46345
rect 31031 46265 31036 46321
rect 31092 46265 31097 46321
rect 40589 46371 40653 46385
rect 40589 46315 40593 46371
rect 40649 46315 40653 46371
rect 40589 46301 40653 46315
rect 31031 46241 31038 46265
rect 31090 46241 31097 46265
rect 31031 46185 31036 46241
rect 31092 46185 31097 46241
rect 31031 46171 31038 46185
rect 31090 46171 31097 46185
rect 31031 46156 31097 46171
rect 10180 46127 10551 46138
rect 344 45843 558 45854
rect 344 44319 361 45843
rect 541 44319 558 45843
rect 344 44308 558 44319
rect 352 41381 512 41393
rect 352 41367 374 41381
rect 490 41367 512 41381
rect 352 39871 364 41367
rect 500 39871 512 41367
rect 352 39857 374 39871
rect 490 39857 512 39871
rect 10180 39867 10211 46127
rect 10519 39867 10551 46127
rect 18245 45744 18309 45758
rect 18245 45688 18249 45744
rect 18305 45688 18309 45744
rect 18245 45674 18309 45688
rect 18791 45744 18855 45758
rect 18791 45688 18795 45744
rect 18851 45688 18855 45744
rect 18791 45674 18855 45688
rect 19337 45735 19401 45749
rect 19337 45679 19341 45735
rect 19397 45679 19401 45735
rect 19337 45665 19401 45679
rect 19882 45734 19946 45748
rect 19882 45678 19886 45734
rect 19942 45678 19946 45734
rect 19882 45664 19946 45678
rect 21513 45722 21577 45736
rect 21513 45666 21517 45722
rect 21573 45666 21577 45722
rect 21513 45652 21577 45666
rect 22056 45719 22120 45733
rect 22056 45663 22060 45719
rect 22116 45663 22120 45719
rect 22056 45649 22120 45663
rect 22598 45718 22662 45732
rect 22598 45662 22602 45718
rect 22658 45662 22662 45718
rect 22598 45648 22662 45662
rect 23145 45723 23209 45737
rect 23145 45667 23149 45723
rect 23205 45667 23209 45723
rect 23145 45653 23209 45667
rect 25863 45734 25927 45748
rect 25863 45678 25867 45734
rect 25923 45678 25927 45734
rect 25863 45664 25927 45678
rect 26406 45738 26470 45752
rect 26406 45682 26410 45738
rect 26466 45682 26470 45738
rect 26406 45668 26470 45682
rect 26948 45732 27012 45746
rect 26948 45676 26952 45732
rect 27008 45676 27012 45732
rect 26948 45662 27012 45676
rect 27505 45723 27569 45737
rect 27505 45667 27509 45723
rect 27565 45667 27569 45723
rect 27505 45653 27569 45667
rect 29129 45734 29193 45748
rect 29129 45678 29133 45734
rect 29189 45678 29193 45734
rect 29129 45664 29193 45678
rect 29673 45727 29737 45741
rect 29673 45671 29677 45727
rect 29733 45671 29737 45727
rect 29673 45657 29737 45671
rect 30223 45731 30287 45745
rect 30223 45675 30227 45731
rect 30283 45675 30287 45731
rect 30223 45661 30287 45675
rect 30756 45731 30820 45745
rect 30756 45675 30760 45731
rect 30816 45675 30820 45731
rect 30756 45661 30820 45675
rect 39557 44887 39621 44901
rect 39557 44831 39561 44887
rect 39617 44831 39621 44887
rect 39557 44817 39621 44831
rect 40595 44830 40647 46301
rect 41146 45815 41210 45829
rect 41146 45759 41150 45815
rect 41206 45759 41210 45815
rect 41146 45745 41210 45759
rect 40988 44987 41052 45001
rect 40988 44931 40992 44987
rect 41048 44931 41052 44987
rect 40988 44917 41052 44931
rect 39557 44697 39621 44711
rect 39557 44641 39561 44697
rect 39617 44641 39621 44697
rect 39557 44627 39621 44641
rect 39557 43737 39621 43751
rect 39557 43681 39561 43737
rect 39617 43681 39621 43737
rect 39557 43667 39621 43681
rect 40595 43680 40647 44778
rect 40995 44819 41047 44917
rect 40894 44762 40946 44772
rect 40995 44757 41047 44767
rect 41152 44823 41204 45745
rect 44754 45068 45306 45084
rect 44754 45012 44762 45068
rect 44818 45066 44842 45068
rect 44898 45066 44922 45068
rect 44978 45066 45002 45068
rect 45058 45066 45082 45068
rect 45138 45066 45162 45068
rect 45218 45066 45242 45068
rect 44832 45014 44842 45066
rect 44898 45014 44908 45066
rect 45152 45014 45162 45066
rect 45218 45014 45228 45066
rect 44818 45012 44842 45014
rect 44898 45012 44922 45014
rect 44978 45012 45002 45014
rect 45058 45012 45082 45014
rect 45138 45012 45162 45014
rect 45218 45012 45242 45014
rect 45298 45012 45306 45068
rect 44754 44997 45306 45012
rect 40894 44617 40946 44710
rect 40888 44603 40952 44617
rect 40888 44547 40892 44603
rect 40948 44547 40952 44603
rect 40888 44533 40952 44547
rect 40988 43837 41052 43851
rect 40988 43781 40992 43837
rect 41048 43781 41052 43837
rect 40988 43767 41052 43781
rect 40595 43618 40647 43628
rect 40995 43669 41047 43767
rect 40894 43612 40946 43622
rect 39557 43547 39621 43561
rect 39557 43491 39561 43547
rect 39617 43491 39621 43547
rect 39557 43477 39621 43491
rect 40995 43607 41047 43617
rect 41152 43673 41204 44771
rect 46294 44929 46530 44949
rect 46294 44713 46304 44929
rect 46520 44713 46530 44929
rect 46294 44693 46530 44713
rect 41516 44522 41874 44537
rect 41516 44520 41547 44522
rect 41603 44520 41627 44522
rect 41683 44520 41707 44522
rect 41763 44520 41787 44522
rect 41843 44520 41874 44522
rect 41516 44468 41541 44520
rect 41603 44468 41605 44520
rect 41785 44468 41787 44520
rect 41849 44468 41874 44520
rect 41516 44466 41547 44468
rect 41603 44466 41627 44468
rect 41683 44466 41707 44468
rect 41763 44466 41787 44468
rect 41843 44466 41874 44468
rect 41516 44452 41874 44466
rect 44766 43917 45293 43935
rect 44766 43915 44801 43917
rect 44857 43915 44881 43917
rect 44937 43915 44961 43917
rect 45017 43915 45041 43917
rect 45097 43915 45121 43917
rect 45177 43915 45201 43917
rect 45257 43915 45293 43917
rect 44766 43863 44779 43915
rect 44959 43863 44961 43915
rect 45023 43863 45035 43915
rect 45097 43863 45099 43915
rect 45279 43863 45293 43915
rect 44766 43861 44801 43863
rect 44857 43861 44881 43863
rect 44937 43861 44961 43863
rect 45017 43861 45041 43863
rect 45097 43861 45121 43863
rect 45177 43861 45201 43863
rect 45257 43861 45293 43863
rect 44766 43844 45293 43861
rect 41152 43611 41204 43621
rect 46282 43778 46518 43798
rect 40894 43467 40946 43560
rect 46282 43562 46292 43778
rect 46508 43562 46518 43778
rect 46282 43542 46518 43562
rect 40888 43453 40952 43467
rect 40888 43397 40892 43453
rect 40948 43397 40952 43453
rect 40888 43383 40952 43397
rect 41514 43372 41872 43387
rect 41514 43370 41545 43372
rect 41601 43370 41625 43372
rect 41681 43370 41705 43372
rect 41761 43370 41785 43372
rect 41841 43370 41872 43372
rect 41514 43318 41539 43370
rect 41601 43318 41603 43370
rect 41783 43318 41785 43370
rect 41847 43318 41872 43370
rect 41514 43316 41545 43318
rect 41601 43316 41625 43318
rect 41681 43316 41705 43318
rect 41761 43316 41785 43318
rect 41841 43316 41872 43318
rect 41514 43302 41872 43316
rect 40589 42681 40653 42695
rect 40589 42625 40593 42681
rect 40649 42625 40653 42681
rect 40589 42611 40653 42625
rect 39557 41197 39621 41211
rect 39557 41141 39561 41197
rect 39617 41141 39621 41197
rect 39557 41127 39621 41141
rect 40595 41140 40647 42611
rect 41146 42125 41210 42139
rect 41146 42069 41150 42125
rect 41206 42069 41210 42125
rect 41146 42055 41210 42069
rect 40988 41297 41052 41311
rect 40988 41241 40992 41297
rect 41048 41241 41052 41297
rect 40988 41227 41052 41241
rect 39557 41007 39621 41021
rect 39557 40951 39561 41007
rect 39617 40951 39621 41007
rect 39557 40937 39621 40951
rect 10180 39857 10551 39867
rect 39557 39927 39621 39941
rect 39557 39871 39561 39927
rect 39617 39871 39621 39927
rect 39557 39857 39621 39871
rect 40595 39870 40647 41088
rect 40995 41129 41047 41227
rect 40894 41072 40946 41082
rect 40995 41067 41047 41077
rect 41152 41133 41204 42055
rect 44756 41375 45283 41393
rect 44756 41373 44791 41375
rect 44847 41373 44871 41375
rect 44927 41373 44951 41375
rect 45007 41373 45031 41375
rect 45087 41373 45111 41375
rect 45167 41373 45191 41375
rect 45247 41373 45283 41375
rect 44756 41321 44769 41373
rect 44949 41321 44951 41373
rect 45013 41321 45025 41373
rect 45087 41321 45089 41373
rect 45269 41321 45283 41373
rect 44756 41319 44791 41321
rect 44847 41319 44871 41321
rect 44927 41319 44951 41321
rect 45007 41319 45031 41321
rect 45087 41319 45111 41321
rect 45167 41319 45191 41321
rect 45247 41319 45283 41321
rect 44756 41302 45283 41319
rect 40894 40927 40946 41020
rect 40888 40913 40952 40927
rect 40888 40857 40892 40913
rect 40948 40857 40952 40913
rect 40888 40843 40952 40857
rect 40988 40027 41052 40041
rect 40988 39971 40992 40027
rect 41048 39971 41052 40027
rect 40988 39957 41052 39971
rect -5924 39809 -5722 39820
rect -5684 39846 -148 39856
rect -5684 39824 -5662 39846
rect -170 39824 -148 39846
rect 352 39845 512 39857
rect -6989 39747 -6983 39799
rect -6931 39747 -6919 39799
rect -6867 39747 -6861 39799
rect -6989 39731 -6861 39747
rect -27077 39671 -27062 39727
rect -27006 39671 -26990 39727
rect -27077 39669 -26990 39671
rect -27077 39647 -27060 39669
rect -27008 39647 -26990 39669
rect -5684 39688 -5664 39824
rect -168 39688 -148 39824
rect 40595 39808 40647 39818
rect 40995 39859 41047 39957
rect 40894 39802 40946 39812
rect -5684 39666 -5662 39688
rect -170 39666 -148 39688
rect 39557 39737 39621 39751
rect 39557 39681 39561 39737
rect 39617 39681 39621 39737
rect 39557 39667 39621 39681
rect 40995 39797 41047 39807
rect 41152 39863 41204 41081
rect 46140 41246 46376 41266
rect 46140 41030 46150 41246
rect 46366 41030 46376 41246
rect 46140 41010 46376 41030
rect 41432 40831 41790 40846
rect 41432 40829 41463 40831
rect 41519 40829 41543 40831
rect 41599 40829 41623 40831
rect 41679 40829 41703 40831
rect 41759 40829 41790 40831
rect 41432 40777 41457 40829
rect 41519 40777 41521 40829
rect 41701 40777 41703 40829
rect 41765 40777 41790 40829
rect 41432 40775 41463 40777
rect 41519 40775 41543 40777
rect 41599 40775 41623 40777
rect 41679 40775 41703 40777
rect 41759 40775 41790 40777
rect 41432 40761 41790 40775
rect 44756 40105 45283 40123
rect 44756 40103 44791 40105
rect 44847 40103 44871 40105
rect 44927 40103 44951 40105
rect 45007 40103 45031 40105
rect 45087 40103 45111 40105
rect 45167 40103 45191 40105
rect 45247 40103 45283 40105
rect 44756 40051 44769 40103
rect 44949 40051 44951 40103
rect 45013 40051 45025 40103
rect 45087 40051 45089 40103
rect 45269 40051 45283 40103
rect 44756 40049 44791 40051
rect 44847 40049 44871 40051
rect 44927 40049 44951 40051
rect 45007 40049 45031 40051
rect 45087 40049 45111 40051
rect 45167 40049 45191 40051
rect 45247 40049 45283 40051
rect 44756 40032 45283 40049
rect 41152 39801 41204 39811
rect 46111 39956 46347 39976
rect -5684 39656 -148 39666
rect 40894 39657 40946 39750
rect 46111 39740 46121 39956
rect 46337 39740 46347 39956
rect 46111 39720 46347 39740
rect -27077 39591 -27062 39647
rect -27006 39591 -26990 39647
rect -27077 39567 -27060 39591
rect -27008 39567 -26990 39591
rect 40888 39643 40952 39657
rect 40888 39587 40892 39643
rect 40948 39587 40952 39643
rect 40888 39573 40952 39587
rect -27077 39511 -27062 39567
rect -27006 39511 -26990 39567
rect 41430 39562 41788 39577
rect 41430 39560 41461 39562
rect 41517 39560 41541 39562
rect 41597 39560 41621 39562
rect 41677 39560 41701 39562
rect 41757 39560 41788 39562
rect -27077 39489 -27060 39511
rect -27008 39489 -26990 39511
rect -27077 39466 -26990 39489
rect -18883 39520 -18807 39547
rect -18883 39498 -18871 39520
rect -18819 39498 -18807 39520
rect -18883 39442 -18873 39498
rect -18817 39442 -18807 39498
rect 41430 39508 41455 39560
rect 41517 39508 41519 39560
rect 41699 39508 41701 39560
rect 41763 39508 41788 39560
rect 41430 39506 41461 39508
rect 41517 39506 41541 39508
rect 41597 39506 41621 39508
rect 41677 39506 41701 39508
rect 41757 39506 41788 39508
rect 41430 39492 41788 39506
rect -18883 39418 -18871 39442
rect -18819 39418 -18807 39442
rect -18883 39362 -18873 39418
rect -18817 39362 -18807 39418
rect -18883 39340 -18871 39362
rect -18819 39340 -18807 39362
rect -18883 39338 -18807 39340
rect -18883 39282 -18873 39338
rect -18817 39282 -18807 39338
rect -18883 39276 -18871 39282
rect -18819 39276 -18807 39282
rect -18883 39264 -18807 39276
rect -18883 39258 -18871 39264
rect -18819 39258 -18807 39264
rect -18883 39202 -18873 39258
rect -18817 39202 -18807 39258
rect -18883 39200 -18807 39202
rect -18883 39178 -18871 39200
rect -18819 39178 -18807 39200
rect -31812 39150 -31748 39176
rect -31812 39144 -31806 39150
rect -31754 39144 -31748 39150
rect -31812 39088 -31808 39144
rect -31752 39088 -31748 39144
rect -31812 39086 -31748 39088
rect -31812 39064 -31806 39086
rect -31754 39064 -31748 39086
rect -31812 39008 -31808 39064
rect -31752 39008 -31748 39064
rect -31812 38984 -31806 39008
rect -31754 38984 -31748 39008
rect -31812 38928 -31808 38984
rect -31752 38928 -31748 38984
rect -31812 38906 -31806 38928
rect -31754 38906 -31748 38928
rect -31812 38904 -31748 38906
rect -31812 38848 -31808 38904
rect -31752 38848 -31748 38904
rect -31812 38842 -31806 38848
rect -31754 38842 -31748 38848
rect -31812 38817 -31748 38842
rect -27082 39118 -26998 39130
rect -27082 39104 -27066 39118
rect -27014 39104 -26998 39118
rect -27082 39048 -27068 39104
rect -27012 39048 -26998 39104
rect -27082 39024 -27066 39048
rect -27014 39024 -26998 39048
rect -27082 38968 -27068 39024
rect -27012 38968 -26998 39024
rect -27082 38944 -27066 38968
rect -27014 38944 -26998 38968
rect -27082 38888 -27068 38944
rect -27012 38888 -26998 38944
rect -27082 38874 -27066 38888
rect -27014 38874 -26998 38888
rect -27082 38864 -26998 38874
rect -27082 38808 -27068 38864
rect -27012 38808 -26998 38864
rect -27082 38798 -26998 38808
rect -27082 38784 -27066 38798
rect -27014 38784 -26998 38798
rect -27082 38728 -27068 38784
rect -27012 38728 -26998 38784
rect -27082 38704 -27066 38728
rect -27014 38704 -26998 38728
rect -27082 38648 -27068 38704
rect -27012 38648 -26998 38704
rect -27082 38624 -27066 38648
rect -27014 38624 -26998 38648
rect -31811 38605 -31747 38623
rect -31811 38549 -31807 38605
rect -31751 38549 -31747 38605
rect -31811 38543 -31805 38549
rect -31753 38543 -31747 38549
rect -31811 38531 -31747 38543
rect -31811 38525 -31805 38531
rect -31753 38525 -31747 38531
rect -31811 38469 -31807 38525
rect -31751 38469 -31747 38525
rect -31811 38467 -31747 38469
rect -31811 38445 -31805 38467
rect -31753 38445 -31747 38467
rect -31811 38389 -31807 38445
rect -31751 38389 -31747 38445
rect -27082 38568 -27068 38624
rect -27012 38568 -26998 38624
rect -27082 38554 -27066 38568
rect -27014 38554 -26998 38568
rect -27082 38544 -26998 38554
rect -27082 38488 -27068 38544
rect -27012 38488 -26998 38544
rect -27082 38478 -26998 38488
rect -27082 38464 -27066 38478
rect -27014 38464 -26998 38478
rect -31811 38365 -31805 38389
rect -31753 38365 -31747 38389
rect -31811 38309 -31807 38365
rect -31751 38309 -31747 38365
rect -29614 38409 -29150 38423
rect -29614 38353 -29610 38409
rect -29554 38407 -29530 38409
rect -29474 38407 -29450 38409
rect -29394 38407 -29370 38409
rect -29314 38407 -29290 38409
rect -29234 38407 -29210 38409
rect -29548 38355 -29536 38407
rect -29474 38355 -29472 38407
rect -29292 38355 -29290 38407
rect -29228 38355 -29216 38407
rect -29554 38353 -29530 38355
rect -29474 38353 -29450 38355
rect -29394 38353 -29370 38355
rect -29314 38353 -29290 38355
rect -29234 38353 -29210 38355
rect -29154 38353 -29150 38409
rect -29614 38339 -29150 38353
rect -27082 38408 -27068 38464
rect -27012 38408 -26998 38464
rect -27082 38384 -27066 38408
rect -27014 38384 -26998 38408
rect -31811 38287 -31805 38309
rect -31753 38287 -31747 38309
rect -31811 38285 -31747 38287
rect -31811 38229 -31807 38285
rect -31751 38229 -31747 38285
rect -27082 38328 -27068 38384
rect -27012 38328 -26998 38384
rect -27082 38304 -27066 38328
rect -27014 38304 -26998 38328
rect -31030 38256 -30901 38266
rect -31811 38223 -31805 38229
rect -31753 38223 -31747 38229
rect -31811 38211 -31747 38223
rect -31811 38205 -31805 38211
rect -31753 38205 -31747 38211
rect -31811 38149 -31807 38205
rect -31751 38149 -31747 38205
rect -31047 38250 -30885 38256
rect -31047 38198 -31024 38250
rect -30972 38198 -30960 38250
rect -30908 38198 -30885 38250
rect -27082 38248 -27068 38304
rect -27012 38248 -26998 38304
rect -27082 38234 -27066 38248
rect -27014 38234 -26998 38248
rect -27082 38222 -26998 38234
rect -18883 39122 -18873 39178
rect -18817 39122 -18807 39178
rect -18883 39098 -18871 39122
rect -18819 39098 -18807 39122
rect -18883 39042 -18873 39098
rect -18817 39042 -18807 39098
rect -18883 39020 -18871 39042
rect -18819 39020 -18807 39042
rect -18883 39018 -18807 39020
rect -18883 38962 -18873 39018
rect -18817 38962 -18807 39018
rect 7082 39210 7318 39220
rect 12542 39210 12778 39220
rect 7082 39182 12778 39210
rect 7082 39002 7110 39182
rect 7290 39002 12570 39182
rect 12750 39002 12778 39182
rect 7082 38974 12778 39002
rect 7082 38964 7318 38974
rect 12542 38964 12778 38974
rect -18883 38956 -18871 38962
rect -18819 38956 -18807 38962
rect -18883 38944 -18807 38956
rect -18883 38938 -18871 38944
rect -18819 38938 -18807 38944
rect -18883 38882 -18873 38938
rect -18817 38882 -18807 38938
rect -18883 38880 -18807 38882
rect -18883 38858 -18871 38880
rect -18819 38858 -18807 38880
rect -18883 38802 -18873 38858
rect -18817 38802 -18807 38858
rect 1473 38874 1537 38888
rect 1473 38818 1477 38874
rect 1533 38818 1537 38874
rect 1473 38804 1537 38818
rect 2513 38869 2595 38891
rect 2513 38813 2526 38869
rect 2582 38813 2595 38869
rect -18883 38778 -18871 38802
rect -18819 38778 -18807 38802
rect -18883 38722 -18873 38778
rect -18817 38722 -18807 38778
rect -18883 38700 -18871 38722
rect -18819 38700 -18807 38722
rect -18883 38698 -18807 38700
rect -18883 38642 -18873 38698
rect -18817 38642 -18807 38698
rect -18883 38636 -18871 38642
rect -18819 38636 -18807 38642
rect -18883 38624 -18807 38636
rect 2513 38799 2528 38813
rect 2580 38799 2595 38813
rect 2513 38789 2595 38799
rect 2513 38733 2526 38789
rect 2582 38733 2595 38789
rect 2513 38723 2595 38733
rect 2513 38709 2528 38723
rect 2580 38709 2595 38723
rect 2513 38653 2526 38709
rect 2582 38653 2595 38709
rect 2513 38632 2595 38653
rect -18883 38618 -18871 38624
rect -18819 38618 -18807 38624
rect -18883 38562 -18873 38618
rect -18817 38562 -18807 38618
rect 93 38566 157 38576
rect 1230 38566 1294 38576
rect -18883 38560 -18807 38562
rect -18883 38538 -18871 38560
rect -18819 38538 -18807 38560
rect -18883 38482 -18873 38538
rect -18817 38482 -18807 38538
rect 87 38560 1294 38566
rect 87 38508 99 38560
rect 151 38508 1236 38560
rect 1288 38508 1294 38560
rect 87 38502 1294 38508
rect 93 38492 157 38502
rect 1230 38492 1294 38502
rect 2626 38568 2690 38578
rect 5361 38568 5425 38578
rect 2626 38562 5425 38568
rect 2626 38510 2632 38562
rect 2684 38510 5367 38562
rect 5419 38510 5425 38562
rect 2626 38504 5425 38510
rect 2626 38494 2690 38504
rect 5361 38494 5425 38504
rect -18883 38458 -18871 38482
rect -18819 38458 -18807 38482
rect -18883 38402 -18873 38458
rect -18817 38402 -18807 38458
rect -18883 38380 -18871 38402
rect -18819 38380 -18807 38402
rect -18883 38378 -18807 38380
rect -18883 38322 -18873 38378
rect -18817 38322 -18807 38378
rect -18883 38316 -18871 38322
rect -18819 38316 -18807 38322
rect -18883 38304 -18807 38316
rect -18883 38298 -18871 38304
rect -18819 38298 -18807 38304
rect -18883 38242 -18873 38298
rect -18817 38242 -18807 38298
rect -18883 38240 -18807 38242
rect -31047 38192 -30885 38198
rect -18883 38218 -18871 38240
rect -18819 38218 -18807 38240
rect -31811 38131 -31747 38149
rect -35518 37558 -35282 37578
rect -35518 37342 -35508 37558
rect -35292 37342 -35282 37558
rect -35518 37322 -35282 37342
rect -31030 27923 -30901 38192
rect -18883 38162 -18873 38218
rect -18817 38162 -18807 38218
rect -18883 38138 -18871 38162
rect -18819 38138 -18807 38162
rect -18883 38082 -18873 38138
rect -18817 38082 -18807 38138
rect -18883 38060 -18871 38082
rect -18819 38060 -18807 38082
rect 2515 38396 2614 38430
rect 2515 38340 2536 38396
rect 2592 38340 2614 38396
rect 2515 38330 2614 38340
rect 2515 38316 2538 38330
rect 2590 38316 2614 38330
rect 2515 38260 2536 38316
rect 2592 38260 2614 38316
rect 2515 38236 2538 38260
rect 2590 38236 2614 38260
rect 2515 38180 2536 38236
rect 2592 38180 2614 38236
rect 2515 38156 2538 38180
rect 2590 38156 2614 38180
rect 2515 38100 2536 38156
rect 2592 38100 2614 38156
rect 2515 38086 2538 38100
rect 2590 38086 2614 38100
rect -18883 38058 -18807 38060
rect -18883 38002 -18873 38058
rect -18817 38002 -18807 38058
rect -18883 37996 -18871 38002
rect -18819 37996 -18807 38002
rect -18883 37984 -18807 37996
rect 1996 38065 2060 38079
rect 1996 38009 2000 38065
rect 2056 38009 2060 38065
rect 1996 37995 2060 38009
rect 2515 38076 2614 38086
rect 5361 38155 5425 38165
rect 7236 38155 7300 38165
rect 5361 38149 7300 38155
rect 5361 38097 5367 38149
rect 5419 38097 7242 38149
rect 7294 38097 7300 38149
rect 5361 38091 7300 38097
rect 5361 38081 5425 38091
rect 7236 38081 7300 38091
rect 2515 38020 2536 38076
rect 2592 38020 2614 38076
rect 2515 37986 2614 38020
rect -18883 37978 -18871 37984
rect -18819 37978 -18807 37984
rect -18883 37922 -18873 37978
rect -18817 37922 -18807 37978
rect -18883 37920 -18807 37922
rect -18883 37898 -18871 37920
rect -18819 37898 -18807 37920
rect -18883 37842 -18873 37898
rect -18817 37842 -18807 37898
rect -18883 37818 -18871 37842
rect -18819 37818 -18807 37842
rect -18883 37762 -18873 37818
rect -18817 37762 -18807 37818
rect -18883 37740 -18871 37762
rect -18819 37740 -18807 37762
rect -18883 37738 -18807 37740
rect -18883 37682 -18873 37738
rect -18817 37682 -18807 37738
rect -18883 37676 -18871 37682
rect -18819 37676 -18807 37682
rect -18883 37664 -18807 37676
rect -18883 37658 -18871 37664
rect -18819 37658 -18807 37664
rect -18883 37602 -18873 37658
rect -18817 37602 -18807 37658
rect -18883 37600 -18807 37602
rect -18883 37578 -18871 37600
rect -18819 37578 -18807 37600
rect -18883 37522 -18873 37578
rect -18817 37522 -18807 37578
rect 93 37651 157 37661
rect 3427 37651 3491 37661
rect 9428 37651 9492 37661
rect 93 37645 9492 37651
rect 93 37593 99 37645
rect 151 37593 3433 37645
rect 3485 37593 9434 37645
rect 9486 37593 9492 37645
rect 93 37587 9492 37593
rect 93 37577 157 37587
rect 3427 37577 3491 37587
rect 9428 37577 9492 37587
rect -18883 37498 -18871 37522
rect -18819 37498 -18807 37522
rect -30199 37475 -30070 37496
rect -30217 37469 -30055 37475
rect -30217 37417 -30193 37469
rect -30141 37417 -30129 37469
rect -30077 37417 -30055 37469
rect -30217 37411 -30055 37417
rect -18883 37442 -18873 37498
rect -18817 37442 -18807 37498
rect -18883 37420 -18871 37442
rect -18819 37420 -18807 37442
rect -18883 37418 -18807 37420
rect -30199 29281 -30070 37411
rect -27079 37351 -26995 37363
rect -27079 37337 -27063 37351
rect -27011 37337 -26995 37351
rect -29652 37319 -29143 37333
rect -29652 37317 -29626 37319
rect -29570 37317 -29546 37319
rect -29490 37317 -29466 37319
rect -29410 37317 -29386 37319
rect -29330 37317 -29306 37319
rect -29250 37317 -29226 37319
rect -29170 37317 -29143 37319
rect -29652 37265 -29648 37317
rect -29468 37265 -29466 37317
rect -29404 37265 -29392 37317
rect -29330 37265 -29328 37317
rect -29148 37265 -29143 37317
rect -29652 37263 -29626 37265
rect -29570 37263 -29546 37265
rect -29490 37263 -29466 37265
rect -29410 37263 -29386 37265
rect -29330 37263 -29306 37265
rect -29250 37263 -29226 37265
rect -29170 37263 -29143 37265
rect -29652 37249 -29143 37263
rect -27079 37281 -27065 37337
rect -27009 37281 -26995 37337
rect -27079 37257 -27063 37281
rect -27011 37257 -26995 37281
rect -27079 37201 -27065 37257
rect -27009 37201 -26995 37257
rect -27079 37177 -27063 37201
rect -27011 37177 -26995 37201
rect -27079 37121 -27065 37177
rect -27009 37121 -26995 37177
rect -27079 37107 -27063 37121
rect -27011 37107 -26995 37121
rect -27079 37097 -26995 37107
rect -27079 37041 -27065 37097
rect -27009 37041 -26995 37097
rect -27079 37031 -26995 37041
rect -27079 37017 -27063 37031
rect -27011 37017 -26995 37031
rect -27079 36961 -27065 37017
rect -27009 36961 -26995 37017
rect -27079 36937 -27063 36961
rect -27011 36937 -26995 36961
rect -27079 36881 -27065 36937
rect -27009 36881 -26995 36937
rect -27079 36857 -27063 36881
rect -27011 36857 -26995 36881
rect -27079 36801 -27065 36857
rect -27009 36801 -26995 36857
rect -27079 36787 -27063 36801
rect -27011 36787 -26995 36801
rect -27079 36777 -26995 36787
rect -27079 36721 -27065 36777
rect -27009 36721 -26995 36777
rect -27079 36711 -26995 36721
rect -27079 36697 -27063 36711
rect -27011 36697 -26995 36711
rect -27079 36641 -27065 36697
rect -27009 36641 -26995 36697
rect -27079 36617 -27063 36641
rect -27011 36617 -26995 36641
rect -27079 36561 -27065 36617
rect -27009 36561 -26995 36617
rect -27079 36537 -27063 36561
rect -27011 36537 -26995 36561
rect -27079 36481 -27065 36537
rect -27009 36481 -26995 36537
rect -27079 36467 -27063 36481
rect -27011 36467 -26995 36481
rect -27079 36455 -26995 36467
rect -18883 37362 -18873 37418
rect -18817 37362 -18807 37418
rect -18883 37356 -18871 37362
rect -18819 37356 -18807 37362
rect -18883 37344 -18807 37356
rect -18883 37338 -18871 37344
rect -18819 37338 -18807 37344
rect -18883 37282 -18873 37338
rect -18817 37282 -18807 37338
rect -18883 37280 -18807 37282
rect -18883 37258 -18871 37280
rect -18819 37258 -18807 37280
rect -18883 37202 -18873 37258
rect -18817 37202 -18807 37258
rect -18883 37178 -18871 37202
rect -18819 37178 -18807 37202
rect -18883 37122 -18873 37178
rect -18817 37122 -18807 37178
rect 2644 37207 2708 37217
rect 5429 37207 5493 37217
rect 6701 37207 6765 37217
rect 2644 37201 6765 37207
rect 2168 37145 2232 37159
rect -18883 37100 -18871 37122
rect -18819 37100 -18807 37122
rect -18883 37098 -18807 37100
rect -18883 37042 -18873 37098
rect -18817 37042 -18807 37098
rect 1473 37125 1537 37139
rect 1473 37069 1477 37125
rect 1533 37069 1537 37125
rect 1473 37055 1537 37069
rect 2168 37131 2174 37145
rect 2226 37131 2232 37145
rect 2644 37149 2650 37201
rect 2702 37149 5435 37201
rect 5487 37149 6707 37201
rect 6759 37149 6765 37201
rect 2644 37143 6765 37149
rect 2644 37133 2708 37143
rect 5429 37133 5493 37143
rect 6701 37133 6765 37143
rect 2168 37075 2172 37131
rect 2228 37075 2232 37131
rect -18883 37036 -18871 37042
rect -18819 37036 -18807 37042
rect -18883 37024 -18807 37036
rect -18883 37018 -18871 37024
rect -18819 37018 -18807 37024
rect -18883 36962 -18873 37018
rect -18817 36962 -18807 37018
rect -18883 36960 -18807 36962
rect -18883 36938 -18871 36960
rect -18819 36938 -18807 36960
rect -18883 36882 -18873 36938
rect -18817 36882 -18807 36938
rect 2168 37051 2174 37075
rect 2226 37051 2232 37075
rect 2168 36995 2172 37051
rect 2228 36995 2232 37051
rect 2168 36971 2174 36995
rect 2226 36971 2232 36995
rect 2168 36915 2172 36971
rect 2228 36915 2232 36971
rect 2168 36901 2174 36915
rect 2226 36901 2232 36915
rect 2168 36888 2232 36901
rect -18883 36858 -18871 36882
rect -18819 36858 -18807 36882
rect -18883 36802 -18873 36858
rect -18817 36802 -18807 36858
rect 93 36816 157 36826
rect 883 36816 947 36826
rect -18883 36780 -18871 36802
rect -18819 36780 -18807 36802
rect -18883 36778 -18807 36780
rect -18883 36722 -18873 36778
rect -18817 36722 -18807 36778
rect 90 36810 947 36816
rect 90 36758 99 36810
rect 151 36758 889 36810
rect 941 36758 947 36810
rect 90 36752 947 36758
rect 93 36742 157 36752
rect 883 36742 947 36752
rect -18883 36716 -18871 36722
rect -18819 36716 -18807 36722
rect -18883 36704 -18807 36716
rect -18883 36698 -18871 36704
rect -18819 36698 -18807 36704
rect -18883 36642 -18873 36698
rect -18817 36642 -18807 36698
rect -18883 36640 -18807 36642
rect -18883 36618 -18871 36640
rect -18819 36618 -18807 36640
rect -18883 36562 -18873 36618
rect -18817 36562 -18807 36618
rect -18883 36538 -18871 36562
rect -18819 36538 -18807 36562
rect -18883 36482 -18873 36538
rect -18817 36482 -18807 36538
rect -18883 36460 -18871 36482
rect -18819 36460 -18807 36482
rect -18883 36458 -18807 36460
rect -18883 36402 -18873 36458
rect -18817 36402 -18807 36458
rect -18883 36396 -18871 36402
rect -18819 36396 -18807 36402
rect -18883 36384 -18807 36396
rect -18883 36378 -18871 36384
rect -18819 36378 -18807 36384
rect -18883 36322 -18873 36378
rect -18817 36322 -18807 36378
rect 2169 36647 2233 36678
rect 2169 36591 2173 36647
rect 2229 36591 2233 36647
rect 6345 36593 6409 36607
rect 6345 36591 6349 36593
rect 2169 36581 2233 36591
rect 2169 36567 2175 36581
rect 2227 36567 2233 36581
rect 2169 36511 2173 36567
rect 2229 36511 2233 36567
rect 2169 36487 2175 36511
rect 2227 36487 2233 36511
rect 2169 36431 2173 36487
rect 2229 36431 2233 36487
rect 2169 36407 2175 36431
rect 2227 36407 2233 36431
rect 2169 36351 2173 36407
rect 2229 36351 2233 36407
rect 2169 36337 2175 36351
rect 2227 36337 2233 36351
rect -18883 36320 -18807 36322
rect -18883 36298 -18871 36320
rect -18819 36298 -18807 36320
rect -18883 36242 -18873 36298
rect -18817 36242 -18807 36298
rect 1996 36315 2060 36329
rect 1996 36259 2000 36315
rect 2056 36259 2060 36315
rect 1996 36245 2060 36259
rect 2169 36327 2233 36337
rect 2169 36271 2173 36327
rect 2229 36271 2233 36327
rect -18883 36218 -18871 36242
rect -18819 36218 -18807 36242
rect 2169 36240 2233 36271
rect 4938 36539 6349 36591
rect -27077 36142 -26996 36170
rect -27077 36120 -27063 36142
rect -27011 36120 -26996 36142
rect -27077 36064 -27065 36120
rect -27009 36064 -26996 36120
rect -18883 36162 -18873 36218
rect -18817 36162 -18807 36218
rect -18883 36140 -18871 36162
rect -18819 36140 -18807 36162
rect -18883 36114 -18807 36140
rect -27077 36040 -27063 36064
rect -27011 36040 -26996 36064
rect -27077 35984 -27065 36040
rect -27009 35984 -26996 36040
rect 2938 36087 3343 36098
rect 2938 36031 2952 36087
rect 3008 36085 3032 36087
rect 3088 36085 3112 36087
rect 3168 36085 3192 36087
rect 3248 36085 3272 36087
rect 3008 36033 3018 36085
rect 3262 36033 3272 36085
rect 3008 36031 3032 36033
rect 3088 36031 3112 36033
rect 3168 36031 3192 36033
rect 3248 36031 3272 36033
rect 3328 36031 3343 36087
rect 2938 36020 3343 36031
rect 3582 36090 3811 36104
rect 3582 36034 3588 36090
rect 3644 36088 3668 36090
rect 3724 36088 3748 36090
rect 3658 36036 3668 36088
rect 3724 36036 3734 36088
rect 3644 36034 3668 36036
rect 3724 36034 3748 36036
rect 3804 36034 3811 36090
rect 3582 36020 3811 36034
rect -27077 35962 -27063 35984
rect -27011 35962 -26996 35984
rect -27077 35960 -26996 35962
rect -27077 35904 -27065 35960
rect -27009 35904 -26996 35960
rect -27077 35898 -27063 35904
rect -27011 35898 -26996 35904
rect -27077 35886 -26996 35898
rect -27077 35880 -27063 35886
rect -27011 35880 -26996 35886
rect -27077 35824 -27065 35880
rect -27009 35824 -26996 35880
rect 4938 35863 4990 36539
rect 6345 36537 6349 36539
rect 6405 36591 6409 36593
rect 6405 36539 7804 36591
rect 6405 36537 6409 36539
rect 6345 36523 6409 36537
rect 6345 36249 6409 36263
rect 6345 36247 6349 36249
rect 5990 36195 6349 36247
rect 5055 36089 5351 36114
rect 5111 36087 5135 36089
rect 5191 36087 5215 36089
rect 5271 36087 5295 36089
rect 5133 36035 5135 36087
rect 5197 36035 5209 36087
rect 5271 36035 5273 36087
rect 5111 36033 5135 36035
rect 5191 36033 5215 36035
rect 5271 36033 5295 36035
rect 5055 36008 5351 36033
rect 5574 36090 5801 36107
rect 5574 36034 5579 36090
rect 5635 36088 5659 36090
rect 5715 36088 5739 36090
rect 5649 36036 5659 36088
rect 5715 36036 5725 36088
rect 5635 36034 5659 36036
rect 5715 36034 5739 36036
rect 5795 36034 5801 36090
rect 5574 36017 5801 36034
rect 5990 35969 6042 36195
rect 6345 36193 6349 36195
rect 6405 36247 6409 36249
rect 6405 36195 6740 36247
rect 6405 36193 6409 36195
rect 6345 36179 6409 36193
rect 5747 35917 6042 35969
rect 6688 35969 6740 36195
rect 6936 36082 7157 36099
rect 6936 36026 6938 36082
rect 6994 36080 7018 36082
rect 7074 36080 7098 36082
rect 7008 36028 7018 36080
rect 7074 36028 7084 36080
rect 6994 36026 7018 36028
rect 7074 36026 7098 36028
rect 7154 36026 7157 36082
rect 6936 36010 7157 36026
rect 7383 36089 7681 36104
rect 7383 36033 7384 36089
rect 7440 36087 7464 36089
rect 7520 36087 7544 36089
rect 7600 36087 7624 36089
rect 7462 36035 7464 36087
rect 7526 36035 7538 36087
rect 7600 36035 7602 36087
rect 7440 36033 7464 36035
rect 7520 36033 7544 36035
rect 7600 36033 7624 36035
rect 7680 36033 7681 36089
rect 7383 36018 7681 36033
rect 6688 35917 6989 35969
rect 7752 35941 7804 36539
rect 8921 36088 9348 36103
rect 8921 36032 8946 36088
rect 9002 36086 9026 36088
rect 9082 36086 9106 36088
rect 9162 36086 9186 36088
rect 9242 36086 9266 36088
rect 9002 36034 9012 36086
rect 9256 36034 9266 36086
rect 9002 36032 9026 36034
rect 9082 36032 9106 36034
rect 9162 36032 9186 36034
rect 9242 36032 9266 36034
rect 9322 36032 9348 36088
rect 8921 36018 9348 36032
rect 9575 36085 9802 36101
rect 9575 36029 9580 36085
rect 9636 36083 9660 36085
rect 9716 36083 9740 36085
rect 9650 36031 9660 36083
rect 9716 36031 9726 36083
rect 9636 36029 9660 36031
rect 9716 36029 9740 36031
rect 9796 36029 9802 36085
rect 9575 36013 9802 36029
rect -27077 35822 -26996 35824
rect -27077 35800 -27063 35822
rect -27011 35800 -26996 35822
rect -27077 35744 -27065 35800
rect -27009 35744 -26996 35800
rect -27077 35720 -27063 35744
rect -27011 35720 -26996 35744
rect -27077 35664 -27065 35720
rect -27009 35664 -26996 35720
rect -27077 35642 -27063 35664
rect -27011 35642 -26996 35664
rect -27077 35640 -26996 35642
rect -27077 35584 -27065 35640
rect -27009 35584 -26996 35640
rect -27077 35578 -27063 35584
rect -27011 35578 -26996 35584
rect -27077 35566 -26996 35578
rect -27077 35560 -27063 35566
rect -27011 35560 -26996 35566
rect -27077 35504 -27065 35560
rect -27009 35504 -26996 35560
rect -27077 35502 -26996 35504
rect -27077 35480 -27063 35502
rect -27011 35480 -26996 35502
rect -27077 35424 -27065 35480
rect -27009 35424 -26996 35480
rect -27077 35400 -27063 35424
rect -27011 35400 -26996 35424
rect -27077 35344 -27065 35400
rect -27009 35344 -26996 35400
rect -27077 35322 -27063 35344
rect -27011 35322 -26996 35344
rect -27077 35320 -26996 35322
rect -27077 35264 -27065 35320
rect -27009 35264 -26996 35320
rect -27077 35258 -27063 35264
rect -27011 35258 -26996 35264
rect -27077 35246 -26996 35258
rect -27077 35240 -27063 35246
rect -27011 35240 -26996 35246
rect -27077 35184 -27065 35240
rect -27009 35184 -26996 35240
rect -27077 35182 -26996 35184
rect -27077 35160 -27063 35182
rect -27011 35160 -26996 35182
rect -27077 35104 -27065 35160
rect -27009 35104 -26996 35160
rect -27077 35080 -27063 35104
rect -27011 35080 -26996 35104
rect -27077 35024 -27065 35080
rect -27009 35024 -26996 35080
rect -27077 35002 -27063 35024
rect -27011 35002 -26996 35024
rect -27077 34975 -26996 35002
rect 5430 35014 5494 35030
rect 5430 34962 5436 35014
rect 5488 34962 5494 35014
rect -27079 34682 -27000 34701
rect -27079 34626 -27068 34682
rect -27012 34626 -27000 34682
rect -27079 34612 -27066 34626
rect -27014 34612 -27000 34626
rect -27079 34602 -27000 34612
rect -9369 34672 -9305 34686
rect -9369 34616 -9365 34672
rect -9309 34616 -9305 34672
rect -9369 34602 -9305 34616
rect -27079 34546 -27068 34602
rect -27012 34546 -27000 34602
rect -27079 34536 -27000 34546
rect -27079 34522 -27066 34536
rect -27014 34522 -27000 34536
rect -27079 34466 -27068 34522
rect -27012 34466 -27000 34522
rect -27079 34442 -27066 34466
rect -27014 34442 -27000 34466
rect -27079 34386 -27068 34442
rect -27012 34386 -27000 34442
rect -27079 34362 -27066 34386
rect -27014 34362 -27000 34386
rect -27079 34306 -27068 34362
rect -27012 34306 -27000 34362
rect -27079 34292 -27066 34306
rect -27014 34292 -27000 34306
rect -27079 34282 -27000 34292
rect -27079 34226 -27068 34282
rect -27012 34226 -27000 34282
rect -27079 34216 -27000 34226
rect -27079 34202 -27066 34216
rect -27014 34202 -27000 34216
rect -27079 34146 -27068 34202
rect -27012 34146 -27000 34202
rect -27079 34122 -27066 34146
rect -27014 34122 -27000 34146
rect 2938 34183 2990 34704
rect 5430 34419 5494 34962
rect 5430 34367 5436 34419
rect 5488 34367 5494 34419
rect 5430 34351 5494 34367
rect 7242 35012 7306 35028
rect 7242 34960 7248 35012
rect 7300 34960 7306 35012
rect 7242 34419 7306 34960
rect 7242 34367 7248 34419
rect 7300 34367 7306 34419
rect 7242 34351 7306 34367
rect 5932 34191 5996 34205
rect 5932 34183 5936 34191
rect 2938 34135 5936 34183
rect 5992 34183 5996 34191
rect 8938 34183 8990 34790
rect 5992 34135 8990 34183
rect 2938 34131 8990 34135
rect -27079 34066 -27068 34122
rect -27012 34066 -27000 34122
rect 5932 34121 5996 34131
rect -27079 34042 -27066 34066
rect -27014 34042 -27000 34066
rect -27079 33986 -27068 34042
rect -27012 33986 -27000 34042
rect -27079 33972 -27066 33986
rect -27014 33972 -27000 33986
rect -27079 33962 -27000 33972
rect -27079 33906 -27068 33962
rect -27012 33906 -27000 33962
rect -27079 33896 -27000 33906
rect -27079 33882 -27066 33896
rect -27014 33882 -27000 33896
rect -27079 33826 -27068 33882
rect -27012 33826 -27000 33882
rect -27079 33802 -27066 33826
rect -27014 33802 -27000 33826
rect -27079 33746 -27068 33802
rect -27012 33746 -27000 33802
rect 3745 33850 3797 33860
rect 6738 33850 6802 33860
rect 9745 33850 9797 33860
rect 3797 33846 9745 33850
rect 3797 33798 6742 33846
rect 3745 33788 3797 33798
rect 6738 33790 6742 33798
rect 6798 33798 9745 33846
rect 9797 33798 9798 33850
rect 6798 33790 6802 33798
rect 6738 33776 6802 33790
rect 9745 33788 9797 33798
rect -27079 33722 -27066 33746
rect -27014 33722 -27000 33746
rect -27079 33666 -27068 33722
rect -27012 33666 -27000 33722
rect -27079 33652 -27066 33666
rect -27014 33652 -27000 33666
rect -27079 33642 -27000 33652
rect -27079 33586 -27068 33642
rect -27012 33586 -27000 33642
rect -27079 33576 -27000 33586
rect -27079 33562 -27066 33576
rect -27014 33562 -27000 33576
rect -27079 33506 -27068 33562
rect -27012 33506 -27000 33562
rect -27079 33488 -27000 33506
rect -21518 33547 -21454 33561
rect -21518 33491 -21514 33547
rect -21458 33491 -21454 33547
rect -21518 33477 -21454 33491
rect 5430 33555 5494 33574
rect 5430 33503 5436 33555
rect 5488 33503 5494 33555
rect -6948 33175 -6884 33189
rect -6948 33119 -6944 33175
rect -6888 33119 -6884 33175
rect -6948 33105 -6884 33119
rect -27084 32882 -27005 32909
rect -27084 32860 -27071 32882
rect -27019 32860 -27005 32882
rect -27084 32804 -27073 32860
rect -27017 32804 -27005 32860
rect -27084 32780 -27071 32804
rect -27019 32780 -27005 32804
rect -27084 32724 -27073 32780
rect -27017 32724 -27005 32780
rect -27084 32702 -27071 32724
rect -27019 32702 -27005 32724
rect -27084 32700 -27005 32702
rect -27084 32644 -27073 32700
rect -27017 32644 -27005 32700
rect -27084 32638 -27071 32644
rect -27019 32638 -27005 32644
rect -27084 32626 -27005 32638
rect -27084 32620 -27071 32626
rect -27019 32620 -27005 32626
rect -27084 32564 -27073 32620
rect -27017 32564 -27005 32620
rect -27084 32562 -27005 32564
rect -27084 32540 -27071 32562
rect -27019 32540 -27005 32562
rect -27084 32484 -27073 32540
rect -27017 32484 -27005 32540
rect -27084 32460 -27071 32484
rect -27019 32460 -27005 32484
rect -27084 32404 -27073 32460
rect -27017 32404 -27005 32460
rect -27084 32382 -27071 32404
rect -27019 32382 -27005 32404
rect -27084 32355 -27005 32382
rect 5317 32345 5381 32355
rect 5430 32345 5494 33503
rect 7428 33563 7492 33579
rect 7428 33511 7434 33563
rect 7486 33511 7492 33563
rect 7428 32362 7492 33511
rect 5317 32341 5494 32345
rect 5317 32285 5321 32341
rect 5377 32285 5494 32341
rect 5317 32281 5494 32285
rect 7364 32348 7492 32362
rect 7364 32292 7368 32348
rect 7424 32292 7492 32348
rect 7364 32288 7492 32292
rect 5317 32271 5381 32281
rect 7364 32278 7428 32288
rect -6989 31807 8057 31840
rect -6989 31805 7969 31807
rect -6989 31753 -6983 31805
rect -6931 31753 -6919 31805
rect -6867 31753 7969 31805
rect -6989 31751 7969 31753
rect 8025 31751 8057 31807
rect -6989 31712 8057 31751
rect 4354 30428 4418 30442
rect 4354 30372 4358 30428
rect 4414 30372 4418 30428
rect 4354 30358 4418 30372
rect 8328 30433 8392 30447
rect 8328 30377 8332 30433
rect 8388 30377 8392 30433
rect 8328 30363 8392 30377
rect -9347 30315 2453 30338
rect -9397 30305 2453 30315
rect 3326 30305 3390 30315
rect -9397 30301 3390 30305
rect -9397 30299 3330 30301
rect -9397 30247 -9391 30299
rect -9339 30247 -9327 30299
rect -9275 30247 3330 30299
rect -9397 30245 3330 30247
rect 3386 30245 3390 30301
rect -9397 30241 3390 30245
rect -9397 30231 2453 30241
rect 3326 30231 3390 30241
rect -9347 30210 2453 30231
rect -12693 29748 -12629 29762
rect -12693 29692 -12689 29748
rect -12633 29692 -12629 29748
rect -12693 29678 -12629 29692
rect 1913 29752 1977 29762
rect 16721 29752 16785 29762
rect 1913 29748 16785 29752
rect 1913 29692 1917 29748
rect 1973 29692 16725 29748
rect 16781 29692 16785 29748
rect 1913 29688 16785 29692
rect 1913 29678 1977 29688
rect 16721 29678 16785 29688
rect -13469 29325 -13405 29339
rect -30199 29165 -30193 29281
rect -30077 29165 -30070 29281
rect -30199 29149 -30070 29165
rect -18523 29281 -18394 29298
rect -18523 29165 -18517 29281
rect -18401 29165 -18394 29281
rect -13469 29269 -13465 29325
rect -13409 29269 -13405 29325
rect -13469 29255 -13405 29269
rect 1913 29329 1977 29339
rect 17412 29329 17476 29339
rect 1913 29325 17476 29329
rect 1913 29269 1917 29325
rect 1973 29269 17416 29325
rect 17472 29269 17476 29325
rect 1913 29265 17476 29269
rect 1913 29255 1977 29265
rect 17412 29255 17476 29265
rect -31030 27807 -31024 27923
rect -30908 27807 -30901 27923
rect -31030 27791 -30901 27807
rect -19383 27923 -19254 27940
rect -19383 27807 -19377 27923
rect -19261 27807 -19254 27923
rect -38190 26590 -34856 26621
rect -38190 26588 -38151 26590
rect -38095 26588 -38071 26590
rect -38015 26588 -37991 26590
rect -37935 26588 -37911 26590
rect -37855 26588 -37831 26590
rect -37775 26588 -37751 26590
rect -37695 26588 -37671 26590
rect -37615 26588 -37591 26590
rect -37535 26588 -37511 26590
rect -37455 26588 -37431 26590
rect -37375 26588 -37351 26590
rect -37295 26588 -37271 26590
rect -37215 26588 -37191 26590
rect -37135 26588 -37111 26590
rect -37055 26588 -37031 26590
rect -36975 26588 -36951 26590
rect -36895 26588 -36871 26590
rect -36815 26588 -36791 26590
rect -36735 26588 -36711 26590
rect -36655 26588 -36631 26590
rect -36575 26588 -36551 26590
rect -36495 26588 -36471 26590
rect -36415 26588 -36391 26590
rect -36335 26588 -36311 26590
rect -36255 26588 -36231 26590
rect -36175 26588 -36151 26590
rect -36095 26588 -36071 26590
rect -36015 26588 -35991 26590
rect -35935 26588 -35911 26590
rect -35855 26588 -35831 26590
rect -35775 26588 -35751 26590
rect -35695 26588 -35671 26590
rect -35615 26588 -35591 26590
rect -35535 26588 -35511 26590
rect -35455 26588 -35431 26590
rect -35375 26588 -35351 26590
rect -35295 26588 -35271 26590
rect -35215 26588 -35191 26590
rect -35135 26588 -35111 26590
rect -35055 26588 -35031 26590
rect -34975 26588 -34951 26590
rect -34895 26588 -34856 26590
rect -38190 26536 -38181 26588
rect -38001 26536 -37991 26588
rect -37935 26536 -37925 26588
rect -37681 26536 -37671 26588
rect -37615 26536 -37605 26588
rect -37361 26536 -37351 26588
rect -37295 26536 -37285 26588
rect -37041 26536 -37031 26588
rect -36975 26536 -36965 26588
rect -36721 26536 -36711 26588
rect -36655 26536 -36645 26588
rect -36401 26536 -36391 26588
rect -36335 26536 -36325 26588
rect -36081 26536 -36071 26588
rect -36015 26536 -36005 26588
rect -35761 26536 -35751 26588
rect -35695 26536 -35685 26588
rect -35441 26536 -35431 26588
rect -35375 26536 -35365 26588
rect -35121 26536 -35111 26588
rect -35055 26536 -35045 26588
rect -34865 26536 -34856 26588
rect -38190 26534 -38151 26536
rect -38095 26534 -38071 26536
rect -38015 26534 -37991 26536
rect -37935 26534 -37911 26536
rect -37855 26534 -37831 26536
rect -37775 26534 -37751 26536
rect -37695 26534 -37671 26536
rect -37615 26534 -37591 26536
rect -37535 26534 -37511 26536
rect -37455 26534 -37431 26536
rect -37375 26534 -37351 26536
rect -37295 26534 -37271 26536
rect -37215 26534 -37191 26536
rect -37135 26534 -37111 26536
rect -37055 26534 -37031 26536
rect -36975 26534 -36951 26536
rect -36895 26534 -36871 26536
rect -36815 26534 -36791 26536
rect -36735 26534 -36711 26536
rect -36655 26534 -36631 26536
rect -36575 26534 -36551 26536
rect -36495 26534 -36471 26536
rect -36415 26534 -36391 26536
rect -36335 26534 -36311 26536
rect -36255 26534 -36231 26536
rect -36175 26534 -36151 26536
rect -36095 26534 -36071 26536
rect -36015 26534 -35991 26536
rect -35935 26534 -35911 26536
rect -35855 26534 -35831 26536
rect -35775 26534 -35751 26536
rect -35695 26534 -35671 26536
rect -35615 26534 -35591 26536
rect -35535 26534 -35511 26536
rect -35455 26534 -35431 26536
rect -35375 26534 -35351 26536
rect -35295 26534 -35271 26536
rect -35215 26534 -35191 26536
rect -35135 26534 -35111 26536
rect -35055 26534 -35031 26536
rect -34975 26534 -34951 26536
rect -34895 26534 -34856 26536
rect -38190 26504 -34856 26534
rect -19383 26015 -19254 27807
rect -18523 27609 -18394 29165
rect 7960 28842 8024 28856
rect 1951 28808 2079 28818
rect 4701 28808 4765 28818
rect 1951 28804 4765 28808
rect 1951 28802 4705 28804
rect 1951 28750 1957 28802
rect 2009 28750 2021 28802
rect 2073 28750 4705 28802
rect 1951 28748 4705 28750
rect 4761 28748 4765 28804
rect 7960 28786 7964 28842
rect 8020 28786 8024 28842
rect 7960 28772 8024 28786
rect 1951 28744 4765 28748
rect 1951 28734 2079 28744
rect 4701 28734 4765 28744
rect -6086 28602 -5958 28633
rect -6086 28550 -6080 28602
rect -6028 28550 -6016 28602
rect -5964 28550 -5958 28602
rect -15712 28089 -15613 28108
rect -15712 28059 -15689 28089
rect -15637 28059 -15613 28089
rect -15712 28003 -15691 28059
rect -15635 28003 -15613 28059
rect -15712 27979 -15689 28003
rect -15637 27979 -15613 28003
rect -15712 27923 -15691 27979
rect -15635 27923 -15613 27979
rect -15712 27909 -15689 27923
rect -15637 27909 -15613 27923
rect -15712 27899 -15613 27909
rect -15712 27843 -15691 27899
rect -15635 27843 -15613 27899
rect -15712 27833 -15613 27843
rect -15712 27819 -15689 27833
rect -15637 27819 -15613 27833
rect -15712 27763 -15691 27819
rect -15635 27763 -15613 27819
rect -15712 27739 -15689 27763
rect -15637 27739 -15613 27763
rect -15712 27683 -15691 27739
rect -15635 27683 -15613 27739
rect -17635 27638 -17507 27654
rect -18523 27569 -18246 27609
rect -18523 27517 -18320 27569
rect -18268 27517 -18246 27569
rect -18523 27480 -18246 27517
rect -17635 27522 -17629 27638
rect -17513 27522 -17507 27638
rect -15712 27653 -15689 27683
rect -15637 27653 -15613 27683
rect -15712 27635 -15613 27653
rect -13983 28066 -13931 28076
rect -17635 27506 -17507 27522
rect -14906 27571 -14854 27581
rect -18326 27098 -18262 27108
rect -18326 27092 -17257 27098
rect -18326 27040 -18320 27092
rect -18268 27040 -17257 27092
rect -18326 27034 -17257 27040
rect -14906 27083 -14854 27519
rect -18326 27024 -18262 27034
rect -18881 26760 -18817 26770
rect -17256 26760 -17192 26770
rect -18881 26754 -17192 26760
rect -18881 26702 -18875 26754
rect -18823 26702 -17250 26754
rect -17198 26702 -17192 26754
rect -18881 26696 -17192 26702
rect -18881 26686 -18817 26696
rect -17256 26686 -17192 26696
rect -17635 26409 -17507 26425
rect -17635 26293 -17629 26409
rect -17513 26293 -17507 26409
rect -17635 26277 -17507 26293
rect -15725 26270 -15636 26291
rect -15725 26214 -15709 26270
rect -15653 26214 -15636 26270
rect -15725 26200 -15707 26214
rect -15655 26200 -15636 26214
rect -15725 26190 -15636 26200
rect -15725 26134 -15709 26190
rect -15653 26134 -15636 26190
rect -15725 26124 -15636 26134
rect -15725 26110 -15707 26124
rect -15655 26110 -15636 26124
rect -15725 26054 -15709 26110
rect -15653 26054 -15636 26110
rect -15725 26034 -15636 26054
rect -19383 25971 -18816 26015
rect -19383 25919 -18876 25971
rect -18824 25919 -18816 25971
rect -19383 25886 -18816 25919
rect -14906 25967 -14854 27031
rect -14906 25905 -14854 25915
rect -14404 27259 -14352 27269
rect -14404 25659 -14352 27207
rect -13983 26466 -13931 28014
rect -12389 28061 -12316 28086
rect -12389 28005 -12381 28061
rect -12325 28005 -12316 28061
rect -12389 27995 -12316 28005
rect -12389 27981 -12379 27995
rect -12327 27981 -12316 27995
rect -12389 27925 -12381 27981
rect -12325 27925 -12316 27981
rect -12389 27901 -12379 27925
rect -12327 27901 -12316 27925
rect -12389 27845 -12381 27901
rect -12325 27845 -12316 27901
rect -12389 27821 -12379 27845
rect -12327 27821 -12316 27845
rect -12389 27765 -12381 27821
rect -12325 27765 -12316 27821
rect -12389 27751 -12379 27765
rect -12327 27751 -12316 27765
rect -12389 27741 -12316 27751
rect -12389 27685 -12381 27741
rect -12325 27685 -12316 27741
rect -12389 27660 -12316 27685
rect -12394 27420 -12297 27437
rect -12394 27364 -12374 27420
rect -12318 27364 -12297 27420
rect -12394 27350 -12372 27364
rect -12320 27350 -12297 27364
rect -12394 27340 -12297 27350
rect -12394 27284 -12374 27340
rect -12318 27284 -12297 27340
rect -12394 27274 -12297 27284
rect -12394 27260 -12372 27274
rect -12320 27260 -12297 27274
rect -12394 27204 -12374 27260
rect -12318 27204 -12297 27260
rect -12394 27188 -12297 27204
rect -10016 26582 -9888 26598
rect -10016 26530 -10010 26582
rect -9958 26530 -9946 26582
rect -9894 26530 -9888 26582
rect -13983 25674 -13931 26414
rect -12396 26459 -12301 26496
rect -12396 26403 -12377 26459
rect -12321 26403 -12301 26459
rect -12396 26393 -12301 26403
rect -12396 26379 -12375 26393
rect -12323 26379 -12301 26393
rect -12396 26323 -12377 26379
rect -12321 26323 -12301 26379
rect -12396 26299 -12375 26323
rect -12323 26299 -12301 26323
rect -12396 26243 -12377 26299
rect -12321 26243 -12301 26299
rect -12396 26219 -12375 26243
rect -12323 26219 -12301 26243
rect -12396 26163 -12377 26219
rect -12321 26163 -12301 26219
rect -12396 26149 -12375 26163
rect -12323 26149 -12301 26163
rect -12396 26139 -12301 26149
rect -12396 26083 -12377 26139
rect -12321 26083 -12301 26139
rect -12396 26047 -12301 26083
rect -12384 25821 -12321 25833
rect -12384 25765 -12381 25821
rect -12325 25765 -12321 25821
rect -12384 25751 -12379 25765
rect -12327 25751 -12321 25765
rect -12384 25741 -12321 25751
rect -12384 25685 -12381 25741
rect -12325 25685 -12321 25741
rect -12384 25675 -12321 25685
rect -25551 25527 -24848 25579
rect -25449 25476 -25369 25492
rect -25449 25420 -25437 25476
rect -25381 25420 -25369 25476
rect -25449 25398 -25435 25420
rect -25383 25398 -25369 25420
rect -25449 25396 -25369 25398
rect -25449 25340 -25437 25396
rect -25381 25340 -25369 25396
rect -25449 25334 -25435 25340
rect -25383 25334 -25369 25340
rect -25449 25322 -25369 25334
rect -25449 25316 -25435 25322
rect -25383 25316 -25369 25322
rect -25449 25260 -25437 25316
rect -25381 25260 -25369 25316
rect -25449 25258 -25369 25260
rect -25449 25236 -25435 25258
rect -25383 25236 -25369 25258
rect -40593 25161 -40357 25181
rect -25449 25180 -25437 25236
rect -25381 25180 -25369 25236
rect -25449 25165 -25369 25180
rect -40593 24945 -40583 25161
rect -40367 24945 -40357 25161
rect -40593 24925 -40357 24945
rect -32991 25106 -32863 25122
rect -32991 24990 -32985 25106
rect -32869 24990 -32863 25106
rect -38182 23582 -34852 23615
rect -38182 23580 -38145 23582
rect -38089 23580 -38065 23582
rect -38009 23580 -37985 23582
rect -37929 23580 -37905 23582
rect -37849 23580 -37825 23582
rect -37769 23580 -37745 23582
rect -37689 23580 -37665 23582
rect -37609 23580 -37585 23582
rect -37529 23580 -37505 23582
rect -37449 23580 -37425 23582
rect -37369 23580 -37345 23582
rect -37289 23580 -37265 23582
rect -37209 23580 -37185 23582
rect -37129 23580 -37105 23582
rect -37049 23580 -37025 23582
rect -36969 23580 -36945 23582
rect -36889 23580 -36865 23582
rect -36809 23580 -36785 23582
rect -36729 23580 -36705 23582
rect -36649 23580 -36625 23582
rect -36569 23580 -36545 23582
rect -36489 23580 -36465 23582
rect -36409 23580 -36385 23582
rect -36329 23580 -36305 23582
rect -36249 23580 -36225 23582
rect -36169 23580 -36145 23582
rect -36089 23580 -36065 23582
rect -36009 23580 -35985 23582
rect -35929 23580 -35905 23582
rect -35849 23580 -35825 23582
rect -35769 23580 -35745 23582
rect -35689 23580 -35665 23582
rect -35609 23580 -35585 23582
rect -35529 23580 -35505 23582
rect -35449 23580 -35425 23582
rect -35369 23580 -35345 23582
rect -35289 23580 -35265 23582
rect -35209 23580 -35185 23582
rect -35129 23580 -35105 23582
rect -35049 23580 -35025 23582
rect -34969 23580 -34945 23582
rect -34889 23580 -34852 23582
rect -38182 23528 -38175 23580
rect -37995 23528 -37985 23580
rect -37929 23528 -37919 23580
rect -37675 23528 -37665 23580
rect -37609 23528 -37599 23580
rect -37355 23528 -37345 23580
rect -37289 23528 -37279 23580
rect -37035 23528 -37025 23580
rect -36969 23528 -36959 23580
rect -36715 23528 -36705 23580
rect -36649 23528 -36639 23580
rect -36395 23528 -36385 23580
rect -36329 23528 -36319 23580
rect -36075 23528 -36065 23580
rect -36009 23528 -35999 23580
rect -35755 23528 -35745 23580
rect -35689 23528 -35679 23580
rect -35435 23528 -35425 23580
rect -35369 23528 -35359 23580
rect -35115 23528 -35105 23580
rect -35049 23528 -35039 23580
rect -34859 23528 -34852 23580
rect -38182 23526 -38145 23528
rect -38089 23526 -38065 23528
rect -38009 23526 -37985 23528
rect -37929 23526 -37905 23528
rect -37849 23526 -37825 23528
rect -37769 23526 -37745 23528
rect -37689 23526 -37665 23528
rect -37609 23526 -37585 23528
rect -37529 23526 -37505 23528
rect -37449 23526 -37425 23528
rect -37369 23526 -37345 23528
rect -37289 23526 -37265 23528
rect -37209 23526 -37185 23528
rect -37129 23526 -37105 23528
rect -37049 23526 -37025 23528
rect -36969 23526 -36945 23528
rect -36889 23526 -36865 23528
rect -36809 23526 -36785 23528
rect -36729 23526 -36705 23528
rect -36649 23526 -36625 23528
rect -36569 23526 -36545 23528
rect -36489 23526 -36465 23528
rect -36409 23526 -36385 23528
rect -36329 23526 -36305 23528
rect -36249 23526 -36225 23528
rect -36169 23526 -36145 23528
rect -36089 23526 -36065 23528
rect -36009 23526 -35985 23528
rect -35929 23526 -35905 23528
rect -35849 23526 -35825 23528
rect -35769 23526 -35745 23528
rect -35689 23526 -35665 23528
rect -35609 23526 -35585 23528
rect -35529 23526 -35505 23528
rect -35449 23526 -35425 23528
rect -35369 23526 -35345 23528
rect -35289 23526 -35265 23528
rect -35209 23526 -35185 23528
rect -35129 23526 -35105 23528
rect -35049 23526 -35025 23528
rect -34969 23526 -34945 23528
rect -34889 23526 -34852 23528
rect -38182 23493 -34852 23526
rect -38168 19054 -34861 19075
rect -38168 18998 -38143 19054
rect -38087 19052 -38063 19054
rect -38007 19052 -37983 19054
rect -37927 19052 -37903 19054
rect -37847 19052 -37823 19054
rect -37767 19052 -37743 19054
rect -37687 19052 -37663 19054
rect -37607 19052 -37583 19054
rect -37527 19052 -37503 19054
rect -37447 19052 -37423 19054
rect -37367 19052 -37343 19054
rect -37287 19052 -37263 19054
rect -37207 19052 -37183 19054
rect -37127 19052 -37103 19054
rect -37047 19052 -37023 19054
rect -36967 19052 -36943 19054
rect -36887 19052 -36863 19054
rect -36807 19052 -36783 19054
rect -36727 19052 -36703 19054
rect -36647 19052 -36623 19054
rect -36567 19052 -36543 19054
rect -36487 19052 -36463 19054
rect -36407 19052 -36383 19054
rect -36327 19052 -36303 19054
rect -36247 19052 -36223 19054
rect -36167 19052 -36143 19054
rect -36087 19052 -36063 19054
rect -36007 19052 -35983 19054
rect -35927 19052 -35903 19054
rect -35847 19052 -35823 19054
rect -35767 19052 -35743 19054
rect -35687 19052 -35663 19054
rect -35607 19052 -35583 19054
rect -35527 19052 -35503 19054
rect -35447 19052 -35423 19054
rect -35367 19052 -35343 19054
rect -35287 19052 -35263 19054
rect -35207 19052 -35183 19054
rect -35127 19052 -35103 19054
rect -35047 19052 -35023 19054
rect -34967 19052 -34943 19054
rect -38087 19000 -38077 19052
rect -37833 19000 -37823 19052
rect -37767 19000 -37757 19052
rect -37513 19000 -37503 19052
rect -37447 19000 -37437 19052
rect -37193 19000 -37183 19052
rect -37127 19000 -37117 19052
rect -36873 19000 -36863 19052
rect -36807 19000 -36797 19052
rect -36553 19000 -36543 19052
rect -36487 19000 -36477 19052
rect -36233 19000 -36223 19052
rect -36167 19000 -36157 19052
rect -35913 19000 -35903 19052
rect -35847 19000 -35837 19052
rect -35593 19000 -35583 19052
rect -35527 19000 -35517 19052
rect -35273 19000 -35263 19052
rect -35207 19000 -35197 19052
rect -34953 19000 -34943 19052
rect -38087 18998 -38063 19000
rect -38007 18998 -37983 19000
rect -37927 18998 -37903 19000
rect -37847 18998 -37823 19000
rect -37767 18998 -37743 19000
rect -37687 18998 -37663 19000
rect -37607 18998 -37583 19000
rect -37527 18998 -37503 19000
rect -37447 18998 -37423 19000
rect -37367 18998 -37343 19000
rect -37287 18998 -37263 19000
rect -37207 18998 -37183 19000
rect -37127 18998 -37103 19000
rect -37047 18998 -37023 19000
rect -36967 18998 -36943 19000
rect -36887 18998 -36863 19000
rect -36807 18998 -36783 19000
rect -36727 18998 -36703 19000
rect -36647 18998 -36623 19000
rect -36567 18998 -36543 19000
rect -36487 18998 -36463 19000
rect -36407 18998 -36383 19000
rect -36327 18998 -36303 19000
rect -36247 18998 -36223 19000
rect -36167 18998 -36143 19000
rect -36087 18998 -36063 19000
rect -36007 18998 -35983 19000
rect -35927 18998 -35903 19000
rect -35847 18998 -35823 19000
rect -35767 18998 -35743 19000
rect -35687 18998 -35663 19000
rect -35607 18998 -35583 19000
rect -35527 18998 -35503 19000
rect -35447 18998 -35423 19000
rect -35367 18998 -35343 19000
rect -35287 18998 -35263 19000
rect -35207 18998 -35183 19000
rect -35127 18998 -35103 19000
rect -35047 18998 -35023 19000
rect -34967 18998 -34943 19000
rect -34887 18998 -34861 19054
rect -38168 18977 -34861 18998
rect -40596 17620 -40360 17640
rect -40596 17404 -40586 17620
rect -40370 17404 -40360 17620
rect -40596 17384 -40360 17404
rect -38174 16059 -34852 16085
rect -38174 16057 -38141 16059
rect -38085 16057 -38061 16059
rect -38005 16057 -37981 16059
rect -37925 16057 -37901 16059
rect -37845 16057 -37821 16059
rect -37765 16057 -37741 16059
rect -37685 16057 -37661 16059
rect -37605 16057 -37581 16059
rect -37525 16057 -37501 16059
rect -37445 16057 -37421 16059
rect -37365 16057 -37341 16059
rect -37285 16057 -37261 16059
rect -37205 16057 -37181 16059
rect -37125 16057 -37101 16059
rect -37045 16057 -37021 16059
rect -36965 16057 -36941 16059
rect -36885 16057 -36861 16059
rect -36805 16057 -36781 16059
rect -36725 16057 -36701 16059
rect -36645 16057 -36621 16059
rect -36565 16057 -36541 16059
rect -36485 16057 -36461 16059
rect -36405 16057 -36381 16059
rect -36325 16057 -36301 16059
rect -36245 16057 -36221 16059
rect -36165 16057 -36141 16059
rect -36085 16057 -36061 16059
rect -36005 16057 -35981 16059
rect -35925 16057 -35901 16059
rect -35845 16057 -35821 16059
rect -35765 16057 -35741 16059
rect -35685 16057 -35661 16059
rect -35605 16057 -35581 16059
rect -35525 16057 -35501 16059
rect -35445 16057 -35421 16059
rect -35365 16057 -35341 16059
rect -35285 16057 -35261 16059
rect -35205 16057 -35181 16059
rect -35125 16057 -35101 16059
rect -35045 16057 -35021 16059
rect -34965 16057 -34941 16059
rect -34885 16057 -34852 16059
rect -38174 16005 -38171 16057
rect -37991 16005 -37981 16057
rect -37925 16005 -37915 16057
rect -37671 16005 -37661 16057
rect -37605 16005 -37595 16057
rect -37351 16005 -37341 16057
rect -37285 16005 -37275 16057
rect -37031 16005 -37021 16057
rect -36965 16005 -36955 16057
rect -36711 16005 -36701 16057
rect -36645 16005 -36635 16057
rect -36391 16005 -36381 16057
rect -36325 16005 -36315 16057
rect -36071 16005 -36061 16057
rect -36005 16005 -35995 16057
rect -35751 16005 -35741 16057
rect -35685 16005 -35675 16057
rect -35431 16005 -35421 16057
rect -35365 16005 -35355 16057
rect -35111 16005 -35101 16057
rect -35045 16005 -35035 16057
rect -34855 16005 -34852 16057
rect -38174 16003 -38141 16005
rect -38085 16003 -38061 16005
rect -38005 16003 -37981 16005
rect -37925 16003 -37901 16005
rect -37845 16003 -37821 16005
rect -37765 16003 -37741 16005
rect -37685 16003 -37661 16005
rect -37605 16003 -37581 16005
rect -37525 16003 -37501 16005
rect -37445 16003 -37421 16005
rect -37365 16003 -37341 16005
rect -37285 16003 -37261 16005
rect -37205 16003 -37181 16005
rect -37125 16003 -37101 16005
rect -37045 16003 -37021 16005
rect -36965 16003 -36941 16005
rect -36885 16003 -36861 16005
rect -36805 16003 -36781 16005
rect -36725 16003 -36701 16005
rect -36645 16003 -36621 16005
rect -36565 16003 -36541 16005
rect -36485 16003 -36461 16005
rect -36405 16003 -36381 16005
rect -36325 16003 -36301 16005
rect -36245 16003 -36221 16005
rect -36165 16003 -36141 16005
rect -36085 16003 -36061 16005
rect -36005 16003 -35981 16005
rect -35925 16003 -35901 16005
rect -35845 16003 -35821 16005
rect -35765 16003 -35741 16005
rect -35685 16003 -35661 16005
rect -35605 16003 -35581 16005
rect -35525 16003 -35501 16005
rect -35445 16003 -35421 16005
rect -35365 16003 -35341 16005
rect -35285 16003 -35261 16005
rect -35205 16003 -35181 16005
rect -35125 16003 -35101 16005
rect -35045 16003 -35021 16005
rect -34965 16003 -34941 16005
rect -34885 16003 -34852 16005
rect -38174 15977 -34852 16003
rect -32991 14096 -32863 24990
rect -25452 24937 -25365 24955
rect -25452 24881 -25437 24937
rect -25381 24881 -25365 24937
rect -25452 24867 -25435 24881
rect -25383 24867 -25365 24881
rect -25452 24857 -25365 24867
rect -25452 24801 -25437 24857
rect -25381 24801 -25365 24857
rect -25452 24791 -25365 24801
rect -25452 24777 -25435 24791
rect -25383 24777 -25365 24791
rect -27178 24719 -26676 24771
rect -25452 24721 -25437 24777
rect -25381 24721 -25365 24777
rect -27178 21000 -27126 24719
rect -25452 24704 -25365 24721
rect -27939 20948 -27126 21000
rect -32991 13980 -32985 14096
rect -32869 13980 -32863 14096
rect -32991 13964 -32863 13980
rect -31130 17576 -31002 17592
rect -31130 17460 -31124 17576
rect -31008 17460 -31002 17576
rect -31130 6331 -31002 17460
rect -27939 15451 -27887 20948
rect -27178 17229 -27126 20948
rect -24900 21808 -24848 25527
rect -15727 25420 -15632 25457
rect -15727 25364 -15708 25420
rect -15652 25364 -15632 25420
rect -15727 25354 -15632 25364
rect -15727 25340 -15706 25354
rect -15654 25340 -15632 25354
rect -15727 25284 -15708 25340
rect -15652 25284 -15632 25340
rect -15727 25260 -15706 25284
rect -15654 25260 -15632 25284
rect -15727 25204 -15708 25260
rect -15652 25204 -15632 25260
rect -15727 25180 -15706 25204
rect -15654 25180 -15632 25204
rect -15727 25124 -15708 25180
rect -15652 25124 -15632 25180
rect -15727 25110 -15706 25124
rect -15654 25110 -15632 25124
rect -15727 25100 -15632 25110
rect -15727 25044 -15708 25100
rect -15652 25044 -15632 25100
rect -17635 24996 -17507 25012
rect -15727 25008 -15632 25044
rect -17635 24880 -17629 24996
rect -17513 24880 -17507 24996
rect -14404 24882 -14352 25607
rect -13989 25660 -13925 25674
rect -13989 25604 -13985 25660
rect -13929 25604 -13925 25660
rect -13989 25590 -13925 25604
rect -12384 25661 -12379 25675
rect -12327 25661 -12321 25675
rect -12384 25605 -12381 25661
rect -12325 25605 -12321 25661
rect -12384 25594 -12321 25605
rect -17635 24864 -17507 24880
rect -14410 24868 -14346 24882
rect -14410 24812 -14406 24868
rect -14350 24812 -14346 24868
rect -14410 24798 -14346 24812
rect -13983 24866 -13931 25590
rect -18326 24458 -18262 24467
rect -18326 24451 -17271 24458
rect -18326 24399 -18320 24451
rect -18268 24399 -17271 24451
rect -18326 24394 -17271 24399
rect -14908 24441 -14856 24451
rect -18326 24383 -18262 24394
rect -18881 24118 -18817 24128
rect -17263 24118 -17199 24128
rect -18881 24112 -17199 24118
rect -18881 24060 -18875 24112
rect -18823 24060 -17257 24112
rect -17205 24060 -17199 24112
rect -18881 24054 -17199 24060
rect -18881 24044 -18817 24054
rect -17263 24044 -17199 24054
rect -17635 23767 -17507 23783
rect -17635 23651 -17629 23767
rect -17513 23651 -17507 23767
rect -17635 23635 -17507 23651
rect -15725 23629 -15658 23647
rect -15725 23573 -15720 23629
rect -15664 23573 -15658 23629
rect -15725 23559 -15718 23573
rect -15666 23559 -15658 23573
rect -15725 23549 -15658 23559
rect -15725 23493 -15720 23549
rect -15664 23493 -15658 23549
rect -15725 23483 -15658 23493
rect -15725 23469 -15718 23483
rect -15666 23469 -15658 23483
rect -15725 23413 -15720 23469
rect -15664 23413 -15658 23469
rect -15725 23395 -15658 23413
rect -14908 22771 -14856 24389
rect -14908 22713 -14856 22719
rect -14404 24059 -14352 24798
rect -14404 22459 -14352 24007
rect -13983 23266 -13931 24814
rect -12393 24707 -12328 24722
rect -12393 24693 -12387 24707
rect -12335 24693 -12328 24707
rect -12393 24637 -12389 24693
rect -12333 24637 -12328 24693
rect -12393 24613 -12387 24637
rect -12335 24613 -12328 24637
rect -12393 24557 -12389 24613
rect -12333 24557 -12328 24613
rect -12393 24533 -12387 24557
rect -12335 24533 -12328 24557
rect -12393 24477 -12389 24533
rect -12333 24477 -12328 24533
rect -12393 24463 -12387 24477
rect -12335 24463 -12328 24477
rect -12393 24448 -12328 24463
rect -12398 24229 -12316 24249
rect -12398 24173 -12385 24229
rect -12329 24173 -12316 24229
rect -12398 24159 -12383 24173
rect -12331 24159 -12316 24173
rect -12398 24149 -12316 24159
rect -12398 24093 -12385 24149
rect -12329 24093 -12316 24149
rect -12398 24083 -12316 24093
rect -12398 24069 -12383 24083
rect -12331 24069 -12316 24083
rect -12398 24013 -12385 24069
rect -12329 24013 -12316 24069
rect -12398 23993 -12316 24013
rect -13983 23203 -13931 23214
rect -12389 23255 -12319 23287
rect -12389 23199 -12382 23255
rect -12326 23199 -12319 23255
rect -12389 23189 -12319 23199
rect -12389 23175 -12380 23189
rect -12328 23175 -12319 23189
rect -12389 23119 -12382 23175
rect -12326 23119 -12319 23175
rect -12389 23095 -12380 23119
rect -12328 23095 -12319 23119
rect -12389 23039 -12382 23095
rect -12326 23039 -12319 23095
rect -12389 23015 -12380 23039
rect -12328 23015 -12319 23039
rect -12389 22959 -12382 23015
rect -12326 22959 -12319 23015
rect -12389 22945 -12380 22959
rect -12328 22945 -12319 22959
rect -12389 22935 -12319 22945
rect -12389 22879 -12382 22935
rect -12326 22879 -12319 22935
rect -12389 22847 -12319 22879
rect -11601 22770 -11473 22786
rect -11601 22718 -11595 22770
rect -11543 22718 -11531 22770
rect -11479 22718 -11473 22770
rect -14404 22397 -14352 22407
rect -12391 22619 -12323 22634
rect -12391 22563 -12385 22619
rect -12329 22563 -12323 22619
rect -12391 22549 -12383 22563
rect -12331 22549 -12323 22563
rect -12391 22539 -12323 22549
rect -12391 22483 -12385 22539
rect -12329 22483 -12323 22539
rect -12391 22473 -12323 22483
rect -12391 22459 -12383 22473
rect -12331 22459 -12323 22473
rect -12391 22403 -12385 22459
rect -12329 22403 -12323 22459
rect -12391 22389 -12323 22403
rect -11601 21851 -11473 22718
rect -24900 21756 -24087 21808
rect -24900 18038 -24848 21756
rect -25557 17986 -24848 18038
rect -25452 17896 -25387 17932
rect -25452 17882 -25446 17896
rect -25394 17882 -25387 17896
rect -25452 17826 -25448 17882
rect -25392 17826 -25387 17882
rect -25452 17802 -25446 17826
rect -25394 17802 -25387 17826
rect -25452 17746 -25448 17802
rect -25392 17746 -25387 17802
rect -25452 17722 -25446 17746
rect -25394 17722 -25387 17746
rect -25452 17666 -25448 17722
rect -25392 17666 -25387 17722
rect -25452 17652 -25446 17666
rect -25394 17652 -25387 17666
rect -25452 17617 -25387 17652
rect -25450 17394 -25378 17414
rect -25450 17338 -25442 17394
rect -25386 17338 -25378 17394
rect -25450 17324 -25440 17338
rect -25388 17324 -25378 17338
rect -25450 17314 -25378 17324
rect -25450 17258 -25442 17314
rect -25386 17258 -25378 17314
rect -25450 17248 -25378 17258
rect -25450 17234 -25440 17248
rect -25388 17234 -25378 17248
rect -27178 17177 -26752 17229
rect -25450 17178 -25442 17234
rect -25386 17178 -25378 17234
rect -25450 17159 -25378 17178
rect -24139 16259 -24087 21756
rect -24191 16245 -24087 16259
rect -24191 16189 -24166 16245
rect -24110 16189 -24087 16245
rect -24191 16175 -24087 16189
rect -27939 15437 -27835 15451
rect -27939 15381 -27916 15437
rect -27860 15381 -27835 15437
rect -27939 15367 -27835 15381
rect -27939 9871 -27887 15367
rect -25572 14514 -24916 14562
rect -25575 14513 -24916 14514
rect -25572 14510 -24916 14513
rect -25517 14423 -25444 14456
rect -25517 14409 -25507 14423
rect -25455 14409 -25444 14423
rect -25517 14353 -25509 14409
rect -25453 14353 -25444 14409
rect -25517 14329 -25507 14353
rect -25455 14329 -25444 14353
rect -25517 14273 -25509 14329
rect -25453 14273 -25444 14329
rect -25517 14249 -25507 14273
rect -25455 14249 -25444 14273
rect -25517 14193 -25509 14249
rect -25453 14193 -25444 14249
rect -25517 14179 -25507 14193
rect -25455 14179 -25444 14193
rect -25517 14147 -25444 14179
rect -25518 13915 -25446 13935
rect -25518 13859 -25510 13915
rect -25454 13859 -25446 13915
rect -25518 13845 -25508 13859
rect -25456 13845 -25446 13859
rect -25518 13835 -25446 13845
rect -25518 13779 -25510 13835
rect -25454 13779 -25446 13835
rect -25518 13769 -25446 13779
rect -25518 13755 -25508 13769
rect -25456 13755 -25446 13769
rect -27246 13723 -26815 13755
rect -27246 13714 -26812 13723
rect -27246 13703 -26815 13714
rect -27246 9871 -27194 13703
rect -25518 13699 -25510 13755
rect -25454 13699 -25446 13755
rect -25518 13680 -25446 13699
rect -27939 9819 -27194 9871
rect -31130 6215 -31124 6331
rect -31008 6215 -31002 6331
rect -31130 6199 -31002 6215
rect -27246 5987 -27194 9819
rect -24968 10677 -24916 14510
rect -24139 10677 -24087 16175
rect -16781 21723 -11473 21851
rect -18223 14069 -18159 14083
rect -18223 14013 -18219 14069
rect -18163 14013 -18159 14069
rect -18223 13999 -18159 14013
rect -24968 10625 -24087 10677
rect -24968 6793 -24916 10625
rect -16781 7603 -16653 21723
rect -10016 21076 -9888 26530
rect -6086 21665 -5958 28550
rect 3399 28595 3463 28605
rect 4328 28595 4392 28605
rect 3399 28591 4398 28595
rect 3399 28589 4332 28591
rect 3399 28537 3405 28589
rect 3457 28537 4332 28589
rect 3399 28535 4332 28537
rect 4388 28535 4398 28591
rect 3399 28531 4398 28535
rect 8338 28592 8402 28602
rect 9399 28592 9463 28602
rect 8338 28588 9473 28592
rect 8338 28532 8342 28588
rect 8398 28586 9473 28588
rect 8398 28534 9405 28586
rect 9457 28534 9473 28586
rect 8398 28532 9473 28534
rect 3399 28521 3463 28531
rect 4328 28521 4392 28531
rect 8338 28528 9473 28532
rect 8338 28518 8402 28528
rect 9399 28518 9463 28528
rect -5279 27532 -5215 27542
rect -5279 27528 19935 27532
rect -5279 27472 -5275 27528
rect -5219 27472 19935 27528
rect -5279 27468 19935 27472
rect -5279 27458 -5215 27468
rect -3918 26855 -3854 26865
rect -3918 26851 17577 26855
rect -3918 26795 -3914 26851
rect -3858 26795 17577 26851
rect -3918 26791 17577 26795
rect -3918 26781 -3854 26791
rect 1952 25820 2080 25830
rect 7960 25820 8024 25830
rect 1952 25814 8024 25820
rect 1952 25762 1958 25814
rect 2010 25762 2022 25814
rect 2074 25762 7966 25814
rect 8018 25762 8024 25814
rect 1952 25756 8024 25762
rect 1952 25746 2080 25756
rect 7960 25746 8024 25756
rect -6086 21613 -6080 21665
rect -6028 21613 -6016 21665
rect -5964 21613 -5958 21665
rect -6086 21597 -5958 21613
rect -3501 25408 -3373 25433
rect -3501 25356 -3495 25408
rect -3443 25356 -3431 25408
rect -3379 25356 -3373 25408
rect -14184 20948 -9888 21076
rect -14184 15366 -14056 20948
rect -3501 20803 -3373 25356
rect 17513 24802 17577 26791
rect 19871 26005 19935 27468
rect 19871 25949 19875 26005
rect 19931 25949 19935 26005
rect 19871 25935 19935 25949
rect 19873 25594 19937 25608
rect 19873 25538 19877 25594
rect 19933 25538 19937 25594
rect 19873 24802 19937 25538
rect 17513 24738 19937 24802
rect 5715 24578 5783 24604
rect 5715 24522 5721 24578
rect 5777 24522 5783 24578
rect 5715 24512 5783 24522
rect 7068 24588 7132 24602
rect 7068 24532 7072 24588
rect 7128 24532 7132 24588
rect 7068 24518 7132 24532
rect 5715 24498 5723 24512
rect 5775 24498 5783 24512
rect 5715 24442 5721 24498
rect 5777 24442 5783 24498
rect 5715 24418 5723 24442
rect 5775 24418 5783 24442
rect 5715 24362 5721 24418
rect 5777 24362 5783 24418
rect 5715 24338 5723 24362
rect 5775 24338 5783 24362
rect 5715 24282 5721 24338
rect 5777 24282 5783 24338
rect 5715 24268 5723 24282
rect 5775 24268 5783 24282
rect 5715 24258 5783 24268
rect 5715 24202 5721 24258
rect 5777 24202 5783 24258
rect 5715 24176 5783 24202
rect 42856 24147 46190 24184
rect 42856 24145 42895 24147
rect 42951 24145 42975 24147
rect 43031 24145 43055 24147
rect 43111 24145 43135 24147
rect 43191 24145 43215 24147
rect 43271 24145 43295 24147
rect 43351 24145 43375 24147
rect 43431 24145 43455 24147
rect 43511 24145 43535 24147
rect 43591 24145 43615 24147
rect 43671 24145 43695 24147
rect 43751 24145 43775 24147
rect 43831 24145 43855 24147
rect 43911 24145 43935 24147
rect 43991 24145 44015 24147
rect 44071 24145 44095 24147
rect 44151 24145 44175 24147
rect 44231 24145 44255 24147
rect 44311 24145 44335 24147
rect 44391 24145 44415 24147
rect 44471 24145 44495 24147
rect 44551 24145 44575 24147
rect 44631 24145 44655 24147
rect 44711 24145 44735 24147
rect 44791 24145 44815 24147
rect 44871 24145 44895 24147
rect 44951 24145 44975 24147
rect 45031 24145 45055 24147
rect 45111 24145 45135 24147
rect 45191 24145 45215 24147
rect 45271 24145 45295 24147
rect 45351 24145 45375 24147
rect 45431 24145 45455 24147
rect 45511 24145 45535 24147
rect 45591 24145 45615 24147
rect 45671 24145 45695 24147
rect 45751 24145 45775 24147
rect 45831 24145 45855 24147
rect 45911 24145 45935 24147
rect 45991 24145 46015 24147
rect 46071 24145 46095 24147
rect 46151 24145 46190 24147
rect 3399 24097 3463 24109
rect 5643 24097 5707 24107
rect 3399 24095 5707 24097
rect 3399 24043 3405 24095
rect 3457 24091 5707 24095
rect 3457 24043 5649 24091
rect 3399 24039 5649 24043
rect 5701 24039 5707 24091
rect 3399 24033 5707 24039
rect 3399 24027 3463 24033
rect 5643 24023 5707 24033
rect 7017 24101 7081 24111
rect 9399 24101 9463 24111
rect 7017 24095 9467 24101
rect 7017 24043 7023 24095
rect 7075 24043 9405 24095
rect 9457 24043 9467 24095
rect 42856 24093 42865 24145
rect 43045 24093 43055 24145
rect 43111 24093 43121 24145
rect 43365 24093 43375 24145
rect 43431 24093 43441 24145
rect 43685 24093 43695 24145
rect 43751 24093 43761 24145
rect 44005 24093 44015 24145
rect 44071 24093 44081 24145
rect 44325 24093 44335 24145
rect 44391 24093 44401 24145
rect 44645 24093 44655 24145
rect 44711 24093 44721 24145
rect 44965 24093 44975 24145
rect 45031 24093 45041 24145
rect 45285 24093 45295 24145
rect 45351 24093 45361 24145
rect 45605 24093 45615 24145
rect 45671 24093 45681 24145
rect 45925 24093 45935 24145
rect 45991 24093 46001 24145
rect 46181 24093 46190 24145
rect 42856 24091 42895 24093
rect 42951 24091 42975 24093
rect 43031 24091 43055 24093
rect 43111 24091 43135 24093
rect 43191 24091 43215 24093
rect 43271 24091 43295 24093
rect 43351 24091 43375 24093
rect 43431 24091 43455 24093
rect 43511 24091 43535 24093
rect 43591 24091 43615 24093
rect 43671 24091 43695 24093
rect 43751 24091 43775 24093
rect 43831 24091 43855 24093
rect 43911 24091 43935 24093
rect 43991 24091 44015 24093
rect 44071 24091 44095 24093
rect 44151 24091 44175 24093
rect 44231 24091 44255 24093
rect 44311 24091 44335 24093
rect 44391 24091 44415 24093
rect 44471 24091 44495 24093
rect 44551 24091 44575 24093
rect 44631 24091 44655 24093
rect 44711 24091 44735 24093
rect 44791 24091 44815 24093
rect 44871 24091 44895 24093
rect 44951 24091 44975 24093
rect 45031 24091 45055 24093
rect 45111 24091 45135 24093
rect 45191 24091 45215 24093
rect 45271 24091 45295 24093
rect 45351 24091 45375 24093
rect 45431 24091 45455 24093
rect 45511 24091 45535 24093
rect 45591 24091 45615 24093
rect 45671 24091 45695 24093
rect 45751 24091 45775 24093
rect 45831 24091 45855 24093
rect 45911 24091 45935 24093
rect 45991 24091 46015 24093
rect 46071 24091 46095 24093
rect 46151 24091 46190 24093
rect 42856 24055 46190 24091
rect 7017 24037 9467 24043
rect 7017 24027 7081 24037
rect 9399 24027 9463 24037
rect 36066 24014 36130 24028
rect 36066 24012 36070 24014
rect 35939 23960 36070 24012
rect 36066 23958 36070 23960
rect 36126 23958 36130 24014
rect 36066 23944 36130 23958
rect 35152 23862 35216 23876
rect 35152 23806 35156 23862
rect 35212 23806 35216 23862
rect 35152 23792 35216 23806
rect 7091 23648 7155 23782
rect 7091 23592 7095 23648
rect 7151 23592 7155 23648
rect 39346 23711 39420 23724
rect 39346 23655 39355 23711
rect 39411 23655 39420 23711
rect 39346 23641 39357 23655
rect 39409 23641 39420 23655
rect 39346 23631 39420 23641
rect 7091 23578 7155 23592
rect 37819 23609 37892 23621
rect 37819 23579 37829 23609
rect 37881 23579 37892 23609
rect 37819 23523 37827 23579
rect 37883 23523 37892 23579
rect 37819 23493 37829 23523
rect 37881 23493 37892 23523
rect 37819 23482 37892 23493
rect 39346 23575 39355 23631
rect 39411 23575 39420 23631
rect 39346 23565 39420 23575
rect 39346 23551 39357 23565
rect 39409 23551 39420 23565
rect 39346 23495 39355 23551
rect 39411 23495 39420 23551
rect 39346 23483 39420 23495
rect 8787 23329 8943 23366
rect 8787 23273 8797 23329
rect 8853 23327 8877 23329
rect 8859 23275 8871 23327
rect 8853 23273 8877 23275
rect 8933 23273 8943 23329
rect 8787 23236 8943 23273
rect 37819 23192 37905 23204
rect 37819 23178 37836 23192
rect 37888 23178 37905 23192
rect 37819 23122 37834 23178
rect 37890 23122 37905 23178
rect 37819 23098 37836 23122
rect 37888 23098 37905 23122
rect 2550 23059 2614 23073
rect 2550 23003 2554 23059
rect 2610 23003 2614 23059
rect 2550 22989 2614 23003
rect 10202 23059 10266 23073
rect 10202 23003 10206 23059
rect 10262 23003 10266 23059
rect 10202 22989 10266 23003
rect 37819 23042 37834 23098
rect 37890 23042 37905 23098
rect 37819 23018 37836 23042
rect 37888 23018 37905 23042
rect 37819 22962 37834 23018
rect 37890 22962 37905 23018
rect 37819 22948 37836 22962
rect 37888 22948 37905 22962
rect 37819 22936 37905 22948
rect 39335 23198 39421 23210
rect 39335 23184 39352 23198
rect 39404 23184 39421 23198
rect 39335 23128 39350 23184
rect 39406 23128 39421 23184
rect 39335 23104 39352 23128
rect 39404 23104 39421 23128
rect 39335 23048 39350 23104
rect 39406 23048 39421 23104
rect 39335 23024 39352 23048
rect 39404 23024 39421 23048
rect 39335 22968 39350 23024
rect 39406 22968 39421 23024
rect 39335 22954 39352 22968
rect 39404 22954 39421 22968
rect 39335 22942 39421 22954
rect 35100 22790 35280 22800
rect 35760 22727 36021 22740
rect 35760 22725 35782 22727
rect 35838 22725 35862 22727
rect 35918 22725 35942 22727
rect 35998 22725 36021 22727
rect 35760 22673 35768 22725
rect 36012 22673 36021 22725
rect 35760 22671 35782 22673
rect 35838 22671 35862 22673
rect 35918 22671 35942 22673
rect 35998 22671 36021 22673
rect 35760 22658 36021 22671
rect 47556 22724 47792 22744
rect 35100 22600 35280 22610
rect 47556 22508 47566 22724
rect 47782 22508 47792 22724
rect 47556 22488 47792 22508
rect 39346 22385 39420 22398
rect 39346 22329 39355 22385
rect 39411 22329 39420 22385
rect 39346 22315 39357 22329
rect 39409 22315 39420 22329
rect 39346 22305 39420 22315
rect 37826 22273 37896 22290
rect 37826 22243 37835 22273
rect 37887 22243 37896 22273
rect 37826 22187 37833 22243
rect 37889 22187 37896 22243
rect 37826 22157 37835 22187
rect 37887 22157 37896 22187
rect 39346 22249 39355 22305
rect 39411 22249 39420 22305
rect 39346 22239 39420 22249
rect 39346 22225 39357 22239
rect 39409 22225 39420 22239
rect 39346 22169 39355 22225
rect 39411 22169 39420 22225
rect 39346 22157 39420 22169
rect 37826 22141 37896 22157
rect 4397 22037 4449 22047
rect -3501 20751 -3495 20803
rect -3443 20751 -3431 20803
rect -3379 20751 -3373 20803
rect -3501 20735 -3373 20751
rect -971 21621 -907 21635
rect -971 21565 -967 21621
rect -911 21565 -907 21621
rect -971 20711 -907 21565
rect 2910 21612 2962 22014
rect 3779 21985 4397 22037
rect 4397 21975 4449 21985
rect 8228 22037 8280 22047
rect 8280 21985 9098 22037
rect 8228 21975 8280 21985
rect 6312 21635 6364 21664
rect 6307 21621 6371 21635
rect 6307 21612 6311 21621
rect 2910 21565 6311 21612
rect 6367 21612 6371 21621
rect 9905 21612 9957 22096
rect 6367 21565 9957 21612
rect 37814 21812 37899 21833
rect 37814 21790 37830 21812
rect 37882 21790 37899 21812
rect 37814 21734 37828 21790
rect 37884 21734 37899 21790
rect 37814 21710 37830 21734
rect 37882 21710 37899 21734
rect 37814 21654 37828 21710
rect 37884 21654 37899 21710
rect 37814 21632 37830 21654
rect 37882 21632 37899 21654
rect 37814 21611 37899 21632
rect 39341 21832 39427 21844
rect 39341 21818 39358 21832
rect 39410 21818 39427 21832
rect 39341 21762 39356 21818
rect 39412 21762 39427 21818
rect 39341 21738 39358 21762
rect 39410 21738 39427 21762
rect 39341 21682 39356 21738
rect 39412 21682 39427 21738
rect 39341 21658 39358 21682
rect 39410 21658 39427 21682
rect 39341 21602 39356 21658
rect 39412 21602 39427 21658
rect 2910 21560 9957 21565
rect 35152 21581 35216 21595
rect 6307 21551 6371 21560
rect 35152 21525 35156 21581
rect 35212 21525 35216 21581
rect 39341 21588 39358 21602
rect 39410 21588 39427 21602
rect 39341 21576 39427 21588
rect 35152 21511 35216 21525
rect 35477 21375 35541 21389
rect 35477 21373 35481 21375
rect 35475 21321 35481 21373
rect 35477 21319 35481 21321
rect 35537 21373 35541 21375
rect 35939 21373 35991 21544
rect 35537 21321 35991 21373
rect 35537 21319 35541 21321
rect 35477 21305 35541 21319
rect 42854 21151 46188 21188
rect 42854 21149 42893 21151
rect 42949 21149 42973 21151
rect 43029 21149 43053 21151
rect 43109 21149 43133 21151
rect 43189 21149 43213 21151
rect 43269 21149 43293 21151
rect 43349 21149 43373 21151
rect 43429 21149 43453 21151
rect 43509 21149 43533 21151
rect 43589 21149 43613 21151
rect 43669 21149 43693 21151
rect 43749 21149 43773 21151
rect 43829 21149 43853 21151
rect 43909 21149 43933 21151
rect 43989 21149 44013 21151
rect 44069 21149 44093 21151
rect 44149 21149 44173 21151
rect 44229 21149 44253 21151
rect 44309 21149 44333 21151
rect 44389 21149 44413 21151
rect 44469 21149 44493 21151
rect 44549 21149 44573 21151
rect 44629 21149 44653 21151
rect 44709 21149 44733 21151
rect 44789 21149 44813 21151
rect 44869 21149 44893 21151
rect 44949 21149 44973 21151
rect 45029 21149 45053 21151
rect 45109 21149 45133 21151
rect 45189 21149 45213 21151
rect 45269 21149 45293 21151
rect 45349 21149 45373 21151
rect 45429 21149 45453 21151
rect 45509 21149 45533 21151
rect 45589 21149 45613 21151
rect 45669 21149 45693 21151
rect 45749 21149 45773 21151
rect 45829 21149 45853 21151
rect 45909 21149 45933 21151
rect 45989 21149 46013 21151
rect 46069 21149 46093 21151
rect 46149 21149 46188 21151
rect 42854 21097 42863 21149
rect 43043 21097 43053 21149
rect 43109 21097 43119 21149
rect 43363 21097 43373 21149
rect 43429 21097 43439 21149
rect 43683 21097 43693 21149
rect 43749 21097 43759 21149
rect 44003 21097 44013 21149
rect 44069 21097 44079 21149
rect 44323 21097 44333 21149
rect 44389 21097 44399 21149
rect 44643 21097 44653 21149
rect 44709 21097 44719 21149
rect 44963 21097 44973 21149
rect 45029 21097 45039 21149
rect 45283 21097 45293 21149
rect 45349 21097 45359 21149
rect 45603 21097 45613 21149
rect 45669 21097 45679 21149
rect 45923 21097 45933 21149
rect 45989 21097 45999 21149
rect 46179 21097 46188 21149
rect 42854 21095 42893 21097
rect 42949 21095 42973 21097
rect 43029 21095 43053 21097
rect 43109 21095 43133 21097
rect 43189 21095 43213 21097
rect 43269 21095 43293 21097
rect 43349 21095 43373 21097
rect 43429 21095 43453 21097
rect 43509 21095 43533 21097
rect 43589 21095 43613 21097
rect 43669 21095 43693 21097
rect 43749 21095 43773 21097
rect 43829 21095 43853 21097
rect 43909 21095 43933 21097
rect 43989 21095 44013 21097
rect 44069 21095 44093 21097
rect 44149 21095 44173 21097
rect 44229 21095 44253 21097
rect 44309 21095 44333 21097
rect 44389 21095 44413 21097
rect 44469 21095 44493 21097
rect 44549 21095 44573 21097
rect 44629 21095 44653 21097
rect 44709 21095 44733 21097
rect 44789 21095 44813 21097
rect 44869 21095 44893 21097
rect 44949 21095 44973 21097
rect 45029 21095 45053 21097
rect 45109 21095 45133 21097
rect 45189 21095 45213 21097
rect 45269 21095 45293 21097
rect 45349 21095 45373 21097
rect 45429 21095 45453 21097
rect 45509 21095 45533 21097
rect 45589 21095 45613 21097
rect 45669 21095 45693 21097
rect 45749 21095 45773 21097
rect 45829 21095 45853 21097
rect 45909 21095 45933 21097
rect 45989 21095 46013 21097
rect 46069 21095 46093 21097
rect 46149 21095 46188 21097
rect 42854 21059 46188 21095
rect 14688 21023 14752 21037
rect 6312 20967 6364 20997
rect 14688 20967 14692 21023
rect 14748 20967 14752 21023
rect 4397 20945 4449 20955
rect 6310 20953 6374 20967
rect 6310 20945 6314 20953
rect 4387 20893 4397 20945
rect 4449 20897 6314 20945
rect 6370 20945 6374 20953
rect 8228 20945 8280 20955
rect 14688 20953 14752 20967
rect 6370 20897 8228 20945
rect 4449 20893 8228 20897
rect 8280 20893 8290 20945
rect 4397 20883 4449 20893
rect 6310 20883 6374 20893
rect 8228 20883 8280 20893
rect -971 20655 -967 20711
rect -911 20655 -907 20711
rect -971 20641 -907 20655
rect 23670 20216 23734 20226
rect 22767 20210 23734 20216
rect 22767 20158 23676 20210
rect 23728 20158 23734 20210
rect 22767 20152 23734 20158
rect -444 20109 -380 20119
rect 5394 20109 5458 20119
rect 9394 20109 9458 20119
rect 12373 20109 12501 20121
rect -14184 15310 -14148 15366
rect -14092 15310 -14056 15366
rect -14184 15264 -14056 15310
rect -10970 20105 12512 20109
rect -10970 20103 12379 20105
rect -10970 20051 -438 20103
rect -386 20051 5400 20103
rect 5452 20051 9400 20103
rect 9452 20051 12379 20103
rect -10970 20039 12379 20051
rect -10970 19987 -438 20039
rect -386 19987 5400 20039
rect 5452 19987 9400 20039
rect 9452 19989 12379 20039
rect 12495 19989 12512 20105
rect 9452 19987 12512 19989
rect -10970 19981 12512 19987
rect -13064 14137 -13000 14151
rect -13064 14081 -13060 14137
rect -13004 14081 -13000 14137
rect -13064 14067 -13000 14081
rect -10970 10219 -10842 19981
rect -444 19971 -380 19981
rect 5394 19971 5458 19981
rect 9394 19971 9458 19981
rect 12373 19973 12501 19981
rect 51 19509 115 19523
rect 51 19453 55 19509
rect 111 19453 115 19509
rect -756 19208 -692 19222
rect -756 19152 -752 19208
rect -696 19152 -692 19208
rect -756 19049 -692 19152
rect 51 19051 115 19453
rect 1684 19410 1748 19420
rect 7394 19410 7458 19420
rect 11295 19410 11423 19422
rect 1684 19406 11452 19410
rect 1684 19404 11301 19406
rect 1684 19352 1690 19404
rect 1742 19352 7400 19404
rect 7452 19352 11301 19404
rect 1684 19340 11301 19352
rect 1684 19288 1690 19340
rect 1742 19288 3401 19340
rect 3453 19288 7400 19340
rect 7452 19290 11301 19340
rect 11417 19290 11452 19406
rect 7452 19288 11452 19290
rect 1684 19282 11452 19288
rect 14687 19323 14751 19337
rect 1684 19272 1748 19282
rect 3395 19272 3459 19282
rect 7394 19272 7458 19282
rect 11295 19274 11423 19282
rect 14687 19267 14691 19323
rect 14747 19267 14751 19323
rect 14687 19253 14751 19267
rect 4857 19168 5194 19183
rect 4857 19158 4877 19168
rect 5173 19158 5194 19168
rect 3061 19102 3125 19116
rect 3061 19046 3065 19102
rect 3121 19046 3125 19102
rect 3061 19032 3125 19046
rect 4857 19042 4871 19158
rect 5179 19042 5194 19158
rect 4857 19032 4877 19042
rect 5173 19032 5194 19042
rect 7085 19102 7149 19116
rect 7085 19046 7089 19102
rect 7145 19046 7149 19102
rect 7085 19032 7149 19046
rect 8981 19102 9045 19116
rect 8981 19046 8985 19102
rect 9041 19046 9045 19102
rect 8981 19032 9045 19046
rect 10232 19054 10296 19068
rect 4857 19017 5194 19032
rect 10232 18998 10236 19054
rect 10292 18998 10296 19054
rect 10232 18984 10296 18998
rect 20971 19062 21035 19072
rect 22767 19062 22831 20152
rect 23670 20142 23734 20152
rect 23689 19378 23753 19392
rect 23689 19322 23693 19378
rect 23749 19322 23753 19378
rect 23689 19308 23753 19322
rect 20971 19058 22831 19062
rect 20971 19002 20975 19058
rect 21031 19002 22831 19058
rect 20971 18998 22831 19002
rect 20971 18988 21035 18998
rect 5707 18906 5771 18920
rect 5707 18850 5711 18906
rect 5767 18850 5771 18906
rect 5707 18836 5771 18850
rect 7706 18906 7770 18920
rect 7706 18850 7710 18906
rect 7766 18850 7770 18906
rect 7706 18836 7770 18850
rect 8280 18714 8344 18728
rect 4899 18647 4963 18661
rect 4899 18591 4903 18647
rect 4959 18591 4963 18647
rect 4899 18577 4963 18591
rect 6897 18647 6961 18661
rect 6897 18591 6901 18647
rect 6957 18591 6961 18647
rect 8280 18658 8284 18714
rect 8340 18658 8344 18714
rect 8280 18644 8344 18658
rect 13574 18684 13638 18698
rect 13574 18628 13578 18684
rect 13634 18628 13638 18684
rect 13574 18614 13638 18628
rect 6897 18577 6961 18591
rect 22767 18428 22831 18998
rect 23658 18428 23722 18438
rect 22767 18422 23722 18428
rect 22767 18370 23664 18422
rect 23716 18370 23722 18422
rect 22767 18364 23722 18370
rect 23658 18354 23722 18364
rect 3707 18308 3771 18322
rect 3707 18252 3711 18308
rect 3767 18252 3771 18308
rect 3707 18238 3771 18252
rect 9706 18308 9770 18322
rect 9706 18252 9710 18308
rect 9766 18252 9770 18308
rect 9706 18238 9770 18252
rect 2898 18027 2962 18041
rect 2898 17971 2902 18027
rect 2958 17971 2962 18027
rect 2898 17957 2962 17971
rect 8899 18027 8963 18041
rect 8899 17971 8903 18027
rect 8959 17971 8963 18027
rect 8899 17957 8963 17971
rect 233 17768 297 17782
rect 233 17712 237 17768
rect 293 17712 297 17768
rect 233 17698 297 17712
rect 14689 17538 14753 17552
rect -821 17521 -757 17535
rect -821 17465 -817 17521
rect -761 17465 -757 17521
rect 14689 17482 14693 17538
rect 14749 17482 14753 17538
rect 14689 17468 14753 17482
rect 23689 17548 23753 17562
rect 23689 17492 23693 17548
rect 23749 17492 23753 17548
rect 23689 17478 23753 17492
rect -821 17451 -757 17465
rect 7393 17359 7457 17369
rect 9396 17359 9460 17369
rect 13885 17359 13949 17369
rect 7393 17353 13962 17359
rect 7393 17301 7399 17353
rect 7451 17301 9402 17353
rect 9454 17301 13891 17353
rect 13943 17301 13962 17353
rect 4295 17285 4359 17299
rect -445 17221 -381 17231
rect 1684 17221 1748 17231
rect -10479 17215 1748 17221
rect 4295 17229 4299 17285
rect 4355 17229 4359 17285
rect 4295 17215 4359 17229
rect 6227 17285 6291 17299
rect 6227 17229 6231 17285
rect 6287 17229 6291 17285
rect 6227 17215 6291 17229
rect 7393 17289 13962 17301
rect 7393 17237 7399 17289
rect 7451 17237 9402 17289
rect 9454 17237 13891 17289
rect 13943 17237 13962 17289
rect 7393 17231 13962 17237
rect 7393 17221 7457 17231
rect 9396 17221 9460 17231
rect 13885 17221 13949 17231
rect -10479 17163 -439 17215
rect -387 17163 1690 17215
rect 1742 17163 1748 17215
rect -10479 17153 1748 17163
rect -10479 17097 -10412 17153
rect -10356 17151 1748 17153
rect -10356 17099 -439 17151
rect -387 17099 1690 17151
rect 1742 17099 1748 17151
rect -10356 17097 1748 17099
rect -10479 17092 1748 17097
rect -10416 17083 -10352 17092
rect -445 17083 -381 17092
rect 1684 17083 1748 17092
rect 13603 17083 13667 17093
rect 14690 17083 14754 17093
rect 13603 17079 14754 17083
rect 13603 17023 13607 17079
rect 13663 17077 14754 17079
rect 13663 17025 14696 17077
rect 14748 17025 14754 17077
rect 13663 17023 14754 17025
rect 13603 17019 14754 17023
rect 13603 17009 13667 17019
rect 14690 17009 14754 17019
rect 3393 16866 3457 16876
rect 5393 16866 5457 16876
rect 13277 16866 13341 16876
rect 3393 16860 13351 16866
rect 3393 16808 3399 16860
rect 3451 16808 5399 16860
rect 5451 16808 13283 16860
rect 13335 16808 13351 16860
rect 3393 16796 13351 16808
rect 3393 16744 3399 16796
rect 3451 16744 5399 16796
rect 5451 16744 13283 16796
rect 13335 16744 13351 16796
rect 3393 16738 13351 16744
rect 3393 16728 3457 16738
rect 5393 16728 5457 16738
rect 13277 16728 13341 16738
rect 251 16432 11139 16456
rect -10415 16288 -10351 16298
rect -3926 16288 -3862 16298
rect -10415 16284 -3862 16288
rect -10415 16228 -10411 16284
rect -10355 16282 -3862 16284
rect -10355 16230 -3920 16282
rect -3868 16230 -3862 16282
rect -10355 16228 -3862 16230
rect 251 16252 261 16432
rect 11129 16252 11139 16432
rect 251 16228 11139 16252
rect -10415 16224 -3862 16228
rect -10415 16214 -10351 16224
rect -3926 16214 -3862 16224
rect -5786 15704 -5722 15718
rect -5786 15648 -5782 15704
rect -5726 15648 -5722 15704
rect -5786 15634 -5722 15648
rect -3914 15135 -3862 16214
rect 28 16162 187 16199
rect -3008 15450 -2944 15464
rect -3008 15394 -3004 15450
rect -2948 15394 -2944 15450
rect -3008 15380 -2944 15394
rect -5026 14663 -4390 14715
rect -5026 14411 -4974 14663
rect -4902 14431 -4832 14456
rect -4902 14409 -4893 14431
rect -4841 14409 -4832 14431
rect -4902 14353 -4895 14409
rect -4839 14353 -4832 14409
rect -4902 14329 -4893 14353
rect -4841 14329 -4832 14353
rect -4902 14273 -4895 14329
rect -4839 14273 -4832 14329
rect -4902 14251 -4893 14273
rect -4841 14251 -4832 14273
rect -4902 14226 -4832 14251
rect -6544 14135 -6480 14151
rect -6544 14083 -6538 14135
rect -6486 14083 -6480 14135
rect -6544 12886 -6480 14083
rect -4917 13974 -4833 14008
rect -4917 13960 -4901 13974
rect -4849 13960 -4833 13974
rect -4917 13904 -4903 13960
rect -4847 13904 -4833 13960
rect -4917 13880 -4901 13904
rect -4849 13880 -4833 13904
rect -4917 13824 -4903 13880
rect -4847 13824 -4833 13880
rect -4917 13800 -4901 13824
rect -4849 13800 -4833 13824
rect -4917 13744 -4903 13800
rect -4847 13744 -4833 13800
rect -4917 13730 -4901 13744
rect -4849 13730 -4833 13744
rect -4917 13696 -4833 13730
rect -5006 13597 -4731 13649
rect -6544 12834 -6538 12886
rect -6486 12834 -6480 12886
rect -6544 12818 -6480 12834
rect -5851 12886 -5787 12902
rect -5851 12834 -5845 12886
rect -5793 12834 -5787 12886
rect -5851 12213 -5787 12834
rect -5851 12161 -5845 12213
rect -5793 12161 -5787 12213
rect -5851 12145 -5787 12161
rect -5845 10943 -5793 10953
rect -6411 10890 -6103 10942
rect -6411 10701 -6359 10890
rect -6162 10823 -5937 10843
rect -6162 10767 -6158 10823
rect -6102 10821 -6078 10823
rect -6022 10821 -5998 10823
rect -6088 10769 -6078 10821
rect -6022 10769 -6012 10821
rect -6102 10767 -6078 10769
rect -6022 10767 -5998 10769
rect -5942 10767 -5937 10823
rect -6162 10748 -5937 10767
rect -6411 10649 -6104 10701
rect -10970 10163 -10966 10219
rect -10910 10163 -10842 10219
rect -10970 10139 -10842 10163
rect -6156 10214 -6104 10649
rect -5845 10412 -5793 10891
rect -5707 10822 -5401 10848
rect -5707 10766 -5702 10822
rect -5646 10820 -5622 10822
rect -5566 10820 -5542 10822
rect -5486 10820 -5462 10822
rect -5624 10768 -5622 10820
rect -5560 10768 -5548 10820
rect -5486 10768 -5484 10820
rect -5646 10766 -5622 10768
rect -5566 10766 -5542 10768
rect -5486 10766 -5462 10768
rect -5406 10766 -5401 10822
rect -5707 10741 -5401 10766
rect -5845 10401 -5792 10412
rect -5793 10349 -5792 10401
rect -5845 10339 -5792 10349
rect -6156 10200 -6092 10214
rect -6156 10144 -6152 10200
rect -6096 10144 -6092 10200
rect -6156 10130 -6092 10144
rect -6156 9717 -6104 10130
rect -6383 9665 -6104 9717
rect -6383 9453 -6331 9665
rect -6167 9580 -5929 9602
rect -6167 9524 -6156 9580
rect -6100 9578 -6076 9580
rect -6020 9578 -5996 9580
rect -6086 9526 -6076 9578
rect -6020 9526 -6010 9578
rect -6100 9524 -6076 9526
rect -6020 9524 -5996 9526
rect -5940 9524 -5929 9580
rect -6167 9503 -5929 9524
rect -6383 9401 -6110 9453
rect -5845 9452 -5793 10339
rect -5348 10214 -5296 10935
rect -4783 10243 -4731 13597
rect -4442 10243 -4390 14663
rect -3914 14139 -3862 15083
rect -678 15136 -626 15146
rect -3144 14980 -3061 15008
rect -3144 14966 -3129 14980
rect -3077 14966 -3061 14980
rect -3144 14910 -3131 14966
rect -3075 14910 -3061 14966
rect -3144 14886 -3129 14910
rect -3077 14886 -3061 14910
rect -3144 14830 -3131 14886
rect -3075 14830 -3061 14886
rect -3144 14806 -3129 14830
rect -3077 14806 -3061 14830
rect -3144 14750 -3131 14806
rect -3075 14750 -3061 14806
rect -3144 14736 -3129 14750
rect -3077 14736 -3061 14750
rect -3144 14709 -3061 14736
rect -3023 14640 -2959 14654
rect -3023 14584 -3019 14640
rect -2963 14584 -2959 14640
rect -3023 14570 -2959 14584
rect -3914 12635 -3862 14087
rect -2598 13133 -2534 13147
rect -2598 13077 -2594 13133
rect -2538 13077 -2534 13133
rect -2598 13063 -2534 13077
rect -1808 13117 -1725 13143
rect -1808 13061 -1795 13117
rect -1739 13061 -1725 13117
rect -1808 13051 -1725 13061
rect -1808 13037 -1793 13051
rect -1741 13037 -1725 13051
rect -1808 12981 -1795 13037
rect -1739 12981 -1725 13037
rect -1808 12957 -1793 12981
rect -1741 12957 -1725 12981
rect -1808 12901 -1795 12957
rect -1739 12901 -1725 12957
rect -1808 12877 -1793 12901
rect -1741 12877 -1725 12901
rect -1808 12821 -1795 12877
rect -1739 12821 -1725 12877
rect -1808 12807 -1793 12821
rect -1741 12807 -1725 12821
rect -1808 12797 -1725 12807
rect -1808 12741 -1795 12797
rect -1739 12741 -1725 12797
rect -1808 12716 -1725 12741
rect -5361 10200 -5296 10214
rect -5361 10198 -5357 10200
rect -5363 10146 -5357 10198
rect -5361 10144 -5357 10146
rect -5301 10144 -5296 10200
rect -4789 10229 -4725 10243
rect -4789 10173 -4785 10229
rect -4729 10173 -4725 10229
rect -4789 10159 -4725 10173
rect -4448 10229 -4384 10243
rect -4448 10173 -4444 10229
rect -4388 10173 -4384 10229
rect -4448 10159 -4384 10173
rect -5361 10130 -5296 10144
rect -5708 9580 -5399 9605
rect -5708 9578 -5702 9580
rect -5646 9578 -5622 9580
rect -5566 9578 -5542 9580
rect -5486 9578 -5462 9580
rect -5406 9578 -5399 9580
rect -5646 9526 -5644 9578
rect -5464 9526 -5462 9578
rect -5400 9526 -5399 9578
rect -5708 9524 -5702 9526
rect -5646 9524 -5622 9526
rect -5566 9524 -5542 9526
rect -5486 9524 -5462 9526
rect -5406 9524 -5399 9526
rect -5708 9499 -5399 9524
rect -5348 9406 -5296 10130
rect -5845 9390 -5793 9400
rect -16781 7547 -16745 7603
rect -16689 7547 -16653 7603
rect -5853 8168 -5789 8184
rect -5853 8116 -5847 8168
rect -5795 8116 -5789 8168
rect -16781 7501 -16653 7547
rect -6565 7585 -6501 7601
rect -6565 7533 -6559 7585
rect -6507 7533 -6501 7585
rect -7214 7231 -6751 7253
rect -7214 7015 -7211 7231
rect -6755 7015 -6751 7231
rect -7214 6993 -6751 7015
rect -25628 6741 -24916 6793
rect -25521 6660 -25446 6679
rect -25521 6646 -25510 6660
rect -25458 6646 -25446 6660
rect -25521 6590 -25512 6646
rect -25456 6590 -25446 6646
rect -25521 6566 -25510 6590
rect -25458 6566 -25446 6590
rect -25521 6510 -25512 6566
rect -25456 6510 -25446 6566
rect -25521 6486 -25510 6510
rect -25458 6486 -25446 6510
rect -25521 6430 -25512 6486
rect -25456 6430 -25446 6486
rect -25521 6416 -25510 6430
rect -25458 6416 -25446 6430
rect -25521 6398 -25446 6416
rect -18251 6299 -18187 6313
rect -18251 6243 -18247 6299
rect -18191 6243 -18187 6299
rect -18251 6229 -18187 6243
rect -13075 6309 -13011 6323
rect -13075 6253 -13071 6309
rect -13015 6253 -13011 6309
rect -13075 6239 -13011 6253
rect -6565 6307 -6501 7533
rect -5853 7589 -5789 8116
rect -5853 7537 -5847 7589
rect -5795 7537 -5789 7589
rect -5853 7521 -5789 7537
rect -4783 6803 -4731 10159
rect -5036 6751 -4731 6803
rect -4917 6691 -4836 6705
rect -4917 6635 -4905 6691
rect -4849 6635 -4836 6691
rect -4917 6613 -4903 6635
rect -4851 6613 -4836 6635
rect -4917 6611 -4836 6613
rect -4917 6555 -4905 6611
rect -4849 6555 -4836 6611
rect -4917 6549 -4903 6555
rect -4851 6549 -4836 6555
rect -4917 6537 -4836 6549
rect -4917 6531 -4903 6537
rect -4851 6531 -4836 6537
rect -4917 6475 -4905 6531
rect -4849 6475 -4836 6531
rect -4917 6473 -4836 6475
rect -4917 6451 -4903 6473
rect -4851 6451 -4836 6473
rect -4917 6395 -4905 6451
rect -4849 6395 -4836 6451
rect -4917 6382 -4836 6395
rect -6565 6255 -6559 6307
rect -6507 6255 -6501 6307
rect -6565 6239 -6501 6255
rect -25522 6173 -25447 6184
rect -25522 6159 -25511 6173
rect -25459 6159 -25447 6173
rect -25522 6103 -25513 6159
rect -25457 6103 -25447 6159
rect -25522 6079 -25511 6103
rect -25459 6079 -25447 6103
rect -25522 6023 -25513 6079
rect -25457 6023 -25447 6079
rect -25522 5999 -25511 6023
rect -25459 5999 -25447 6023
rect -27246 5936 -26782 5987
rect -27165 5935 -26782 5936
rect -25522 5943 -25513 5999
rect -25457 5943 -25447 5999
rect -4907 6146 -4841 6173
rect -4907 6124 -4900 6146
rect -4848 6124 -4841 6146
rect -4907 6068 -4902 6124
rect -4846 6068 -4841 6124
rect -4907 6044 -4900 6068
rect -4848 6044 -4841 6068
rect -25522 5929 -25511 5943
rect -25459 5929 -25447 5943
rect -25522 5919 -25447 5929
rect -5029 5826 -4977 5994
rect -4907 5988 -4902 6044
rect -4846 5988 -4841 6044
rect -4907 5966 -4900 5988
rect -4848 5966 -4841 5988
rect -4907 5940 -4841 5966
rect -4442 5826 -4390 10159
rect -3914 9437 -3862 12583
rect -1498 12405 -1434 12419
rect -1498 12349 -1494 12405
rect -1438 12349 -1434 12405
rect -2885 12324 -2821 12338
rect -1498 12335 -1434 12349
rect -2885 12268 -2881 12324
rect -2825 12268 -2821 12324
rect -2885 12254 -2821 12268
rect -1926 11531 -1862 11545
rect -1926 11475 -1922 11531
rect -1866 11475 -1862 11531
rect -1926 11461 -1862 11475
rect -1759 11522 -1693 11539
rect -1759 11466 -1754 11522
rect -1698 11466 -1693 11522
rect -1759 11456 -1693 11466
rect -1759 11442 -1752 11456
rect -1700 11442 -1693 11456
rect -1759 11386 -1754 11442
rect -1698 11386 -1693 11442
rect -1759 11362 -1752 11386
rect -1700 11362 -1693 11386
rect -1759 11306 -1754 11362
rect -1698 11306 -1693 11362
rect -1759 11282 -1752 11306
rect -1700 11282 -1693 11306
rect -1759 11226 -1754 11282
rect -1698 11226 -1693 11282
rect -1759 11212 -1752 11226
rect -1700 11212 -1693 11226
rect -1759 11202 -1693 11212
rect -1759 11146 -1754 11202
rect -1698 11146 -1693 11202
rect -1759 11130 -1693 11146
rect -3914 9375 -3862 9385
rect -3415 11034 -3363 11044
rect -5029 5774 -4390 5826
rect -3415 7835 -3363 10982
rect -1498 10779 -1434 10793
rect -2212 10725 -2148 10739
rect -2212 10669 -2208 10725
rect -2152 10669 -2148 10725
rect -1498 10723 -1494 10779
rect -1438 10723 -1434 10779
rect -1498 10709 -1434 10723
rect -2212 10655 -2148 10669
rect -678 10402 -626 15084
rect -1926 9933 -1862 9947
rect -1926 9877 -1922 9933
rect -1866 9877 -1862 9933
rect -1926 9863 -1862 9877
rect -1759 9919 -1695 9940
rect -1759 9863 -1755 9919
rect -1699 9863 -1695 9919
rect -1759 9853 -1695 9863
rect -1759 9839 -1753 9853
rect -1701 9839 -1695 9853
rect -1759 9783 -1755 9839
rect -1699 9783 -1695 9839
rect -1759 9759 -1753 9783
rect -1701 9759 -1695 9783
rect -1759 9703 -1755 9759
rect -1699 9703 -1695 9759
rect -1759 9679 -1753 9703
rect -1701 9679 -1695 9703
rect -1759 9623 -1755 9679
rect -1699 9623 -1695 9679
rect -1759 9609 -1753 9623
rect -1701 9609 -1695 9623
rect -1759 9599 -1695 9609
rect -1759 9543 -1755 9599
rect -1699 9543 -1695 9599
rect -1759 9522 -1695 9543
rect -1149 9435 -1097 9451
rect -2212 9125 -2148 9139
rect -2212 9069 -2208 9125
rect -2152 9069 -2148 9125
rect -2212 9055 -2148 9069
rect -1498 9121 -1434 9135
rect -1498 9065 -1494 9121
rect -1438 9065 -1434 9121
rect -1498 9051 -1434 9065
rect -2598 8331 -2534 8345
rect -2598 8275 -2594 8331
rect -2538 8275 -2534 8331
rect -2598 8261 -2534 8275
rect -1758 8318 -1690 8340
rect -1758 8262 -1752 8318
rect -1696 8262 -1690 8318
rect -1758 8252 -1690 8262
rect -1758 8238 -1750 8252
rect -1698 8238 -1690 8252
rect -1758 8182 -1752 8238
rect -1696 8182 -1690 8238
rect -1758 8158 -1750 8182
rect -1698 8158 -1690 8182
rect -1758 8102 -1752 8158
rect -1696 8102 -1690 8158
rect -1758 8078 -1750 8102
rect -1698 8078 -1690 8102
rect -1758 8022 -1752 8078
rect -1696 8022 -1690 8078
rect -1758 8008 -1750 8022
rect -1698 8008 -1690 8022
rect -1758 7998 -1690 8008
rect -1758 7942 -1752 7998
rect -1696 7942 -1690 7998
rect -1758 7920 -1690 7942
rect -3415 6310 -3363 7783
rect -1149 7835 -1097 9383
rect -1498 7582 -1434 7596
rect -2885 7523 -2821 7537
rect -2885 7467 -2881 7523
rect -2825 7467 -2821 7523
rect -1498 7526 -1494 7582
rect -1438 7526 -1434 7582
rect -1498 7512 -1434 7526
rect -2885 7453 -2821 7467
rect -1498 7238 -1434 7268
rect -1498 7224 -1492 7238
rect -1440 7224 -1434 7238
rect -1498 7168 -1494 7224
rect -1438 7168 -1434 7224
rect -1498 7144 -1492 7168
rect -1440 7144 -1434 7168
rect -1498 7088 -1494 7144
rect -1438 7088 -1434 7144
rect -1498 7064 -1492 7088
rect -1440 7064 -1434 7088
rect -1498 7008 -1494 7064
rect -1438 7008 -1434 7064
rect -1498 6994 -1492 7008
rect -1440 6994 -1434 7008
rect -1498 6964 -1434 6994
rect -1498 6447 -1434 6461
rect -1498 6391 -1494 6447
rect -1438 6391 -1434 6447
rect -1498 6377 -1434 6391
rect -3415 5723 -3363 6258
rect -3050 6038 -2986 6052
rect -3050 5982 -3046 6038
rect -2990 5982 -2986 6038
rect -3050 5968 -2986 5982
rect -3415 5057 -3363 5671
rect -3193 5558 -3110 5587
rect -3193 5544 -3178 5558
rect -3126 5544 -3110 5558
rect -3193 5488 -3180 5544
rect -3124 5488 -3110 5544
rect -3193 5464 -3178 5488
rect -3126 5464 -3110 5488
rect -3193 5408 -3180 5464
rect -3124 5408 -3110 5464
rect -3193 5384 -3178 5408
rect -3126 5384 -3110 5408
rect -3193 5328 -3180 5384
rect -3124 5328 -3110 5384
rect -3193 5314 -3178 5328
rect -3126 5314 -3110 5328
rect -3193 5286 -3110 5314
rect -3028 5229 -2964 5243
rect -3028 5173 -3024 5229
rect -2968 5173 -2964 5229
rect -3028 5159 -2964 5173
rect -1149 5129 -1097 7783
rect -678 5723 -626 10350
rect -678 5661 -626 5671
rect -279 12637 -227 12647
rect -279 11035 -227 12585
rect -1149 5067 -1097 5077
rect -10766 5047 -10702 5057
rect -3427 5047 -3363 5057
rect -10766 5043 -3363 5047
rect -10766 4987 -10762 5043
rect -10706 5041 -3363 5043
rect -10706 4989 -3421 5041
rect -3369 4989 -3363 5041
rect -10706 4987 -3363 4989
rect -10766 4983 -3363 4987
rect -10766 4973 -10702 4983
rect -3427 4973 -3363 4983
rect -279 3789 -227 10983
rect 28 10666 39 16162
rect 175 10666 187 16162
rect 11239 16173 11399 16194
rect 11239 14437 11251 16173
rect 11387 14437 11399 16173
rect 23686 15784 23750 15798
rect 14665 15707 14771 15743
rect 23686 15728 23690 15784
rect 23746 15728 23750 15784
rect 23686 15714 23750 15728
rect 14665 15651 14690 15707
rect 14746 15651 14771 15707
rect 14665 15616 14771 15651
rect 20928 15492 20992 15506
rect 20928 15436 20932 15492
rect 20988 15436 20992 15492
rect 20928 15422 20992 15436
rect 14690 15224 14754 15238
rect 14690 15168 14694 15224
rect 14750 15168 14754 15224
rect 14690 15154 14754 15168
rect 11239 14416 11399 14437
rect 23686 13993 23750 14007
rect 11257 13946 11384 13964
rect 11257 12998 11262 13946
rect 11378 12998 11384 13946
rect 14685 13961 14749 13975
rect 14685 13905 14689 13961
rect 14745 13905 14749 13961
rect 23686 13937 23690 13993
rect 23746 13937 23750 13993
rect 23686 13923 23750 13937
rect 14685 13891 14749 13905
rect 13636 13528 13700 13538
rect 14690 13528 14754 13538
rect 13636 13524 14754 13528
rect 13636 13468 13640 13524
rect 13696 13522 14754 13524
rect 13696 13470 14696 13522
rect 14748 13470 14754 13522
rect 13696 13468 14754 13470
rect 13636 13464 14754 13468
rect 13636 13454 13700 13464
rect 14690 13454 14754 13464
rect 23685 13006 23749 13016
rect 11257 12980 11384 12998
rect 23094 13000 23749 13006
rect 23094 12948 23691 13000
rect 23743 12948 23749 13000
rect 23094 12942 23749 12948
rect 14702 12176 14766 12190
rect 11243 12110 11398 12139
rect 11243 11334 11252 12110
rect 11388 11334 11398 12110
rect 14702 12120 14706 12176
rect 14762 12120 14766 12176
rect 14702 12106 14766 12120
rect 20985 11906 21049 11916
rect 23094 11906 23158 12942
rect 23685 12932 23749 12942
rect 23691 12186 23755 12200
rect 23691 12130 23695 12186
rect 23751 12130 23755 12186
rect 23691 12116 23755 12130
rect 20968 11902 23753 11906
rect 20968 11846 20989 11902
rect 21045 11846 23753 11902
rect 20968 11842 23753 11846
rect 20985 11832 21049 11842
rect 13699 11676 13763 11686
rect 14692 11676 14756 11686
rect 13699 11672 14756 11676
rect 13699 11616 13703 11672
rect 13759 11670 14756 11672
rect 13759 11618 14698 11670
rect 14750 11618 14756 11670
rect 13759 11616 14756 11618
rect 13699 11612 14756 11616
rect 13699 11602 13763 11612
rect 14692 11602 14756 11612
rect 23689 11513 23753 11842
rect 23689 11461 23695 11513
rect 23747 11461 23753 11513
rect 23689 11445 23753 11461
rect 11243 11306 11398 11334
rect 28 10630 187 10666
rect 6483 10514 11218 10547
rect 6483 10378 6502 10514
rect 11198 10378 11218 10514
rect 6483 10346 11218 10378
rect 14691 10379 14755 10393
rect 14691 10323 14695 10379
rect 14751 10323 14755 10379
rect 14691 10309 14755 10323
rect 23691 10376 23755 10390
rect 23691 10320 23695 10376
rect 23751 10320 23755 10376
rect 23691 10306 23755 10320
rect 5223 9418 5276 9428
rect 24544 9418 24608 9434
rect 5223 9417 24550 9418
rect 5275 9366 24550 9417
rect 24602 9366 24608 9418
rect 5275 9365 24608 9366
rect 5223 9355 5276 9365
rect 24544 9350 24608 9365
rect 36066 9150 36130 9164
rect 23208 7845 23261 7855
rect 17771 7844 23261 7845
rect 17771 7792 23208 7844
rect 23260 7792 23261 7844
rect 17771 7717 17824 7792
rect 23208 7782 23261 7792
rect 12920 7664 17824 7717
rect 25495 7651 25559 9116
rect 35842 9096 36070 9150
rect 35489 8527 35553 8541
rect 35489 8471 35493 8527
rect 35549 8471 35553 8527
rect 35489 8457 35553 8471
rect 35842 8400 35896 9096
rect 36066 9094 36070 9096
rect 36126 9094 36130 9150
rect 36066 9080 36130 9094
rect 36631 8465 36695 8479
rect 35982 8413 36635 8465
rect 36631 8409 36635 8413
rect 36691 8409 36695 8465
rect 36631 8395 36695 8409
rect 35024 8279 35088 8293
rect 35024 8223 35028 8279
rect 35084 8223 35088 8279
rect 35024 8209 35088 8223
rect 40100 8117 40181 8131
rect 40100 8095 40114 8117
rect 40166 8095 40181 8117
rect 38575 8033 38645 8048
rect 38575 7977 38582 8033
rect 38638 7977 38645 8033
rect 38575 7971 38584 7977
rect 38636 7971 38645 7977
rect 38575 7959 38645 7971
rect 38575 7953 38584 7959
rect 38636 7953 38645 7959
rect 38575 7897 38582 7953
rect 38638 7897 38645 7953
rect 40100 8039 40112 8095
rect 40168 8039 40181 8095
rect 40100 8015 40114 8039
rect 40166 8015 40181 8039
rect 40100 7959 40112 8015
rect 40168 7959 40181 8015
rect 40100 7937 40114 7959
rect 40166 7937 40181 7959
rect 40100 7923 40181 7937
rect 36301 7875 36532 7891
rect 38575 7882 38645 7897
rect 36301 7819 36308 7875
rect 36364 7873 36388 7875
rect 36444 7873 36468 7875
rect 36378 7821 36388 7873
rect 36444 7821 36454 7873
rect 36364 7819 36388 7821
rect 36444 7819 36468 7821
rect 36524 7819 36532 7875
rect 36301 7804 36532 7819
rect 33746 7651 33810 7661
rect 25495 7645 33810 7651
rect 25495 7593 33752 7645
rect 33804 7593 33810 7645
rect 25495 7587 33810 7593
rect 33746 7577 33810 7587
rect 38568 7559 38649 7573
rect 38568 7537 38582 7559
rect 38634 7537 38649 7559
rect 38568 7481 38580 7537
rect 38636 7481 38649 7537
rect 38568 7457 38582 7481
rect 38634 7457 38649 7481
rect 38568 7401 38580 7457
rect 38636 7401 38649 7457
rect 38568 7379 38582 7401
rect 38634 7379 38649 7401
rect 38568 7365 38649 7379
rect 40087 7572 40168 7586
rect 40087 7550 40101 7572
rect 40153 7550 40168 7572
rect 40087 7494 40099 7550
rect 40155 7494 40168 7550
rect 40087 7470 40101 7494
rect 40153 7470 40168 7494
rect 40087 7414 40099 7470
rect 40155 7414 40168 7470
rect 40087 7392 40101 7414
rect 40153 7392 40168 7414
rect 40087 7378 40168 7392
rect 36362 7334 36531 7347
rect 36362 7278 36378 7334
rect 36434 7332 36458 7334
rect 36440 7280 36452 7332
rect 36434 7278 36458 7280
rect 36514 7278 36531 7334
rect 36362 7265 36531 7278
rect 35028 7219 35092 7233
rect 35028 7163 35032 7219
rect 35088 7163 35092 7219
rect 35028 7149 35092 7163
rect 42602 7215 45923 7242
rect 42602 7213 42634 7215
rect 42690 7213 42714 7215
rect 42770 7213 42794 7215
rect 42850 7213 42874 7215
rect 42930 7213 42954 7215
rect 43010 7213 43034 7215
rect 43090 7213 43114 7215
rect 43170 7213 43194 7215
rect 43250 7213 43274 7215
rect 43330 7213 43354 7215
rect 43410 7213 43434 7215
rect 43490 7213 43514 7215
rect 43570 7213 43594 7215
rect 43650 7213 43674 7215
rect 43730 7213 43754 7215
rect 43810 7213 43834 7215
rect 43890 7213 43914 7215
rect 43970 7213 43994 7215
rect 44050 7213 44074 7215
rect 44130 7213 44154 7215
rect 44210 7213 44234 7215
rect 44290 7213 44314 7215
rect 44370 7213 44394 7215
rect 44450 7213 44474 7215
rect 44530 7213 44554 7215
rect 44610 7213 44634 7215
rect 44690 7213 44714 7215
rect 44770 7213 44794 7215
rect 44850 7213 44874 7215
rect 44930 7213 44954 7215
rect 45010 7213 45034 7215
rect 45090 7213 45114 7215
rect 45170 7213 45194 7215
rect 45250 7213 45274 7215
rect 45330 7213 45354 7215
rect 45410 7213 45434 7215
rect 45490 7213 45514 7215
rect 45570 7213 45594 7215
rect 45650 7213 45674 7215
rect 45730 7213 45754 7215
rect 45810 7213 45834 7215
rect 45890 7213 45923 7215
rect 42602 7161 42604 7213
rect 42784 7161 42794 7213
rect 42850 7161 42860 7213
rect 43104 7161 43114 7213
rect 43170 7161 43180 7213
rect 43424 7161 43434 7213
rect 43490 7161 43500 7213
rect 43744 7161 43754 7213
rect 43810 7161 43820 7213
rect 44064 7161 44074 7213
rect 44130 7161 44140 7213
rect 44384 7161 44394 7213
rect 44450 7161 44460 7213
rect 44704 7161 44714 7213
rect 44770 7161 44780 7213
rect 45024 7161 45034 7213
rect 45090 7161 45100 7213
rect 45344 7161 45354 7213
rect 45410 7161 45420 7213
rect 45664 7161 45674 7213
rect 45730 7161 45740 7213
rect 45920 7161 45923 7213
rect 42602 7159 42634 7161
rect 42690 7159 42714 7161
rect 42770 7159 42794 7161
rect 42850 7159 42874 7161
rect 42930 7159 42954 7161
rect 43010 7159 43034 7161
rect 43090 7159 43114 7161
rect 43170 7159 43194 7161
rect 43250 7159 43274 7161
rect 43330 7159 43354 7161
rect 43410 7159 43434 7161
rect 43490 7159 43514 7161
rect 43570 7159 43594 7161
rect 43650 7159 43674 7161
rect 43730 7159 43754 7161
rect 43810 7159 43834 7161
rect 43890 7159 43914 7161
rect 43970 7159 43994 7161
rect 44050 7159 44074 7161
rect 44130 7159 44154 7161
rect 44210 7159 44234 7161
rect 44290 7159 44314 7161
rect 44370 7159 44394 7161
rect 44450 7159 44474 7161
rect 44530 7159 44554 7161
rect 44610 7159 44634 7161
rect 44690 7159 44714 7161
rect 44770 7159 44794 7161
rect 44850 7159 44874 7161
rect 44930 7159 44954 7161
rect 45010 7159 45034 7161
rect 45090 7159 45114 7161
rect 45170 7159 45194 7161
rect 45250 7159 45274 7161
rect 45330 7159 45354 7161
rect 45410 7159 45434 7161
rect 45490 7159 45514 7161
rect 45570 7159 45594 7161
rect 45650 7159 45674 7161
rect 45730 7159 45754 7161
rect 45810 7159 45834 7161
rect 45890 7159 45923 7161
rect 42602 7133 45923 7159
rect 35027 6950 35091 6964
rect 35027 6894 35031 6950
rect 35087 6894 35091 6950
rect 35027 6880 35091 6894
rect 36352 6786 36437 6805
rect 36352 6730 36366 6786
rect 36422 6730 36437 6786
rect 36352 6711 36437 6730
rect 40092 6781 40173 6795
rect 40092 6759 40106 6781
rect 40158 6759 40173 6781
rect 38571 6702 38649 6717
rect 38571 6672 38584 6702
rect 38636 6672 38649 6702
rect 38571 6616 38582 6672
rect 38638 6616 38649 6672
rect 38571 6586 38584 6616
rect 38636 6586 38649 6616
rect 40092 6703 40104 6759
rect 40160 6703 40173 6759
rect 40092 6679 40106 6703
rect 40158 6679 40173 6703
rect 40092 6623 40104 6679
rect 40160 6623 40173 6679
rect 40092 6601 40106 6623
rect 40158 6601 40173 6623
rect 40092 6587 40173 6601
rect 38571 6572 38649 6586
rect 24544 6312 24608 6322
rect 33734 6312 33798 6322
rect 24544 6306 33798 6312
rect 24544 6254 24550 6306
rect 24602 6254 33740 6306
rect 33792 6254 33798 6306
rect 24544 6248 33798 6254
rect 24544 6238 24608 6248
rect 33734 6238 33798 6248
rect 36971 6245 37067 6275
rect 36971 6189 36991 6245
rect 37047 6189 37067 6245
rect 36971 6159 37067 6189
rect 38563 6228 38644 6242
rect 38563 6206 38577 6228
rect 38629 6206 38644 6228
rect 38563 6150 38575 6206
rect 38631 6150 38644 6206
rect 38563 6126 38577 6150
rect 38629 6126 38644 6150
rect 38563 6070 38575 6126
rect 38631 6070 38644 6126
rect 38563 6048 38577 6070
rect 38629 6048 38644 6070
rect 38563 6034 38644 6048
rect 40092 6225 40173 6239
rect 40092 6203 40106 6225
rect 40158 6203 40173 6225
rect 40092 6147 40104 6203
rect 40160 6147 40173 6203
rect 40092 6123 40106 6147
rect 40158 6123 40173 6147
rect 40092 6067 40104 6123
rect 40160 6067 40173 6123
rect 40092 6045 40106 6067
rect 40158 6045 40173 6067
rect 40092 6031 40173 6045
rect 35027 5881 35091 5895
rect 35027 5825 35031 5881
rect 35087 5825 35091 5881
rect 35027 5811 35091 5825
rect 47473 5790 47709 5810
rect 35970 5703 36149 5717
rect 35970 5647 35991 5703
rect 36047 5701 36071 5703
rect 36053 5649 36065 5701
rect 36047 5647 36071 5649
rect 36127 5647 36149 5703
rect 35970 5634 36149 5647
rect 47473 5574 47483 5790
rect 47699 5574 47709 5790
rect 35024 5558 35088 5572
rect 35024 5502 35028 5558
rect 35084 5502 35088 5558
rect 47473 5554 47709 5574
rect 35024 5488 35088 5502
rect 40109 5401 40190 5415
rect 40109 5379 40123 5401
rect 40175 5379 40190 5401
rect 38574 5312 38648 5332
rect 38574 5282 38585 5312
rect 38637 5282 38648 5312
rect 38574 5226 38583 5282
rect 38639 5226 38648 5282
rect 38574 5196 38585 5226
rect 38637 5196 38648 5226
rect 40109 5323 40121 5379
rect 40177 5323 40190 5379
rect 40109 5299 40123 5323
rect 40175 5299 40190 5323
rect 40109 5243 40121 5299
rect 40177 5243 40190 5299
rect 40109 5221 40123 5243
rect 40175 5221 40190 5243
rect 40109 5207 40190 5221
rect 38574 5177 38648 5196
rect 36514 5155 36734 5172
rect 36514 5099 36516 5155
rect 36572 5153 36596 5155
rect 36652 5153 36676 5155
rect 36586 5101 36596 5153
rect 36652 5101 36662 5153
rect 36572 5099 36596 5101
rect 36652 5099 36676 5101
rect 36732 5099 36734 5155
rect 36514 5082 36734 5099
rect 23208 4916 23261 4926
rect 33742 4916 33795 4926
rect 23208 4915 33795 4916
rect 23260 4863 33742 4915
rect 33794 4863 33795 4915
rect 23208 4853 23261 4863
rect 33742 4853 33795 4863
rect 38562 4875 38643 4889
rect 38562 4853 38576 4875
rect 38628 4853 38643 4875
rect 38562 4797 38574 4853
rect 38630 4797 38643 4853
rect 38562 4773 38576 4797
rect 38628 4773 38643 4797
rect 38562 4717 38574 4773
rect 38630 4717 38643 4773
rect 38562 4695 38576 4717
rect 38628 4695 38643 4717
rect 38562 4681 38643 4695
rect 40092 4853 40173 4867
rect 40092 4831 40106 4853
rect 40158 4831 40173 4853
rect 40092 4775 40104 4831
rect 40160 4775 40173 4831
rect 40092 4751 40106 4775
rect 40158 4751 40173 4775
rect 40092 4695 40104 4751
rect 40160 4695 40173 4751
rect 40092 4673 40106 4695
rect 40158 4673 40173 4695
rect 40092 4659 40173 4673
rect 36364 4612 36509 4623
rect 36364 4556 36368 4612
rect 36424 4610 36448 4612
rect 36430 4558 36442 4610
rect 36424 4556 36448 4558
rect 36504 4556 36509 4612
rect 36364 4545 36509 4556
rect 35035 4488 35099 4502
rect 35035 4432 35039 4488
rect 35095 4432 35099 4488
rect 35035 4418 35099 4432
rect 42599 4216 45959 4243
rect 35024 4183 35088 4197
rect 35024 4127 35028 4183
rect 35084 4127 35088 4183
rect 42599 4160 42611 4216
rect 42667 4214 42691 4216
rect 42747 4214 42771 4216
rect 42827 4214 42851 4216
rect 42907 4214 42931 4216
rect 42987 4214 43011 4216
rect 43067 4214 43091 4216
rect 43147 4214 43171 4216
rect 43227 4214 43251 4216
rect 43307 4214 43331 4216
rect 43387 4214 43411 4216
rect 43467 4214 43491 4216
rect 43547 4214 43571 4216
rect 43627 4214 43651 4216
rect 43707 4214 43731 4216
rect 43787 4214 43811 4216
rect 43867 4214 43891 4216
rect 43947 4214 43971 4216
rect 44027 4214 44051 4216
rect 44107 4214 44131 4216
rect 44187 4214 44211 4216
rect 44267 4214 44291 4216
rect 44347 4214 44371 4216
rect 44427 4214 44451 4216
rect 44507 4214 44531 4216
rect 44587 4214 44611 4216
rect 44667 4214 44691 4216
rect 44747 4214 44771 4216
rect 44827 4214 44851 4216
rect 44907 4214 44931 4216
rect 44987 4214 45011 4216
rect 45067 4214 45091 4216
rect 45147 4214 45171 4216
rect 45227 4214 45251 4216
rect 45307 4214 45331 4216
rect 45387 4214 45411 4216
rect 45467 4214 45491 4216
rect 45547 4214 45571 4216
rect 45627 4214 45651 4216
rect 45707 4214 45731 4216
rect 45787 4214 45811 4216
rect 45867 4214 45891 4216
rect 42673 4162 42685 4214
rect 42747 4162 42749 4214
rect 42929 4162 42931 4214
rect 42993 4162 43005 4214
rect 43067 4162 43069 4214
rect 43249 4162 43251 4214
rect 43313 4162 43325 4214
rect 43387 4162 43389 4214
rect 43569 4162 43571 4214
rect 43633 4162 43645 4214
rect 43707 4162 43709 4214
rect 43889 4162 43891 4214
rect 43953 4162 43965 4214
rect 44027 4162 44029 4214
rect 44209 4162 44211 4214
rect 44273 4162 44285 4214
rect 44347 4162 44349 4214
rect 44529 4162 44531 4214
rect 44593 4162 44605 4214
rect 44667 4162 44669 4214
rect 44849 4162 44851 4214
rect 44913 4162 44925 4214
rect 44987 4162 44989 4214
rect 45169 4162 45171 4214
rect 45233 4162 45245 4214
rect 45307 4162 45309 4214
rect 45489 4162 45491 4214
rect 45553 4162 45565 4214
rect 45627 4162 45629 4214
rect 45809 4162 45811 4214
rect 45873 4162 45885 4214
rect 42667 4160 42691 4162
rect 42747 4160 42771 4162
rect 42827 4160 42851 4162
rect 42907 4160 42931 4162
rect 42987 4160 43011 4162
rect 43067 4160 43091 4162
rect 43147 4160 43171 4162
rect 43227 4160 43251 4162
rect 43307 4160 43331 4162
rect 43387 4160 43411 4162
rect 43467 4160 43491 4162
rect 43547 4160 43571 4162
rect 43627 4160 43651 4162
rect 43707 4160 43731 4162
rect 43787 4160 43811 4162
rect 43867 4160 43891 4162
rect 43947 4160 43971 4162
rect 44027 4160 44051 4162
rect 44107 4160 44131 4162
rect 44187 4160 44211 4162
rect 44267 4160 44291 4162
rect 44347 4160 44371 4162
rect 44427 4160 44451 4162
rect 44507 4160 44531 4162
rect 44587 4160 44611 4162
rect 44667 4160 44691 4162
rect 44747 4160 44771 4162
rect 44827 4160 44851 4162
rect 44907 4160 44931 4162
rect 44987 4160 45011 4162
rect 45067 4160 45091 4162
rect 45147 4160 45171 4162
rect 45227 4160 45251 4162
rect 45307 4160 45331 4162
rect 45387 4160 45411 4162
rect 45467 4160 45491 4162
rect 45547 4160 45571 4162
rect 45627 4160 45651 4162
rect 45707 4160 45731 4162
rect 45787 4160 45811 4162
rect 45867 4160 45891 4162
rect 45947 4160 45959 4216
rect 42599 4134 45959 4160
rect 35024 4113 35088 4127
rect 36972 4069 37068 4099
rect 36972 4013 36992 4069
rect 37048 4013 37068 4069
rect 36972 3983 37068 4013
rect 40099 4022 40180 4036
rect 40099 4000 40113 4022
rect 40165 4000 40180 4022
rect 40099 3944 40111 4000
rect 40167 3944 40180 4000
rect 38572 3925 38651 3944
rect 38572 3869 38583 3925
rect 38639 3869 38651 3925
rect 38572 3863 38585 3869
rect 38637 3863 38651 3869
rect 38572 3851 38651 3863
rect 38572 3845 38585 3851
rect 38637 3845 38651 3851
rect 38572 3789 38583 3845
rect 38639 3789 38651 3845
rect 40099 3920 40113 3944
rect 40165 3920 40180 3944
rect 40099 3864 40111 3920
rect 40167 3864 40180 3920
rect 40099 3842 40113 3864
rect 40165 3842 40180 3864
rect 40099 3828 40180 3842
rect 38572 3771 38651 3789
rect -279 3727 -227 3737
rect 36359 3523 36486 3541
rect 36359 3521 36394 3523
rect 36450 3521 36486 3523
rect 36359 3469 36364 3521
rect 36480 3469 36486 3521
rect 36359 3467 36394 3469
rect 36450 3467 36486 3469
rect 36359 3449 36486 3467
rect 38565 3475 38646 3489
rect 38565 3453 38579 3475
rect 38631 3453 38646 3475
rect 38565 3397 38577 3453
rect 38633 3397 38646 3453
rect 38565 3373 38579 3397
rect 38631 3373 38646 3397
rect 38565 3317 38577 3373
rect 38633 3317 38646 3373
rect 38565 3295 38579 3317
rect 38631 3295 38646 3317
rect 38565 3281 38646 3295
rect 40089 3469 40170 3483
rect 40089 3447 40103 3469
rect 40155 3447 40170 3469
rect 40089 3391 40101 3447
rect 40157 3391 40170 3447
rect 40089 3367 40103 3391
rect 40155 3367 40170 3391
rect 40089 3311 40101 3367
rect 40157 3311 40170 3367
rect 40089 3289 40103 3311
rect 40155 3289 40170 3311
rect 40089 3275 40170 3289
rect 35031 3118 35095 3132
rect 35031 3062 35035 3118
rect 35091 3062 35095 3118
rect 35031 3048 35095 3062
rect 3670 2688 5404 2741
rect 5351 2407 5404 2688
rect 23432 2407 23485 2417
rect 5351 2406 23485 2407
rect 5351 2354 23432 2406
rect 23484 2354 23485 2406
rect 23432 2344 23485 2354
rect 36066 2210 36130 2224
rect 35842 2156 36070 2210
rect 35489 1587 35553 1601
rect 35489 1531 35493 1587
rect 35549 1531 35553 1587
rect 35489 1517 35553 1531
rect 35842 1460 35896 2156
rect 36066 2154 36070 2156
rect 36126 2154 36130 2210
rect 36066 2140 36130 2154
rect 36631 1525 36695 1539
rect 35982 1473 36635 1525
rect 36631 1469 36635 1473
rect 36691 1469 36695 1525
rect 36631 1455 36695 1469
rect 35024 1339 35088 1353
rect 35024 1283 35028 1339
rect 35084 1283 35088 1339
rect 35024 1269 35088 1283
rect 40100 1177 40181 1191
rect 40100 1155 40114 1177
rect 40166 1155 40181 1177
rect 22589 1097 22642 1107
rect 18808 1096 22642 1097
rect 18808 1044 22589 1096
rect 22641 1044 22642 1096
rect 22589 1034 22642 1044
rect 38575 1093 38645 1108
rect 38575 1037 38582 1093
rect 38638 1037 38645 1093
rect 38575 1031 38584 1037
rect 38636 1031 38645 1037
rect 38575 1019 38645 1031
rect 38575 1013 38584 1019
rect 38636 1013 38645 1019
rect 38575 957 38582 1013
rect 38638 957 38645 1013
rect 40100 1099 40112 1155
rect 40168 1099 40181 1155
rect 40100 1075 40114 1099
rect 40166 1075 40181 1099
rect 40100 1019 40112 1075
rect 40168 1019 40181 1075
rect 40100 997 40114 1019
rect 40166 997 40181 1019
rect 40100 983 40181 997
rect 36301 935 36532 951
rect 38575 942 38645 957
rect 36301 879 36308 935
rect 36364 933 36388 935
rect 36444 933 36468 935
rect 36378 881 36388 933
rect 36444 881 36454 933
rect 36364 879 36388 881
rect 36444 879 36468 881
rect 36524 879 36532 935
rect 36301 864 36532 879
rect 26001 716 26076 726
rect 33730 721 33805 726
rect 33730 716 33810 721
rect 26001 704 33810 716
rect 26001 652 26012 704
rect 26064 652 33741 704
rect 33793 652 33810 704
rect 26001 641 33810 652
rect 26001 631 26076 641
rect 33730 637 33810 641
rect 33730 631 33805 637
rect 38568 619 38649 633
rect 38568 597 38582 619
rect 38634 597 38649 619
rect 38568 541 38580 597
rect 38636 541 38649 597
rect 38568 517 38582 541
rect 38634 517 38649 541
rect 38568 461 38580 517
rect 38636 461 38649 517
rect 38568 439 38582 461
rect 38634 439 38649 461
rect 38568 425 38649 439
rect 40087 632 40168 646
rect 40087 610 40101 632
rect 40153 610 40168 632
rect 40087 554 40099 610
rect 40155 554 40168 610
rect 40087 530 40101 554
rect 40153 530 40168 554
rect 40087 474 40099 530
rect 40155 474 40168 530
rect 40087 452 40101 474
rect 40153 452 40168 474
rect 40087 438 40168 452
rect 36362 394 36531 407
rect 36362 338 36378 394
rect 36434 392 36458 394
rect 36440 340 36452 392
rect 36434 338 36458 340
rect 36514 338 36531 394
rect 36362 325 36531 338
rect 35028 279 35092 293
rect 322 217 21107 242
rect 322 81 326 217
rect 21102 81 21107 217
rect 35028 223 35032 279
rect 35088 223 35092 279
rect 35028 209 35092 223
rect 42599 282 45930 319
rect 42599 280 42636 282
rect 42692 280 42716 282
rect 42772 280 42796 282
rect 42852 280 42876 282
rect 42932 280 42956 282
rect 43012 280 43036 282
rect 43092 280 43116 282
rect 43172 280 43196 282
rect 43252 280 43276 282
rect 43332 280 43356 282
rect 43412 280 43436 282
rect 43492 280 43516 282
rect 43572 280 43596 282
rect 43652 280 43676 282
rect 43732 280 43756 282
rect 43812 280 43836 282
rect 43892 280 43916 282
rect 43972 280 43996 282
rect 44052 280 44076 282
rect 44132 280 44156 282
rect 44212 280 44236 282
rect 44292 280 44316 282
rect 44372 280 44396 282
rect 44452 280 44476 282
rect 44532 280 44556 282
rect 44612 280 44636 282
rect 44692 280 44716 282
rect 44772 280 44796 282
rect 44852 280 44876 282
rect 44932 280 44956 282
rect 45012 280 45036 282
rect 45092 280 45116 282
rect 45172 280 45196 282
rect 45252 280 45276 282
rect 45332 280 45356 282
rect 45412 280 45436 282
rect 45492 280 45516 282
rect 45572 280 45596 282
rect 45652 280 45676 282
rect 45732 280 45756 282
rect 45812 280 45836 282
rect 45892 280 45930 282
rect 42599 228 42606 280
rect 42786 228 42796 280
rect 42852 228 42862 280
rect 43106 228 43116 280
rect 43172 228 43182 280
rect 43426 228 43436 280
rect 43492 228 43502 280
rect 43746 228 43756 280
rect 43812 228 43822 280
rect 44066 228 44076 280
rect 44132 228 44142 280
rect 44386 228 44396 280
rect 44452 228 44462 280
rect 44706 228 44716 280
rect 44772 228 44782 280
rect 45026 228 45036 280
rect 45092 228 45102 280
rect 45346 228 45356 280
rect 45412 228 45422 280
rect 45666 228 45676 280
rect 45732 228 45742 280
rect 45922 228 45930 280
rect 42599 226 42636 228
rect 42692 226 42716 228
rect 42772 226 42796 228
rect 42852 226 42876 228
rect 42932 226 42956 228
rect 43012 226 43036 228
rect 43092 226 43116 228
rect 43172 226 43196 228
rect 43252 226 43276 228
rect 43332 226 43356 228
rect 43412 226 43436 228
rect 43492 226 43516 228
rect 43572 226 43596 228
rect 43652 226 43676 228
rect 43732 226 43756 228
rect 43812 226 43836 228
rect 43892 226 43916 228
rect 43972 226 43996 228
rect 44052 226 44076 228
rect 44132 226 44156 228
rect 44212 226 44236 228
rect 44292 226 44316 228
rect 44372 226 44396 228
rect 44452 226 44476 228
rect 44532 226 44556 228
rect 44612 226 44636 228
rect 44692 226 44716 228
rect 44772 226 44796 228
rect 44852 226 44876 228
rect 44932 226 44956 228
rect 45012 226 45036 228
rect 45092 226 45116 228
rect 45172 226 45196 228
rect 45252 226 45276 228
rect 45332 226 45356 228
rect 45412 226 45436 228
rect 45492 226 45516 228
rect 45572 226 45596 228
rect 45652 226 45676 228
rect 45732 226 45756 228
rect 45812 226 45836 228
rect 45892 226 45930 228
rect 42599 189 45930 226
rect 322 57 21107 81
rect 35027 10 35091 24
rect 35027 -46 35031 10
rect 35087 -46 35091 10
rect 35027 -60 35091 -46
rect 36352 -154 36437 -135
rect 36352 -210 36366 -154
rect 36422 -210 36437 -154
rect 36352 -229 36437 -210
rect 40092 -159 40173 -145
rect 40092 -181 40106 -159
rect 40158 -181 40173 -159
rect 38571 -238 38649 -223
rect 38571 -268 38584 -238
rect 38636 -268 38649 -238
rect 38571 -324 38582 -268
rect 38638 -324 38649 -268
rect 38571 -354 38584 -324
rect 38636 -354 38649 -324
rect 40092 -237 40104 -181
rect 40160 -237 40173 -181
rect 40092 -261 40106 -237
rect 40158 -261 40173 -237
rect 40092 -317 40104 -261
rect 40160 -317 40173 -261
rect 40092 -339 40106 -317
rect 40158 -339 40173 -317
rect 40092 -353 40173 -339
rect 38571 -368 38649 -354
rect 33734 -628 33798 -618
rect 23417 -635 33798 -628
rect 23417 -641 33741 -635
rect 23417 -693 23432 -641
rect 23484 -687 33741 -641
rect 33793 -687 33798 -635
rect 23484 -693 33798 -687
rect 23432 -703 23485 -693
rect 33734 -702 33798 -693
rect 36971 -695 37067 -665
rect 33741 -703 33794 -702
rect 36971 -751 36991 -695
rect 37047 -751 37067 -695
rect 36971 -781 37067 -751
rect 38563 -712 38644 -698
rect 38563 -734 38577 -712
rect 38629 -734 38644 -712
rect 38563 -790 38575 -734
rect 38631 -790 38644 -734
rect 38563 -814 38577 -790
rect 38629 -814 38644 -790
rect 38563 -870 38575 -814
rect 38631 -870 38644 -814
rect 38563 -892 38577 -870
rect 38629 -892 38644 -870
rect 38563 -906 38644 -892
rect 40092 -715 40173 -701
rect 40092 -737 40106 -715
rect 40158 -737 40173 -715
rect 40092 -793 40104 -737
rect 40160 -793 40173 -737
rect 40092 -817 40106 -793
rect 40158 -817 40173 -793
rect 40092 -873 40104 -817
rect 40160 -873 40173 -817
rect 40092 -895 40106 -873
rect 40158 -895 40173 -873
rect 40092 -909 40173 -895
rect 35027 -1059 35091 -1045
rect 35027 -1115 35031 -1059
rect 35087 -1115 35091 -1059
rect 35027 -1129 35091 -1115
rect 47489 -1150 47725 -1130
rect 35970 -1237 36149 -1223
rect 35970 -1293 35991 -1237
rect 36047 -1239 36071 -1237
rect 36053 -1291 36065 -1239
rect 36047 -1293 36071 -1291
rect 36127 -1293 36149 -1237
rect 35970 -1306 36149 -1293
rect 47489 -1366 47499 -1150
rect 47715 -1366 47725 -1150
rect 35024 -1382 35088 -1368
rect 35024 -1438 35028 -1382
rect 35084 -1438 35088 -1382
rect 47489 -1386 47725 -1366
rect 35024 -1452 35088 -1438
rect 40109 -1539 40190 -1525
rect 40109 -1561 40123 -1539
rect 40175 -1561 40190 -1539
rect 38574 -1628 38648 -1608
rect 38574 -1658 38585 -1628
rect 38637 -1658 38648 -1628
rect 38574 -1714 38583 -1658
rect 38639 -1714 38648 -1658
rect 38574 -1744 38585 -1714
rect 38637 -1744 38648 -1714
rect 40109 -1617 40121 -1561
rect 40177 -1617 40190 -1561
rect 40109 -1641 40123 -1617
rect 40175 -1641 40190 -1617
rect 40109 -1697 40121 -1641
rect 40177 -1697 40190 -1641
rect 40109 -1719 40123 -1697
rect 40175 -1719 40190 -1697
rect 40109 -1733 40190 -1719
rect 38574 -1763 38648 -1744
rect 36514 -1785 36734 -1768
rect 36514 -1841 36516 -1785
rect 36572 -1787 36596 -1785
rect 36652 -1787 36676 -1785
rect 36586 -1839 36596 -1787
rect 36652 -1839 36662 -1787
rect 36572 -1841 36596 -1839
rect 36652 -1841 36676 -1839
rect 36732 -1841 36734 -1785
rect 36514 -1858 36734 -1841
rect 22589 -2017 22643 -2007
rect 33746 -2017 33806 -2007
rect 22587 -2018 33806 -2017
rect 22587 -2070 22590 -2018
rect 22642 -2021 33806 -2018
rect 22642 -2070 33750 -2021
rect 22587 -2073 33750 -2070
rect 33802 -2073 33806 -2021
rect 22587 -2077 33806 -2073
rect 22589 -2080 22643 -2077
rect 33746 -2087 33806 -2077
rect 38562 -2065 38643 -2051
rect 38562 -2087 38576 -2065
rect 38628 -2087 38643 -2065
rect 38562 -2143 38574 -2087
rect 38630 -2143 38643 -2087
rect 38562 -2167 38576 -2143
rect 38628 -2167 38643 -2143
rect 38562 -2223 38574 -2167
rect 38630 -2223 38643 -2167
rect 38562 -2245 38576 -2223
rect 38628 -2245 38643 -2223
rect 38562 -2259 38643 -2245
rect 40092 -2087 40173 -2073
rect 40092 -2109 40106 -2087
rect 40158 -2109 40173 -2087
rect 40092 -2165 40104 -2109
rect 40160 -2165 40173 -2109
rect 40092 -2189 40106 -2165
rect 40158 -2189 40173 -2165
rect 40092 -2245 40104 -2189
rect 40160 -2245 40173 -2189
rect 40092 -2267 40106 -2245
rect 40158 -2267 40173 -2245
rect 40092 -2281 40173 -2267
rect 36364 -2328 36509 -2317
rect 36364 -2384 36368 -2328
rect 36424 -2330 36448 -2328
rect 36430 -2382 36442 -2330
rect 36424 -2384 36448 -2382
rect 36504 -2384 36509 -2328
rect 36364 -2395 36509 -2384
rect 35035 -2452 35099 -2438
rect 35035 -2508 35039 -2452
rect 35095 -2508 35099 -2452
rect 35035 -2522 35099 -2508
rect 42587 -2724 45933 -2698
rect 35024 -2757 35088 -2743
rect 35024 -2813 35028 -2757
rect 35084 -2813 35088 -2757
rect 42587 -2780 42592 -2724
rect 42648 -2726 42672 -2724
rect 42728 -2726 42752 -2724
rect 42808 -2726 42832 -2724
rect 42888 -2726 42912 -2724
rect 42968 -2726 42992 -2724
rect 43048 -2726 43072 -2724
rect 43128 -2726 43152 -2724
rect 43208 -2726 43232 -2724
rect 43288 -2726 43312 -2724
rect 43368 -2726 43392 -2724
rect 43448 -2726 43472 -2724
rect 43528 -2726 43552 -2724
rect 43608 -2726 43632 -2724
rect 43688 -2726 43712 -2724
rect 43768 -2726 43792 -2724
rect 43848 -2726 43872 -2724
rect 43928 -2726 43952 -2724
rect 44008 -2726 44032 -2724
rect 44088 -2726 44112 -2724
rect 44168 -2726 44192 -2724
rect 44248 -2726 44272 -2724
rect 44328 -2726 44352 -2724
rect 44408 -2726 44432 -2724
rect 44488 -2726 44512 -2724
rect 44568 -2726 44592 -2724
rect 44648 -2726 44672 -2724
rect 44728 -2726 44752 -2724
rect 44808 -2726 44832 -2724
rect 44888 -2726 44912 -2724
rect 44968 -2726 44992 -2724
rect 45048 -2726 45072 -2724
rect 45128 -2726 45152 -2724
rect 45208 -2726 45232 -2724
rect 45288 -2726 45312 -2724
rect 45368 -2726 45392 -2724
rect 45448 -2726 45472 -2724
rect 45528 -2726 45552 -2724
rect 45608 -2726 45632 -2724
rect 45688 -2726 45712 -2724
rect 45768 -2726 45792 -2724
rect 45848 -2726 45872 -2724
rect 42654 -2778 42666 -2726
rect 42728 -2778 42730 -2726
rect 42910 -2778 42912 -2726
rect 42974 -2778 42986 -2726
rect 43048 -2778 43050 -2726
rect 43230 -2778 43232 -2726
rect 43294 -2778 43306 -2726
rect 43368 -2778 43370 -2726
rect 43550 -2778 43552 -2726
rect 43614 -2778 43626 -2726
rect 43688 -2778 43690 -2726
rect 43870 -2778 43872 -2726
rect 43934 -2778 43946 -2726
rect 44008 -2778 44010 -2726
rect 44190 -2778 44192 -2726
rect 44254 -2778 44266 -2726
rect 44328 -2778 44330 -2726
rect 44510 -2778 44512 -2726
rect 44574 -2778 44586 -2726
rect 44648 -2778 44650 -2726
rect 44830 -2778 44832 -2726
rect 44894 -2778 44906 -2726
rect 44968 -2778 44970 -2726
rect 45150 -2778 45152 -2726
rect 45214 -2778 45226 -2726
rect 45288 -2778 45290 -2726
rect 45470 -2778 45472 -2726
rect 45534 -2778 45546 -2726
rect 45608 -2778 45610 -2726
rect 45790 -2778 45792 -2726
rect 45854 -2778 45866 -2726
rect 42648 -2780 42672 -2778
rect 42728 -2780 42752 -2778
rect 42808 -2780 42832 -2778
rect 42888 -2780 42912 -2778
rect 42968 -2780 42992 -2778
rect 43048 -2780 43072 -2778
rect 43128 -2780 43152 -2778
rect 43208 -2780 43232 -2778
rect 43288 -2780 43312 -2778
rect 43368 -2780 43392 -2778
rect 43448 -2780 43472 -2778
rect 43528 -2780 43552 -2778
rect 43608 -2780 43632 -2778
rect 43688 -2780 43712 -2778
rect 43768 -2780 43792 -2778
rect 43848 -2780 43872 -2778
rect 43928 -2780 43952 -2778
rect 44008 -2780 44032 -2778
rect 44088 -2780 44112 -2778
rect 44168 -2780 44192 -2778
rect 44248 -2780 44272 -2778
rect 44328 -2780 44352 -2778
rect 44408 -2780 44432 -2778
rect 44488 -2780 44512 -2778
rect 44568 -2780 44592 -2778
rect 44648 -2780 44672 -2778
rect 44728 -2780 44752 -2778
rect 44808 -2780 44832 -2778
rect 44888 -2780 44912 -2778
rect 44968 -2780 44992 -2778
rect 45048 -2780 45072 -2778
rect 45128 -2780 45152 -2778
rect 45208 -2780 45232 -2778
rect 45288 -2780 45312 -2778
rect 45368 -2780 45392 -2778
rect 45448 -2780 45472 -2778
rect 45528 -2780 45552 -2778
rect 45608 -2780 45632 -2778
rect 45688 -2780 45712 -2778
rect 45768 -2780 45792 -2778
rect 45848 -2780 45872 -2778
rect 45928 -2780 45933 -2724
rect 42587 -2806 45933 -2780
rect 35024 -2827 35088 -2813
rect 36972 -2871 37068 -2841
rect 36972 -2927 36992 -2871
rect 37048 -2927 37068 -2871
rect 36972 -2957 37068 -2927
rect 40099 -2918 40180 -2904
rect 40099 -2940 40113 -2918
rect 40165 -2940 40180 -2918
rect 40099 -2996 40111 -2940
rect 40167 -2996 40180 -2940
rect 38572 -3015 38651 -2996
rect 38572 -3071 38583 -3015
rect 38639 -3071 38651 -3015
rect 38572 -3077 38585 -3071
rect 38637 -3077 38651 -3071
rect 38572 -3089 38651 -3077
rect 38572 -3095 38585 -3089
rect 38637 -3095 38651 -3089
rect 38572 -3151 38583 -3095
rect 38639 -3151 38651 -3095
rect 40099 -3020 40113 -2996
rect 40165 -3020 40180 -2996
rect 40099 -3076 40111 -3020
rect 40167 -3076 40180 -3020
rect 40099 -3098 40113 -3076
rect 40165 -3098 40180 -3076
rect 40099 -3112 40180 -3098
rect 38572 -3169 38651 -3151
rect 36359 -3417 36486 -3399
rect 36359 -3419 36394 -3417
rect 36450 -3419 36486 -3417
rect 36359 -3471 36364 -3419
rect 36480 -3471 36486 -3419
rect 36359 -3473 36394 -3471
rect 36450 -3473 36486 -3471
rect 36359 -3491 36486 -3473
rect 38565 -3465 38646 -3451
rect 38565 -3487 38579 -3465
rect 38631 -3487 38646 -3465
rect 38565 -3543 38577 -3487
rect 38633 -3543 38646 -3487
rect 38565 -3567 38579 -3543
rect 38631 -3567 38646 -3543
rect 38565 -3623 38577 -3567
rect 38633 -3623 38646 -3567
rect 38565 -3645 38579 -3623
rect 38631 -3645 38646 -3623
rect 38565 -3659 38646 -3645
rect 40089 -3471 40170 -3457
rect 40089 -3493 40103 -3471
rect 40155 -3493 40170 -3471
rect 40089 -3549 40101 -3493
rect 40157 -3549 40170 -3493
rect 40089 -3573 40103 -3549
rect 40155 -3573 40170 -3549
rect 40089 -3629 40101 -3573
rect 40157 -3629 40170 -3573
rect 40089 -3651 40103 -3629
rect 40155 -3651 40170 -3629
rect 40089 -3665 40170 -3651
rect 35031 -3822 35095 -3808
rect 35031 -3878 35035 -3822
rect 35091 -3878 35095 -3822
rect 35031 -3892 35095 -3878
rect -3595 -6848 -3503 -6812
rect -3595 -6904 -3577 -6848
rect -3521 -6904 -3503 -6848
rect -3595 -6914 -3503 -6904
rect -3595 -6928 -3575 -6914
rect -3523 -6928 -3503 -6914
rect -3595 -6984 -3577 -6928
rect -3521 -6984 -3503 -6928
rect -3595 -7008 -3575 -6984
rect -3523 -7008 -3503 -6984
rect -3595 -7064 -3577 -7008
rect -3521 -7064 -3503 -7008
rect -3595 -7088 -3575 -7064
rect -3523 -7088 -3503 -7064
rect -3595 -7144 -3577 -7088
rect -3521 -7144 -3503 -7088
rect -3595 -7158 -3575 -7144
rect -3523 -7158 -3503 -7144
rect -3595 -7168 -3503 -7158
rect -3595 -7224 -3577 -7168
rect -3521 -7224 -3503 -7168
rect -3595 -7234 -3503 -7224
rect -3595 -7248 -3575 -7234
rect -3523 -7248 -3503 -7234
rect -3595 -7304 -3577 -7248
rect -3521 -7304 -3503 -7248
rect -3595 -7328 -3575 -7304
rect -3523 -7328 -3503 -7304
rect -3595 -7384 -3577 -7328
rect -3521 -7384 -3503 -7328
rect -3595 -7408 -3575 -7384
rect -3523 -7408 -3503 -7384
rect -3595 -7464 -3577 -7408
rect -3521 -7464 -3503 -7408
rect -3595 -7478 -3575 -7464
rect -3523 -7478 -3503 -7464
rect -3595 -7488 -3503 -7478
rect -3595 -7544 -3577 -7488
rect -3521 -7544 -3503 -7488
rect -3595 -7554 -3503 -7544
rect -3595 -7568 -3575 -7554
rect -3523 -7568 -3503 -7554
rect -3595 -7624 -3577 -7568
rect -3521 -7624 -3503 -7568
rect -3595 -7648 -3575 -7624
rect -3523 -7648 -3503 -7624
rect -3595 -7704 -3577 -7648
rect -3521 -7704 -3503 -7648
rect -3595 -7728 -3575 -7704
rect -3523 -7728 -3503 -7704
rect -3595 -7784 -3577 -7728
rect -3521 -7784 -3503 -7728
rect -3595 -7798 -3575 -7784
rect -3523 -7798 -3503 -7784
rect -3595 -7808 -3503 -7798
rect -3595 -7864 -3577 -7808
rect -3521 -7864 -3503 -7808
rect -3595 -7874 -3503 -7864
rect -3595 -7888 -3575 -7874
rect -3523 -7888 -3503 -7874
rect -3595 -7944 -3577 -7888
rect -3521 -7944 -3503 -7888
rect -3595 -7968 -3575 -7944
rect -3523 -7968 -3503 -7944
rect -3595 -8024 -3577 -7968
rect -3521 -8024 -3503 -7968
rect -3595 -8048 -3575 -8024
rect -3523 -8048 -3503 -8024
rect -3595 -8104 -3577 -8048
rect -3521 -8104 -3503 -8048
rect -3595 -8118 -3575 -8104
rect -3523 -8118 -3503 -8104
rect -3595 -8128 -3503 -8118
rect -3595 -8184 -3577 -8128
rect -3521 -8184 -3503 -8128
rect -3595 -8194 -3503 -8184
rect -3595 -8208 -3575 -8194
rect -3523 -8208 -3503 -8194
rect -3595 -8264 -3577 -8208
rect -3521 -8264 -3503 -8208
rect -3595 -8288 -3575 -8264
rect -3523 -8288 -3503 -8264
rect -3595 -8344 -3577 -8288
rect -3521 -8344 -3503 -8288
rect -3595 -8368 -3575 -8344
rect -3523 -8368 -3503 -8344
rect -3595 -8424 -3577 -8368
rect -3521 -8424 -3503 -8368
rect -3595 -8438 -3575 -8424
rect -3523 -8438 -3503 -8424
rect -3595 -8448 -3503 -8438
rect -3595 -8504 -3577 -8448
rect -3521 -8504 -3503 -8448
rect -3595 -8514 -3503 -8504
rect -3595 -8528 -3575 -8514
rect -3523 -8528 -3503 -8514
rect -3595 -8584 -3577 -8528
rect -3521 -8584 -3503 -8528
rect -3595 -8608 -3575 -8584
rect -3523 -8608 -3503 -8584
rect -3595 -8664 -3577 -8608
rect -3521 -8664 -3503 -8608
rect -3595 -8688 -3575 -8664
rect -3523 -8688 -3503 -8664
rect -3595 -8744 -3577 -8688
rect -3521 -8744 -3503 -8688
rect -3595 -8758 -3575 -8744
rect -3523 -8758 -3503 -8744
rect -3595 -8768 -3503 -8758
rect -3595 -8824 -3577 -8768
rect -3521 -8824 -3503 -8768
rect -3595 -8834 -3503 -8824
rect -3595 -8848 -3575 -8834
rect -3523 -8848 -3503 -8834
rect -3595 -8904 -3577 -8848
rect -3521 -8904 -3503 -8848
rect -3595 -8928 -3575 -8904
rect -3523 -8928 -3503 -8904
rect -3595 -8984 -3577 -8928
rect -3521 -8984 -3503 -8928
rect -3595 -9008 -3575 -8984
rect -3523 -9008 -3503 -8984
rect -3595 -9064 -3577 -9008
rect -3521 -9064 -3503 -9008
rect -3595 -9078 -3575 -9064
rect -3523 -9078 -3503 -9064
rect -3595 -9088 -3503 -9078
rect -3595 -9144 -3577 -9088
rect -3521 -9144 -3503 -9088
rect -3595 -9154 -3503 -9144
rect -3595 -9168 -3575 -9154
rect -3523 -9168 -3503 -9154
rect -3595 -9224 -3577 -9168
rect -3521 -9224 -3503 -9168
rect -3595 -9248 -3575 -9224
rect -3523 -9248 -3503 -9224
rect -3595 -9304 -3577 -9248
rect -3521 -9304 -3503 -9248
rect -3595 -9328 -3575 -9304
rect -3523 -9328 -3503 -9304
rect -3595 -9384 -3577 -9328
rect -3521 -9384 -3503 -9328
rect -3595 -9398 -3575 -9384
rect -3523 -9398 -3503 -9384
rect -3595 -9408 -3503 -9398
rect -3595 -9464 -3577 -9408
rect -3521 -9464 -3503 -9408
rect -3595 -9474 -3503 -9464
rect -3595 -9488 -3575 -9474
rect -3523 -9488 -3503 -9474
rect -3595 -9544 -3577 -9488
rect -3521 -9544 -3503 -9488
rect -3595 -9568 -3575 -9544
rect -3523 -9568 -3503 -9544
rect -3595 -9624 -3577 -9568
rect -3521 -9624 -3503 -9568
rect -3595 -9648 -3575 -9624
rect -3523 -9648 -3503 -9624
rect -3595 -9704 -3577 -9648
rect -3521 -9704 -3503 -9648
rect -3595 -9718 -3575 -9704
rect -3523 -9718 -3503 -9704
rect -3595 -9728 -3503 -9718
rect -3595 -9784 -3577 -9728
rect -3521 -9784 -3503 -9728
rect -3595 -9794 -3503 -9784
rect -3595 -9808 -3575 -9794
rect -3523 -9808 -3503 -9794
rect -3595 -9864 -3577 -9808
rect -3521 -9864 -3503 -9808
rect -3595 -9888 -3575 -9864
rect -3523 -9888 -3503 -9864
rect -3595 -9944 -3577 -9888
rect -3521 -9944 -3503 -9888
rect -3595 -9968 -3575 -9944
rect -3523 -9968 -3503 -9944
rect -3595 -10024 -3577 -9968
rect -3521 -10024 -3503 -9968
rect -3595 -10038 -3575 -10024
rect -3523 -10038 -3503 -10024
rect -3595 -10048 -3503 -10038
rect -3595 -10104 -3577 -10048
rect -3521 -10104 -3503 -10048
rect -3595 -10140 -3503 -10104
rect -600 -6855 -486 -6815
rect -600 -6911 -571 -6855
rect -515 -6911 -486 -6855
rect -600 -6921 -486 -6911
rect -600 -6935 -569 -6921
rect -517 -6935 -486 -6921
rect -600 -6991 -571 -6935
rect -515 -6991 -486 -6935
rect -600 -7015 -569 -6991
rect -517 -7015 -486 -6991
rect -600 -7071 -571 -7015
rect -515 -7071 -486 -7015
rect -600 -7095 -569 -7071
rect -517 -7095 -486 -7071
rect -600 -7151 -571 -7095
rect -515 -7151 -486 -7095
rect -600 -7165 -569 -7151
rect -517 -7165 -486 -7151
rect -600 -7175 -486 -7165
rect -600 -7231 -571 -7175
rect -515 -7231 -486 -7175
rect -600 -7241 -486 -7231
rect -600 -7255 -569 -7241
rect -517 -7255 -486 -7241
rect -600 -7311 -571 -7255
rect -515 -7311 -486 -7255
rect -600 -7335 -569 -7311
rect -517 -7335 -486 -7311
rect -600 -7391 -571 -7335
rect -515 -7391 -486 -7335
rect -600 -7415 -569 -7391
rect -517 -7415 -486 -7391
rect -600 -7471 -571 -7415
rect -515 -7471 -486 -7415
rect -600 -7485 -569 -7471
rect -517 -7485 -486 -7471
rect -600 -7495 -486 -7485
rect -600 -7551 -571 -7495
rect -515 -7551 -486 -7495
rect -600 -7561 -486 -7551
rect -600 -7575 -569 -7561
rect -517 -7575 -486 -7561
rect -600 -7631 -571 -7575
rect -515 -7631 -486 -7575
rect -600 -7655 -569 -7631
rect -517 -7655 -486 -7631
rect -600 -7711 -571 -7655
rect -515 -7711 -486 -7655
rect -600 -7735 -569 -7711
rect -517 -7735 -486 -7711
rect -600 -7791 -571 -7735
rect -515 -7791 -486 -7735
rect -600 -7805 -569 -7791
rect -517 -7805 -486 -7791
rect -600 -7815 -486 -7805
rect -600 -7871 -571 -7815
rect -515 -7871 -486 -7815
rect -600 -7881 -486 -7871
rect -600 -7895 -569 -7881
rect -517 -7895 -486 -7881
rect -600 -7951 -571 -7895
rect -515 -7951 -486 -7895
rect -600 -7975 -569 -7951
rect -517 -7975 -486 -7951
rect -600 -8031 -571 -7975
rect -515 -8031 -486 -7975
rect -600 -8055 -569 -8031
rect -517 -8055 -486 -8031
rect -600 -8111 -571 -8055
rect -515 -8111 -486 -8055
rect -600 -8125 -569 -8111
rect -517 -8125 -486 -8111
rect -600 -8135 -486 -8125
rect -600 -8191 -571 -8135
rect -515 -8191 -486 -8135
rect -600 -8201 -486 -8191
rect -600 -8215 -569 -8201
rect -517 -8215 -486 -8201
rect -600 -8271 -571 -8215
rect -515 -8271 -486 -8215
rect -600 -8295 -569 -8271
rect -517 -8295 -486 -8271
rect -600 -8351 -571 -8295
rect -515 -8351 -486 -8295
rect -600 -8375 -569 -8351
rect -517 -8375 -486 -8351
rect -600 -8431 -571 -8375
rect -515 -8431 -486 -8375
rect -600 -8445 -569 -8431
rect -517 -8445 -486 -8431
rect -600 -8455 -486 -8445
rect -600 -8511 -571 -8455
rect -515 -8511 -486 -8455
rect -600 -8521 -486 -8511
rect -600 -8535 -569 -8521
rect -517 -8535 -486 -8521
rect -600 -8591 -571 -8535
rect -515 -8591 -486 -8535
rect -600 -8615 -569 -8591
rect -517 -8615 -486 -8591
rect -600 -8671 -571 -8615
rect -515 -8671 -486 -8615
rect -600 -8695 -569 -8671
rect -517 -8695 -486 -8671
rect -600 -8751 -571 -8695
rect -515 -8751 -486 -8695
rect -600 -8765 -569 -8751
rect -517 -8765 -486 -8751
rect -600 -8775 -486 -8765
rect -600 -8831 -571 -8775
rect -515 -8831 -486 -8775
rect -600 -8841 -486 -8831
rect -600 -8855 -569 -8841
rect -517 -8855 -486 -8841
rect -600 -8911 -571 -8855
rect -515 -8911 -486 -8855
rect -600 -8935 -569 -8911
rect -517 -8935 -486 -8911
rect -600 -8991 -571 -8935
rect -515 -8991 -486 -8935
rect -600 -9015 -569 -8991
rect -517 -9015 -486 -8991
rect -600 -9071 -571 -9015
rect -515 -9071 -486 -9015
rect -600 -9085 -569 -9071
rect -517 -9085 -486 -9071
rect -600 -9095 -486 -9085
rect -600 -9151 -571 -9095
rect -515 -9151 -486 -9095
rect -600 -9161 -486 -9151
rect -600 -9175 -569 -9161
rect -517 -9175 -486 -9161
rect -600 -9231 -571 -9175
rect -515 -9231 -486 -9175
rect -600 -9255 -569 -9231
rect -517 -9255 -486 -9231
rect -600 -9311 -571 -9255
rect -515 -9311 -486 -9255
rect -600 -9335 -569 -9311
rect -517 -9335 -486 -9311
rect -600 -9391 -571 -9335
rect -515 -9391 -486 -9335
rect -600 -9405 -569 -9391
rect -517 -9405 -486 -9391
rect -600 -9415 -486 -9405
rect -600 -9471 -571 -9415
rect -515 -9471 -486 -9415
rect -600 -9481 -486 -9471
rect -600 -9495 -569 -9481
rect -517 -9495 -486 -9481
rect -600 -9551 -571 -9495
rect -515 -9551 -486 -9495
rect -600 -9575 -569 -9551
rect -517 -9575 -486 -9551
rect -600 -9631 -571 -9575
rect -515 -9631 -486 -9575
rect -600 -9655 -569 -9631
rect -517 -9655 -486 -9631
rect -600 -9711 -571 -9655
rect -515 -9711 -486 -9655
rect -600 -9725 -569 -9711
rect -517 -9725 -486 -9711
rect -600 -9735 -486 -9725
rect -600 -9791 -571 -9735
rect -515 -9791 -486 -9735
rect -600 -9801 -486 -9791
rect -600 -9815 -569 -9801
rect -517 -9815 -486 -9801
rect -600 -9871 -571 -9815
rect -515 -9871 -486 -9815
rect -600 -9895 -569 -9871
rect -517 -9895 -486 -9871
rect -600 -9951 -571 -9895
rect -515 -9951 -486 -9895
rect -600 -9975 -569 -9951
rect -517 -9975 -486 -9951
rect -600 -10031 -571 -9975
rect -515 -10031 -486 -9975
rect -600 -10045 -569 -10031
rect -517 -10045 -486 -10031
rect -600 -10055 -486 -10045
rect -600 -10111 -571 -10055
rect -515 -10111 -486 -10055
rect -600 -10150 -486 -10111
rect -2179 -12092 -1943 -12072
rect -2179 -12308 -2169 -12092
rect -1953 -12308 -1943 -12092
rect -2179 -12328 -1943 -12308
<< via2 >>
rect -15400 78112 -15184 78130
rect -15400 77932 -15382 78112
rect -15382 77932 -15202 78112
rect -15202 77932 -15184 78112
rect -15400 77914 -15184 77932
rect 12616 78083 12832 78101
rect 12616 77903 12634 78083
rect 12634 77903 12814 78083
rect 12814 77903 12832 78083
rect 12616 77885 12832 77903
rect 24666 78084 24882 78102
rect 24666 77904 24684 78084
rect 24684 77904 24864 78084
rect 24864 77904 24882 78084
rect 24666 77886 24882 77904
rect -16827 76666 -16825 76688
rect -16825 76666 -16773 76688
rect -16773 76666 -16771 76688
rect -16827 76654 -16771 76666
rect -16827 76632 -16825 76654
rect -16825 76632 -16773 76654
rect -16773 76632 -16771 76654
rect -16827 76602 -16825 76608
rect -16825 76602 -16773 76608
rect -16773 76602 -16771 76608
rect -16827 76590 -16771 76602
rect -16827 76552 -16825 76590
rect -16825 76552 -16773 76590
rect -16773 76552 -16771 76590
rect -16827 76526 -16771 76528
rect -16827 76474 -16825 76526
rect -16825 76474 -16773 76526
rect -16773 76474 -16771 76526
rect -16827 76472 -16771 76474
rect -16827 76410 -16825 76448
rect -16825 76410 -16773 76448
rect -16773 76410 -16771 76448
rect -16827 76398 -16771 76410
rect -16827 76392 -16825 76398
rect -16825 76392 -16773 76398
rect -16773 76392 -16771 76398
rect -16827 76346 -16825 76368
rect -16825 76346 -16773 76368
rect -16773 76346 -16771 76368
rect -16827 76334 -16771 76346
rect -16827 76312 -16825 76334
rect -16825 76312 -16773 76334
rect -16773 76312 -16771 76334
rect -16827 76282 -16825 76288
rect -16825 76282 -16773 76288
rect -16773 76282 -16771 76288
rect -16827 76270 -16771 76282
rect -16827 76232 -16825 76270
rect -16825 76232 -16773 76270
rect -16773 76232 -16771 76270
rect -16827 76206 -16771 76208
rect -16827 76154 -16825 76206
rect -16825 76154 -16773 76206
rect -16773 76154 -16771 76206
rect -16827 76152 -16771 76154
rect -16827 76090 -16825 76128
rect -16825 76090 -16773 76128
rect -16773 76090 -16771 76128
rect -16827 76078 -16771 76090
rect -16827 76072 -16825 76078
rect -16825 76072 -16773 76078
rect -16773 76072 -16771 76078
rect -16827 76026 -16825 76048
rect -16825 76026 -16773 76048
rect -16773 76026 -16771 76048
rect -16827 76014 -16771 76026
rect -16827 75992 -16825 76014
rect -16825 75992 -16773 76014
rect -16773 75992 -16771 76014
rect -16827 75962 -16825 75968
rect -16825 75962 -16773 75968
rect -16773 75962 -16771 75968
rect -16827 75950 -16771 75962
rect -16827 75912 -16825 75950
rect -16825 75912 -16773 75950
rect -16773 75912 -16771 75950
rect -16827 75886 -16771 75888
rect -16827 75834 -16825 75886
rect -16825 75834 -16773 75886
rect -16773 75834 -16771 75886
rect -16827 75832 -16771 75834
rect -16827 75770 -16825 75808
rect -16825 75770 -16773 75808
rect -16773 75770 -16771 75808
rect -16827 75758 -16771 75770
rect -16827 75752 -16825 75758
rect -16825 75752 -16773 75758
rect -16773 75752 -16771 75758
rect -16827 75706 -16825 75728
rect -16825 75706 -16773 75728
rect -16773 75706 -16771 75728
rect -16827 75694 -16771 75706
rect -16827 75672 -16825 75694
rect -16825 75672 -16773 75694
rect -16773 75672 -16771 75694
rect -16827 75642 -16825 75648
rect -16825 75642 -16773 75648
rect -16773 75642 -16771 75648
rect -16827 75630 -16771 75642
rect -16827 75592 -16825 75630
rect -16825 75592 -16773 75630
rect -16773 75592 -16771 75630
rect -16827 75566 -16771 75568
rect -16827 75514 -16825 75566
rect -16825 75514 -16773 75566
rect -16773 75514 -16771 75566
rect -16827 75512 -16771 75514
rect -16827 75450 -16825 75488
rect -16825 75450 -16773 75488
rect -16773 75450 -16771 75488
rect -16827 75438 -16771 75450
rect -16827 75432 -16825 75438
rect -16825 75432 -16773 75438
rect -16773 75432 -16771 75438
rect -16827 75386 -16825 75408
rect -16825 75386 -16773 75408
rect -16773 75386 -16771 75408
rect -16827 75374 -16771 75386
rect -16827 75352 -16825 75374
rect -16825 75352 -16773 75374
rect -16773 75352 -16771 75374
rect -16827 75322 -16825 75328
rect -16825 75322 -16773 75328
rect -16773 75322 -16771 75328
rect -16827 75310 -16771 75322
rect -16827 75272 -16825 75310
rect -16825 75272 -16773 75310
rect -16773 75272 -16771 75310
rect -16827 75246 -16771 75248
rect -16827 75194 -16825 75246
rect -16825 75194 -16773 75246
rect -16773 75194 -16771 75246
rect -16827 75192 -16771 75194
rect -16827 75130 -16825 75168
rect -16825 75130 -16773 75168
rect -16773 75130 -16771 75168
rect -16827 75118 -16771 75130
rect -16827 75112 -16825 75118
rect -16825 75112 -16773 75118
rect -16773 75112 -16771 75118
rect -16827 75066 -16825 75088
rect -16825 75066 -16773 75088
rect -16773 75066 -16771 75088
rect -16827 75054 -16771 75066
rect -16827 75032 -16825 75054
rect -16825 75032 -16773 75054
rect -16773 75032 -16771 75054
rect -16827 75002 -16825 75008
rect -16825 75002 -16773 75008
rect -16773 75002 -16771 75008
rect -16827 74990 -16771 75002
rect -16827 74952 -16825 74990
rect -16825 74952 -16773 74990
rect -16773 74952 -16771 74990
rect -16827 74926 -16771 74928
rect -16827 74874 -16825 74926
rect -16825 74874 -16773 74926
rect -16773 74874 -16771 74926
rect -16827 74872 -16771 74874
rect -16827 74810 -16825 74848
rect -16825 74810 -16773 74848
rect -16773 74810 -16771 74848
rect -16827 74798 -16771 74810
rect -16827 74792 -16825 74798
rect -16825 74792 -16773 74798
rect -16773 74792 -16771 74798
rect -16827 74746 -16825 74768
rect -16825 74746 -16773 74768
rect -16773 74746 -16771 74768
rect -16827 74734 -16771 74746
rect -16827 74712 -16825 74734
rect -16825 74712 -16773 74734
rect -16773 74712 -16771 74734
rect -16827 74682 -16825 74688
rect -16825 74682 -16773 74688
rect -16773 74682 -16771 74688
rect -16827 74670 -16771 74682
rect -16827 74632 -16825 74670
rect -16825 74632 -16773 74670
rect -16773 74632 -16771 74670
rect -16827 74606 -16771 74608
rect -16827 74554 -16825 74606
rect -16825 74554 -16773 74606
rect -16773 74554 -16771 74606
rect -16827 74552 -16771 74554
rect -16827 74490 -16825 74528
rect -16825 74490 -16773 74528
rect -16773 74490 -16771 74528
rect -16827 74478 -16771 74490
rect -16827 74472 -16825 74478
rect -16825 74472 -16773 74478
rect -16773 74472 -16771 74478
rect -16827 74426 -16825 74448
rect -16825 74426 -16773 74448
rect -16773 74426 -16771 74448
rect -16827 74414 -16771 74426
rect -16827 74392 -16825 74414
rect -16825 74392 -16773 74414
rect -16773 74392 -16771 74414
rect -16827 74362 -16825 74368
rect -16825 74362 -16773 74368
rect -16773 74362 -16771 74368
rect -16827 74350 -16771 74362
rect -16827 74312 -16825 74350
rect -16825 74312 -16773 74350
rect -16773 74312 -16771 74350
rect -16827 74286 -16771 74288
rect -16827 74234 -16825 74286
rect -16825 74234 -16773 74286
rect -16773 74234 -16771 74286
rect -16827 74232 -16771 74234
rect -16827 74170 -16825 74208
rect -16825 74170 -16773 74208
rect -16773 74170 -16771 74208
rect -16827 74158 -16771 74170
rect -16827 74152 -16825 74158
rect -16825 74152 -16773 74158
rect -16773 74152 -16771 74158
rect -16827 74106 -16825 74128
rect -16825 74106 -16773 74128
rect -16773 74106 -16771 74128
rect -16827 74094 -16771 74106
rect -16827 74072 -16825 74094
rect -16825 74072 -16773 74094
rect -16773 74072 -16771 74094
rect -16827 74042 -16825 74048
rect -16825 74042 -16773 74048
rect -16773 74042 -16771 74048
rect -16827 74030 -16771 74042
rect -16827 73992 -16825 74030
rect -16825 73992 -16773 74030
rect -16773 73992 -16771 74030
rect -16827 73966 -16771 73968
rect -16827 73914 -16825 73966
rect -16825 73914 -16773 73966
rect -16773 73914 -16771 73966
rect -16827 73912 -16771 73914
rect -16827 73850 -16825 73888
rect -16825 73850 -16773 73888
rect -16773 73850 -16771 73888
rect -16827 73838 -16771 73850
rect -16827 73832 -16825 73838
rect -16825 73832 -16773 73838
rect -16773 73832 -16771 73838
rect -16827 73786 -16825 73808
rect -16825 73786 -16773 73808
rect -16773 73786 -16771 73808
rect -16827 73774 -16771 73786
rect -16827 73752 -16825 73774
rect -16825 73752 -16773 73774
rect -16773 73752 -16771 73774
rect -16827 73722 -16825 73728
rect -16825 73722 -16773 73728
rect -16773 73722 -16771 73728
rect -16827 73710 -16771 73722
rect -16827 73672 -16825 73710
rect -16825 73672 -16773 73710
rect -16773 73672 -16771 73710
rect -16827 73646 -16771 73648
rect -16827 73594 -16825 73646
rect -16825 73594 -16773 73646
rect -16773 73594 -16771 73646
rect -16827 73592 -16771 73594
rect -16827 73530 -16825 73568
rect -16825 73530 -16773 73568
rect -16773 73530 -16771 73568
rect -16827 73518 -16771 73530
rect -16827 73512 -16825 73518
rect -16825 73512 -16773 73518
rect -16773 73512 -16771 73518
rect -16827 73466 -16825 73488
rect -16825 73466 -16773 73488
rect -16773 73466 -16771 73488
rect -16827 73454 -16771 73466
rect -16827 73432 -16825 73454
rect -16825 73432 -16773 73454
rect -16773 73432 -16771 73454
rect -13826 76672 -13824 76694
rect -13824 76672 -13772 76694
rect -13772 76672 -13770 76694
rect -13826 76660 -13770 76672
rect -13826 76638 -13824 76660
rect -13824 76638 -13772 76660
rect -13772 76638 -13770 76660
rect -13826 76608 -13824 76614
rect -13824 76608 -13772 76614
rect -13772 76608 -13770 76614
rect -13826 76596 -13770 76608
rect -13826 76558 -13824 76596
rect -13824 76558 -13772 76596
rect -13772 76558 -13770 76596
rect -13826 76532 -13770 76534
rect -13826 76480 -13824 76532
rect -13824 76480 -13772 76532
rect -13772 76480 -13770 76532
rect -13826 76478 -13770 76480
rect -13826 76416 -13824 76454
rect -13824 76416 -13772 76454
rect -13772 76416 -13770 76454
rect -13826 76404 -13770 76416
rect -13826 76398 -13824 76404
rect -13824 76398 -13772 76404
rect -13772 76398 -13770 76404
rect -13826 76352 -13824 76374
rect -13824 76352 -13772 76374
rect -13772 76352 -13770 76374
rect -13826 76340 -13770 76352
rect -13826 76318 -13824 76340
rect -13824 76318 -13772 76340
rect -13772 76318 -13770 76340
rect -13826 76288 -13824 76294
rect -13824 76288 -13772 76294
rect -13772 76288 -13770 76294
rect -13826 76276 -13770 76288
rect -13826 76238 -13824 76276
rect -13824 76238 -13772 76276
rect -13772 76238 -13770 76276
rect -13826 76212 -13770 76214
rect -13826 76160 -13824 76212
rect -13824 76160 -13772 76212
rect -13772 76160 -13770 76212
rect -13826 76158 -13770 76160
rect -13826 76096 -13824 76134
rect -13824 76096 -13772 76134
rect -13772 76096 -13770 76134
rect -13826 76084 -13770 76096
rect -13826 76078 -13824 76084
rect -13824 76078 -13772 76084
rect -13772 76078 -13770 76084
rect -13826 76032 -13824 76054
rect -13824 76032 -13772 76054
rect -13772 76032 -13770 76054
rect -13826 76020 -13770 76032
rect -13826 75998 -13824 76020
rect -13824 75998 -13772 76020
rect -13772 75998 -13770 76020
rect -13826 75968 -13824 75974
rect -13824 75968 -13772 75974
rect -13772 75968 -13770 75974
rect -13826 75956 -13770 75968
rect -13826 75918 -13824 75956
rect -13824 75918 -13772 75956
rect -13772 75918 -13770 75956
rect -13826 75892 -13770 75894
rect -13826 75840 -13824 75892
rect -13824 75840 -13772 75892
rect -13772 75840 -13770 75892
rect -13826 75838 -13770 75840
rect -13826 75776 -13824 75814
rect -13824 75776 -13772 75814
rect -13772 75776 -13770 75814
rect -13826 75764 -13770 75776
rect -13826 75758 -13824 75764
rect -13824 75758 -13772 75764
rect -13772 75758 -13770 75764
rect -13826 75712 -13824 75734
rect -13824 75712 -13772 75734
rect -13772 75712 -13770 75734
rect -13826 75700 -13770 75712
rect -13826 75678 -13824 75700
rect -13824 75678 -13772 75700
rect -13772 75678 -13770 75700
rect -13826 75648 -13824 75654
rect -13824 75648 -13772 75654
rect -13772 75648 -13770 75654
rect -13826 75636 -13770 75648
rect -13826 75598 -13824 75636
rect -13824 75598 -13772 75636
rect -13772 75598 -13770 75636
rect -13826 75572 -13770 75574
rect -13826 75520 -13824 75572
rect -13824 75520 -13772 75572
rect -13772 75520 -13770 75572
rect -13826 75518 -13770 75520
rect -13826 75456 -13824 75494
rect -13824 75456 -13772 75494
rect -13772 75456 -13770 75494
rect -13826 75444 -13770 75456
rect -13826 75438 -13824 75444
rect -13824 75438 -13772 75444
rect -13772 75438 -13770 75444
rect -13826 75392 -13824 75414
rect -13824 75392 -13772 75414
rect -13772 75392 -13770 75414
rect -13826 75380 -13770 75392
rect -13826 75358 -13824 75380
rect -13824 75358 -13772 75380
rect -13772 75358 -13770 75380
rect -13826 75328 -13824 75334
rect -13824 75328 -13772 75334
rect -13772 75328 -13770 75334
rect -13826 75316 -13770 75328
rect -13826 75278 -13824 75316
rect -13824 75278 -13772 75316
rect -13772 75278 -13770 75316
rect -13826 75252 -13770 75254
rect -13826 75200 -13824 75252
rect -13824 75200 -13772 75252
rect -13772 75200 -13770 75252
rect -13826 75198 -13770 75200
rect -13826 75136 -13824 75174
rect -13824 75136 -13772 75174
rect -13772 75136 -13770 75174
rect -13826 75124 -13770 75136
rect -13826 75118 -13824 75124
rect -13824 75118 -13772 75124
rect -13772 75118 -13770 75124
rect -13826 75072 -13824 75094
rect -13824 75072 -13772 75094
rect -13772 75072 -13770 75094
rect -13826 75060 -13770 75072
rect -13826 75038 -13824 75060
rect -13824 75038 -13772 75060
rect -13772 75038 -13770 75060
rect -13826 75008 -13824 75014
rect -13824 75008 -13772 75014
rect -13772 75008 -13770 75014
rect -13826 74996 -13770 75008
rect -13826 74958 -13824 74996
rect -13824 74958 -13772 74996
rect -13772 74958 -13770 74996
rect -13826 74932 -13770 74934
rect -13826 74880 -13824 74932
rect -13824 74880 -13772 74932
rect -13772 74880 -13770 74932
rect -13826 74878 -13770 74880
rect -13826 74816 -13824 74854
rect -13824 74816 -13772 74854
rect -13772 74816 -13770 74854
rect -13826 74804 -13770 74816
rect -13826 74798 -13824 74804
rect -13824 74798 -13772 74804
rect -13772 74798 -13770 74804
rect -13826 74752 -13824 74774
rect -13824 74752 -13772 74774
rect -13772 74752 -13770 74774
rect -13826 74740 -13770 74752
rect -13826 74718 -13824 74740
rect -13824 74718 -13772 74740
rect -13772 74718 -13770 74740
rect -13826 74688 -13824 74694
rect -13824 74688 -13772 74694
rect -13772 74688 -13770 74694
rect -13826 74676 -13770 74688
rect -13826 74638 -13824 74676
rect -13824 74638 -13772 74676
rect -13772 74638 -13770 74676
rect -13826 74612 -13770 74614
rect -13826 74560 -13824 74612
rect -13824 74560 -13772 74612
rect -13772 74560 -13770 74612
rect -13826 74558 -13770 74560
rect -13826 74496 -13824 74534
rect -13824 74496 -13772 74534
rect -13772 74496 -13770 74534
rect -13826 74484 -13770 74496
rect -13826 74478 -13824 74484
rect -13824 74478 -13772 74484
rect -13772 74478 -13770 74484
rect -13826 74432 -13824 74454
rect -13824 74432 -13772 74454
rect -13772 74432 -13770 74454
rect -13826 74420 -13770 74432
rect -13826 74398 -13824 74420
rect -13824 74398 -13772 74420
rect -13772 74398 -13770 74420
rect -13826 74368 -13824 74374
rect -13824 74368 -13772 74374
rect -13772 74368 -13770 74374
rect -13826 74356 -13770 74368
rect -13826 74318 -13824 74356
rect -13824 74318 -13772 74356
rect -13772 74318 -13770 74356
rect -13826 74292 -13770 74294
rect -13826 74240 -13824 74292
rect -13824 74240 -13772 74292
rect -13772 74240 -13770 74292
rect -13826 74238 -13770 74240
rect -13826 74176 -13824 74214
rect -13824 74176 -13772 74214
rect -13772 74176 -13770 74214
rect -13826 74164 -13770 74176
rect -13826 74158 -13824 74164
rect -13824 74158 -13772 74164
rect -13772 74158 -13770 74164
rect -13826 74112 -13824 74134
rect -13824 74112 -13772 74134
rect -13772 74112 -13770 74134
rect -13826 74100 -13770 74112
rect -13826 74078 -13824 74100
rect -13824 74078 -13772 74100
rect -13772 74078 -13770 74100
rect -13826 74048 -13824 74054
rect -13824 74048 -13772 74054
rect -13772 74048 -13770 74054
rect -13826 74036 -13770 74048
rect -13826 73998 -13824 74036
rect -13824 73998 -13772 74036
rect -13772 73998 -13770 74036
rect -13826 73972 -13770 73974
rect -13826 73920 -13824 73972
rect -13824 73920 -13772 73972
rect -13772 73920 -13770 73972
rect -13826 73918 -13770 73920
rect -13826 73856 -13824 73894
rect -13824 73856 -13772 73894
rect -13772 73856 -13770 73894
rect -13826 73844 -13770 73856
rect -13826 73838 -13824 73844
rect -13824 73838 -13772 73844
rect -13772 73838 -13770 73844
rect -13826 73792 -13824 73814
rect -13824 73792 -13772 73814
rect -13772 73792 -13770 73814
rect -13826 73780 -13770 73792
rect -13826 73758 -13824 73780
rect -13824 73758 -13772 73780
rect -13772 73758 -13770 73780
rect -13826 73728 -13824 73734
rect -13824 73728 -13772 73734
rect -13772 73728 -13770 73734
rect -13826 73716 -13770 73728
rect -13826 73678 -13824 73716
rect -13824 73678 -13772 73716
rect -13772 73678 -13770 73716
rect -13826 73652 -13770 73654
rect -13826 73600 -13824 73652
rect -13824 73600 -13772 73652
rect -13772 73600 -13770 73652
rect -13826 73598 -13770 73600
rect -13826 73536 -13824 73574
rect -13824 73536 -13772 73574
rect -13772 73536 -13770 73574
rect -13826 73524 -13770 73536
rect -13826 73518 -13824 73524
rect -13824 73518 -13772 73524
rect -13772 73518 -13770 73524
rect -13826 73472 -13824 73494
rect -13824 73472 -13772 73494
rect -13772 73472 -13770 73494
rect -13826 73460 -13770 73472
rect -13826 73438 -13824 73460
rect -13824 73438 -13772 73460
rect -13772 73438 -13770 73460
rect 11179 76720 11235 76730
rect 11179 76674 11235 76720
rect 11179 76594 11235 76650
rect 11179 76514 11235 76570
rect 11179 76434 11235 76490
rect 11179 76354 11235 76410
rect 11179 76274 11235 76330
rect 11179 76194 11235 76250
rect 11179 76114 11235 76170
rect 11179 76034 11235 76090
rect 11179 75954 11235 76010
rect 11179 75874 11235 75930
rect 11179 75794 11235 75850
rect 11179 75714 11235 75770
rect 11179 75634 11235 75690
rect 11179 75554 11235 75610
rect 11179 75474 11235 75530
rect 11179 75394 11235 75450
rect 11179 75314 11235 75370
rect 11179 75234 11235 75290
rect 11179 75154 11235 75210
rect 11179 75074 11235 75130
rect 11179 74994 11235 75050
rect 11179 74914 11235 74970
rect 11179 74834 11235 74890
rect 11179 74754 11235 74810
rect 11179 74674 11235 74730
rect 11179 74594 11235 74650
rect 11179 74514 11235 74570
rect 11179 74434 11235 74490
rect 11179 74354 11235 74410
rect 11179 74274 11235 74330
rect 11179 74194 11235 74250
rect 11179 74114 11235 74170
rect 11179 74034 11235 74090
rect 11179 73954 11235 74010
rect 11179 73874 11235 73930
rect 11179 73794 11235 73850
rect 11179 73714 11235 73770
rect 11179 73634 11235 73690
rect 11179 73554 11235 73610
rect 11179 73474 11235 73530
rect 11179 73404 11235 73450
rect 11179 73394 11235 73404
rect 14180 76733 14236 76743
rect 14180 76687 14236 76733
rect 14180 76607 14236 76663
rect 14180 76527 14236 76583
rect 14180 76447 14236 76503
rect 14180 76367 14236 76423
rect 14180 76287 14236 76343
rect 14180 76207 14236 76263
rect 14180 76127 14236 76183
rect 14180 76047 14236 76103
rect 14180 75967 14236 76023
rect 14180 75887 14236 75943
rect 14180 75807 14236 75863
rect 14180 75727 14236 75783
rect 14180 75647 14236 75703
rect 14180 75567 14236 75623
rect 14180 75487 14236 75543
rect 14180 75407 14236 75463
rect 14180 75327 14236 75383
rect 14180 75247 14236 75303
rect 14180 75167 14236 75223
rect 14180 75087 14236 75143
rect 14180 75007 14236 75063
rect 14180 74927 14236 74983
rect 14180 74847 14236 74903
rect 14180 74767 14236 74823
rect 14180 74687 14236 74743
rect 14180 74607 14236 74663
rect 14180 74527 14236 74583
rect 14180 74447 14236 74503
rect 14180 74367 14236 74423
rect 14180 74287 14236 74343
rect 14180 74207 14236 74263
rect 14180 74127 14236 74183
rect 14180 74047 14236 74103
rect 14180 73967 14236 74023
rect 14180 73887 14236 73943
rect 14180 73807 14236 73863
rect 14180 73727 14236 73783
rect 14180 73647 14236 73703
rect 14180 73567 14236 73623
rect 14180 73487 14236 73543
rect 14180 73417 14236 73463
rect 14180 73407 14236 73417
rect -16660 71796 -16604 71798
rect -16660 71744 -16658 71796
rect -16658 71744 -16606 71796
rect -16606 71744 -16604 71796
rect -16660 71742 -16604 71744
rect -15482 71792 -15426 71794
rect -15482 71740 -15480 71792
rect -15480 71740 -15428 71792
rect -15428 71740 -15426 71792
rect -15482 71738 -15426 71740
rect -15265 71799 -15209 71801
rect -15265 71747 -15263 71799
rect -15263 71747 -15211 71799
rect -15211 71747 -15209 71799
rect -15265 71745 -15209 71747
rect -14131 71796 -14075 71798
rect -14131 71744 -14129 71796
rect -14129 71744 -14077 71796
rect -14077 71744 -14075 71796
rect -14131 71742 -14075 71744
rect -16550 70292 -16494 70294
rect -16550 70240 -16548 70292
rect -16548 70240 -16496 70292
rect -16496 70240 -16494 70292
rect -16550 70238 -16494 70240
rect -15436 70278 -15380 70280
rect -15436 70226 -15434 70278
rect -15434 70226 -15382 70278
rect -15382 70226 -15380 70278
rect -15436 70224 -15380 70226
rect -15223 70279 -15167 70281
rect -15223 70227 -15221 70279
rect -15221 70227 -15169 70279
rect -15169 70227 -15167 70279
rect -15223 70225 -15167 70227
rect -14059 70279 -14003 70281
rect -14059 70227 -14057 70279
rect -14057 70227 -14005 70279
rect -14005 70227 -14003 70279
rect -14059 70225 -14003 70227
rect -16704 68643 -16648 68699
rect -15418 68442 -15416 68488
rect -15416 68442 -15364 68488
rect -15364 68442 -15362 68488
rect -15418 68432 -15362 68442
rect -15418 68378 -15416 68408
rect -15416 68378 -15364 68408
rect -15364 68378 -15362 68408
rect -15418 68366 -15362 68378
rect -15418 68352 -15416 68366
rect -15416 68352 -15364 68366
rect -15364 68352 -15362 68366
rect -15418 68314 -15416 68328
rect -15416 68314 -15364 68328
rect -15364 68314 -15362 68328
rect -15418 68302 -15362 68314
rect -15418 68272 -15416 68302
rect -15416 68272 -15364 68302
rect -15364 68272 -15362 68302
rect -15955 68241 -15899 68251
rect -15955 68195 -15953 68241
rect -15953 68195 -15901 68241
rect -15901 68195 -15899 68241
rect -15955 68125 -15953 68171
rect -15953 68125 -15901 68171
rect -15901 68125 -15899 68171
rect -15955 68115 -15899 68125
rect -15418 68238 -15362 68248
rect -15418 68192 -15416 68238
rect -15416 68192 -15364 68238
rect -15364 68192 -15362 68238
rect -14871 68244 -14815 68254
rect -14871 68198 -14869 68244
rect -14869 68198 -14817 68244
rect -14817 68198 -14815 68244
rect -14871 68128 -14869 68174
rect -14869 68128 -14817 68174
rect -14817 68128 -14815 68174
rect -14871 68118 -14815 68128
rect -14195 68013 -14139 68069
rect -16573 67607 -16517 67609
rect -16573 67555 -16571 67607
rect -16571 67555 -16519 67607
rect -16519 67555 -16517 67607
rect -16573 67553 -16517 67555
rect -15418 67601 -15362 67603
rect -15418 67549 -15416 67601
rect -15416 67549 -15364 67601
rect -15364 67549 -15362 67601
rect -15418 67547 -15362 67549
rect -14300 67612 -14244 67614
rect -14300 67560 -14298 67612
rect -14298 67560 -14246 67612
rect -14246 67560 -14244 67612
rect -14300 67558 -14244 67560
rect 17435 64686 17437 64724
rect 17437 64686 17489 64724
rect 17489 64686 17491 64724
rect 17435 64674 17491 64686
rect 17435 64668 17437 64674
rect 17437 64668 17489 64674
rect 17489 64668 17491 64674
rect 17435 64622 17437 64644
rect 17437 64622 17489 64644
rect 17489 64622 17491 64644
rect 17435 64610 17491 64622
rect 17435 64588 17437 64610
rect 17437 64588 17489 64610
rect 17489 64588 17491 64610
rect 17435 64558 17437 64564
rect 17437 64558 17489 64564
rect 17489 64558 17491 64564
rect 17435 64546 17491 64558
rect 17435 64508 17437 64546
rect 17437 64508 17489 64546
rect 17489 64508 17491 64546
rect 17435 64482 17491 64484
rect 17435 64430 17437 64482
rect 17437 64430 17489 64482
rect 17489 64430 17491 64482
rect 17435 64428 17491 64430
rect 17435 64366 17437 64404
rect 17437 64366 17489 64404
rect 17489 64366 17491 64404
rect 17435 64354 17491 64366
rect 17435 64348 17437 64354
rect 17437 64348 17489 64354
rect 17489 64348 17491 64354
rect 17435 64302 17437 64324
rect 17437 64302 17489 64324
rect 17489 64302 17491 64324
rect 17435 64290 17491 64302
rect 17435 64268 17437 64290
rect 17437 64268 17489 64290
rect 17489 64268 17491 64290
rect 17435 64238 17437 64244
rect 17437 64238 17489 64244
rect 17489 64238 17491 64244
rect 17435 64226 17491 64238
rect 17435 64188 17437 64226
rect 17437 64188 17489 64226
rect 17489 64188 17491 64226
rect 23963 64686 23965 64724
rect 23965 64686 24017 64724
rect 24017 64686 24019 64724
rect 23963 64674 24019 64686
rect 23963 64668 23965 64674
rect 23965 64668 24017 64674
rect 24017 64668 24019 64674
rect 23963 64622 23965 64644
rect 23965 64622 24017 64644
rect 24017 64622 24019 64644
rect 23963 64610 24019 64622
rect 23963 64588 23965 64610
rect 23965 64588 24017 64610
rect 24017 64588 24019 64610
rect 23963 64558 23965 64564
rect 23965 64558 24017 64564
rect 24017 64558 24019 64564
rect 23963 64546 24019 64558
rect 23963 64508 23965 64546
rect 23965 64508 24017 64546
rect 24017 64508 24019 64546
rect 23963 64482 24019 64484
rect 23963 64430 23965 64482
rect 23965 64430 24017 64482
rect 24017 64430 24019 64482
rect 23963 64428 24019 64430
rect 23963 64366 23965 64404
rect 23965 64366 24017 64404
rect 24017 64366 24019 64404
rect 23963 64354 24019 64366
rect 23963 64348 23965 64354
rect 23965 64348 24017 64354
rect 24017 64348 24019 64354
rect 23963 64302 23965 64324
rect 23965 64302 24017 64324
rect 24017 64302 24019 64324
rect 23963 64290 24019 64302
rect 23963 64268 23965 64290
rect 23965 64268 24017 64290
rect 24017 64268 24019 64290
rect 23963 64238 23965 64244
rect 23965 64238 24017 64244
rect 24017 64238 24019 64244
rect 23963 64226 24019 64238
rect 23963 64188 23965 64226
rect 23965 64188 24017 64226
rect 24017 64188 24019 64226
rect 31579 64686 31581 64724
rect 31581 64686 31633 64724
rect 31633 64686 31635 64724
rect 31579 64674 31635 64686
rect 31579 64668 31581 64674
rect 31581 64668 31633 64674
rect 31633 64668 31635 64674
rect 31579 64622 31581 64644
rect 31581 64622 31633 64644
rect 31633 64622 31635 64644
rect 31579 64610 31635 64622
rect 31579 64588 31581 64610
rect 31581 64588 31633 64610
rect 31633 64588 31635 64610
rect 31579 64558 31581 64564
rect 31581 64558 31633 64564
rect 31633 64558 31635 64564
rect 31579 64546 31635 64558
rect 31579 64508 31581 64546
rect 31581 64508 31633 64546
rect 31633 64508 31635 64546
rect 31579 64482 31635 64484
rect 31579 64430 31581 64482
rect 31581 64430 31633 64482
rect 31633 64430 31635 64482
rect 31579 64428 31635 64430
rect 31579 64366 31581 64404
rect 31581 64366 31633 64404
rect 31633 64366 31635 64404
rect 31579 64354 31635 64366
rect 31579 64348 31581 64354
rect 31581 64348 31633 64354
rect 31633 64348 31635 64354
rect 31579 64302 31581 64324
rect 31581 64302 31633 64324
rect 31633 64302 31635 64324
rect 31579 64290 31635 64302
rect 31579 64268 31581 64290
rect 31581 64268 31633 64290
rect 31633 64268 31635 64290
rect 31579 64238 31581 64244
rect 31581 64238 31633 64244
rect 31633 64238 31635 64244
rect 31579 64226 31635 64238
rect 31579 64188 31581 64226
rect 31581 64188 31633 64226
rect 31633 64188 31635 64226
rect -9851 63396 -9795 63398
rect -9771 63396 -9715 63398
rect -9691 63396 -9635 63398
rect -9611 63396 -9555 63398
rect -9531 63396 -9475 63398
rect -9851 63344 -9829 63396
rect -9829 63344 -9817 63396
rect -9817 63344 -9795 63396
rect -9771 63344 -9765 63396
rect -9765 63344 -9753 63396
rect -9753 63344 -9715 63396
rect -9691 63344 -9689 63396
rect -9689 63344 -9637 63396
rect -9637 63344 -9635 63396
rect -9611 63344 -9573 63396
rect -9573 63344 -9561 63396
rect -9561 63344 -9555 63396
rect -9531 63344 -9509 63396
rect -9509 63344 -9497 63396
rect -9497 63344 -9475 63396
rect -9851 63342 -9795 63344
rect -9771 63342 -9715 63344
rect -9691 63342 -9635 63344
rect -9611 63342 -9555 63344
rect -9531 63342 -9475 63344
rect -8040 63398 -7984 63400
rect -7960 63398 -7904 63400
rect -7880 63398 -7824 63400
rect -7800 63398 -7744 63400
rect -7720 63398 -7664 63400
rect -8040 63346 -8018 63398
rect -8018 63346 -8006 63398
rect -8006 63346 -7984 63398
rect -7960 63346 -7954 63398
rect -7954 63346 -7942 63398
rect -7942 63346 -7904 63398
rect -7880 63346 -7878 63398
rect -7878 63346 -7826 63398
rect -7826 63346 -7824 63398
rect -7800 63346 -7762 63398
rect -7762 63346 -7750 63398
rect -7750 63346 -7744 63398
rect -7720 63346 -7698 63398
rect -7698 63346 -7686 63398
rect -7686 63346 -7664 63398
rect -8040 63344 -7984 63346
rect -7960 63344 -7904 63346
rect -7880 63344 -7824 63346
rect -7800 63344 -7744 63346
rect -7720 63344 -7664 63346
rect -6245 63394 -6189 63396
rect -6165 63394 -6109 63396
rect -6085 63394 -6029 63396
rect -6005 63394 -5949 63396
rect -5925 63394 -5869 63396
rect -6245 63342 -6223 63394
rect -6223 63342 -6211 63394
rect -6211 63342 -6189 63394
rect -6165 63342 -6159 63394
rect -6159 63342 -6147 63394
rect -6147 63342 -6109 63394
rect -6085 63342 -6083 63394
rect -6083 63342 -6031 63394
rect -6031 63342 -6029 63394
rect -6005 63342 -5967 63394
rect -5967 63342 -5955 63394
rect -5955 63342 -5949 63394
rect -5925 63342 -5903 63394
rect -5903 63342 -5891 63394
rect -5891 63342 -5869 63394
rect -6245 63340 -6189 63342
rect -6165 63340 -6109 63342
rect -6085 63340 -6029 63342
rect -6005 63340 -5949 63342
rect -5925 63340 -5869 63342
rect -4446 63392 -4390 63394
rect -4366 63392 -4310 63394
rect -4286 63392 -4230 63394
rect -4206 63392 -4150 63394
rect -4126 63392 -4070 63394
rect -4446 63340 -4424 63392
rect -4424 63340 -4412 63392
rect -4412 63340 -4390 63392
rect -4366 63340 -4360 63392
rect -4360 63340 -4348 63392
rect -4348 63340 -4310 63392
rect -4286 63340 -4284 63392
rect -4284 63340 -4232 63392
rect -4232 63340 -4230 63392
rect -4206 63340 -4168 63392
rect -4168 63340 -4156 63392
rect -4156 63340 -4150 63392
rect -4126 63340 -4104 63392
rect -4104 63340 -4092 63392
rect -4092 63340 -4070 63392
rect -4446 63338 -4390 63340
rect -4366 63338 -4310 63340
rect -4286 63338 -4230 63340
rect -4206 63338 -4150 63340
rect -4126 63338 -4070 63340
rect -2655 63396 -2599 63398
rect -2575 63396 -2519 63398
rect -2495 63396 -2439 63398
rect -2415 63396 -2359 63398
rect -2335 63396 -2279 63398
rect -2655 63344 -2633 63396
rect -2633 63344 -2621 63396
rect -2621 63344 -2599 63396
rect -2575 63344 -2569 63396
rect -2569 63344 -2557 63396
rect -2557 63344 -2519 63396
rect -2495 63344 -2493 63396
rect -2493 63344 -2441 63396
rect -2441 63344 -2439 63396
rect -2415 63344 -2377 63396
rect -2377 63344 -2365 63396
rect -2365 63344 -2359 63396
rect -2335 63344 -2313 63396
rect -2313 63344 -2301 63396
rect -2301 63344 -2279 63396
rect -2655 63342 -2599 63344
rect -2575 63342 -2519 63344
rect -2495 63342 -2439 63344
rect -2415 63342 -2359 63344
rect -2335 63342 -2279 63344
rect -853 63392 -797 63394
rect -773 63392 -717 63394
rect -693 63392 -637 63394
rect -613 63392 -557 63394
rect -533 63392 -477 63394
rect -853 63340 -831 63392
rect -831 63340 -819 63392
rect -819 63340 -797 63392
rect -773 63340 -767 63392
rect -767 63340 -755 63392
rect -755 63340 -717 63392
rect -693 63340 -691 63392
rect -691 63340 -639 63392
rect -639 63340 -637 63392
rect -613 63340 -575 63392
rect -575 63340 -563 63392
rect -563 63340 -557 63392
rect -533 63340 -511 63392
rect -511 63340 -499 63392
rect -499 63340 -477 63392
rect -853 63338 -797 63340
rect -773 63338 -717 63340
rect -693 63338 -637 63340
rect -613 63338 -557 63340
rect -533 63338 -477 63340
rect -6927 63176 -6711 63194
rect -6927 62996 -6909 63176
rect -6909 62996 -6729 63176
rect -6729 62996 -6711 63176
rect -6927 62978 -6711 62996
rect 794 63202 1250 63220
rect 794 63022 1250 63202
rect 794 63004 1250 63022
rect 17980 62683 17982 62721
rect 17982 62683 18034 62721
rect 18034 62683 18036 62721
rect 17980 62671 18036 62683
rect 17980 62665 17982 62671
rect 17982 62665 18034 62671
rect 18034 62665 18036 62671
rect 17980 62619 17982 62641
rect 17982 62619 18034 62641
rect 18034 62619 18036 62641
rect 17980 62607 18036 62619
rect 17980 62585 17982 62607
rect 17982 62585 18034 62607
rect 18034 62585 18036 62607
rect 17980 62555 17982 62561
rect 17982 62555 18034 62561
rect 18034 62555 18036 62561
rect 17980 62543 18036 62555
rect 17980 62505 17982 62543
rect 17982 62505 18034 62543
rect 18034 62505 18036 62543
rect 17980 62479 18036 62481
rect 17980 62427 17982 62479
rect 17982 62427 18034 62479
rect 18034 62427 18036 62479
rect 17980 62425 18036 62427
rect 17980 62363 17982 62401
rect 17982 62363 18034 62401
rect 18034 62363 18036 62401
rect 17980 62351 18036 62363
rect 17980 62345 17982 62351
rect 17982 62345 18034 62351
rect 18034 62345 18036 62351
rect 17980 62299 17982 62321
rect 17982 62299 18034 62321
rect 18034 62299 18036 62321
rect 17980 62287 18036 62299
rect 17980 62265 17982 62287
rect 17982 62265 18034 62287
rect 18034 62265 18036 62287
rect 17980 62235 17982 62241
rect 17982 62235 18034 62241
rect 18034 62235 18036 62241
rect 17980 62223 18036 62235
rect 17980 62185 17982 62223
rect 17982 62185 18034 62223
rect 18034 62185 18036 62223
rect 19068 62683 19070 62721
rect 19070 62683 19122 62721
rect 19122 62683 19124 62721
rect 19068 62671 19124 62683
rect 19068 62665 19070 62671
rect 19070 62665 19122 62671
rect 19122 62665 19124 62671
rect 19068 62619 19070 62641
rect 19070 62619 19122 62641
rect 19122 62619 19124 62641
rect 19068 62607 19124 62619
rect 19068 62585 19070 62607
rect 19070 62585 19122 62607
rect 19122 62585 19124 62607
rect 19068 62555 19070 62561
rect 19070 62555 19122 62561
rect 19122 62555 19124 62561
rect 19068 62543 19124 62555
rect 19068 62505 19070 62543
rect 19070 62505 19122 62543
rect 19122 62505 19124 62543
rect 19068 62479 19124 62481
rect 19068 62427 19070 62479
rect 19070 62427 19122 62479
rect 19122 62427 19124 62479
rect 19068 62425 19124 62427
rect 19068 62363 19070 62401
rect 19070 62363 19122 62401
rect 19122 62363 19124 62401
rect 19068 62351 19124 62363
rect 19068 62345 19070 62351
rect 19070 62345 19122 62351
rect 19122 62345 19124 62351
rect 19068 62299 19070 62321
rect 19070 62299 19122 62321
rect 19122 62299 19124 62321
rect 19068 62287 19124 62299
rect 19068 62265 19070 62287
rect 19070 62265 19122 62287
rect 19122 62265 19124 62287
rect 19068 62235 19070 62241
rect 19070 62235 19122 62241
rect 19122 62235 19124 62241
rect 19068 62223 19124 62235
rect 19068 62185 19070 62223
rect 19070 62185 19122 62223
rect 19122 62185 19124 62223
rect 21244 62683 21246 62721
rect 21246 62683 21298 62721
rect 21298 62683 21300 62721
rect 21244 62671 21300 62683
rect 21244 62665 21246 62671
rect 21246 62665 21298 62671
rect 21298 62665 21300 62671
rect 21244 62619 21246 62641
rect 21246 62619 21298 62641
rect 21298 62619 21300 62641
rect 21244 62607 21300 62619
rect 21244 62585 21246 62607
rect 21246 62585 21298 62607
rect 21298 62585 21300 62607
rect 21244 62555 21246 62561
rect 21246 62555 21298 62561
rect 21298 62555 21300 62561
rect 21244 62543 21300 62555
rect 21244 62505 21246 62543
rect 21246 62505 21298 62543
rect 21298 62505 21300 62543
rect 21244 62479 21300 62481
rect 21244 62427 21246 62479
rect 21246 62427 21298 62479
rect 21298 62427 21300 62479
rect 21244 62425 21300 62427
rect 21244 62363 21246 62401
rect 21246 62363 21298 62401
rect 21298 62363 21300 62401
rect 21244 62351 21300 62363
rect 21244 62345 21246 62351
rect 21246 62345 21298 62351
rect 21298 62345 21300 62351
rect 21244 62299 21246 62321
rect 21246 62299 21298 62321
rect 21298 62299 21300 62321
rect 21244 62287 21300 62299
rect 21244 62265 21246 62287
rect 21246 62265 21298 62287
rect 21298 62265 21300 62287
rect 21244 62235 21246 62241
rect 21246 62235 21298 62241
rect 21298 62235 21300 62241
rect 21244 62223 21300 62235
rect 21244 62185 21246 62223
rect 21246 62185 21298 62223
rect 21298 62185 21300 62223
rect 22332 62683 22334 62721
rect 22334 62683 22386 62721
rect 22386 62683 22388 62721
rect 22332 62671 22388 62683
rect 22332 62665 22334 62671
rect 22334 62665 22386 62671
rect 22386 62665 22388 62671
rect 22332 62619 22334 62641
rect 22334 62619 22386 62641
rect 22386 62619 22388 62641
rect 22332 62607 22388 62619
rect 22332 62585 22334 62607
rect 22334 62585 22386 62607
rect 22386 62585 22388 62607
rect 22332 62555 22334 62561
rect 22334 62555 22386 62561
rect 22386 62555 22388 62561
rect 22332 62543 22388 62555
rect 22332 62505 22334 62543
rect 22334 62505 22386 62543
rect 22386 62505 22388 62543
rect 22332 62479 22388 62481
rect 22332 62427 22334 62479
rect 22334 62427 22386 62479
rect 22386 62427 22388 62479
rect 22332 62425 22388 62427
rect 22332 62363 22334 62401
rect 22334 62363 22386 62401
rect 22386 62363 22388 62401
rect 22332 62351 22388 62363
rect 22332 62345 22334 62351
rect 22334 62345 22386 62351
rect 22386 62345 22388 62351
rect 22332 62299 22334 62321
rect 22334 62299 22386 62321
rect 22386 62299 22388 62321
rect 22332 62287 22388 62299
rect 22332 62265 22334 62287
rect 22334 62265 22386 62287
rect 22386 62265 22388 62287
rect 22332 62235 22334 62241
rect 22334 62235 22386 62241
rect 22386 62235 22388 62241
rect 22332 62223 22388 62235
rect 22332 62185 22334 62223
rect 22334 62185 22386 62223
rect 22386 62185 22388 62223
rect 23420 62683 23422 62721
rect 23422 62683 23474 62721
rect 23474 62683 23476 62721
rect 23420 62671 23476 62683
rect 23420 62665 23422 62671
rect 23422 62665 23474 62671
rect 23474 62665 23476 62671
rect 23420 62619 23422 62641
rect 23422 62619 23474 62641
rect 23474 62619 23476 62641
rect 23420 62607 23476 62619
rect 23420 62585 23422 62607
rect 23422 62585 23474 62607
rect 23474 62585 23476 62607
rect 23420 62555 23422 62561
rect 23422 62555 23474 62561
rect 23474 62555 23476 62561
rect 23420 62543 23476 62555
rect 23420 62505 23422 62543
rect 23422 62505 23474 62543
rect 23474 62505 23476 62543
rect 23420 62479 23476 62481
rect 23420 62427 23422 62479
rect 23422 62427 23474 62479
rect 23474 62427 23476 62479
rect 23420 62425 23476 62427
rect 23420 62363 23422 62401
rect 23422 62363 23474 62401
rect 23474 62363 23476 62401
rect 23420 62351 23476 62363
rect 23420 62345 23422 62351
rect 23422 62345 23474 62351
rect 23474 62345 23476 62351
rect 23420 62299 23422 62321
rect 23422 62299 23474 62321
rect 23474 62299 23476 62321
rect 23420 62287 23476 62299
rect 23420 62265 23422 62287
rect 23422 62265 23474 62287
rect 23474 62265 23476 62287
rect 23420 62235 23422 62241
rect 23422 62235 23474 62241
rect 23474 62235 23476 62241
rect 23420 62223 23476 62235
rect 23420 62185 23422 62223
rect 23422 62185 23474 62223
rect 23474 62185 23476 62223
rect 24508 62683 24510 62721
rect 24510 62683 24562 62721
rect 24562 62683 24564 62721
rect 24508 62671 24564 62683
rect 24508 62665 24510 62671
rect 24510 62665 24562 62671
rect 24562 62665 24564 62671
rect 24508 62619 24510 62641
rect 24510 62619 24562 62641
rect 24562 62619 24564 62641
rect 24508 62607 24564 62619
rect 24508 62585 24510 62607
rect 24510 62585 24562 62607
rect 24562 62585 24564 62607
rect 24508 62555 24510 62561
rect 24510 62555 24562 62561
rect 24562 62555 24564 62561
rect 24508 62543 24564 62555
rect 24508 62505 24510 62543
rect 24510 62505 24562 62543
rect 24562 62505 24564 62543
rect 24508 62479 24564 62481
rect 24508 62427 24510 62479
rect 24510 62427 24562 62479
rect 24562 62427 24564 62479
rect 24508 62425 24564 62427
rect 24508 62363 24510 62401
rect 24510 62363 24562 62401
rect 24562 62363 24564 62401
rect 24508 62351 24564 62363
rect 24508 62345 24510 62351
rect 24510 62345 24562 62351
rect 24562 62345 24564 62351
rect 24508 62299 24510 62321
rect 24510 62299 24562 62321
rect 24562 62299 24564 62321
rect 24508 62287 24564 62299
rect 24508 62265 24510 62287
rect 24510 62265 24562 62287
rect 24562 62265 24564 62287
rect 24508 62235 24510 62241
rect 24510 62235 24562 62241
rect 24562 62235 24564 62241
rect 24508 62223 24564 62235
rect 24508 62185 24510 62223
rect 24510 62185 24562 62223
rect 24562 62185 24564 62223
rect 25596 62683 25598 62721
rect 25598 62683 25650 62721
rect 25650 62683 25652 62721
rect 25596 62671 25652 62683
rect 25596 62665 25598 62671
rect 25598 62665 25650 62671
rect 25650 62665 25652 62671
rect 25596 62619 25598 62641
rect 25598 62619 25650 62641
rect 25650 62619 25652 62641
rect 25596 62607 25652 62619
rect 25596 62585 25598 62607
rect 25598 62585 25650 62607
rect 25650 62585 25652 62607
rect 25596 62555 25598 62561
rect 25598 62555 25650 62561
rect 25650 62555 25652 62561
rect 25596 62543 25652 62555
rect 25596 62505 25598 62543
rect 25598 62505 25650 62543
rect 25650 62505 25652 62543
rect 25596 62479 25652 62481
rect 25596 62427 25598 62479
rect 25598 62427 25650 62479
rect 25650 62427 25652 62479
rect 25596 62425 25652 62427
rect 25596 62363 25598 62401
rect 25598 62363 25650 62401
rect 25650 62363 25652 62401
rect 25596 62351 25652 62363
rect 25596 62345 25598 62351
rect 25598 62345 25650 62351
rect 25650 62345 25652 62351
rect 25596 62299 25598 62321
rect 25598 62299 25650 62321
rect 25650 62299 25652 62321
rect 25596 62287 25652 62299
rect 25596 62265 25598 62287
rect 25598 62265 25650 62287
rect 25650 62265 25652 62287
rect 25596 62235 25598 62241
rect 25598 62235 25650 62241
rect 25650 62235 25652 62241
rect 25596 62223 25652 62235
rect 25596 62185 25598 62223
rect 25598 62185 25650 62223
rect 25650 62185 25652 62223
rect 26684 62683 26686 62721
rect 26686 62683 26738 62721
rect 26738 62683 26740 62721
rect 26684 62671 26740 62683
rect 26684 62665 26686 62671
rect 26686 62665 26738 62671
rect 26738 62665 26740 62671
rect 26684 62619 26686 62641
rect 26686 62619 26738 62641
rect 26738 62619 26740 62641
rect 26684 62607 26740 62619
rect 26684 62585 26686 62607
rect 26686 62585 26738 62607
rect 26738 62585 26740 62607
rect 26684 62555 26686 62561
rect 26686 62555 26738 62561
rect 26738 62555 26740 62561
rect 26684 62543 26740 62555
rect 26684 62505 26686 62543
rect 26686 62505 26738 62543
rect 26738 62505 26740 62543
rect 26684 62479 26740 62481
rect 26684 62427 26686 62479
rect 26686 62427 26738 62479
rect 26738 62427 26740 62479
rect 26684 62425 26740 62427
rect 26684 62363 26686 62401
rect 26686 62363 26738 62401
rect 26738 62363 26740 62401
rect 26684 62351 26740 62363
rect 26684 62345 26686 62351
rect 26686 62345 26738 62351
rect 26738 62345 26740 62351
rect 26684 62299 26686 62321
rect 26686 62299 26738 62321
rect 26738 62299 26740 62321
rect 26684 62287 26740 62299
rect 26684 62265 26686 62287
rect 26686 62265 26738 62287
rect 26738 62265 26740 62287
rect 26684 62235 26686 62241
rect 26686 62235 26738 62241
rect 26738 62235 26740 62241
rect 26684 62223 26740 62235
rect 26684 62185 26686 62223
rect 26686 62185 26738 62223
rect 26738 62185 26740 62223
rect 28860 62683 28862 62721
rect 28862 62683 28914 62721
rect 28914 62683 28916 62721
rect 28860 62671 28916 62683
rect 28860 62665 28862 62671
rect 28862 62665 28914 62671
rect 28914 62665 28916 62671
rect 28860 62619 28862 62641
rect 28862 62619 28914 62641
rect 28914 62619 28916 62641
rect 28860 62607 28916 62619
rect 28860 62585 28862 62607
rect 28862 62585 28914 62607
rect 28914 62585 28916 62607
rect 28860 62555 28862 62561
rect 28862 62555 28914 62561
rect 28914 62555 28916 62561
rect 28860 62543 28916 62555
rect 28860 62505 28862 62543
rect 28862 62505 28914 62543
rect 28914 62505 28916 62543
rect 28860 62479 28916 62481
rect 28860 62427 28862 62479
rect 28862 62427 28914 62479
rect 28914 62427 28916 62479
rect 28860 62425 28916 62427
rect 28860 62363 28862 62401
rect 28862 62363 28914 62401
rect 28914 62363 28916 62401
rect 28860 62351 28916 62363
rect 28860 62345 28862 62351
rect 28862 62345 28914 62351
rect 28914 62345 28916 62351
rect 28860 62299 28862 62321
rect 28862 62299 28914 62321
rect 28914 62299 28916 62321
rect 28860 62287 28916 62299
rect 28860 62265 28862 62287
rect 28862 62265 28914 62287
rect 28914 62265 28916 62287
rect 28860 62235 28862 62241
rect 28862 62235 28914 62241
rect 28914 62235 28916 62241
rect 28860 62223 28916 62235
rect 28860 62185 28862 62223
rect 28862 62185 28914 62223
rect 28914 62185 28916 62223
rect 29948 62683 29950 62721
rect 29950 62683 30002 62721
rect 30002 62683 30004 62721
rect 29948 62671 30004 62683
rect 29948 62665 29950 62671
rect 29950 62665 30002 62671
rect 30002 62665 30004 62671
rect 29948 62619 29950 62641
rect 29950 62619 30002 62641
rect 30002 62619 30004 62641
rect 29948 62607 30004 62619
rect 29948 62585 29950 62607
rect 29950 62585 30002 62607
rect 30002 62585 30004 62607
rect 29948 62555 29950 62561
rect 29950 62555 30002 62561
rect 30002 62555 30004 62561
rect 29948 62543 30004 62555
rect 29948 62505 29950 62543
rect 29950 62505 30002 62543
rect 30002 62505 30004 62543
rect 29948 62479 30004 62481
rect 29948 62427 29950 62479
rect 29950 62427 30002 62479
rect 30002 62427 30004 62479
rect 29948 62425 30004 62427
rect 29948 62363 29950 62401
rect 29950 62363 30002 62401
rect 30002 62363 30004 62401
rect 29948 62351 30004 62363
rect 29948 62345 29950 62351
rect 29950 62345 30002 62351
rect 30002 62345 30004 62351
rect 29948 62299 29950 62321
rect 29950 62299 30002 62321
rect 30002 62299 30004 62321
rect 29948 62287 30004 62299
rect 29948 62265 29950 62287
rect 29950 62265 30002 62287
rect 30002 62265 30004 62287
rect 29948 62235 29950 62241
rect 29950 62235 30002 62241
rect 30002 62235 30004 62241
rect 29948 62223 30004 62235
rect 29948 62185 29950 62223
rect 29950 62185 30002 62223
rect 30002 62185 30004 62223
rect 31036 62683 31038 62721
rect 31038 62683 31090 62721
rect 31090 62683 31092 62721
rect 31036 62671 31092 62683
rect 31036 62665 31038 62671
rect 31038 62665 31090 62671
rect 31090 62665 31092 62671
rect 31036 62619 31038 62641
rect 31038 62619 31090 62641
rect 31090 62619 31092 62641
rect 31036 62607 31092 62619
rect 31036 62585 31038 62607
rect 31038 62585 31090 62607
rect 31090 62585 31092 62607
rect 31036 62555 31038 62561
rect 31038 62555 31090 62561
rect 31090 62555 31092 62561
rect 31036 62543 31092 62555
rect 31036 62505 31038 62543
rect 31038 62505 31090 62543
rect 31090 62505 31092 62543
rect 31036 62479 31092 62481
rect 31036 62427 31038 62479
rect 31038 62427 31090 62479
rect 31090 62427 31092 62479
rect 31036 62425 31092 62427
rect 31036 62363 31038 62401
rect 31038 62363 31090 62401
rect 31090 62363 31092 62401
rect 31036 62351 31092 62363
rect 31036 62345 31038 62351
rect 31038 62345 31090 62351
rect 31090 62345 31092 62351
rect 31036 62299 31038 62321
rect 31038 62299 31090 62321
rect 31090 62299 31092 62321
rect 31036 62287 31092 62299
rect 31036 62265 31038 62287
rect 31038 62265 31090 62287
rect 31090 62265 31092 62287
rect 31036 62235 31038 62241
rect 31038 62235 31090 62241
rect 31090 62235 31092 62241
rect 31036 62223 31092 62235
rect 31036 62185 31038 62223
rect 31038 62185 31090 62223
rect 31090 62185 31092 62223
rect -8553 54589 -8497 54591
rect -8553 54537 -8551 54589
rect -8551 54537 -8499 54589
rect -8499 54537 -8497 54589
rect -8553 54535 -8497 54537
rect -6862 54590 -6806 54592
rect -6862 54538 -6860 54590
rect -6860 54538 -6808 54590
rect -6808 54538 -6806 54590
rect -6862 54536 -6806 54538
rect -5157 54589 -5101 54591
rect -5157 54537 -5155 54589
rect -5155 54537 -5103 54589
rect -5103 54537 -5101 54589
rect -5157 54535 -5101 54537
rect -3361 54589 -3305 54591
rect -3361 54537 -3359 54589
rect -3359 54537 -3307 54589
rect -3307 54537 -3305 54589
rect -3361 54535 -3305 54537
rect -1532 54589 -1476 54591
rect -1532 54537 -1530 54589
rect -1530 54537 -1478 54589
rect -1478 54537 -1476 54589
rect -1532 54535 -1476 54537
rect -9691 54397 -9635 54399
rect -9611 54397 -9555 54399
rect -9531 54397 -9475 54399
rect -9691 54345 -9673 54397
rect -9673 54345 -9635 54397
rect -9611 54345 -9609 54397
rect -9609 54345 -9557 54397
rect -9557 54345 -9555 54397
rect -9531 54345 -9493 54397
rect -9493 54345 -9475 54397
rect -9691 54343 -9635 54345
rect -9611 54343 -9555 54345
rect -9531 54343 -9475 54345
rect -7896 54396 -7840 54398
rect -7816 54396 -7760 54398
rect -7736 54396 -7680 54398
rect -7896 54344 -7878 54396
rect -7878 54344 -7840 54396
rect -7816 54344 -7814 54396
rect -7814 54344 -7762 54396
rect -7762 54344 -7760 54396
rect -7736 54344 -7698 54396
rect -7698 54344 -7680 54396
rect -7896 54342 -7840 54344
rect -7816 54342 -7760 54344
rect -7736 54342 -7680 54344
rect -6096 54398 -6040 54400
rect -6016 54398 -5960 54400
rect -5936 54398 -5880 54400
rect -6096 54346 -6078 54398
rect -6078 54346 -6040 54398
rect -6016 54346 -6014 54398
rect -6014 54346 -5962 54398
rect -5962 54346 -5960 54398
rect -5936 54346 -5898 54398
rect -5898 54346 -5880 54398
rect -6096 54344 -6040 54346
rect -6016 54344 -5960 54346
rect -5936 54344 -5880 54346
rect -4298 54397 -4242 54399
rect -4218 54397 -4162 54399
rect -4138 54397 -4082 54399
rect -4298 54345 -4280 54397
rect -4280 54345 -4242 54397
rect -4218 54345 -4216 54397
rect -4216 54345 -4164 54397
rect -4164 54345 -4162 54397
rect -4138 54345 -4100 54397
rect -4100 54345 -4082 54397
rect -4298 54343 -4242 54345
rect -4218 54343 -4162 54345
rect -4138 54343 -4082 54345
rect -2500 54398 -2444 54400
rect -2420 54398 -2364 54400
rect -2340 54398 -2284 54400
rect -2500 54346 -2482 54398
rect -2482 54346 -2444 54398
rect -2420 54346 -2418 54398
rect -2418 54346 -2366 54398
rect -2366 54346 -2364 54398
rect -2340 54346 -2302 54398
rect -2302 54346 -2284 54398
rect -2500 54344 -2444 54346
rect -2420 54344 -2364 54346
rect -2340 54344 -2284 54346
rect -697 54397 -641 54399
rect -617 54397 -561 54399
rect -537 54397 -481 54399
rect -697 54345 -679 54397
rect -679 54345 -641 54397
rect -617 54345 -615 54397
rect -615 54345 -563 54397
rect -563 54345 -561 54397
rect -537 54345 -499 54397
rect -499 54345 -481 54397
rect -697 54343 -641 54345
rect -617 54343 -561 54345
rect -537 54343 -481 54345
rect 180 54398 236 54400
rect 180 54346 182 54398
rect 182 54346 234 54398
rect 234 54346 236 54398
rect 180 54344 236 54346
rect -8840 51221 -8784 51239
rect -8840 51183 -8838 51221
rect -8838 51183 -8786 51221
rect -8786 51183 -8784 51221
rect -7718 51187 -7662 51243
rect -8840 51157 -8784 51159
rect -8840 51105 -8838 51157
rect -8838 51105 -8786 51157
rect -8786 51105 -8784 51157
rect -8840 51103 -8784 51105
rect -8840 51041 -8838 51079
rect -8838 51041 -8786 51079
rect -8786 51041 -8784 51079
rect -8840 51023 -8784 51041
rect -27046 49714 -26990 49716
rect -26966 49714 -26910 49716
rect -26886 49714 -26830 49716
rect -26806 49714 -26750 49716
rect -27046 49662 -27000 49714
rect -27000 49662 -26990 49714
rect -26966 49662 -26936 49714
rect -26936 49662 -26924 49714
rect -26924 49662 -26910 49714
rect -26886 49662 -26872 49714
rect -26872 49662 -26860 49714
rect -26860 49662 -26830 49714
rect -26806 49662 -26796 49714
rect -26796 49662 -26750 49714
rect -27046 49660 -26990 49662
rect -26966 49660 -26910 49662
rect -26886 49660 -26830 49662
rect -26806 49660 -26750 49662
rect -26391 49407 -26335 49409
rect -26311 49407 -26255 49409
rect -26231 49407 -26175 49409
rect -26391 49355 -26353 49407
rect -26353 49355 -26341 49407
rect -26341 49355 -26335 49407
rect -26311 49355 -26289 49407
rect -26289 49355 -26277 49407
rect -26277 49355 -26255 49407
rect -26231 49355 -26225 49407
rect -26225 49355 -26213 49407
rect -26213 49355 -26175 49407
rect -26391 49353 -26335 49355
rect -26311 49353 -26255 49355
rect -26231 49353 -26175 49355
rect -26056 49418 -26000 49420
rect -26056 49366 -26054 49418
rect -26054 49366 -26002 49418
rect -26002 49366 -26000 49418
rect -26056 49364 -26000 49366
rect -25960 49172 -25904 49174
rect -25880 49172 -25824 49174
rect -25800 49172 -25744 49174
rect -25720 49172 -25664 49174
rect -25960 49120 -25914 49172
rect -25914 49120 -25904 49172
rect -25880 49120 -25850 49172
rect -25850 49120 -25838 49172
rect -25838 49120 -25824 49172
rect -25800 49120 -25786 49172
rect -25786 49120 -25774 49172
rect -25774 49120 -25744 49172
rect -25720 49120 -25710 49172
rect -25710 49120 -25664 49172
rect -25960 49118 -25904 49120
rect -25880 49118 -25824 49120
rect -25800 49118 -25744 49120
rect -25720 49118 -25664 49120
rect -27067 43244 -27065 43274
rect -27065 43244 -27013 43274
rect -27013 43244 -27011 43274
rect -27067 43232 -27011 43244
rect -27067 43218 -27065 43232
rect -27065 43218 -27013 43232
rect -27013 43218 -27011 43232
rect -27067 43180 -27065 43194
rect -27065 43180 -27013 43194
rect -27013 43180 -27011 43194
rect -27067 43168 -27011 43180
rect -27067 43138 -27065 43168
rect -27065 43138 -27013 43168
rect -27013 43138 -27011 43168
rect -27067 43104 -27011 43114
rect -27067 43058 -27065 43104
rect -27065 43058 -27013 43104
rect -27013 43058 -27011 43104
rect -27067 42988 -27065 43034
rect -27065 42988 -27013 43034
rect -27013 42988 -27011 43034
rect -27067 42978 -27011 42988
rect -13465 43055 -13409 43057
rect -13465 43003 -13463 43055
rect -13463 43003 -13411 43055
rect -13411 43003 -13409 43055
rect -13465 43001 -13409 43003
rect -27067 42924 -27065 42954
rect -27065 42924 -27013 42954
rect -27013 42924 -27011 42954
rect -27067 42912 -27011 42924
rect -27067 42898 -27065 42912
rect -27065 42898 -27013 42912
rect -27013 42898 -27011 42912
rect -27067 42860 -27065 42874
rect -27065 42860 -27013 42874
rect -27013 42860 -27011 42874
rect -27067 42848 -27011 42860
rect -27067 42818 -27065 42848
rect -27065 42818 -27013 42848
rect -27013 42818 -27011 42848
rect -12689 42392 -12633 42394
rect -12689 42340 -12687 42392
rect -12687 42340 -12635 42392
rect -12635 42340 -12633 42392
rect -12689 42338 -12633 42340
rect -27067 42103 -27065 42133
rect -27065 42103 -27013 42133
rect -27013 42103 -27011 42133
rect -27067 42091 -27011 42103
rect -27067 42077 -27065 42091
rect -27065 42077 -27013 42091
rect -27013 42077 -27011 42091
rect -21471 42103 -21415 42159
rect -27067 42039 -27065 42053
rect -27065 42039 -27013 42053
rect -27013 42039 -27011 42053
rect -27067 42027 -27011 42039
rect -27067 41997 -27065 42027
rect -27065 41997 -27013 42027
rect -27013 41997 -27011 42027
rect -27067 41963 -27011 41973
rect -27067 41917 -27065 41963
rect -27065 41917 -27013 41963
rect -27013 41917 -27011 41963
rect -27067 41847 -27065 41893
rect -27065 41847 -27013 41893
rect -27013 41847 -27011 41893
rect -27067 41837 -27011 41847
rect -27067 41783 -27065 41813
rect -27065 41783 -27013 41813
rect -27013 41783 -27011 41813
rect -27067 41771 -27011 41783
rect -27067 41757 -27065 41771
rect -27065 41757 -27013 41771
rect -27013 41757 -27011 41771
rect -27067 41719 -27065 41733
rect -27065 41719 -27013 41733
rect -27013 41719 -27011 41733
rect -27067 41707 -27011 41719
rect -27067 41677 -27065 41707
rect -27065 41677 -27013 41707
rect -27013 41677 -27011 41707
rect -27067 41643 -27011 41653
rect -27067 41597 -27065 41643
rect -27065 41597 -27013 41643
rect -27013 41597 -27011 41643
rect -27067 41527 -27065 41573
rect -27065 41527 -27013 41573
rect -27013 41527 -27011 41573
rect -27067 41517 -27011 41527
rect -27067 41463 -27065 41493
rect -27065 41463 -27013 41493
rect -27013 41463 -27011 41493
rect -27067 41451 -27011 41463
rect -27067 41437 -27065 41451
rect -27065 41437 -27013 41451
rect -27013 41437 -27011 41451
rect -27067 41399 -27065 41413
rect -27065 41399 -27013 41413
rect -27013 41399 -27011 41413
rect -27067 41387 -27011 41399
rect -27067 41357 -27065 41387
rect -27065 41357 -27013 41387
rect -27013 41357 -27011 41387
rect -27067 41323 -27011 41333
rect -27067 41277 -27065 41323
rect -27065 41277 -27013 41323
rect -27013 41277 -27011 41323
rect -27067 41207 -27065 41253
rect -27065 41207 -27013 41253
rect -27013 41207 -27011 41253
rect -27067 41197 -27011 41207
rect -27067 41143 -27065 41173
rect -27065 41143 -27013 41173
rect -27013 41143 -27011 41173
rect -27067 41131 -27011 41143
rect -27067 41117 -27065 41131
rect -27065 41117 -27013 41131
rect -27013 41117 -27011 41131
rect -27067 41079 -27065 41093
rect -27065 41079 -27013 41093
rect -27013 41079 -27011 41093
rect -27067 41067 -27011 41079
rect -27067 41037 -27065 41067
rect -27065 41037 -27013 41067
rect -27013 41037 -27011 41067
rect -27062 40577 -27060 40607
rect -27060 40577 -27008 40607
rect -27008 40577 -27006 40607
rect -27062 40565 -27006 40577
rect -27062 40551 -27060 40565
rect -27060 40551 -27008 40565
rect -27008 40551 -27006 40565
rect -27062 40513 -27060 40527
rect -27060 40513 -27008 40527
rect -27008 40513 -27006 40527
rect -27062 40501 -27006 40513
rect -27062 40471 -27060 40501
rect -27060 40471 -27008 40501
rect -27008 40471 -27006 40501
rect -27062 40437 -27006 40447
rect -27062 40391 -27060 40437
rect -27060 40391 -27008 40437
rect -27008 40391 -27006 40437
rect -27062 40321 -27060 40367
rect -27060 40321 -27008 40367
rect -27008 40321 -27006 40367
rect -27062 40311 -27006 40321
rect -27062 40257 -27060 40287
rect -27060 40257 -27008 40287
rect -27008 40257 -27006 40287
rect -27062 40245 -27006 40257
rect -27062 40231 -27060 40245
rect -27060 40231 -27008 40245
rect -27008 40231 -27006 40245
rect -27062 40193 -27060 40207
rect -27060 40193 -27008 40207
rect -27008 40193 -27006 40207
rect -27062 40181 -27006 40193
rect -27062 40151 -27060 40181
rect -27060 40151 -27008 40181
rect -27008 40151 -27006 40181
rect -27062 40117 -27006 40127
rect -27062 40071 -27060 40117
rect -27060 40071 -27008 40117
rect -27008 40071 -27006 40117
rect -27062 40001 -27060 40047
rect -27060 40001 -27008 40047
rect -27008 40001 -27006 40047
rect -27062 39991 -27006 40001
rect -27062 39937 -27060 39967
rect -27060 39937 -27008 39967
rect -27008 39937 -27006 39967
rect -27062 39925 -27006 39937
rect -27062 39911 -27060 39925
rect -27060 39911 -27008 39925
rect -27008 39911 -27006 39925
rect -27062 39873 -27060 39887
rect -27060 39873 -27008 39887
rect -27008 39873 -27006 39887
rect -27062 39861 -27006 39873
rect -27062 39831 -27060 39861
rect -27060 39831 -27008 39861
rect -27008 39831 -27006 39861
rect -27062 39797 -27006 39807
rect -27062 39751 -27060 39797
rect -27060 39751 -27008 39797
rect -27008 39751 -27006 39797
rect 365 53146 375 60802
rect 375 53146 491 60802
rect 491 53146 501 60802
rect 10216 60812 10512 60814
rect -8855 50770 -8799 50772
rect -8855 50718 -8853 50770
rect -8853 50718 -8801 50770
rect -8801 50718 -8799 50770
rect -8855 50716 -8799 50718
rect -8855 50654 -8853 50692
rect -8853 50654 -8801 50692
rect -8801 50654 -8799 50692
rect -8855 50642 -8799 50654
rect -8855 50636 -8853 50642
rect -8853 50636 -8801 50642
rect -8801 50636 -8799 50642
rect -8855 50590 -8853 50612
rect -8853 50590 -8801 50612
rect -8801 50590 -8799 50612
rect -8855 50578 -8799 50590
rect -8855 50556 -8853 50578
rect -8853 50556 -8801 50578
rect -8801 50556 -8799 50578
rect -8855 50526 -8853 50532
rect -8853 50526 -8801 50532
rect -8801 50526 -8799 50532
rect -8855 50514 -8799 50526
rect -8855 50476 -8853 50514
rect -8853 50476 -8801 50514
rect -8801 50476 -8799 50514
rect -8855 50450 -8799 50452
rect -8855 50398 -8853 50450
rect -8853 50398 -8801 50450
rect -8801 50398 -8799 50450
rect -8855 50396 -8799 50398
rect -8476 50381 -8420 50437
rect -5656 50906 -3920 51042
rect -3337 51043 -2561 51053
rect -3337 50927 -2561 51043
rect -3337 50917 -2561 50927
rect -1638 51033 -782 51043
rect -1638 50917 -782 51033
rect -1638 50907 -782 50917
rect -47 50761 89 50771
rect -5908 50714 -5772 50716
rect -5908 47782 -5772 50714
rect -5908 47780 -5772 47782
rect -47 47765 89 50761
rect -47 47755 89 47765
rect 10216 47640 10512 60812
rect 17435 60686 17437 60724
rect 17437 60686 17489 60724
rect 17489 60686 17491 60724
rect 17435 60674 17491 60686
rect 17435 60668 17437 60674
rect 17437 60668 17489 60674
rect 17489 60668 17491 60674
rect 17435 60622 17437 60644
rect 17437 60622 17489 60644
rect 17489 60622 17491 60644
rect 17435 60610 17491 60622
rect 17435 60588 17437 60610
rect 17437 60588 17489 60610
rect 17489 60588 17491 60610
rect 17435 60558 17437 60564
rect 17437 60558 17489 60564
rect 17489 60558 17491 60564
rect 17435 60546 17491 60558
rect 17435 60508 17437 60546
rect 17437 60508 17489 60546
rect 17489 60508 17491 60546
rect 17435 60482 17491 60484
rect 17435 60430 17437 60482
rect 17437 60430 17489 60482
rect 17489 60430 17491 60482
rect 17435 60428 17491 60430
rect 17435 60366 17437 60404
rect 17437 60366 17489 60404
rect 17489 60366 17491 60404
rect 17435 60354 17491 60366
rect 17435 60348 17437 60354
rect 17437 60348 17489 60354
rect 17489 60348 17491 60354
rect 17435 60302 17437 60324
rect 17437 60302 17489 60324
rect 17489 60302 17491 60324
rect 17435 60290 17491 60302
rect 17435 60268 17437 60290
rect 17437 60268 17489 60290
rect 17489 60268 17491 60290
rect 17435 60238 17437 60244
rect 17437 60238 17489 60244
rect 17489 60238 17491 60244
rect 17435 60226 17491 60238
rect 17435 60188 17437 60226
rect 17437 60188 17489 60226
rect 17489 60188 17491 60226
rect 18523 60686 18525 60724
rect 18525 60686 18577 60724
rect 18577 60686 18579 60724
rect 18523 60674 18579 60686
rect 18523 60668 18525 60674
rect 18525 60668 18577 60674
rect 18577 60668 18579 60674
rect 18523 60622 18525 60644
rect 18525 60622 18577 60644
rect 18577 60622 18579 60644
rect 18523 60610 18579 60622
rect 18523 60588 18525 60610
rect 18525 60588 18577 60610
rect 18577 60588 18579 60610
rect 18523 60558 18525 60564
rect 18525 60558 18577 60564
rect 18577 60558 18579 60564
rect 18523 60546 18579 60558
rect 18523 60508 18525 60546
rect 18525 60508 18577 60546
rect 18577 60508 18579 60546
rect 18523 60482 18579 60484
rect 18523 60430 18525 60482
rect 18525 60430 18577 60482
rect 18577 60430 18579 60482
rect 18523 60428 18579 60430
rect 18523 60366 18525 60404
rect 18525 60366 18577 60404
rect 18577 60366 18579 60404
rect 18523 60354 18579 60366
rect 18523 60348 18525 60354
rect 18525 60348 18577 60354
rect 18577 60348 18579 60354
rect 18523 60302 18525 60324
rect 18525 60302 18577 60324
rect 18577 60302 18579 60324
rect 18523 60290 18579 60302
rect 18523 60268 18525 60290
rect 18525 60268 18577 60290
rect 18577 60268 18579 60290
rect 18523 60238 18525 60244
rect 18525 60238 18577 60244
rect 18577 60238 18579 60244
rect 18523 60226 18579 60238
rect 18523 60188 18525 60226
rect 18525 60188 18577 60226
rect 18577 60188 18579 60226
rect 19611 60686 19613 60724
rect 19613 60686 19665 60724
rect 19665 60686 19667 60724
rect 19611 60674 19667 60686
rect 19611 60668 19613 60674
rect 19613 60668 19665 60674
rect 19665 60668 19667 60674
rect 19611 60622 19613 60644
rect 19613 60622 19665 60644
rect 19665 60622 19667 60644
rect 19611 60610 19667 60622
rect 19611 60588 19613 60610
rect 19613 60588 19665 60610
rect 19665 60588 19667 60610
rect 19611 60558 19613 60564
rect 19613 60558 19665 60564
rect 19665 60558 19667 60564
rect 19611 60546 19667 60558
rect 19611 60508 19613 60546
rect 19613 60508 19665 60546
rect 19665 60508 19667 60546
rect 19611 60482 19667 60484
rect 19611 60430 19613 60482
rect 19613 60430 19665 60482
rect 19665 60430 19667 60482
rect 19611 60428 19667 60430
rect 19611 60366 19613 60404
rect 19613 60366 19665 60404
rect 19665 60366 19667 60404
rect 19611 60354 19667 60366
rect 19611 60348 19613 60354
rect 19613 60348 19665 60354
rect 19665 60348 19667 60354
rect 19611 60302 19613 60324
rect 19613 60302 19665 60324
rect 19665 60302 19667 60324
rect 19611 60290 19667 60302
rect 19611 60268 19613 60290
rect 19613 60268 19665 60290
rect 19665 60268 19667 60290
rect 19611 60238 19613 60244
rect 19613 60238 19665 60244
rect 19665 60238 19667 60244
rect 19611 60226 19667 60238
rect 19611 60188 19613 60226
rect 19613 60188 19665 60226
rect 19665 60188 19667 60226
rect 20699 60686 20701 60724
rect 20701 60686 20753 60724
rect 20753 60686 20755 60724
rect 20699 60674 20755 60686
rect 20699 60668 20701 60674
rect 20701 60668 20753 60674
rect 20753 60668 20755 60674
rect 20699 60622 20701 60644
rect 20701 60622 20753 60644
rect 20753 60622 20755 60644
rect 20699 60610 20755 60622
rect 20699 60588 20701 60610
rect 20701 60588 20753 60610
rect 20753 60588 20755 60610
rect 20699 60558 20701 60564
rect 20701 60558 20753 60564
rect 20753 60558 20755 60564
rect 20699 60546 20755 60558
rect 20699 60508 20701 60546
rect 20701 60508 20753 60546
rect 20753 60508 20755 60546
rect 20699 60482 20755 60484
rect 20699 60430 20701 60482
rect 20701 60430 20753 60482
rect 20753 60430 20755 60482
rect 20699 60428 20755 60430
rect 20699 60366 20701 60404
rect 20701 60366 20753 60404
rect 20753 60366 20755 60404
rect 20699 60354 20755 60366
rect 20699 60348 20701 60354
rect 20701 60348 20753 60354
rect 20753 60348 20755 60354
rect 20699 60302 20701 60324
rect 20701 60302 20753 60324
rect 20753 60302 20755 60324
rect 20699 60290 20755 60302
rect 20699 60268 20701 60290
rect 20701 60268 20753 60290
rect 20753 60268 20755 60290
rect 20699 60238 20701 60244
rect 20701 60238 20753 60244
rect 20753 60238 20755 60244
rect 20699 60226 20755 60238
rect 20699 60188 20701 60226
rect 20701 60188 20753 60226
rect 20753 60188 20755 60226
rect 21787 60686 21789 60724
rect 21789 60686 21841 60724
rect 21841 60686 21843 60724
rect 21787 60674 21843 60686
rect 21787 60668 21789 60674
rect 21789 60668 21841 60674
rect 21841 60668 21843 60674
rect 21787 60622 21789 60644
rect 21789 60622 21841 60644
rect 21841 60622 21843 60644
rect 21787 60610 21843 60622
rect 21787 60588 21789 60610
rect 21789 60588 21841 60610
rect 21841 60588 21843 60610
rect 21787 60558 21789 60564
rect 21789 60558 21841 60564
rect 21841 60558 21843 60564
rect 21787 60546 21843 60558
rect 21787 60508 21789 60546
rect 21789 60508 21841 60546
rect 21841 60508 21843 60546
rect 21787 60482 21843 60484
rect 21787 60430 21789 60482
rect 21789 60430 21841 60482
rect 21841 60430 21843 60482
rect 21787 60428 21843 60430
rect 21787 60366 21789 60404
rect 21789 60366 21841 60404
rect 21841 60366 21843 60404
rect 21787 60354 21843 60366
rect 21787 60348 21789 60354
rect 21789 60348 21841 60354
rect 21841 60348 21843 60354
rect 21787 60302 21789 60324
rect 21789 60302 21841 60324
rect 21841 60302 21843 60324
rect 21787 60290 21843 60302
rect 21787 60268 21789 60290
rect 21789 60268 21841 60290
rect 21841 60268 21843 60290
rect 21787 60238 21789 60244
rect 21789 60238 21841 60244
rect 21841 60238 21843 60244
rect 21787 60226 21843 60238
rect 21787 60188 21789 60226
rect 21789 60188 21841 60226
rect 21841 60188 21843 60226
rect 22875 60686 22877 60724
rect 22877 60686 22929 60724
rect 22929 60686 22931 60724
rect 22875 60674 22931 60686
rect 22875 60668 22877 60674
rect 22877 60668 22929 60674
rect 22929 60668 22931 60674
rect 22875 60622 22877 60644
rect 22877 60622 22929 60644
rect 22929 60622 22931 60644
rect 22875 60610 22931 60622
rect 22875 60588 22877 60610
rect 22877 60588 22929 60610
rect 22929 60588 22931 60610
rect 22875 60558 22877 60564
rect 22877 60558 22929 60564
rect 22929 60558 22931 60564
rect 22875 60546 22931 60558
rect 22875 60508 22877 60546
rect 22877 60508 22929 60546
rect 22929 60508 22931 60546
rect 22875 60482 22931 60484
rect 22875 60430 22877 60482
rect 22877 60430 22929 60482
rect 22929 60430 22931 60482
rect 22875 60428 22931 60430
rect 22875 60366 22877 60404
rect 22877 60366 22929 60404
rect 22929 60366 22931 60404
rect 22875 60354 22931 60366
rect 22875 60348 22877 60354
rect 22877 60348 22929 60354
rect 22929 60348 22931 60354
rect 22875 60302 22877 60324
rect 22877 60302 22929 60324
rect 22929 60302 22931 60324
rect 22875 60290 22931 60302
rect 22875 60268 22877 60290
rect 22877 60268 22929 60290
rect 22929 60268 22931 60290
rect 22875 60238 22877 60244
rect 22877 60238 22929 60244
rect 22929 60238 22931 60244
rect 22875 60226 22931 60238
rect 22875 60188 22877 60226
rect 22877 60188 22929 60226
rect 22929 60188 22931 60226
rect 23963 60686 23965 60724
rect 23965 60686 24017 60724
rect 24017 60686 24019 60724
rect 23963 60674 24019 60686
rect 23963 60668 23965 60674
rect 23965 60668 24017 60674
rect 24017 60668 24019 60674
rect 23963 60622 23965 60644
rect 23965 60622 24017 60644
rect 24017 60622 24019 60644
rect 23963 60610 24019 60622
rect 23963 60588 23965 60610
rect 23965 60588 24017 60610
rect 24017 60588 24019 60610
rect 23963 60558 23965 60564
rect 23965 60558 24017 60564
rect 24017 60558 24019 60564
rect 23963 60546 24019 60558
rect 23963 60508 23965 60546
rect 23965 60508 24017 60546
rect 24017 60508 24019 60546
rect 23963 60482 24019 60484
rect 23963 60430 23965 60482
rect 23965 60430 24017 60482
rect 24017 60430 24019 60482
rect 23963 60428 24019 60430
rect 23963 60366 23965 60404
rect 23965 60366 24017 60404
rect 24017 60366 24019 60404
rect 23963 60354 24019 60366
rect 23963 60348 23965 60354
rect 23965 60348 24017 60354
rect 24017 60348 24019 60354
rect 23963 60302 23965 60324
rect 23965 60302 24017 60324
rect 24017 60302 24019 60324
rect 23963 60290 24019 60302
rect 23963 60268 23965 60290
rect 23965 60268 24017 60290
rect 24017 60268 24019 60290
rect 23963 60238 23965 60244
rect 23965 60238 24017 60244
rect 24017 60238 24019 60244
rect 23963 60226 24019 60238
rect 23963 60188 23965 60226
rect 23965 60188 24017 60226
rect 24017 60188 24019 60226
rect 25051 60686 25053 60724
rect 25053 60686 25105 60724
rect 25105 60686 25107 60724
rect 25051 60674 25107 60686
rect 25051 60668 25053 60674
rect 25053 60668 25105 60674
rect 25105 60668 25107 60674
rect 25051 60622 25053 60644
rect 25053 60622 25105 60644
rect 25105 60622 25107 60644
rect 25051 60610 25107 60622
rect 25051 60588 25053 60610
rect 25053 60588 25105 60610
rect 25105 60588 25107 60610
rect 25051 60558 25053 60564
rect 25053 60558 25105 60564
rect 25105 60558 25107 60564
rect 25051 60546 25107 60558
rect 25051 60508 25053 60546
rect 25053 60508 25105 60546
rect 25105 60508 25107 60546
rect 25051 60482 25107 60484
rect 25051 60430 25053 60482
rect 25053 60430 25105 60482
rect 25105 60430 25107 60482
rect 25051 60428 25107 60430
rect 25051 60366 25053 60404
rect 25053 60366 25105 60404
rect 25105 60366 25107 60404
rect 25051 60354 25107 60366
rect 25051 60348 25053 60354
rect 25053 60348 25105 60354
rect 25105 60348 25107 60354
rect 25051 60302 25053 60324
rect 25053 60302 25105 60324
rect 25105 60302 25107 60324
rect 25051 60290 25107 60302
rect 25051 60268 25053 60290
rect 25053 60268 25105 60290
rect 25105 60268 25107 60290
rect 25051 60238 25053 60244
rect 25053 60238 25105 60244
rect 25105 60238 25107 60244
rect 25051 60226 25107 60238
rect 25051 60188 25053 60226
rect 25053 60188 25105 60226
rect 25105 60188 25107 60226
rect 26139 60686 26141 60724
rect 26141 60686 26193 60724
rect 26193 60686 26195 60724
rect 26139 60674 26195 60686
rect 26139 60668 26141 60674
rect 26141 60668 26193 60674
rect 26193 60668 26195 60674
rect 26139 60622 26141 60644
rect 26141 60622 26193 60644
rect 26193 60622 26195 60644
rect 26139 60610 26195 60622
rect 26139 60588 26141 60610
rect 26141 60588 26193 60610
rect 26193 60588 26195 60610
rect 26139 60558 26141 60564
rect 26141 60558 26193 60564
rect 26193 60558 26195 60564
rect 26139 60546 26195 60558
rect 26139 60508 26141 60546
rect 26141 60508 26193 60546
rect 26193 60508 26195 60546
rect 26139 60482 26195 60484
rect 26139 60430 26141 60482
rect 26141 60430 26193 60482
rect 26193 60430 26195 60482
rect 26139 60428 26195 60430
rect 26139 60366 26141 60404
rect 26141 60366 26193 60404
rect 26193 60366 26195 60404
rect 26139 60354 26195 60366
rect 26139 60348 26141 60354
rect 26141 60348 26193 60354
rect 26193 60348 26195 60354
rect 26139 60302 26141 60324
rect 26141 60302 26193 60324
rect 26193 60302 26195 60324
rect 26139 60290 26195 60302
rect 26139 60268 26141 60290
rect 26141 60268 26193 60290
rect 26193 60268 26195 60290
rect 26139 60238 26141 60244
rect 26141 60238 26193 60244
rect 26193 60238 26195 60244
rect 26139 60226 26195 60238
rect 26139 60188 26141 60226
rect 26141 60188 26193 60226
rect 26193 60188 26195 60226
rect 27227 60686 27229 60724
rect 27229 60686 27281 60724
rect 27281 60686 27283 60724
rect 27227 60674 27283 60686
rect 27227 60668 27229 60674
rect 27229 60668 27281 60674
rect 27281 60668 27283 60674
rect 27227 60622 27229 60644
rect 27229 60622 27281 60644
rect 27281 60622 27283 60644
rect 27227 60610 27283 60622
rect 27227 60588 27229 60610
rect 27229 60588 27281 60610
rect 27281 60588 27283 60610
rect 27227 60558 27229 60564
rect 27229 60558 27281 60564
rect 27281 60558 27283 60564
rect 27227 60546 27283 60558
rect 27227 60508 27229 60546
rect 27229 60508 27281 60546
rect 27281 60508 27283 60546
rect 27227 60482 27283 60484
rect 27227 60430 27229 60482
rect 27229 60430 27281 60482
rect 27281 60430 27283 60482
rect 27227 60428 27283 60430
rect 27227 60366 27229 60404
rect 27229 60366 27281 60404
rect 27281 60366 27283 60404
rect 27227 60354 27283 60366
rect 27227 60348 27229 60354
rect 27229 60348 27281 60354
rect 27281 60348 27283 60354
rect 27227 60302 27229 60324
rect 27229 60302 27281 60324
rect 27281 60302 27283 60324
rect 27227 60290 27283 60302
rect 27227 60268 27229 60290
rect 27229 60268 27281 60290
rect 27281 60268 27283 60290
rect 27227 60238 27229 60244
rect 27229 60238 27281 60244
rect 27281 60238 27283 60244
rect 27227 60226 27283 60238
rect 27227 60188 27229 60226
rect 27229 60188 27281 60226
rect 27281 60188 27283 60226
rect 28315 60686 28317 60724
rect 28317 60686 28369 60724
rect 28369 60686 28371 60724
rect 28315 60674 28371 60686
rect 28315 60668 28317 60674
rect 28317 60668 28369 60674
rect 28369 60668 28371 60674
rect 28315 60622 28317 60644
rect 28317 60622 28369 60644
rect 28369 60622 28371 60644
rect 28315 60610 28371 60622
rect 28315 60588 28317 60610
rect 28317 60588 28369 60610
rect 28369 60588 28371 60610
rect 28315 60558 28317 60564
rect 28317 60558 28369 60564
rect 28369 60558 28371 60564
rect 28315 60546 28371 60558
rect 28315 60508 28317 60546
rect 28317 60508 28369 60546
rect 28369 60508 28371 60546
rect 28315 60482 28371 60484
rect 28315 60430 28317 60482
rect 28317 60430 28369 60482
rect 28369 60430 28371 60482
rect 28315 60428 28371 60430
rect 28315 60366 28317 60404
rect 28317 60366 28369 60404
rect 28369 60366 28371 60404
rect 28315 60354 28371 60366
rect 28315 60348 28317 60354
rect 28317 60348 28369 60354
rect 28369 60348 28371 60354
rect 28315 60302 28317 60324
rect 28317 60302 28369 60324
rect 28369 60302 28371 60324
rect 28315 60290 28371 60302
rect 28315 60268 28317 60290
rect 28317 60268 28369 60290
rect 28369 60268 28371 60290
rect 28315 60238 28317 60244
rect 28317 60238 28369 60244
rect 28369 60238 28371 60244
rect 28315 60226 28371 60238
rect 28315 60188 28317 60226
rect 28317 60188 28369 60226
rect 28369 60188 28371 60226
rect 29403 60686 29405 60724
rect 29405 60686 29457 60724
rect 29457 60686 29459 60724
rect 29403 60674 29459 60686
rect 29403 60668 29405 60674
rect 29405 60668 29457 60674
rect 29457 60668 29459 60674
rect 29403 60622 29405 60644
rect 29405 60622 29457 60644
rect 29457 60622 29459 60644
rect 29403 60610 29459 60622
rect 29403 60588 29405 60610
rect 29405 60588 29457 60610
rect 29457 60588 29459 60610
rect 29403 60558 29405 60564
rect 29405 60558 29457 60564
rect 29457 60558 29459 60564
rect 29403 60546 29459 60558
rect 29403 60508 29405 60546
rect 29405 60508 29457 60546
rect 29457 60508 29459 60546
rect 29403 60482 29459 60484
rect 29403 60430 29405 60482
rect 29405 60430 29457 60482
rect 29457 60430 29459 60482
rect 29403 60428 29459 60430
rect 29403 60366 29405 60404
rect 29405 60366 29457 60404
rect 29457 60366 29459 60404
rect 29403 60354 29459 60366
rect 29403 60348 29405 60354
rect 29405 60348 29457 60354
rect 29457 60348 29459 60354
rect 29403 60302 29405 60324
rect 29405 60302 29457 60324
rect 29457 60302 29459 60324
rect 29403 60290 29459 60302
rect 29403 60268 29405 60290
rect 29405 60268 29457 60290
rect 29457 60268 29459 60290
rect 29403 60238 29405 60244
rect 29405 60238 29457 60244
rect 29457 60238 29459 60244
rect 29403 60226 29459 60238
rect 29403 60188 29405 60226
rect 29405 60188 29457 60226
rect 29457 60188 29459 60226
rect 30491 60686 30493 60724
rect 30493 60686 30545 60724
rect 30545 60686 30547 60724
rect 30491 60674 30547 60686
rect 30491 60668 30493 60674
rect 30493 60668 30545 60674
rect 30545 60668 30547 60674
rect 30491 60622 30493 60644
rect 30493 60622 30545 60644
rect 30545 60622 30547 60644
rect 30491 60610 30547 60622
rect 30491 60588 30493 60610
rect 30493 60588 30545 60610
rect 30545 60588 30547 60610
rect 30491 60558 30493 60564
rect 30493 60558 30545 60564
rect 30545 60558 30547 60564
rect 30491 60546 30547 60558
rect 30491 60508 30493 60546
rect 30493 60508 30545 60546
rect 30545 60508 30547 60546
rect 30491 60482 30547 60484
rect 30491 60430 30493 60482
rect 30493 60430 30545 60482
rect 30545 60430 30547 60482
rect 30491 60428 30547 60430
rect 30491 60366 30493 60404
rect 30493 60366 30545 60404
rect 30545 60366 30547 60404
rect 30491 60354 30547 60366
rect 30491 60348 30493 60354
rect 30493 60348 30545 60354
rect 30545 60348 30547 60354
rect 30491 60302 30493 60324
rect 30493 60302 30545 60324
rect 30545 60302 30547 60324
rect 30491 60290 30547 60302
rect 30491 60268 30493 60290
rect 30493 60268 30545 60290
rect 30545 60268 30547 60290
rect 30491 60238 30493 60244
rect 30493 60238 30545 60244
rect 30545 60238 30547 60244
rect 30491 60226 30547 60238
rect 30491 60188 30493 60226
rect 30493 60188 30545 60226
rect 30545 60188 30547 60226
rect 31579 60686 31581 60724
rect 31581 60686 31633 60724
rect 31633 60686 31635 60724
rect 31579 60674 31635 60686
rect 31579 60668 31581 60674
rect 31581 60668 31633 60674
rect 31633 60668 31635 60674
rect 31579 60622 31581 60644
rect 31581 60622 31633 60644
rect 31633 60622 31635 60644
rect 31579 60610 31635 60622
rect 31579 60588 31581 60610
rect 31581 60588 31633 60610
rect 31633 60588 31635 60610
rect 31579 60558 31581 60564
rect 31581 60558 31633 60564
rect 31633 60558 31635 60564
rect 31579 60546 31635 60558
rect 31579 60508 31581 60546
rect 31581 60508 31633 60546
rect 31633 60508 31635 60546
rect 31579 60482 31635 60484
rect 31579 60430 31581 60482
rect 31581 60430 31633 60482
rect 31633 60430 31635 60482
rect 31579 60428 31635 60430
rect 31579 60366 31581 60404
rect 31581 60366 31633 60404
rect 31633 60366 31635 60404
rect 31579 60354 31635 60366
rect 31579 60348 31581 60354
rect 31581 60348 31633 60354
rect 31633 60348 31635 60354
rect 31579 60302 31581 60324
rect 31581 60302 31633 60324
rect 31633 60302 31635 60324
rect 31579 60290 31635 60302
rect 31579 60268 31581 60290
rect 31581 60268 31633 60290
rect 31633 60268 31635 60290
rect 31579 60238 31581 60244
rect 31581 60238 31633 60244
rect 31633 60238 31635 60244
rect 31579 60226 31635 60238
rect 31579 60188 31581 60226
rect 31581 60188 31633 60226
rect 31633 60188 31635 60226
rect 17980 58683 17982 58721
rect 17982 58683 18034 58721
rect 18034 58683 18036 58721
rect 17980 58671 18036 58683
rect 17980 58665 17982 58671
rect 17982 58665 18034 58671
rect 18034 58665 18036 58671
rect 17980 58619 17982 58641
rect 17982 58619 18034 58641
rect 18034 58619 18036 58641
rect 17980 58607 18036 58619
rect 17980 58585 17982 58607
rect 17982 58585 18034 58607
rect 18034 58585 18036 58607
rect 17980 58555 17982 58561
rect 17982 58555 18034 58561
rect 18034 58555 18036 58561
rect 17980 58543 18036 58555
rect 17980 58505 17982 58543
rect 17982 58505 18034 58543
rect 18034 58505 18036 58543
rect 17980 58479 18036 58481
rect 17980 58427 17982 58479
rect 17982 58427 18034 58479
rect 18034 58427 18036 58479
rect 17980 58425 18036 58427
rect 17980 58363 17982 58401
rect 17982 58363 18034 58401
rect 18034 58363 18036 58401
rect 17980 58351 18036 58363
rect 17980 58345 17982 58351
rect 17982 58345 18034 58351
rect 18034 58345 18036 58351
rect 17980 58299 17982 58321
rect 17982 58299 18034 58321
rect 18034 58299 18036 58321
rect 17980 58287 18036 58299
rect 17980 58265 17982 58287
rect 17982 58265 18034 58287
rect 18034 58265 18036 58287
rect 17980 58235 17982 58241
rect 17982 58235 18034 58241
rect 18034 58235 18036 58241
rect 17980 58223 18036 58235
rect 17980 58185 17982 58223
rect 17982 58185 18034 58223
rect 18034 58185 18036 58223
rect 19068 58683 19070 58721
rect 19070 58683 19122 58721
rect 19122 58683 19124 58721
rect 19068 58671 19124 58683
rect 19068 58665 19070 58671
rect 19070 58665 19122 58671
rect 19122 58665 19124 58671
rect 19068 58619 19070 58641
rect 19070 58619 19122 58641
rect 19122 58619 19124 58641
rect 19068 58607 19124 58619
rect 19068 58585 19070 58607
rect 19070 58585 19122 58607
rect 19122 58585 19124 58607
rect 19068 58555 19070 58561
rect 19070 58555 19122 58561
rect 19122 58555 19124 58561
rect 19068 58543 19124 58555
rect 19068 58505 19070 58543
rect 19070 58505 19122 58543
rect 19122 58505 19124 58543
rect 19068 58479 19124 58481
rect 19068 58427 19070 58479
rect 19070 58427 19122 58479
rect 19122 58427 19124 58479
rect 19068 58425 19124 58427
rect 19068 58363 19070 58401
rect 19070 58363 19122 58401
rect 19122 58363 19124 58401
rect 19068 58351 19124 58363
rect 19068 58345 19070 58351
rect 19070 58345 19122 58351
rect 19122 58345 19124 58351
rect 19068 58299 19070 58321
rect 19070 58299 19122 58321
rect 19122 58299 19124 58321
rect 19068 58287 19124 58299
rect 19068 58265 19070 58287
rect 19070 58265 19122 58287
rect 19122 58265 19124 58287
rect 19068 58235 19070 58241
rect 19070 58235 19122 58241
rect 19122 58235 19124 58241
rect 19068 58223 19124 58235
rect 19068 58185 19070 58223
rect 19070 58185 19122 58223
rect 19122 58185 19124 58223
rect 20156 58683 20158 58721
rect 20158 58683 20210 58721
rect 20210 58683 20212 58721
rect 20156 58671 20212 58683
rect 20156 58665 20158 58671
rect 20158 58665 20210 58671
rect 20210 58665 20212 58671
rect 20156 58619 20158 58641
rect 20158 58619 20210 58641
rect 20210 58619 20212 58641
rect 20156 58607 20212 58619
rect 20156 58585 20158 58607
rect 20158 58585 20210 58607
rect 20210 58585 20212 58607
rect 20156 58555 20158 58561
rect 20158 58555 20210 58561
rect 20210 58555 20212 58561
rect 20156 58543 20212 58555
rect 20156 58505 20158 58543
rect 20158 58505 20210 58543
rect 20210 58505 20212 58543
rect 20156 58479 20212 58481
rect 20156 58427 20158 58479
rect 20158 58427 20210 58479
rect 20210 58427 20212 58479
rect 20156 58425 20212 58427
rect 20156 58363 20158 58401
rect 20158 58363 20210 58401
rect 20210 58363 20212 58401
rect 20156 58351 20212 58363
rect 20156 58345 20158 58351
rect 20158 58345 20210 58351
rect 20210 58345 20212 58351
rect 20156 58299 20158 58321
rect 20158 58299 20210 58321
rect 20210 58299 20212 58321
rect 20156 58287 20212 58299
rect 20156 58265 20158 58287
rect 20158 58265 20210 58287
rect 20210 58265 20212 58287
rect 20156 58235 20158 58241
rect 20158 58235 20210 58241
rect 20210 58235 20212 58241
rect 20156 58223 20212 58235
rect 20156 58185 20158 58223
rect 20158 58185 20210 58223
rect 20210 58185 20212 58223
rect 21244 58683 21246 58721
rect 21246 58683 21298 58721
rect 21298 58683 21300 58721
rect 21244 58671 21300 58683
rect 21244 58665 21246 58671
rect 21246 58665 21298 58671
rect 21298 58665 21300 58671
rect 21244 58619 21246 58641
rect 21246 58619 21298 58641
rect 21298 58619 21300 58641
rect 21244 58607 21300 58619
rect 21244 58585 21246 58607
rect 21246 58585 21298 58607
rect 21298 58585 21300 58607
rect 21244 58555 21246 58561
rect 21246 58555 21298 58561
rect 21298 58555 21300 58561
rect 21244 58543 21300 58555
rect 21244 58505 21246 58543
rect 21246 58505 21298 58543
rect 21298 58505 21300 58543
rect 21244 58479 21300 58481
rect 21244 58427 21246 58479
rect 21246 58427 21298 58479
rect 21298 58427 21300 58479
rect 21244 58425 21300 58427
rect 21244 58363 21246 58401
rect 21246 58363 21298 58401
rect 21298 58363 21300 58401
rect 21244 58351 21300 58363
rect 21244 58345 21246 58351
rect 21246 58345 21298 58351
rect 21298 58345 21300 58351
rect 21244 58299 21246 58321
rect 21246 58299 21298 58321
rect 21298 58299 21300 58321
rect 21244 58287 21300 58299
rect 21244 58265 21246 58287
rect 21246 58265 21298 58287
rect 21298 58265 21300 58287
rect 21244 58235 21246 58241
rect 21246 58235 21298 58241
rect 21298 58235 21300 58241
rect 21244 58223 21300 58235
rect 21244 58185 21246 58223
rect 21246 58185 21298 58223
rect 21298 58185 21300 58223
rect 22332 58683 22334 58721
rect 22334 58683 22386 58721
rect 22386 58683 22388 58721
rect 22332 58671 22388 58683
rect 22332 58665 22334 58671
rect 22334 58665 22386 58671
rect 22386 58665 22388 58671
rect 22332 58619 22334 58641
rect 22334 58619 22386 58641
rect 22386 58619 22388 58641
rect 22332 58607 22388 58619
rect 22332 58585 22334 58607
rect 22334 58585 22386 58607
rect 22386 58585 22388 58607
rect 22332 58555 22334 58561
rect 22334 58555 22386 58561
rect 22386 58555 22388 58561
rect 22332 58543 22388 58555
rect 22332 58505 22334 58543
rect 22334 58505 22386 58543
rect 22386 58505 22388 58543
rect 22332 58479 22388 58481
rect 22332 58427 22334 58479
rect 22334 58427 22386 58479
rect 22386 58427 22388 58479
rect 22332 58425 22388 58427
rect 22332 58363 22334 58401
rect 22334 58363 22386 58401
rect 22386 58363 22388 58401
rect 22332 58351 22388 58363
rect 22332 58345 22334 58351
rect 22334 58345 22386 58351
rect 22386 58345 22388 58351
rect 22332 58299 22334 58321
rect 22334 58299 22386 58321
rect 22386 58299 22388 58321
rect 22332 58287 22388 58299
rect 22332 58265 22334 58287
rect 22334 58265 22386 58287
rect 22386 58265 22388 58287
rect 22332 58235 22334 58241
rect 22334 58235 22386 58241
rect 22386 58235 22388 58241
rect 22332 58223 22388 58235
rect 22332 58185 22334 58223
rect 22334 58185 22386 58223
rect 22386 58185 22388 58223
rect 23420 58683 23422 58721
rect 23422 58683 23474 58721
rect 23474 58683 23476 58721
rect 23420 58671 23476 58683
rect 23420 58665 23422 58671
rect 23422 58665 23474 58671
rect 23474 58665 23476 58671
rect 23420 58619 23422 58641
rect 23422 58619 23474 58641
rect 23474 58619 23476 58641
rect 23420 58607 23476 58619
rect 23420 58585 23422 58607
rect 23422 58585 23474 58607
rect 23474 58585 23476 58607
rect 23420 58555 23422 58561
rect 23422 58555 23474 58561
rect 23474 58555 23476 58561
rect 23420 58543 23476 58555
rect 23420 58505 23422 58543
rect 23422 58505 23474 58543
rect 23474 58505 23476 58543
rect 23420 58479 23476 58481
rect 23420 58427 23422 58479
rect 23422 58427 23474 58479
rect 23474 58427 23476 58479
rect 23420 58425 23476 58427
rect 23420 58363 23422 58401
rect 23422 58363 23474 58401
rect 23474 58363 23476 58401
rect 23420 58351 23476 58363
rect 23420 58345 23422 58351
rect 23422 58345 23474 58351
rect 23474 58345 23476 58351
rect 23420 58299 23422 58321
rect 23422 58299 23474 58321
rect 23474 58299 23476 58321
rect 23420 58287 23476 58299
rect 23420 58265 23422 58287
rect 23422 58265 23474 58287
rect 23474 58265 23476 58287
rect 23420 58235 23422 58241
rect 23422 58235 23474 58241
rect 23474 58235 23476 58241
rect 23420 58223 23476 58235
rect 23420 58185 23422 58223
rect 23422 58185 23474 58223
rect 23474 58185 23476 58223
rect 24508 58683 24510 58721
rect 24510 58683 24562 58721
rect 24562 58683 24564 58721
rect 24508 58671 24564 58683
rect 24508 58665 24510 58671
rect 24510 58665 24562 58671
rect 24562 58665 24564 58671
rect 24508 58619 24510 58641
rect 24510 58619 24562 58641
rect 24562 58619 24564 58641
rect 24508 58607 24564 58619
rect 24508 58585 24510 58607
rect 24510 58585 24562 58607
rect 24562 58585 24564 58607
rect 24508 58555 24510 58561
rect 24510 58555 24562 58561
rect 24562 58555 24564 58561
rect 24508 58543 24564 58555
rect 24508 58505 24510 58543
rect 24510 58505 24562 58543
rect 24562 58505 24564 58543
rect 24508 58479 24564 58481
rect 24508 58427 24510 58479
rect 24510 58427 24562 58479
rect 24562 58427 24564 58479
rect 24508 58425 24564 58427
rect 24508 58363 24510 58401
rect 24510 58363 24562 58401
rect 24562 58363 24564 58401
rect 24508 58351 24564 58363
rect 24508 58345 24510 58351
rect 24510 58345 24562 58351
rect 24562 58345 24564 58351
rect 24508 58299 24510 58321
rect 24510 58299 24562 58321
rect 24562 58299 24564 58321
rect 24508 58287 24564 58299
rect 24508 58265 24510 58287
rect 24510 58265 24562 58287
rect 24562 58265 24564 58287
rect 24508 58235 24510 58241
rect 24510 58235 24562 58241
rect 24562 58235 24564 58241
rect 24508 58223 24564 58235
rect 24508 58185 24510 58223
rect 24510 58185 24562 58223
rect 24562 58185 24564 58223
rect 25596 58683 25598 58721
rect 25598 58683 25650 58721
rect 25650 58683 25652 58721
rect 25596 58671 25652 58683
rect 25596 58665 25598 58671
rect 25598 58665 25650 58671
rect 25650 58665 25652 58671
rect 25596 58619 25598 58641
rect 25598 58619 25650 58641
rect 25650 58619 25652 58641
rect 25596 58607 25652 58619
rect 25596 58585 25598 58607
rect 25598 58585 25650 58607
rect 25650 58585 25652 58607
rect 25596 58555 25598 58561
rect 25598 58555 25650 58561
rect 25650 58555 25652 58561
rect 25596 58543 25652 58555
rect 25596 58505 25598 58543
rect 25598 58505 25650 58543
rect 25650 58505 25652 58543
rect 25596 58479 25652 58481
rect 25596 58427 25598 58479
rect 25598 58427 25650 58479
rect 25650 58427 25652 58479
rect 25596 58425 25652 58427
rect 25596 58363 25598 58401
rect 25598 58363 25650 58401
rect 25650 58363 25652 58401
rect 25596 58351 25652 58363
rect 25596 58345 25598 58351
rect 25598 58345 25650 58351
rect 25650 58345 25652 58351
rect 25596 58299 25598 58321
rect 25598 58299 25650 58321
rect 25650 58299 25652 58321
rect 25596 58287 25652 58299
rect 25596 58265 25598 58287
rect 25598 58265 25650 58287
rect 25650 58265 25652 58287
rect 25596 58235 25598 58241
rect 25598 58235 25650 58241
rect 25650 58235 25652 58241
rect 25596 58223 25652 58235
rect 25596 58185 25598 58223
rect 25598 58185 25650 58223
rect 25650 58185 25652 58223
rect 26684 58683 26686 58721
rect 26686 58683 26738 58721
rect 26738 58683 26740 58721
rect 26684 58671 26740 58683
rect 26684 58665 26686 58671
rect 26686 58665 26738 58671
rect 26738 58665 26740 58671
rect 26684 58619 26686 58641
rect 26686 58619 26738 58641
rect 26738 58619 26740 58641
rect 26684 58607 26740 58619
rect 26684 58585 26686 58607
rect 26686 58585 26738 58607
rect 26738 58585 26740 58607
rect 26684 58555 26686 58561
rect 26686 58555 26738 58561
rect 26738 58555 26740 58561
rect 26684 58543 26740 58555
rect 26684 58505 26686 58543
rect 26686 58505 26738 58543
rect 26738 58505 26740 58543
rect 26684 58479 26740 58481
rect 26684 58427 26686 58479
rect 26686 58427 26738 58479
rect 26738 58427 26740 58479
rect 26684 58425 26740 58427
rect 26684 58363 26686 58401
rect 26686 58363 26738 58401
rect 26738 58363 26740 58401
rect 26684 58351 26740 58363
rect 26684 58345 26686 58351
rect 26686 58345 26738 58351
rect 26738 58345 26740 58351
rect 26684 58299 26686 58321
rect 26686 58299 26738 58321
rect 26738 58299 26740 58321
rect 26684 58287 26740 58299
rect 26684 58265 26686 58287
rect 26686 58265 26738 58287
rect 26738 58265 26740 58287
rect 26684 58235 26686 58241
rect 26686 58235 26738 58241
rect 26738 58235 26740 58241
rect 26684 58223 26740 58235
rect 26684 58185 26686 58223
rect 26686 58185 26738 58223
rect 26738 58185 26740 58223
rect 27772 58683 27774 58721
rect 27774 58683 27826 58721
rect 27826 58683 27828 58721
rect 27772 58671 27828 58683
rect 27772 58665 27774 58671
rect 27774 58665 27826 58671
rect 27826 58665 27828 58671
rect 27772 58619 27774 58641
rect 27774 58619 27826 58641
rect 27826 58619 27828 58641
rect 27772 58607 27828 58619
rect 27772 58585 27774 58607
rect 27774 58585 27826 58607
rect 27826 58585 27828 58607
rect 27772 58555 27774 58561
rect 27774 58555 27826 58561
rect 27826 58555 27828 58561
rect 27772 58543 27828 58555
rect 27772 58505 27774 58543
rect 27774 58505 27826 58543
rect 27826 58505 27828 58543
rect 27772 58479 27828 58481
rect 27772 58427 27774 58479
rect 27774 58427 27826 58479
rect 27826 58427 27828 58479
rect 27772 58425 27828 58427
rect 27772 58363 27774 58401
rect 27774 58363 27826 58401
rect 27826 58363 27828 58401
rect 27772 58351 27828 58363
rect 27772 58345 27774 58351
rect 27774 58345 27826 58351
rect 27826 58345 27828 58351
rect 27772 58299 27774 58321
rect 27774 58299 27826 58321
rect 27826 58299 27828 58321
rect 27772 58287 27828 58299
rect 27772 58265 27774 58287
rect 27774 58265 27826 58287
rect 27826 58265 27828 58287
rect 27772 58235 27774 58241
rect 27774 58235 27826 58241
rect 27826 58235 27828 58241
rect 27772 58223 27828 58235
rect 27772 58185 27774 58223
rect 27774 58185 27826 58223
rect 27826 58185 27828 58223
rect 28860 58683 28862 58721
rect 28862 58683 28914 58721
rect 28914 58683 28916 58721
rect 28860 58671 28916 58683
rect 28860 58665 28862 58671
rect 28862 58665 28914 58671
rect 28914 58665 28916 58671
rect 28860 58619 28862 58641
rect 28862 58619 28914 58641
rect 28914 58619 28916 58641
rect 28860 58607 28916 58619
rect 28860 58585 28862 58607
rect 28862 58585 28914 58607
rect 28914 58585 28916 58607
rect 28860 58555 28862 58561
rect 28862 58555 28914 58561
rect 28914 58555 28916 58561
rect 28860 58543 28916 58555
rect 28860 58505 28862 58543
rect 28862 58505 28914 58543
rect 28914 58505 28916 58543
rect 28860 58479 28916 58481
rect 28860 58427 28862 58479
rect 28862 58427 28914 58479
rect 28914 58427 28916 58479
rect 28860 58425 28916 58427
rect 28860 58363 28862 58401
rect 28862 58363 28914 58401
rect 28914 58363 28916 58401
rect 28860 58351 28916 58363
rect 28860 58345 28862 58351
rect 28862 58345 28914 58351
rect 28914 58345 28916 58351
rect 28860 58299 28862 58321
rect 28862 58299 28914 58321
rect 28914 58299 28916 58321
rect 28860 58287 28916 58299
rect 28860 58265 28862 58287
rect 28862 58265 28914 58287
rect 28914 58265 28916 58287
rect 28860 58235 28862 58241
rect 28862 58235 28914 58241
rect 28914 58235 28916 58241
rect 28860 58223 28916 58235
rect 28860 58185 28862 58223
rect 28862 58185 28914 58223
rect 28914 58185 28916 58223
rect 29948 58683 29950 58721
rect 29950 58683 30002 58721
rect 30002 58683 30004 58721
rect 29948 58671 30004 58683
rect 29948 58665 29950 58671
rect 29950 58665 30002 58671
rect 30002 58665 30004 58671
rect 29948 58619 29950 58641
rect 29950 58619 30002 58641
rect 30002 58619 30004 58641
rect 29948 58607 30004 58619
rect 29948 58585 29950 58607
rect 29950 58585 30002 58607
rect 30002 58585 30004 58607
rect 29948 58555 29950 58561
rect 29950 58555 30002 58561
rect 30002 58555 30004 58561
rect 29948 58543 30004 58555
rect 29948 58505 29950 58543
rect 29950 58505 30002 58543
rect 30002 58505 30004 58543
rect 29948 58479 30004 58481
rect 29948 58427 29950 58479
rect 29950 58427 30002 58479
rect 30002 58427 30004 58479
rect 29948 58425 30004 58427
rect 29948 58363 29950 58401
rect 29950 58363 30002 58401
rect 30002 58363 30004 58401
rect 29948 58351 30004 58363
rect 29948 58345 29950 58351
rect 29950 58345 30002 58351
rect 30002 58345 30004 58351
rect 29948 58299 29950 58321
rect 29950 58299 30002 58321
rect 30002 58299 30004 58321
rect 29948 58287 30004 58299
rect 29948 58265 29950 58287
rect 29950 58265 30002 58287
rect 30002 58265 30004 58287
rect 29948 58235 29950 58241
rect 29950 58235 30002 58241
rect 30002 58235 30004 58241
rect 29948 58223 30004 58235
rect 29948 58185 29950 58223
rect 29950 58185 30002 58223
rect 30002 58185 30004 58223
rect 31036 58683 31038 58721
rect 31038 58683 31090 58721
rect 31090 58683 31092 58721
rect 31036 58671 31092 58683
rect 31036 58665 31038 58671
rect 31038 58665 31090 58671
rect 31090 58665 31092 58671
rect 31036 58619 31038 58641
rect 31038 58619 31090 58641
rect 31090 58619 31092 58641
rect 31036 58607 31092 58619
rect 31036 58585 31038 58607
rect 31038 58585 31090 58607
rect 31090 58585 31092 58607
rect 31036 58555 31038 58561
rect 31038 58555 31090 58561
rect 31090 58555 31092 58561
rect 31036 58543 31092 58555
rect 31036 58505 31038 58543
rect 31038 58505 31090 58543
rect 31090 58505 31092 58543
rect 31036 58479 31092 58481
rect 31036 58427 31038 58479
rect 31038 58427 31090 58479
rect 31090 58427 31092 58479
rect 31036 58425 31092 58427
rect 31036 58363 31038 58401
rect 31038 58363 31090 58401
rect 31090 58363 31092 58401
rect 31036 58351 31092 58363
rect 31036 58345 31038 58351
rect 31038 58345 31090 58351
rect 31090 58345 31092 58351
rect 31036 58299 31038 58321
rect 31038 58299 31090 58321
rect 31090 58299 31092 58321
rect 31036 58287 31092 58299
rect 31036 58265 31038 58287
rect 31038 58265 31090 58287
rect 31090 58265 31092 58287
rect 31036 58235 31038 58241
rect 31038 58235 31090 58241
rect 31090 58235 31092 58241
rect 31036 58223 31092 58235
rect 31036 58185 31038 58223
rect 31038 58185 31090 58223
rect 31090 58185 31092 58223
rect 17435 56686 17437 56724
rect 17437 56686 17489 56724
rect 17489 56686 17491 56724
rect 17435 56674 17491 56686
rect 17435 56668 17437 56674
rect 17437 56668 17489 56674
rect 17489 56668 17491 56674
rect 17435 56622 17437 56644
rect 17437 56622 17489 56644
rect 17489 56622 17491 56644
rect 17435 56610 17491 56622
rect 17435 56588 17437 56610
rect 17437 56588 17489 56610
rect 17489 56588 17491 56610
rect 17435 56558 17437 56564
rect 17437 56558 17489 56564
rect 17489 56558 17491 56564
rect 17435 56546 17491 56558
rect 17435 56508 17437 56546
rect 17437 56508 17489 56546
rect 17489 56508 17491 56546
rect 17435 56482 17491 56484
rect 17435 56430 17437 56482
rect 17437 56430 17489 56482
rect 17489 56430 17491 56482
rect 17435 56428 17491 56430
rect 17435 56366 17437 56404
rect 17437 56366 17489 56404
rect 17489 56366 17491 56404
rect 17435 56354 17491 56366
rect 17435 56348 17437 56354
rect 17437 56348 17489 56354
rect 17489 56348 17491 56354
rect 17435 56302 17437 56324
rect 17437 56302 17489 56324
rect 17489 56302 17491 56324
rect 17435 56290 17491 56302
rect 17435 56268 17437 56290
rect 17437 56268 17489 56290
rect 17489 56268 17491 56290
rect 17435 56238 17437 56244
rect 17437 56238 17489 56244
rect 17489 56238 17491 56244
rect 17435 56226 17491 56238
rect 17435 56188 17437 56226
rect 17437 56188 17489 56226
rect 17489 56188 17491 56226
rect 18523 56686 18525 56724
rect 18525 56686 18577 56724
rect 18577 56686 18579 56724
rect 18523 56674 18579 56686
rect 18523 56668 18525 56674
rect 18525 56668 18577 56674
rect 18577 56668 18579 56674
rect 18523 56622 18525 56644
rect 18525 56622 18577 56644
rect 18577 56622 18579 56644
rect 18523 56610 18579 56622
rect 18523 56588 18525 56610
rect 18525 56588 18577 56610
rect 18577 56588 18579 56610
rect 18523 56558 18525 56564
rect 18525 56558 18577 56564
rect 18577 56558 18579 56564
rect 18523 56546 18579 56558
rect 18523 56508 18525 56546
rect 18525 56508 18577 56546
rect 18577 56508 18579 56546
rect 18523 56482 18579 56484
rect 18523 56430 18525 56482
rect 18525 56430 18577 56482
rect 18577 56430 18579 56482
rect 18523 56428 18579 56430
rect 18523 56366 18525 56404
rect 18525 56366 18577 56404
rect 18577 56366 18579 56404
rect 18523 56354 18579 56366
rect 18523 56348 18525 56354
rect 18525 56348 18577 56354
rect 18577 56348 18579 56354
rect 18523 56302 18525 56324
rect 18525 56302 18577 56324
rect 18577 56302 18579 56324
rect 18523 56290 18579 56302
rect 18523 56268 18525 56290
rect 18525 56268 18577 56290
rect 18577 56268 18579 56290
rect 18523 56238 18525 56244
rect 18525 56238 18577 56244
rect 18577 56238 18579 56244
rect 18523 56226 18579 56238
rect 18523 56188 18525 56226
rect 18525 56188 18577 56226
rect 18577 56188 18579 56226
rect 19611 56686 19613 56724
rect 19613 56686 19665 56724
rect 19665 56686 19667 56724
rect 19611 56674 19667 56686
rect 19611 56668 19613 56674
rect 19613 56668 19665 56674
rect 19665 56668 19667 56674
rect 19611 56622 19613 56644
rect 19613 56622 19665 56644
rect 19665 56622 19667 56644
rect 19611 56610 19667 56622
rect 19611 56588 19613 56610
rect 19613 56588 19665 56610
rect 19665 56588 19667 56610
rect 19611 56558 19613 56564
rect 19613 56558 19665 56564
rect 19665 56558 19667 56564
rect 19611 56546 19667 56558
rect 19611 56508 19613 56546
rect 19613 56508 19665 56546
rect 19665 56508 19667 56546
rect 19611 56482 19667 56484
rect 19611 56430 19613 56482
rect 19613 56430 19665 56482
rect 19665 56430 19667 56482
rect 19611 56428 19667 56430
rect 19611 56366 19613 56404
rect 19613 56366 19665 56404
rect 19665 56366 19667 56404
rect 19611 56354 19667 56366
rect 19611 56348 19613 56354
rect 19613 56348 19665 56354
rect 19665 56348 19667 56354
rect 19611 56302 19613 56324
rect 19613 56302 19665 56324
rect 19665 56302 19667 56324
rect 19611 56290 19667 56302
rect 19611 56268 19613 56290
rect 19613 56268 19665 56290
rect 19665 56268 19667 56290
rect 19611 56238 19613 56244
rect 19613 56238 19665 56244
rect 19665 56238 19667 56244
rect 19611 56226 19667 56238
rect 19611 56188 19613 56226
rect 19613 56188 19665 56226
rect 19665 56188 19667 56226
rect 20699 56686 20701 56724
rect 20701 56686 20753 56724
rect 20753 56686 20755 56724
rect 20699 56674 20755 56686
rect 20699 56668 20701 56674
rect 20701 56668 20753 56674
rect 20753 56668 20755 56674
rect 20699 56622 20701 56644
rect 20701 56622 20753 56644
rect 20753 56622 20755 56644
rect 20699 56610 20755 56622
rect 20699 56588 20701 56610
rect 20701 56588 20753 56610
rect 20753 56588 20755 56610
rect 20699 56558 20701 56564
rect 20701 56558 20753 56564
rect 20753 56558 20755 56564
rect 20699 56546 20755 56558
rect 20699 56508 20701 56546
rect 20701 56508 20753 56546
rect 20753 56508 20755 56546
rect 20699 56482 20755 56484
rect 20699 56430 20701 56482
rect 20701 56430 20753 56482
rect 20753 56430 20755 56482
rect 20699 56428 20755 56430
rect 20699 56366 20701 56404
rect 20701 56366 20753 56404
rect 20753 56366 20755 56404
rect 20699 56354 20755 56366
rect 20699 56348 20701 56354
rect 20701 56348 20753 56354
rect 20753 56348 20755 56354
rect 20699 56302 20701 56324
rect 20701 56302 20753 56324
rect 20753 56302 20755 56324
rect 20699 56290 20755 56302
rect 20699 56268 20701 56290
rect 20701 56268 20753 56290
rect 20753 56268 20755 56290
rect 20699 56238 20701 56244
rect 20701 56238 20753 56244
rect 20753 56238 20755 56244
rect 20699 56226 20755 56238
rect 20699 56188 20701 56226
rect 20701 56188 20753 56226
rect 20753 56188 20755 56226
rect 21787 56686 21789 56724
rect 21789 56686 21841 56724
rect 21841 56686 21843 56724
rect 21787 56674 21843 56686
rect 21787 56668 21789 56674
rect 21789 56668 21841 56674
rect 21841 56668 21843 56674
rect 21787 56622 21789 56644
rect 21789 56622 21841 56644
rect 21841 56622 21843 56644
rect 21787 56610 21843 56622
rect 21787 56588 21789 56610
rect 21789 56588 21841 56610
rect 21841 56588 21843 56610
rect 21787 56558 21789 56564
rect 21789 56558 21841 56564
rect 21841 56558 21843 56564
rect 21787 56546 21843 56558
rect 21787 56508 21789 56546
rect 21789 56508 21841 56546
rect 21841 56508 21843 56546
rect 21787 56482 21843 56484
rect 21787 56430 21789 56482
rect 21789 56430 21841 56482
rect 21841 56430 21843 56482
rect 21787 56428 21843 56430
rect 21787 56366 21789 56404
rect 21789 56366 21841 56404
rect 21841 56366 21843 56404
rect 21787 56354 21843 56366
rect 21787 56348 21789 56354
rect 21789 56348 21841 56354
rect 21841 56348 21843 56354
rect 21787 56302 21789 56324
rect 21789 56302 21841 56324
rect 21841 56302 21843 56324
rect 21787 56290 21843 56302
rect 21787 56268 21789 56290
rect 21789 56268 21841 56290
rect 21841 56268 21843 56290
rect 21787 56238 21789 56244
rect 21789 56238 21841 56244
rect 21841 56238 21843 56244
rect 21787 56226 21843 56238
rect 21787 56188 21789 56226
rect 21789 56188 21841 56226
rect 21841 56188 21843 56226
rect 22875 56686 22877 56724
rect 22877 56686 22929 56724
rect 22929 56686 22931 56724
rect 22875 56674 22931 56686
rect 22875 56668 22877 56674
rect 22877 56668 22929 56674
rect 22929 56668 22931 56674
rect 22875 56622 22877 56644
rect 22877 56622 22929 56644
rect 22929 56622 22931 56644
rect 22875 56610 22931 56622
rect 22875 56588 22877 56610
rect 22877 56588 22929 56610
rect 22929 56588 22931 56610
rect 22875 56558 22877 56564
rect 22877 56558 22929 56564
rect 22929 56558 22931 56564
rect 22875 56546 22931 56558
rect 22875 56508 22877 56546
rect 22877 56508 22929 56546
rect 22929 56508 22931 56546
rect 22875 56482 22931 56484
rect 22875 56430 22877 56482
rect 22877 56430 22929 56482
rect 22929 56430 22931 56482
rect 22875 56428 22931 56430
rect 22875 56366 22877 56404
rect 22877 56366 22929 56404
rect 22929 56366 22931 56404
rect 22875 56354 22931 56366
rect 22875 56348 22877 56354
rect 22877 56348 22929 56354
rect 22929 56348 22931 56354
rect 22875 56302 22877 56324
rect 22877 56302 22929 56324
rect 22929 56302 22931 56324
rect 22875 56290 22931 56302
rect 22875 56268 22877 56290
rect 22877 56268 22929 56290
rect 22929 56268 22931 56290
rect 22875 56238 22877 56244
rect 22877 56238 22929 56244
rect 22929 56238 22931 56244
rect 22875 56226 22931 56238
rect 22875 56188 22877 56226
rect 22877 56188 22929 56226
rect 22929 56188 22931 56226
rect 23963 56686 23965 56724
rect 23965 56686 24017 56724
rect 24017 56686 24019 56724
rect 23963 56674 24019 56686
rect 23963 56668 23965 56674
rect 23965 56668 24017 56674
rect 24017 56668 24019 56674
rect 23963 56622 23965 56644
rect 23965 56622 24017 56644
rect 24017 56622 24019 56644
rect 23963 56610 24019 56622
rect 23963 56588 23965 56610
rect 23965 56588 24017 56610
rect 24017 56588 24019 56610
rect 23963 56558 23965 56564
rect 23965 56558 24017 56564
rect 24017 56558 24019 56564
rect 23963 56546 24019 56558
rect 23963 56508 23965 56546
rect 23965 56508 24017 56546
rect 24017 56508 24019 56546
rect 23963 56482 24019 56484
rect 23963 56430 23965 56482
rect 23965 56430 24017 56482
rect 24017 56430 24019 56482
rect 23963 56428 24019 56430
rect 23963 56366 23965 56404
rect 23965 56366 24017 56404
rect 24017 56366 24019 56404
rect 23963 56354 24019 56366
rect 23963 56348 23965 56354
rect 23965 56348 24017 56354
rect 24017 56348 24019 56354
rect 23963 56302 23965 56324
rect 23965 56302 24017 56324
rect 24017 56302 24019 56324
rect 23963 56290 24019 56302
rect 23963 56268 23965 56290
rect 23965 56268 24017 56290
rect 24017 56268 24019 56290
rect 23963 56238 23965 56244
rect 23965 56238 24017 56244
rect 24017 56238 24019 56244
rect 23963 56226 24019 56238
rect 23963 56188 23965 56226
rect 23965 56188 24017 56226
rect 24017 56188 24019 56226
rect 25051 56686 25053 56724
rect 25053 56686 25105 56724
rect 25105 56686 25107 56724
rect 25051 56674 25107 56686
rect 25051 56668 25053 56674
rect 25053 56668 25105 56674
rect 25105 56668 25107 56674
rect 25051 56622 25053 56644
rect 25053 56622 25105 56644
rect 25105 56622 25107 56644
rect 25051 56610 25107 56622
rect 25051 56588 25053 56610
rect 25053 56588 25105 56610
rect 25105 56588 25107 56610
rect 25051 56558 25053 56564
rect 25053 56558 25105 56564
rect 25105 56558 25107 56564
rect 25051 56546 25107 56558
rect 25051 56508 25053 56546
rect 25053 56508 25105 56546
rect 25105 56508 25107 56546
rect 25051 56482 25107 56484
rect 25051 56430 25053 56482
rect 25053 56430 25105 56482
rect 25105 56430 25107 56482
rect 25051 56428 25107 56430
rect 25051 56366 25053 56404
rect 25053 56366 25105 56404
rect 25105 56366 25107 56404
rect 25051 56354 25107 56366
rect 25051 56348 25053 56354
rect 25053 56348 25105 56354
rect 25105 56348 25107 56354
rect 25051 56302 25053 56324
rect 25053 56302 25105 56324
rect 25105 56302 25107 56324
rect 25051 56290 25107 56302
rect 25051 56268 25053 56290
rect 25053 56268 25105 56290
rect 25105 56268 25107 56290
rect 25051 56238 25053 56244
rect 25053 56238 25105 56244
rect 25105 56238 25107 56244
rect 25051 56226 25107 56238
rect 25051 56188 25053 56226
rect 25053 56188 25105 56226
rect 25105 56188 25107 56226
rect 26139 56686 26141 56724
rect 26141 56686 26193 56724
rect 26193 56686 26195 56724
rect 26139 56674 26195 56686
rect 26139 56668 26141 56674
rect 26141 56668 26193 56674
rect 26193 56668 26195 56674
rect 26139 56622 26141 56644
rect 26141 56622 26193 56644
rect 26193 56622 26195 56644
rect 26139 56610 26195 56622
rect 26139 56588 26141 56610
rect 26141 56588 26193 56610
rect 26193 56588 26195 56610
rect 26139 56558 26141 56564
rect 26141 56558 26193 56564
rect 26193 56558 26195 56564
rect 26139 56546 26195 56558
rect 26139 56508 26141 56546
rect 26141 56508 26193 56546
rect 26193 56508 26195 56546
rect 26139 56482 26195 56484
rect 26139 56430 26141 56482
rect 26141 56430 26193 56482
rect 26193 56430 26195 56482
rect 26139 56428 26195 56430
rect 26139 56366 26141 56404
rect 26141 56366 26193 56404
rect 26193 56366 26195 56404
rect 26139 56354 26195 56366
rect 26139 56348 26141 56354
rect 26141 56348 26193 56354
rect 26193 56348 26195 56354
rect 26139 56302 26141 56324
rect 26141 56302 26193 56324
rect 26193 56302 26195 56324
rect 26139 56290 26195 56302
rect 26139 56268 26141 56290
rect 26141 56268 26193 56290
rect 26193 56268 26195 56290
rect 26139 56238 26141 56244
rect 26141 56238 26193 56244
rect 26193 56238 26195 56244
rect 26139 56226 26195 56238
rect 26139 56188 26141 56226
rect 26141 56188 26193 56226
rect 26193 56188 26195 56226
rect 27227 56686 27229 56724
rect 27229 56686 27281 56724
rect 27281 56686 27283 56724
rect 27227 56674 27283 56686
rect 27227 56668 27229 56674
rect 27229 56668 27281 56674
rect 27281 56668 27283 56674
rect 27227 56622 27229 56644
rect 27229 56622 27281 56644
rect 27281 56622 27283 56644
rect 27227 56610 27283 56622
rect 27227 56588 27229 56610
rect 27229 56588 27281 56610
rect 27281 56588 27283 56610
rect 27227 56558 27229 56564
rect 27229 56558 27281 56564
rect 27281 56558 27283 56564
rect 27227 56546 27283 56558
rect 27227 56508 27229 56546
rect 27229 56508 27281 56546
rect 27281 56508 27283 56546
rect 27227 56482 27283 56484
rect 27227 56430 27229 56482
rect 27229 56430 27281 56482
rect 27281 56430 27283 56482
rect 27227 56428 27283 56430
rect 27227 56366 27229 56404
rect 27229 56366 27281 56404
rect 27281 56366 27283 56404
rect 27227 56354 27283 56366
rect 27227 56348 27229 56354
rect 27229 56348 27281 56354
rect 27281 56348 27283 56354
rect 27227 56302 27229 56324
rect 27229 56302 27281 56324
rect 27281 56302 27283 56324
rect 27227 56290 27283 56302
rect 27227 56268 27229 56290
rect 27229 56268 27281 56290
rect 27281 56268 27283 56290
rect 27227 56238 27229 56244
rect 27229 56238 27281 56244
rect 27281 56238 27283 56244
rect 27227 56226 27283 56238
rect 27227 56188 27229 56226
rect 27229 56188 27281 56226
rect 27281 56188 27283 56226
rect 28315 56686 28317 56724
rect 28317 56686 28369 56724
rect 28369 56686 28371 56724
rect 28315 56674 28371 56686
rect 28315 56668 28317 56674
rect 28317 56668 28369 56674
rect 28369 56668 28371 56674
rect 28315 56622 28317 56644
rect 28317 56622 28369 56644
rect 28369 56622 28371 56644
rect 28315 56610 28371 56622
rect 28315 56588 28317 56610
rect 28317 56588 28369 56610
rect 28369 56588 28371 56610
rect 28315 56558 28317 56564
rect 28317 56558 28369 56564
rect 28369 56558 28371 56564
rect 28315 56546 28371 56558
rect 28315 56508 28317 56546
rect 28317 56508 28369 56546
rect 28369 56508 28371 56546
rect 28315 56482 28371 56484
rect 28315 56430 28317 56482
rect 28317 56430 28369 56482
rect 28369 56430 28371 56482
rect 28315 56428 28371 56430
rect 28315 56366 28317 56404
rect 28317 56366 28369 56404
rect 28369 56366 28371 56404
rect 28315 56354 28371 56366
rect 28315 56348 28317 56354
rect 28317 56348 28369 56354
rect 28369 56348 28371 56354
rect 28315 56302 28317 56324
rect 28317 56302 28369 56324
rect 28369 56302 28371 56324
rect 28315 56290 28371 56302
rect 28315 56268 28317 56290
rect 28317 56268 28369 56290
rect 28369 56268 28371 56290
rect 28315 56238 28317 56244
rect 28317 56238 28369 56244
rect 28369 56238 28371 56244
rect 28315 56226 28371 56238
rect 28315 56188 28317 56226
rect 28317 56188 28369 56226
rect 28369 56188 28371 56226
rect 29403 56686 29405 56724
rect 29405 56686 29457 56724
rect 29457 56686 29459 56724
rect 29403 56674 29459 56686
rect 29403 56668 29405 56674
rect 29405 56668 29457 56674
rect 29457 56668 29459 56674
rect 29403 56622 29405 56644
rect 29405 56622 29457 56644
rect 29457 56622 29459 56644
rect 29403 56610 29459 56622
rect 29403 56588 29405 56610
rect 29405 56588 29457 56610
rect 29457 56588 29459 56610
rect 29403 56558 29405 56564
rect 29405 56558 29457 56564
rect 29457 56558 29459 56564
rect 29403 56546 29459 56558
rect 29403 56508 29405 56546
rect 29405 56508 29457 56546
rect 29457 56508 29459 56546
rect 29403 56482 29459 56484
rect 29403 56430 29405 56482
rect 29405 56430 29457 56482
rect 29457 56430 29459 56482
rect 29403 56428 29459 56430
rect 29403 56366 29405 56404
rect 29405 56366 29457 56404
rect 29457 56366 29459 56404
rect 29403 56354 29459 56366
rect 29403 56348 29405 56354
rect 29405 56348 29457 56354
rect 29457 56348 29459 56354
rect 29403 56302 29405 56324
rect 29405 56302 29457 56324
rect 29457 56302 29459 56324
rect 29403 56290 29459 56302
rect 29403 56268 29405 56290
rect 29405 56268 29457 56290
rect 29457 56268 29459 56290
rect 29403 56238 29405 56244
rect 29405 56238 29457 56244
rect 29457 56238 29459 56244
rect 29403 56226 29459 56238
rect 29403 56188 29405 56226
rect 29405 56188 29457 56226
rect 29457 56188 29459 56226
rect 30491 56686 30493 56724
rect 30493 56686 30545 56724
rect 30545 56686 30547 56724
rect 30491 56674 30547 56686
rect 30491 56668 30493 56674
rect 30493 56668 30545 56674
rect 30545 56668 30547 56674
rect 30491 56622 30493 56644
rect 30493 56622 30545 56644
rect 30545 56622 30547 56644
rect 30491 56610 30547 56622
rect 30491 56588 30493 56610
rect 30493 56588 30545 56610
rect 30545 56588 30547 56610
rect 30491 56558 30493 56564
rect 30493 56558 30545 56564
rect 30545 56558 30547 56564
rect 30491 56546 30547 56558
rect 30491 56508 30493 56546
rect 30493 56508 30545 56546
rect 30545 56508 30547 56546
rect 30491 56482 30547 56484
rect 30491 56430 30493 56482
rect 30493 56430 30545 56482
rect 30545 56430 30547 56482
rect 30491 56428 30547 56430
rect 30491 56366 30493 56404
rect 30493 56366 30545 56404
rect 30545 56366 30547 56404
rect 30491 56354 30547 56366
rect 30491 56348 30493 56354
rect 30493 56348 30545 56354
rect 30545 56348 30547 56354
rect 30491 56302 30493 56324
rect 30493 56302 30545 56324
rect 30545 56302 30547 56324
rect 30491 56290 30547 56302
rect 30491 56268 30493 56290
rect 30493 56268 30545 56290
rect 30545 56268 30547 56290
rect 30491 56238 30493 56244
rect 30493 56238 30545 56244
rect 30545 56238 30547 56244
rect 30491 56226 30547 56238
rect 30491 56188 30493 56226
rect 30493 56188 30545 56226
rect 30545 56188 30547 56226
rect 31579 56686 31581 56724
rect 31581 56686 31633 56724
rect 31633 56686 31635 56724
rect 31579 56674 31635 56686
rect 31579 56668 31581 56674
rect 31581 56668 31633 56674
rect 31633 56668 31635 56674
rect 31579 56622 31581 56644
rect 31581 56622 31633 56644
rect 31633 56622 31635 56644
rect 31579 56610 31635 56622
rect 31579 56588 31581 56610
rect 31581 56588 31633 56610
rect 31633 56588 31635 56610
rect 31579 56558 31581 56564
rect 31581 56558 31633 56564
rect 31633 56558 31635 56564
rect 31579 56546 31635 56558
rect 31579 56508 31581 56546
rect 31581 56508 31633 56546
rect 31633 56508 31635 56546
rect 31579 56482 31635 56484
rect 31579 56430 31581 56482
rect 31581 56430 31633 56482
rect 31633 56430 31635 56482
rect 31579 56428 31635 56430
rect 31579 56366 31581 56404
rect 31581 56366 31633 56404
rect 31633 56366 31635 56404
rect 31579 56354 31635 56366
rect 31579 56348 31581 56354
rect 31581 56348 31633 56354
rect 31633 56348 31635 56354
rect 31579 56302 31581 56324
rect 31581 56302 31633 56324
rect 31633 56302 31635 56324
rect 31579 56290 31635 56302
rect 31579 56268 31581 56290
rect 31581 56268 31633 56290
rect 31633 56268 31635 56290
rect 31579 56238 31581 56244
rect 31581 56238 31633 56244
rect 31633 56238 31635 56244
rect 31579 56226 31635 56238
rect 31579 56188 31581 56226
rect 31581 56188 31633 56226
rect 31633 56188 31635 56226
rect 17980 54683 17982 54721
rect 17982 54683 18034 54721
rect 18034 54683 18036 54721
rect 17980 54671 18036 54683
rect 17980 54665 17982 54671
rect 17982 54665 18034 54671
rect 18034 54665 18036 54671
rect 17980 54619 17982 54641
rect 17982 54619 18034 54641
rect 18034 54619 18036 54641
rect 17980 54607 18036 54619
rect 17980 54585 17982 54607
rect 17982 54585 18034 54607
rect 18034 54585 18036 54607
rect 17980 54555 17982 54561
rect 17982 54555 18034 54561
rect 18034 54555 18036 54561
rect 17980 54543 18036 54555
rect 17980 54505 17982 54543
rect 17982 54505 18034 54543
rect 18034 54505 18036 54543
rect 17980 54479 18036 54481
rect 17980 54427 17982 54479
rect 17982 54427 18034 54479
rect 18034 54427 18036 54479
rect 17980 54425 18036 54427
rect 17980 54363 17982 54401
rect 17982 54363 18034 54401
rect 18034 54363 18036 54401
rect 17980 54351 18036 54363
rect 17980 54345 17982 54351
rect 17982 54345 18034 54351
rect 18034 54345 18036 54351
rect 17980 54299 17982 54321
rect 17982 54299 18034 54321
rect 18034 54299 18036 54321
rect 17980 54287 18036 54299
rect 17980 54265 17982 54287
rect 17982 54265 18034 54287
rect 18034 54265 18036 54287
rect 17980 54235 17982 54241
rect 17982 54235 18034 54241
rect 18034 54235 18036 54241
rect 17980 54223 18036 54235
rect 17980 54185 17982 54223
rect 17982 54185 18034 54223
rect 18034 54185 18036 54223
rect 19068 54683 19070 54721
rect 19070 54683 19122 54721
rect 19122 54683 19124 54721
rect 19068 54671 19124 54683
rect 19068 54665 19070 54671
rect 19070 54665 19122 54671
rect 19122 54665 19124 54671
rect 19068 54619 19070 54641
rect 19070 54619 19122 54641
rect 19122 54619 19124 54641
rect 19068 54607 19124 54619
rect 19068 54585 19070 54607
rect 19070 54585 19122 54607
rect 19122 54585 19124 54607
rect 19068 54555 19070 54561
rect 19070 54555 19122 54561
rect 19122 54555 19124 54561
rect 19068 54543 19124 54555
rect 19068 54505 19070 54543
rect 19070 54505 19122 54543
rect 19122 54505 19124 54543
rect 19068 54479 19124 54481
rect 19068 54427 19070 54479
rect 19070 54427 19122 54479
rect 19122 54427 19124 54479
rect 19068 54425 19124 54427
rect 19068 54363 19070 54401
rect 19070 54363 19122 54401
rect 19122 54363 19124 54401
rect 19068 54351 19124 54363
rect 19068 54345 19070 54351
rect 19070 54345 19122 54351
rect 19122 54345 19124 54351
rect 19068 54299 19070 54321
rect 19070 54299 19122 54321
rect 19122 54299 19124 54321
rect 19068 54287 19124 54299
rect 19068 54265 19070 54287
rect 19070 54265 19122 54287
rect 19122 54265 19124 54287
rect 19068 54235 19070 54241
rect 19070 54235 19122 54241
rect 19122 54235 19124 54241
rect 19068 54223 19124 54235
rect 19068 54185 19070 54223
rect 19070 54185 19122 54223
rect 19122 54185 19124 54223
rect 20156 54683 20158 54721
rect 20158 54683 20210 54721
rect 20210 54683 20212 54721
rect 20156 54671 20212 54683
rect 20156 54665 20158 54671
rect 20158 54665 20210 54671
rect 20210 54665 20212 54671
rect 20156 54619 20158 54641
rect 20158 54619 20210 54641
rect 20210 54619 20212 54641
rect 20156 54607 20212 54619
rect 20156 54585 20158 54607
rect 20158 54585 20210 54607
rect 20210 54585 20212 54607
rect 20156 54555 20158 54561
rect 20158 54555 20210 54561
rect 20210 54555 20212 54561
rect 20156 54543 20212 54555
rect 20156 54505 20158 54543
rect 20158 54505 20210 54543
rect 20210 54505 20212 54543
rect 20156 54479 20212 54481
rect 20156 54427 20158 54479
rect 20158 54427 20210 54479
rect 20210 54427 20212 54479
rect 20156 54425 20212 54427
rect 20156 54363 20158 54401
rect 20158 54363 20210 54401
rect 20210 54363 20212 54401
rect 20156 54351 20212 54363
rect 20156 54345 20158 54351
rect 20158 54345 20210 54351
rect 20210 54345 20212 54351
rect 20156 54299 20158 54321
rect 20158 54299 20210 54321
rect 20210 54299 20212 54321
rect 20156 54287 20212 54299
rect 20156 54265 20158 54287
rect 20158 54265 20210 54287
rect 20210 54265 20212 54287
rect 20156 54235 20158 54241
rect 20158 54235 20210 54241
rect 20210 54235 20212 54241
rect 20156 54223 20212 54235
rect 20156 54185 20158 54223
rect 20158 54185 20210 54223
rect 20210 54185 20212 54223
rect 21244 54683 21246 54721
rect 21246 54683 21298 54721
rect 21298 54683 21300 54721
rect 21244 54671 21300 54683
rect 21244 54665 21246 54671
rect 21246 54665 21298 54671
rect 21298 54665 21300 54671
rect 21244 54619 21246 54641
rect 21246 54619 21298 54641
rect 21298 54619 21300 54641
rect 21244 54607 21300 54619
rect 21244 54585 21246 54607
rect 21246 54585 21298 54607
rect 21298 54585 21300 54607
rect 21244 54555 21246 54561
rect 21246 54555 21298 54561
rect 21298 54555 21300 54561
rect 21244 54543 21300 54555
rect 21244 54505 21246 54543
rect 21246 54505 21298 54543
rect 21298 54505 21300 54543
rect 21244 54479 21300 54481
rect 21244 54427 21246 54479
rect 21246 54427 21298 54479
rect 21298 54427 21300 54479
rect 21244 54425 21300 54427
rect 21244 54363 21246 54401
rect 21246 54363 21298 54401
rect 21298 54363 21300 54401
rect 21244 54351 21300 54363
rect 21244 54345 21246 54351
rect 21246 54345 21298 54351
rect 21298 54345 21300 54351
rect 21244 54299 21246 54321
rect 21246 54299 21298 54321
rect 21298 54299 21300 54321
rect 21244 54287 21300 54299
rect 21244 54265 21246 54287
rect 21246 54265 21298 54287
rect 21298 54265 21300 54287
rect 21244 54235 21246 54241
rect 21246 54235 21298 54241
rect 21298 54235 21300 54241
rect 21244 54223 21300 54235
rect 21244 54185 21246 54223
rect 21246 54185 21298 54223
rect 21298 54185 21300 54223
rect 22332 54683 22334 54721
rect 22334 54683 22386 54721
rect 22386 54683 22388 54721
rect 22332 54671 22388 54683
rect 22332 54665 22334 54671
rect 22334 54665 22386 54671
rect 22386 54665 22388 54671
rect 22332 54619 22334 54641
rect 22334 54619 22386 54641
rect 22386 54619 22388 54641
rect 22332 54607 22388 54619
rect 22332 54585 22334 54607
rect 22334 54585 22386 54607
rect 22386 54585 22388 54607
rect 22332 54555 22334 54561
rect 22334 54555 22386 54561
rect 22386 54555 22388 54561
rect 22332 54543 22388 54555
rect 22332 54505 22334 54543
rect 22334 54505 22386 54543
rect 22386 54505 22388 54543
rect 22332 54479 22388 54481
rect 22332 54427 22334 54479
rect 22334 54427 22386 54479
rect 22386 54427 22388 54479
rect 22332 54425 22388 54427
rect 22332 54363 22334 54401
rect 22334 54363 22386 54401
rect 22386 54363 22388 54401
rect 22332 54351 22388 54363
rect 22332 54345 22334 54351
rect 22334 54345 22386 54351
rect 22386 54345 22388 54351
rect 22332 54299 22334 54321
rect 22334 54299 22386 54321
rect 22386 54299 22388 54321
rect 22332 54287 22388 54299
rect 22332 54265 22334 54287
rect 22334 54265 22386 54287
rect 22386 54265 22388 54287
rect 22332 54235 22334 54241
rect 22334 54235 22386 54241
rect 22386 54235 22388 54241
rect 22332 54223 22388 54235
rect 22332 54185 22334 54223
rect 22334 54185 22386 54223
rect 22386 54185 22388 54223
rect 23420 54683 23422 54721
rect 23422 54683 23474 54721
rect 23474 54683 23476 54721
rect 23420 54671 23476 54683
rect 23420 54665 23422 54671
rect 23422 54665 23474 54671
rect 23474 54665 23476 54671
rect 23420 54619 23422 54641
rect 23422 54619 23474 54641
rect 23474 54619 23476 54641
rect 23420 54607 23476 54619
rect 23420 54585 23422 54607
rect 23422 54585 23474 54607
rect 23474 54585 23476 54607
rect 23420 54555 23422 54561
rect 23422 54555 23474 54561
rect 23474 54555 23476 54561
rect 23420 54543 23476 54555
rect 23420 54505 23422 54543
rect 23422 54505 23474 54543
rect 23474 54505 23476 54543
rect 23420 54479 23476 54481
rect 23420 54427 23422 54479
rect 23422 54427 23474 54479
rect 23474 54427 23476 54479
rect 23420 54425 23476 54427
rect 23420 54363 23422 54401
rect 23422 54363 23474 54401
rect 23474 54363 23476 54401
rect 23420 54351 23476 54363
rect 23420 54345 23422 54351
rect 23422 54345 23474 54351
rect 23474 54345 23476 54351
rect 23420 54299 23422 54321
rect 23422 54299 23474 54321
rect 23474 54299 23476 54321
rect 23420 54287 23476 54299
rect 23420 54265 23422 54287
rect 23422 54265 23474 54287
rect 23474 54265 23476 54287
rect 23420 54235 23422 54241
rect 23422 54235 23474 54241
rect 23474 54235 23476 54241
rect 23420 54223 23476 54235
rect 23420 54185 23422 54223
rect 23422 54185 23474 54223
rect 23474 54185 23476 54223
rect 24508 54683 24510 54721
rect 24510 54683 24562 54721
rect 24562 54683 24564 54721
rect 24508 54671 24564 54683
rect 24508 54665 24510 54671
rect 24510 54665 24562 54671
rect 24562 54665 24564 54671
rect 24508 54619 24510 54641
rect 24510 54619 24562 54641
rect 24562 54619 24564 54641
rect 24508 54607 24564 54619
rect 24508 54585 24510 54607
rect 24510 54585 24562 54607
rect 24562 54585 24564 54607
rect 24508 54555 24510 54561
rect 24510 54555 24562 54561
rect 24562 54555 24564 54561
rect 24508 54543 24564 54555
rect 24508 54505 24510 54543
rect 24510 54505 24562 54543
rect 24562 54505 24564 54543
rect 24508 54479 24564 54481
rect 24508 54427 24510 54479
rect 24510 54427 24562 54479
rect 24562 54427 24564 54479
rect 24508 54425 24564 54427
rect 24508 54363 24510 54401
rect 24510 54363 24562 54401
rect 24562 54363 24564 54401
rect 24508 54351 24564 54363
rect 24508 54345 24510 54351
rect 24510 54345 24562 54351
rect 24562 54345 24564 54351
rect 24508 54299 24510 54321
rect 24510 54299 24562 54321
rect 24562 54299 24564 54321
rect 24508 54287 24564 54299
rect 24508 54265 24510 54287
rect 24510 54265 24562 54287
rect 24562 54265 24564 54287
rect 24508 54235 24510 54241
rect 24510 54235 24562 54241
rect 24562 54235 24564 54241
rect 24508 54223 24564 54235
rect 24508 54185 24510 54223
rect 24510 54185 24562 54223
rect 24562 54185 24564 54223
rect 25596 54683 25598 54721
rect 25598 54683 25650 54721
rect 25650 54683 25652 54721
rect 25596 54671 25652 54683
rect 25596 54665 25598 54671
rect 25598 54665 25650 54671
rect 25650 54665 25652 54671
rect 25596 54619 25598 54641
rect 25598 54619 25650 54641
rect 25650 54619 25652 54641
rect 25596 54607 25652 54619
rect 25596 54585 25598 54607
rect 25598 54585 25650 54607
rect 25650 54585 25652 54607
rect 25596 54555 25598 54561
rect 25598 54555 25650 54561
rect 25650 54555 25652 54561
rect 25596 54543 25652 54555
rect 25596 54505 25598 54543
rect 25598 54505 25650 54543
rect 25650 54505 25652 54543
rect 25596 54479 25652 54481
rect 25596 54427 25598 54479
rect 25598 54427 25650 54479
rect 25650 54427 25652 54479
rect 25596 54425 25652 54427
rect 25596 54363 25598 54401
rect 25598 54363 25650 54401
rect 25650 54363 25652 54401
rect 25596 54351 25652 54363
rect 25596 54345 25598 54351
rect 25598 54345 25650 54351
rect 25650 54345 25652 54351
rect 25596 54299 25598 54321
rect 25598 54299 25650 54321
rect 25650 54299 25652 54321
rect 25596 54287 25652 54299
rect 25596 54265 25598 54287
rect 25598 54265 25650 54287
rect 25650 54265 25652 54287
rect 25596 54235 25598 54241
rect 25598 54235 25650 54241
rect 25650 54235 25652 54241
rect 25596 54223 25652 54235
rect 25596 54185 25598 54223
rect 25598 54185 25650 54223
rect 25650 54185 25652 54223
rect 26684 54683 26686 54721
rect 26686 54683 26738 54721
rect 26738 54683 26740 54721
rect 26684 54671 26740 54683
rect 26684 54665 26686 54671
rect 26686 54665 26738 54671
rect 26738 54665 26740 54671
rect 26684 54619 26686 54641
rect 26686 54619 26738 54641
rect 26738 54619 26740 54641
rect 26684 54607 26740 54619
rect 26684 54585 26686 54607
rect 26686 54585 26738 54607
rect 26738 54585 26740 54607
rect 26684 54555 26686 54561
rect 26686 54555 26738 54561
rect 26738 54555 26740 54561
rect 26684 54543 26740 54555
rect 26684 54505 26686 54543
rect 26686 54505 26738 54543
rect 26738 54505 26740 54543
rect 26684 54479 26740 54481
rect 26684 54427 26686 54479
rect 26686 54427 26738 54479
rect 26738 54427 26740 54479
rect 26684 54425 26740 54427
rect 26684 54363 26686 54401
rect 26686 54363 26738 54401
rect 26738 54363 26740 54401
rect 26684 54351 26740 54363
rect 26684 54345 26686 54351
rect 26686 54345 26738 54351
rect 26738 54345 26740 54351
rect 26684 54299 26686 54321
rect 26686 54299 26738 54321
rect 26738 54299 26740 54321
rect 26684 54287 26740 54299
rect 26684 54265 26686 54287
rect 26686 54265 26738 54287
rect 26738 54265 26740 54287
rect 26684 54235 26686 54241
rect 26686 54235 26738 54241
rect 26738 54235 26740 54241
rect 26684 54223 26740 54235
rect 26684 54185 26686 54223
rect 26686 54185 26738 54223
rect 26738 54185 26740 54223
rect 27772 54683 27774 54721
rect 27774 54683 27826 54721
rect 27826 54683 27828 54721
rect 27772 54671 27828 54683
rect 27772 54665 27774 54671
rect 27774 54665 27826 54671
rect 27826 54665 27828 54671
rect 27772 54619 27774 54641
rect 27774 54619 27826 54641
rect 27826 54619 27828 54641
rect 27772 54607 27828 54619
rect 27772 54585 27774 54607
rect 27774 54585 27826 54607
rect 27826 54585 27828 54607
rect 27772 54555 27774 54561
rect 27774 54555 27826 54561
rect 27826 54555 27828 54561
rect 27772 54543 27828 54555
rect 27772 54505 27774 54543
rect 27774 54505 27826 54543
rect 27826 54505 27828 54543
rect 27772 54479 27828 54481
rect 27772 54427 27774 54479
rect 27774 54427 27826 54479
rect 27826 54427 27828 54479
rect 27772 54425 27828 54427
rect 27772 54363 27774 54401
rect 27774 54363 27826 54401
rect 27826 54363 27828 54401
rect 27772 54351 27828 54363
rect 27772 54345 27774 54351
rect 27774 54345 27826 54351
rect 27826 54345 27828 54351
rect 27772 54299 27774 54321
rect 27774 54299 27826 54321
rect 27826 54299 27828 54321
rect 27772 54287 27828 54299
rect 27772 54265 27774 54287
rect 27774 54265 27826 54287
rect 27826 54265 27828 54287
rect 27772 54235 27774 54241
rect 27774 54235 27826 54241
rect 27826 54235 27828 54241
rect 27772 54223 27828 54235
rect 27772 54185 27774 54223
rect 27774 54185 27826 54223
rect 27826 54185 27828 54223
rect 28860 54683 28862 54721
rect 28862 54683 28914 54721
rect 28914 54683 28916 54721
rect 28860 54671 28916 54683
rect 28860 54665 28862 54671
rect 28862 54665 28914 54671
rect 28914 54665 28916 54671
rect 28860 54619 28862 54641
rect 28862 54619 28914 54641
rect 28914 54619 28916 54641
rect 28860 54607 28916 54619
rect 28860 54585 28862 54607
rect 28862 54585 28914 54607
rect 28914 54585 28916 54607
rect 28860 54555 28862 54561
rect 28862 54555 28914 54561
rect 28914 54555 28916 54561
rect 28860 54543 28916 54555
rect 28860 54505 28862 54543
rect 28862 54505 28914 54543
rect 28914 54505 28916 54543
rect 28860 54479 28916 54481
rect 28860 54427 28862 54479
rect 28862 54427 28914 54479
rect 28914 54427 28916 54479
rect 28860 54425 28916 54427
rect 28860 54363 28862 54401
rect 28862 54363 28914 54401
rect 28914 54363 28916 54401
rect 28860 54351 28916 54363
rect 28860 54345 28862 54351
rect 28862 54345 28914 54351
rect 28914 54345 28916 54351
rect 28860 54299 28862 54321
rect 28862 54299 28914 54321
rect 28914 54299 28916 54321
rect 28860 54287 28916 54299
rect 28860 54265 28862 54287
rect 28862 54265 28914 54287
rect 28914 54265 28916 54287
rect 28860 54235 28862 54241
rect 28862 54235 28914 54241
rect 28914 54235 28916 54241
rect 28860 54223 28916 54235
rect 28860 54185 28862 54223
rect 28862 54185 28914 54223
rect 28914 54185 28916 54223
rect 29948 54683 29950 54721
rect 29950 54683 30002 54721
rect 30002 54683 30004 54721
rect 29948 54671 30004 54683
rect 29948 54665 29950 54671
rect 29950 54665 30002 54671
rect 30002 54665 30004 54671
rect 29948 54619 29950 54641
rect 29950 54619 30002 54641
rect 30002 54619 30004 54641
rect 29948 54607 30004 54619
rect 29948 54585 29950 54607
rect 29950 54585 30002 54607
rect 30002 54585 30004 54607
rect 29948 54555 29950 54561
rect 29950 54555 30002 54561
rect 30002 54555 30004 54561
rect 29948 54543 30004 54555
rect 29948 54505 29950 54543
rect 29950 54505 30002 54543
rect 30002 54505 30004 54543
rect 29948 54479 30004 54481
rect 29948 54427 29950 54479
rect 29950 54427 30002 54479
rect 30002 54427 30004 54479
rect 29948 54425 30004 54427
rect 29948 54363 29950 54401
rect 29950 54363 30002 54401
rect 30002 54363 30004 54401
rect 29948 54351 30004 54363
rect 29948 54345 29950 54351
rect 29950 54345 30002 54351
rect 30002 54345 30004 54351
rect 29948 54299 29950 54321
rect 29950 54299 30002 54321
rect 30002 54299 30004 54321
rect 29948 54287 30004 54299
rect 29948 54265 29950 54287
rect 29950 54265 30002 54287
rect 30002 54265 30004 54287
rect 29948 54235 29950 54241
rect 29950 54235 30002 54241
rect 30002 54235 30004 54241
rect 29948 54223 30004 54235
rect 29948 54185 29950 54223
rect 29950 54185 30002 54223
rect 30002 54185 30004 54223
rect 31036 54683 31038 54721
rect 31038 54683 31090 54721
rect 31090 54683 31092 54721
rect 31036 54671 31092 54683
rect 31036 54665 31038 54671
rect 31038 54665 31090 54671
rect 31090 54665 31092 54671
rect 31036 54619 31038 54641
rect 31038 54619 31090 54641
rect 31090 54619 31092 54641
rect 31036 54607 31092 54619
rect 31036 54585 31038 54607
rect 31038 54585 31090 54607
rect 31090 54585 31092 54607
rect 31036 54555 31038 54561
rect 31038 54555 31090 54561
rect 31090 54555 31092 54561
rect 31036 54543 31092 54555
rect 31036 54505 31038 54543
rect 31038 54505 31090 54543
rect 31090 54505 31092 54543
rect 31036 54479 31092 54481
rect 31036 54427 31038 54479
rect 31038 54427 31090 54479
rect 31090 54427 31092 54479
rect 31036 54425 31092 54427
rect 31036 54363 31038 54401
rect 31038 54363 31090 54401
rect 31090 54363 31092 54401
rect 31036 54351 31092 54363
rect 31036 54345 31038 54351
rect 31038 54345 31090 54351
rect 31090 54345 31092 54351
rect 31036 54299 31038 54321
rect 31038 54299 31090 54321
rect 31090 54299 31092 54321
rect 31036 54287 31092 54299
rect 31036 54265 31038 54287
rect 31038 54265 31090 54287
rect 31090 54265 31092 54287
rect 31036 54235 31038 54241
rect 31038 54235 31090 54241
rect 31090 54235 31092 54241
rect 31036 54223 31092 54235
rect 31036 54185 31038 54223
rect 31038 54185 31090 54223
rect 31090 54185 31092 54223
rect 17435 52686 17437 52724
rect 17437 52686 17489 52724
rect 17489 52686 17491 52724
rect 17435 52674 17491 52686
rect 17435 52668 17437 52674
rect 17437 52668 17489 52674
rect 17489 52668 17491 52674
rect 17435 52622 17437 52644
rect 17437 52622 17489 52644
rect 17489 52622 17491 52644
rect 17435 52610 17491 52622
rect 17435 52588 17437 52610
rect 17437 52588 17489 52610
rect 17489 52588 17491 52610
rect 17435 52558 17437 52564
rect 17437 52558 17489 52564
rect 17489 52558 17491 52564
rect 17435 52546 17491 52558
rect 17435 52508 17437 52546
rect 17437 52508 17489 52546
rect 17489 52508 17491 52546
rect 17435 52482 17491 52484
rect 17435 52430 17437 52482
rect 17437 52430 17489 52482
rect 17489 52430 17491 52482
rect 17435 52428 17491 52430
rect 17435 52366 17437 52404
rect 17437 52366 17489 52404
rect 17489 52366 17491 52404
rect 17435 52354 17491 52366
rect 17435 52348 17437 52354
rect 17437 52348 17489 52354
rect 17489 52348 17491 52354
rect 17435 52302 17437 52324
rect 17437 52302 17489 52324
rect 17489 52302 17491 52324
rect 17435 52290 17491 52302
rect 17435 52268 17437 52290
rect 17437 52268 17489 52290
rect 17489 52268 17491 52290
rect 17435 52238 17437 52244
rect 17437 52238 17489 52244
rect 17489 52238 17491 52244
rect 17435 52226 17491 52238
rect 17435 52188 17437 52226
rect 17437 52188 17489 52226
rect 17489 52188 17491 52226
rect 18523 52686 18525 52724
rect 18525 52686 18577 52724
rect 18577 52686 18579 52724
rect 18523 52674 18579 52686
rect 18523 52668 18525 52674
rect 18525 52668 18577 52674
rect 18577 52668 18579 52674
rect 18523 52622 18525 52644
rect 18525 52622 18577 52644
rect 18577 52622 18579 52644
rect 18523 52610 18579 52622
rect 18523 52588 18525 52610
rect 18525 52588 18577 52610
rect 18577 52588 18579 52610
rect 18523 52558 18525 52564
rect 18525 52558 18577 52564
rect 18577 52558 18579 52564
rect 18523 52546 18579 52558
rect 18523 52508 18525 52546
rect 18525 52508 18577 52546
rect 18577 52508 18579 52546
rect 18523 52482 18579 52484
rect 18523 52430 18525 52482
rect 18525 52430 18577 52482
rect 18577 52430 18579 52482
rect 18523 52428 18579 52430
rect 18523 52366 18525 52404
rect 18525 52366 18577 52404
rect 18577 52366 18579 52404
rect 18523 52354 18579 52366
rect 18523 52348 18525 52354
rect 18525 52348 18577 52354
rect 18577 52348 18579 52354
rect 18523 52302 18525 52324
rect 18525 52302 18577 52324
rect 18577 52302 18579 52324
rect 18523 52290 18579 52302
rect 18523 52268 18525 52290
rect 18525 52268 18577 52290
rect 18577 52268 18579 52290
rect 18523 52238 18525 52244
rect 18525 52238 18577 52244
rect 18577 52238 18579 52244
rect 18523 52226 18579 52238
rect 18523 52188 18525 52226
rect 18525 52188 18577 52226
rect 18577 52188 18579 52226
rect 19611 52686 19613 52724
rect 19613 52686 19665 52724
rect 19665 52686 19667 52724
rect 19611 52674 19667 52686
rect 19611 52668 19613 52674
rect 19613 52668 19665 52674
rect 19665 52668 19667 52674
rect 19611 52622 19613 52644
rect 19613 52622 19665 52644
rect 19665 52622 19667 52644
rect 19611 52610 19667 52622
rect 19611 52588 19613 52610
rect 19613 52588 19665 52610
rect 19665 52588 19667 52610
rect 19611 52558 19613 52564
rect 19613 52558 19665 52564
rect 19665 52558 19667 52564
rect 19611 52546 19667 52558
rect 19611 52508 19613 52546
rect 19613 52508 19665 52546
rect 19665 52508 19667 52546
rect 19611 52482 19667 52484
rect 19611 52430 19613 52482
rect 19613 52430 19665 52482
rect 19665 52430 19667 52482
rect 19611 52428 19667 52430
rect 19611 52366 19613 52404
rect 19613 52366 19665 52404
rect 19665 52366 19667 52404
rect 19611 52354 19667 52366
rect 19611 52348 19613 52354
rect 19613 52348 19665 52354
rect 19665 52348 19667 52354
rect 19611 52302 19613 52324
rect 19613 52302 19665 52324
rect 19665 52302 19667 52324
rect 19611 52290 19667 52302
rect 19611 52268 19613 52290
rect 19613 52268 19665 52290
rect 19665 52268 19667 52290
rect 19611 52238 19613 52244
rect 19613 52238 19665 52244
rect 19665 52238 19667 52244
rect 19611 52226 19667 52238
rect 19611 52188 19613 52226
rect 19613 52188 19665 52226
rect 19665 52188 19667 52226
rect 20699 52686 20701 52724
rect 20701 52686 20753 52724
rect 20753 52686 20755 52724
rect 20699 52674 20755 52686
rect 20699 52668 20701 52674
rect 20701 52668 20753 52674
rect 20753 52668 20755 52674
rect 20699 52622 20701 52644
rect 20701 52622 20753 52644
rect 20753 52622 20755 52644
rect 20699 52610 20755 52622
rect 20699 52588 20701 52610
rect 20701 52588 20753 52610
rect 20753 52588 20755 52610
rect 20699 52558 20701 52564
rect 20701 52558 20753 52564
rect 20753 52558 20755 52564
rect 20699 52546 20755 52558
rect 20699 52508 20701 52546
rect 20701 52508 20753 52546
rect 20753 52508 20755 52546
rect 20699 52482 20755 52484
rect 20699 52430 20701 52482
rect 20701 52430 20753 52482
rect 20753 52430 20755 52482
rect 20699 52428 20755 52430
rect 20699 52366 20701 52404
rect 20701 52366 20753 52404
rect 20753 52366 20755 52404
rect 20699 52354 20755 52366
rect 20699 52348 20701 52354
rect 20701 52348 20753 52354
rect 20753 52348 20755 52354
rect 20699 52302 20701 52324
rect 20701 52302 20753 52324
rect 20753 52302 20755 52324
rect 20699 52290 20755 52302
rect 20699 52268 20701 52290
rect 20701 52268 20753 52290
rect 20753 52268 20755 52290
rect 20699 52238 20701 52244
rect 20701 52238 20753 52244
rect 20753 52238 20755 52244
rect 20699 52226 20755 52238
rect 20699 52188 20701 52226
rect 20701 52188 20753 52226
rect 20753 52188 20755 52226
rect 21787 52686 21789 52724
rect 21789 52686 21841 52724
rect 21841 52686 21843 52724
rect 21787 52674 21843 52686
rect 21787 52668 21789 52674
rect 21789 52668 21841 52674
rect 21841 52668 21843 52674
rect 21787 52622 21789 52644
rect 21789 52622 21841 52644
rect 21841 52622 21843 52644
rect 21787 52610 21843 52622
rect 21787 52588 21789 52610
rect 21789 52588 21841 52610
rect 21841 52588 21843 52610
rect 21787 52558 21789 52564
rect 21789 52558 21841 52564
rect 21841 52558 21843 52564
rect 21787 52546 21843 52558
rect 21787 52508 21789 52546
rect 21789 52508 21841 52546
rect 21841 52508 21843 52546
rect 21787 52482 21843 52484
rect 21787 52430 21789 52482
rect 21789 52430 21841 52482
rect 21841 52430 21843 52482
rect 21787 52428 21843 52430
rect 21787 52366 21789 52404
rect 21789 52366 21841 52404
rect 21841 52366 21843 52404
rect 21787 52354 21843 52366
rect 21787 52348 21789 52354
rect 21789 52348 21841 52354
rect 21841 52348 21843 52354
rect 21787 52302 21789 52324
rect 21789 52302 21841 52324
rect 21841 52302 21843 52324
rect 21787 52290 21843 52302
rect 21787 52268 21789 52290
rect 21789 52268 21841 52290
rect 21841 52268 21843 52290
rect 21787 52238 21789 52244
rect 21789 52238 21841 52244
rect 21841 52238 21843 52244
rect 21787 52226 21843 52238
rect 21787 52188 21789 52226
rect 21789 52188 21841 52226
rect 21841 52188 21843 52226
rect 22875 52686 22877 52724
rect 22877 52686 22929 52724
rect 22929 52686 22931 52724
rect 22875 52674 22931 52686
rect 22875 52668 22877 52674
rect 22877 52668 22929 52674
rect 22929 52668 22931 52674
rect 22875 52622 22877 52644
rect 22877 52622 22929 52644
rect 22929 52622 22931 52644
rect 22875 52610 22931 52622
rect 22875 52588 22877 52610
rect 22877 52588 22929 52610
rect 22929 52588 22931 52610
rect 22875 52558 22877 52564
rect 22877 52558 22929 52564
rect 22929 52558 22931 52564
rect 22875 52546 22931 52558
rect 22875 52508 22877 52546
rect 22877 52508 22929 52546
rect 22929 52508 22931 52546
rect 22875 52482 22931 52484
rect 22875 52430 22877 52482
rect 22877 52430 22929 52482
rect 22929 52430 22931 52482
rect 22875 52428 22931 52430
rect 22875 52366 22877 52404
rect 22877 52366 22929 52404
rect 22929 52366 22931 52404
rect 22875 52354 22931 52366
rect 22875 52348 22877 52354
rect 22877 52348 22929 52354
rect 22929 52348 22931 52354
rect 22875 52302 22877 52324
rect 22877 52302 22929 52324
rect 22929 52302 22931 52324
rect 22875 52290 22931 52302
rect 22875 52268 22877 52290
rect 22877 52268 22929 52290
rect 22929 52268 22931 52290
rect 22875 52238 22877 52244
rect 22877 52238 22929 52244
rect 22929 52238 22931 52244
rect 22875 52226 22931 52238
rect 22875 52188 22877 52226
rect 22877 52188 22929 52226
rect 22929 52188 22931 52226
rect 23963 52686 23965 52724
rect 23965 52686 24017 52724
rect 24017 52686 24019 52724
rect 23963 52674 24019 52686
rect 23963 52668 23965 52674
rect 23965 52668 24017 52674
rect 24017 52668 24019 52674
rect 23963 52622 23965 52644
rect 23965 52622 24017 52644
rect 24017 52622 24019 52644
rect 23963 52610 24019 52622
rect 23963 52588 23965 52610
rect 23965 52588 24017 52610
rect 24017 52588 24019 52610
rect 23963 52558 23965 52564
rect 23965 52558 24017 52564
rect 24017 52558 24019 52564
rect 23963 52546 24019 52558
rect 23963 52508 23965 52546
rect 23965 52508 24017 52546
rect 24017 52508 24019 52546
rect 23963 52482 24019 52484
rect 23963 52430 23965 52482
rect 23965 52430 24017 52482
rect 24017 52430 24019 52482
rect 23963 52428 24019 52430
rect 23963 52366 23965 52404
rect 23965 52366 24017 52404
rect 24017 52366 24019 52404
rect 23963 52354 24019 52366
rect 23963 52348 23965 52354
rect 23965 52348 24017 52354
rect 24017 52348 24019 52354
rect 23963 52302 23965 52324
rect 23965 52302 24017 52324
rect 24017 52302 24019 52324
rect 23963 52290 24019 52302
rect 23963 52268 23965 52290
rect 23965 52268 24017 52290
rect 24017 52268 24019 52290
rect 23963 52238 23965 52244
rect 23965 52238 24017 52244
rect 24017 52238 24019 52244
rect 23963 52226 24019 52238
rect 23963 52188 23965 52226
rect 23965 52188 24017 52226
rect 24017 52188 24019 52226
rect 25051 52686 25053 52724
rect 25053 52686 25105 52724
rect 25105 52686 25107 52724
rect 25051 52674 25107 52686
rect 25051 52668 25053 52674
rect 25053 52668 25105 52674
rect 25105 52668 25107 52674
rect 25051 52622 25053 52644
rect 25053 52622 25105 52644
rect 25105 52622 25107 52644
rect 25051 52610 25107 52622
rect 25051 52588 25053 52610
rect 25053 52588 25105 52610
rect 25105 52588 25107 52610
rect 25051 52558 25053 52564
rect 25053 52558 25105 52564
rect 25105 52558 25107 52564
rect 25051 52546 25107 52558
rect 25051 52508 25053 52546
rect 25053 52508 25105 52546
rect 25105 52508 25107 52546
rect 25051 52482 25107 52484
rect 25051 52430 25053 52482
rect 25053 52430 25105 52482
rect 25105 52430 25107 52482
rect 25051 52428 25107 52430
rect 25051 52366 25053 52404
rect 25053 52366 25105 52404
rect 25105 52366 25107 52404
rect 25051 52354 25107 52366
rect 25051 52348 25053 52354
rect 25053 52348 25105 52354
rect 25105 52348 25107 52354
rect 25051 52302 25053 52324
rect 25053 52302 25105 52324
rect 25105 52302 25107 52324
rect 25051 52290 25107 52302
rect 25051 52268 25053 52290
rect 25053 52268 25105 52290
rect 25105 52268 25107 52290
rect 25051 52238 25053 52244
rect 25053 52238 25105 52244
rect 25105 52238 25107 52244
rect 25051 52226 25107 52238
rect 25051 52188 25053 52226
rect 25053 52188 25105 52226
rect 25105 52188 25107 52226
rect 26139 52686 26141 52724
rect 26141 52686 26193 52724
rect 26193 52686 26195 52724
rect 26139 52674 26195 52686
rect 26139 52668 26141 52674
rect 26141 52668 26193 52674
rect 26193 52668 26195 52674
rect 26139 52622 26141 52644
rect 26141 52622 26193 52644
rect 26193 52622 26195 52644
rect 26139 52610 26195 52622
rect 26139 52588 26141 52610
rect 26141 52588 26193 52610
rect 26193 52588 26195 52610
rect 26139 52558 26141 52564
rect 26141 52558 26193 52564
rect 26193 52558 26195 52564
rect 26139 52546 26195 52558
rect 26139 52508 26141 52546
rect 26141 52508 26193 52546
rect 26193 52508 26195 52546
rect 26139 52482 26195 52484
rect 26139 52430 26141 52482
rect 26141 52430 26193 52482
rect 26193 52430 26195 52482
rect 26139 52428 26195 52430
rect 26139 52366 26141 52404
rect 26141 52366 26193 52404
rect 26193 52366 26195 52404
rect 26139 52354 26195 52366
rect 26139 52348 26141 52354
rect 26141 52348 26193 52354
rect 26193 52348 26195 52354
rect 26139 52302 26141 52324
rect 26141 52302 26193 52324
rect 26193 52302 26195 52324
rect 26139 52290 26195 52302
rect 26139 52268 26141 52290
rect 26141 52268 26193 52290
rect 26193 52268 26195 52290
rect 26139 52238 26141 52244
rect 26141 52238 26193 52244
rect 26193 52238 26195 52244
rect 26139 52226 26195 52238
rect 26139 52188 26141 52226
rect 26141 52188 26193 52226
rect 26193 52188 26195 52226
rect 27227 52686 27229 52724
rect 27229 52686 27281 52724
rect 27281 52686 27283 52724
rect 27227 52674 27283 52686
rect 27227 52668 27229 52674
rect 27229 52668 27281 52674
rect 27281 52668 27283 52674
rect 27227 52622 27229 52644
rect 27229 52622 27281 52644
rect 27281 52622 27283 52644
rect 27227 52610 27283 52622
rect 27227 52588 27229 52610
rect 27229 52588 27281 52610
rect 27281 52588 27283 52610
rect 27227 52558 27229 52564
rect 27229 52558 27281 52564
rect 27281 52558 27283 52564
rect 27227 52546 27283 52558
rect 27227 52508 27229 52546
rect 27229 52508 27281 52546
rect 27281 52508 27283 52546
rect 27227 52482 27283 52484
rect 27227 52430 27229 52482
rect 27229 52430 27281 52482
rect 27281 52430 27283 52482
rect 27227 52428 27283 52430
rect 27227 52366 27229 52404
rect 27229 52366 27281 52404
rect 27281 52366 27283 52404
rect 27227 52354 27283 52366
rect 27227 52348 27229 52354
rect 27229 52348 27281 52354
rect 27281 52348 27283 52354
rect 27227 52302 27229 52324
rect 27229 52302 27281 52324
rect 27281 52302 27283 52324
rect 27227 52290 27283 52302
rect 27227 52268 27229 52290
rect 27229 52268 27281 52290
rect 27281 52268 27283 52290
rect 27227 52238 27229 52244
rect 27229 52238 27281 52244
rect 27281 52238 27283 52244
rect 27227 52226 27283 52238
rect 27227 52188 27229 52226
rect 27229 52188 27281 52226
rect 27281 52188 27283 52226
rect 28315 52686 28317 52724
rect 28317 52686 28369 52724
rect 28369 52686 28371 52724
rect 28315 52674 28371 52686
rect 28315 52668 28317 52674
rect 28317 52668 28369 52674
rect 28369 52668 28371 52674
rect 28315 52622 28317 52644
rect 28317 52622 28369 52644
rect 28369 52622 28371 52644
rect 28315 52610 28371 52622
rect 28315 52588 28317 52610
rect 28317 52588 28369 52610
rect 28369 52588 28371 52610
rect 28315 52558 28317 52564
rect 28317 52558 28369 52564
rect 28369 52558 28371 52564
rect 28315 52546 28371 52558
rect 28315 52508 28317 52546
rect 28317 52508 28369 52546
rect 28369 52508 28371 52546
rect 28315 52482 28371 52484
rect 28315 52430 28317 52482
rect 28317 52430 28369 52482
rect 28369 52430 28371 52482
rect 28315 52428 28371 52430
rect 28315 52366 28317 52404
rect 28317 52366 28369 52404
rect 28369 52366 28371 52404
rect 28315 52354 28371 52366
rect 28315 52348 28317 52354
rect 28317 52348 28369 52354
rect 28369 52348 28371 52354
rect 28315 52302 28317 52324
rect 28317 52302 28369 52324
rect 28369 52302 28371 52324
rect 28315 52290 28371 52302
rect 28315 52268 28317 52290
rect 28317 52268 28369 52290
rect 28369 52268 28371 52290
rect 28315 52238 28317 52244
rect 28317 52238 28369 52244
rect 28369 52238 28371 52244
rect 28315 52226 28371 52238
rect 28315 52188 28317 52226
rect 28317 52188 28369 52226
rect 28369 52188 28371 52226
rect 29403 52686 29405 52724
rect 29405 52686 29457 52724
rect 29457 52686 29459 52724
rect 29403 52674 29459 52686
rect 29403 52668 29405 52674
rect 29405 52668 29457 52674
rect 29457 52668 29459 52674
rect 29403 52622 29405 52644
rect 29405 52622 29457 52644
rect 29457 52622 29459 52644
rect 29403 52610 29459 52622
rect 29403 52588 29405 52610
rect 29405 52588 29457 52610
rect 29457 52588 29459 52610
rect 29403 52558 29405 52564
rect 29405 52558 29457 52564
rect 29457 52558 29459 52564
rect 29403 52546 29459 52558
rect 29403 52508 29405 52546
rect 29405 52508 29457 52546
rect 29457 52508 29459 52546
rect 29403 52482 29459 52484
rect 29403 52430 29405 52482
rect 29405 52430 29457 52482
rect 29457 52430 29459 52482
rect 29403 52428 29459 52430
rect 29403 52366 29405 52404
rect 29405 52366 29457 52404
rect 29457 52366 29459 52404
rect 29403 52354 29459 52366
rect 29403 52348 29405 52354
rect 29405 52348 29457 52354
rect 29457 52348 29459 52354
rect 29403 52302 29405 52324
rect 29405 52302 29457 52324
rect 29457 52302 29459 52324
rect 29403 52290 29459 52302
rect 29403 52268 29405 52290
rect 29405 52268 29457 52290
rect 29457 52268 29459 52290
rect 29403 52238 29405 52244
rect 29405 52238 29457 52244
rect 29457 52238 29459 52244
rect 29403 52226 29459 52238
rect 29403 52188 29405 52226
rect 29405 52188 29457 52226
rect 29457 52188 29459 52226
rect 30491 52686 30493 52724
rect 30493 52686 30545 52724
rect 30545 52686 30547 52724
rect 30491 52674 30547 52686
rect 30491 52668 30493 52674
rect 30493 52668 30545 52674
rect 30545 52668 30547 52674
rect 30491 52622 30493 52644
rect 30493 52622 30545 52644
rect 30545 52622 30547 52644
rect 30491 52610 30547 52622
rect 30491 52588 30493 52610
rect 30493 52588 30545 52610
rect 30545 52588 30547 52610
rect 30491 52558 30493 52564
rect 30493 52558 30545 52564
rect 30545 52558 30547 52564
rect 30491 52546 30547 52558
rect 30491 52508 30493 52546
rect 30493 52508 30545 52546
rect 30545 52508 30547 52546
rect 30491 52482 30547 52484
rect 30491 52430 30493 52482
rect 30493 52430 30545 52482
rect 30545 52430 30547 52482
rect 30491 52428 30547 52430
rect 30491 52366 30493 52404
rect 30493 52366 30545 52404
rect 30545 52366 30547 52404
rect 30491 52354 30547 52366
rect 30491 52348 30493 52354
rect 30493 52348 30545 52354
rect 30545 52348 30547 52354
rect 30491 52302 30493 52324
rect 30493 52302 30545 52324
rect 30545 52302 30547 52324
rect 30491 52290 30547 52302
rect 30491 52268 30493 52290
rect 30493 52268 30545 52290
rect 30545 52268 30547 52290
rect 30491 52238 30493 52244
rect 30493 52238 30545 52244
rect 30545 52238 30547 52244
rect 30491 52226 30547 52238
rect 30491 52188 30493 52226
rect 30493 52188 30545 52226
rect 30545 52188 30547 52226
rect 31579 52686 31581 52724
rect 31581 52686 31633 52724
rect 31633 52686 31635 52724
rect 31579 52674 31635 52686
rect 31579 52668 31581 52674
rect 31581 52668 31633 52674
rect 31633 52668 31635 52674
rect 31579 52622 31581 52644
rect 31581 52622 31633 52644
rect 31633 52622 31635 52644
rect 31579 52610 31635 52622
rect 31579 52588 31581 52610
rect 31581 52588 31633 52610
rect 31633 52588 31635 52610
rect 31579 52558 31581 52564
rect 31581 52558 31633 52564
rect 31633 52558 31635 52564
rect 31579 52546 31635 52558
rect 31579 52508 31581 52546
rect 31581 52508 31633 52546
rect 31633 52508 31635 52546
rect 31579 52482 31635 52484
rect 31579 52430 31581 52482
rect 31581 52430 31633 52482
rect 31633 52430 31635 52482
rect 31579 52428 31635 52430
rect 31579 52366 31581 52404
rect 31581 52366 31633 52404
rect 31633 52366 31635 52404
rect 31579 52354 31635 52366
rect 31579 52348 31581 52354
rect 31581 52348 31633 52354
rect 31633 52348 31635 52354
rect 31579 52302 31581 52324
rect 31581 52302 31633 52324
rect 31633 52302 31635 52324
rect 31579 52290 31635 52302
rect 31579 52268 31581 52290
rect 31581 52268 31633 52290
rect 31633 52268 31635 52290
rect 31579 52238 31581 52244
rect 31581 52238 31633 52244
rect 31633 52238 31635 52244
rect 31579 52226 31635 52238
rect 31579 52188 31581 52226
rect 31581 52188 31633 52226
rect 31633 52188 31635 52226
rect 17980 50683 17982 50721
rect 17982 50683 18034 50721
rect 18034 50683 18036 50721
rect 17980 50671 18036 50683
rect 17980 50665 17982 50671
rect 17982 50665 18034 50671
rect 18034 50665 18036 50671
rect 17980 50619 17982 50641
rect 17982 50619 18034 50641
rect 18034 50619 18036 50641
rect 17980 50607 18036 50619
rect 17980 50585 17982 50607
rect 17982 50585 18034 50607
rect 18034 50585 18036 50607
rect 17980 50555 17982 50561
rect 17982 50555 18034 50561
rect 18034 50555 18036 50561
rect 17980 50543 18036 50555
rect 17980 50505 17982 50543
rect 17982 50505 18034 50543
rect 18034 50505 18036 50543
rect 17980 50479 18036 50481
rect 17980 50427 17982 50479
rect 17982 50427 18034 50479
rect 18034 50427 18036 50479
rect 17980 50425 18036 50427
rect 17980 50363 17982 50401
rect 17982 50363 18034 50401
rect 18034 50363 18036 50401
rect 17980 50351 18036 50363
rect 17980 50345 17982 50351
rect 17982 50345 18034 50351
rect 18034 50345 18036 50351
rect 17980 50299 17982 50321
rect 17982 50299 18034 50321
rect 18034 50299 18036 50321
rect 17980 50287 18036 50299
rect 17980 50265 17982 50287
rect 17982 50265 18034 50287
rect 18034 50265 18036 50287
rect 17980 50235 17982 50241
rect 17982 50235 18034 50241
rect 18034 50235 18036 50241
rect 17980 50223 18036 50235
rect 17980 50185 17982 50223
rect 17982 50185 18034 50223
rect 18034 50185 18036 50223
rect 20156 50683 20158 50721
rect 20158 50683 20210 50721
rect 20210 50683 20212 50721
rect 20156 50671 20212 50683
rect 20156 50665 20158 50671
rect 20158 50665 20210 50671
rect 20210 50665 20212 50671
rect 20156 50619 20158 50641
rect 20158 50619 20210 50641
rect 20210 50619 20212 50641
rect 20156 50607 20212 50619
rect 20156 50585 20158 50607
rect 20158 50585 20210 50607
rect 20210 50585 20212 50607
rect 20156 50555 20158 50561
rect 20158 50555 20210 50561
rect 20210 50555 20212 50561
rect 20156 50543 20212 50555
rect 20156 50505 20158 50543
rect 20158 50505 20210 50543
rect 20210 50505 20212 50543
rect 20156 50479 20212 50481
rect 20156 50427 20158 50479
rect 20158 50427 20210 50479
rect 20210 50427 20212 50479
rect 20156 50425 20212 50427
rect 20156 50363 20158 50401
rect 20158 50363 20210 50401
rect 20210 50363 20212 50401
rect 20156 50351 20212 50363
rect 20156 50345 20158 50351
rect 20158 50345 20210 50351
rect 20210 50345 20212 50351
rect 20156 50299 20158 50321
rect 20158 50299 20210 50321
rect 20210 50299 20212 50321
rect 20156 50287 20212 50299
rect 20156 50265 20158 50287
rect 20158 50265 20210 50287
rect 20210 50265 20212 50287
rect 20156 50235 20158 50241
rect 20158 50235 20210 50241
rect 20210 50235 20212 50241
rect 20156 50223 20212 50235
rect 20156 50185 20158 50223
rect 20158 50185 20210 50223
rect 20210 50185 20212 50223
rect 21244 50683 21246 50721
rect 21246 50683 21298 50721
rect 21298 50683 21300 50721
rect 21244 50671 21300 50683
rect 21244 50665 21246 50671
rect 21246 50665 21298 50671
rect 21298 50665 21300 50671
rect 21244 50619 21246 50641
rect 21246 50619 21298 50641
rect 21298 50619 21300 50641
rect 21244 50607 21300 50619
rect 21244 50585 21246 50607
rect 21246 50585 21298 50607
rect 21298 50585 21300 50607
rect 21244 50555 21246 50561
rect 21246 50555 21298 50561
rect 21298 50555 21300 50561
rect 21244 50543 21300 50555
rect 21244 50505 21246 50543
rect 21246 50505 21298 50543
rect 21298 50505 21300 50543
rect 21244 50479 21300 50481
rect 21244 50427 21246 50479
rect 21246 50427 21298 50479
rect 21298 50427 21300 50479
rect 21244 50425 21300 50427
rect 21244 50363 21246 50401
rect 21246 50363 21298 50401
rect 21298 50363 21300 50401
rect 21244 50351 21300 50363
rect 21244 50345 21246 50351
rect 21246 50345 21298 50351
rect 21298 50345 21300 50351
rect 21244 50299 21246 50321
rect 21246 50299 21298 50321
rect 21298 50299 21300 50321
rect 21244 50287 21300 50299
rect 21244 50265 21246 50287
rect 21246 50265 21298 50287
rect 21298 50265 21300 50287
rect 21244 50235 21246 50241
rect 21246 50235 21298 50241
rect 21298 50235 21300 50241
rect 21244 50223 21300 50235
rect 21244 50185 21246 50223
rect 21246 50185 21298 50223
rect 21298 50185 21300 50223
rect 23420 50683 23422 50721
rect 23422 50683 23474 50721
rect 23474 50683 23476 50721
rect 23420 50671 23476 50683
rect 23420 50665 23422 50671
rect 23422 50665 23474 50671
rect 23474 50665 23476 50671
rect 23420 50619 23422 50641
rect 23422 50619 23474 50641
rect 23474 50619 23476 50641
rect 23420 50607 23476 50619
rect 23420 50585 23422 50607
rect 23422 50585 23474 50607
rect 23474 50585 23476 50607
rect 23420 50555 23422 50561
rect 23422 50555 23474 50561
rect 23474 50555 23476 50561
rect 23420 50543 23476 50555
rect 23420 50505 23422 50543
rect 23422 50505 23474 50543
rect 23474 50505 23476 50543
rect 23420 50479 23476 50481
rect 23420 50427 23422 50479
rect 23422 50427 23474 50479
rect 23474 50427 23476 50479
rect 23420 50425 23476 50427
rect 23420 50363 23422 50401
rect 23422 50363 23474 50401
rect 23474 50363 23476 50401
rect 23420 50351 23476 50363
rect 23420 50345 23422 50351
rect 23422 50345 23474 50351
rect 23474 50345 23476 50351
rect 23420 50299 23422 50321
rect 23422 50299 23474 50321
rect 23474 50299 23476 50321
rect 23420 50287 23476 50299
rect 23420 50265 23422 50287
rect 23422 50265 23474 50287
rect 23474 50265 23476 50287
rect 23420 50235 23422 50241
rect 23422 50235 23474 50241
rect 23474 50235 23476 50241
rect 23420 50223 23476 50235
rect 23420 50185 23422 50223
rect 23422 50185 23474 50223
rect 23474 50185 23476 50223
rect 24508 50683 24510 50721
rect 24510 50683 24562 50721
rect 24562 50683 24564 50721
rect 24508 50671 24564 50683
rect 24508 50665 24510 50671
rect 24510 50665 24562 50671
rect 24562 50665 24564 50671
rect 24508 50619 24510 50641
rect 24510 50619 24562 50641
rect 24562 50619 24564 50641
rect 24508 50607 24564 50619
rect 24508 50585 24510 50607
rect 24510 50585 24562 50607
rect 24562 50585 24564 50607
rect 24508 50555 24510 50561
rect 24510 50555 24562 50561
rect 24562 50555 24564 50561
rect 24508 50543 24564 50555
rect 24508 50505 24510 50543
rect 24510 50505 24562 50543
rect 24562 50505 24564 50543
rect 24508 50479 24564 50481
rect 24508 50427 24510 50479
rect 24510 50427 24562 50479
rect 24562 50427 24564 50479
rect 24508 50425 24564 50427
rect 24508 50363 24510 50401
rect 24510 50363 24562 50401
rect 24562 50363 24564 50401
rect 24508 50351 24564 50363
rect 24508 50345 24510 50351
rect 24510 50345 24562 50351
rect 24562 50345 24564 50351
rect 24508 50299 24510 50321
rect 24510 50299 24562 50321
rect 24562 50299 24564 50321
rect 24508 50287 24564 50299
rect 24508 50265 24510 50287
rect 24510 50265 24562 50287
rect 24562 50265 24564 50287
rect 24508 50235 24510 50241
rect 24510 50235 24562 50241
rect 24562 50235 24564 50241
rect 24508 50223 24564 50235
rect 24508 50185 24510 50223
rect 24510 50185 24562 50223
rect 24562 50185 24564 50223
rect 25596 50683 25598 50721
rect 25598 50683 25650 50721
rect 25650 50683 25652 50721
rect 25596 50671 25652 50683
rect 25596 50665 25598 50671
rect 25598 50665 25650 50671
rect 25650 50665 25652 50671
rect 25596 50619 25598 50641
rect 25598 50619 25650 50641
rect 25650 50619 25652 50641
rect 25596 50607 25652 50619
rect 25596 50585 25598 50607
rect 25598 50585 25650 50607
rect 25650 50585 25652 50607
rect 25596 50555 25598 50561
rect 25598 50555 25650 50561
rect 25650 50555 25652 50561
rect 25596 50543 25652 50555
rect 25596 50505 25598 50543
rect 25598 50505 25650 50543
rect 25650 50505 25652 50543
rect 25596 50479 25652 50481
rect 25596 50427 25598 50479
rect 25598 50427 25650 50479
rect 25650 50427 25652 50479
rect 25596 50425 25652 50427
rect 25596 50363 25598 50401
rect 25598 50363 25650 50401
rect 25650 50363 25652 50401
rect 25596 50351 25652 50363
rect 25596 50345 25598 50351
rect 25598 50345 25650 50351
rect 25650 50345 25652 50351
rect 25596 50299 25598 50321
rect 25598 50299 25650 50321
rect 25650 50299 25652 50321
rect 25596 50287 25652 50299
rect 25596 50265 25598 50287
rect 25598 50265 25650 50287
rect 25650 50265 25652 50287
rect 25596 50235 25598 50241
rect 25598 50235 25650 50241
rect 25650 50235 25652 50241
rect 25596 50223 25652 50235
rect 25596 50185 25598 50223
rect 25598 50185 25650 50223
rect 25650 50185 25652 50223
rect 27772 50683 27774 50721
rect 27774 50683 27826 50721
rect 27826 50683 27828 50721
rect 27772 50671 27828 50683
rect 27772 50665 27774 50671
rect 27774 50665 27826 50671
rect 27826 50665 27828 50671
rect 27772 50619 27774 50641
rect 27774 50619 27826 50641
rect 27826 50619 27828 50641
rect 27772 50607 27828 50619
rect 27772 50585 27774 50607
rect 27774 50585 27826 50607
rect 27826 50585 27828 50607
rect 27772 50555 27774 50561
rect 27774 50555 27826 50561
rect 27826 50555 27828 50561
rect 27772 50543 27828 50555
rect 27772 50505 27774 50543
rect 27774 50505 27826 50543
rect 27826 50505 27828 50543
rect 27772 50479 27828 50481
rect 27772 50427 27774 50479
rect 27774 50427 27826 50479
rect 27826 50427 27828 50479
rect 27772 50425 27828 50427
rect 27772 50363 27774 50401
rect 27774 50363 27826 50401
rect 27826 50363 27828 50401
rect 27772 50351 27828 50363
rect 27772 50345 27774 50351
rect 27774 50345 27826 50351
rect 27826 50345 27828 50351
rect 27772 50299 27774 50321
rect 27774 50299 27826 50321
rect 27826 50299 27828 50321
rect 27772 50287 27828 50299
rect 27772 50265 27774 50287
rect 27774 50265 27826 50287
rect 27826 50265 27828 50287
rect 27772 50235 27774 50241
rect 27774 50235 27826 50241
rect 27826 50235 27828 50241
rect 27772 50223 27828 50235
rect 27772 50185 27774 50223
rect 27774 50185 27826 50223
rect 27826 50185 27828 50223
rect 28860 50683 28862 50721
rect 28862 50683 28914 50721
rect 28914 50683 28916 50721
rect 28860 50671 28916 50683
rect 28860 50665 28862 50671
rect 28862 50665 28914 50671
rect 28914 50665 28916 50671
rect 28860 50619 28862 50641
rect 28862 50619 28914 50641
rect 28914 50619 28916 50641
rect 28860 50607 28916 50619
rect 28860 50585 28862 50607
rect 28862 50585 28914 50607
rect 28914 50585 28916 50607
rect 28860 50555 28862 50561
rect 28862 50555 28914 50561
rect 28914 50555 28916 50561
rect 28860 50543 28916 50555
rect 28860 50505 28862 50543
rect 28862 50505 28914 50543
rect 28914 50505 28916 50543
rect 28860 50479 28916 50481
rect 28860 50427 28862 50479
rect 28862 50427 28914 50479
rect 28914 50427 28916 50479
rect 28860 50425 28916 50427
rect 28860 50363 28862 50401
rect 28862 50363 28914 50401
rect 28914 50363 28916 50401
rect 28860 50351 28916 50363
rect 28860 50345 28862 50351
rect 28862 50345 28914 50351
rect 28914 50345 28916 50351
rect 28860 50299 28862 50321
rect 28862 50299 28914 50321
rect 28914 50299 28916 50321
rect 28860 50287 28916 50299
rect 28860 50265 28862 50287
rect 28862 50265 28914 50287
rect 28914 50265 28916 50287
rect 28860 50235 28862 50241
rect 28862 50235 28914 50241
rect 28914 50235 28916 50241
rect 28860 50223 28916 50235
rect 28860 50185 28862 50223
rect 28862 50185 28914 50223
rect 28914 50185 28916 50223
rect 31036 50683 31038 50721
rect 31038 50683 31090 50721
rect 31090 50683 31092 50721
rect 31036 50671 31092 50683
rect 31036 50665 31038 50671
rect 31038 50665 31090 50671
rect 31090 50665 31092 50671
rect 31036 50619 31038 50641
rect 31038 50619 31090 50641
rect 31090 50619 31092 50641
rect 31036 50607 31092 50619
rect 31036 50585 31038 50607
rect 31038 50585 31090 50607
rect 31090 50585 31092 50607
rect 31036 50555 31038 50561
rect 31038 50555 31090 50561
rect 31090 50555 31092 50561
rect 31036 50543 31092 50555
rect 31036 50505 31038 50543
rect 31038 50505 31090 50543
rect 31090 50505 31092 50543
rect 31036 50479 31092 50481
rect 31036 50427 31038 50479
rect 31038 50427 31090 50479
rect 31090 50427 31092 50479
rect 31036 50425 31092 50427
rect 31036 50363 31038 50401
rect 31038 50363 31090 50401
rect 31090 50363 31092 50401
rect 31036 50351 31092 50363
rect 31036 50345 31038 50351
rect 31038 50345 31090 50351
rect 31090 50345 31092 50351
rect 31036 50299 31038 50321
rect 31038 50299 31090 50321
rect 31090 50299 31092 50321
rect 31036 50287 31092 50299
rect 31036 50265 31038 50287
rect 31038 50265 31090 50287
rect 31090 50265 31092 50287
rect 31036 50235 31038 50241
rect 31038 50235 31090 50241
rect 31090 50235 31092 50241
rect 31036 50223 31092 50235
rect 31036 50185 31038 50223
rect 31038 50185 31090 50223
rect 31090 50185 31092 50223
rect 17435 48686 17437 48724
rect 17437 48686 17489 48724
rect 17489 48686 17491 48724
rect 17435 48674 17491 48686
rect 17435 48668 17437 48674
rect 17437 48668 17489 48674
rect 17489 48668 17491 48674
rect 17435 48622 17437 48644
rect 17437 48622 17489 48644
rect 17489 48622 17491 48644
rect 17435 48610 17491 48622
rect 17435 48588 17437 48610
rect 17437 48588 17489 48610
rect 17489 48588 17491 48610
rect 17435 48558 17437 48564
rect 17437 48558 17489 48564
rect 17489 48558 17491 48564
rect 17435 48546 17491 48558
rect 17435 48508 17437 48546
rect 17437 48508 17489 48546
rect 17489 48508 17491 48546
rect 17435 48482 17491 48484
rect 17435 48430 17437 48482
rect 17437 48430 17489 48482
rect 17489 48430 17491 48482
rect 17435 48428 17491 48430
rect 17435 48366 17437 48404
rect 17437 48366 17489 48404
rect 17489 48366 17491 48404
rect 17435 48354 17491 48366
rect 17435 48348 17437 48354
rect 17437 48348 17489 48354
rect 17489 48348 17491 48354
rect 17435 48302 17437 48324
rect 17437 48302 17489 48324
rect 17489 48302 17491 48324
rect 17435 48290 17491 48302
rect 17435 48268 17437 48290
rect 17437 48268 17489 48290
rect 17489 48268 17491 48290
rect 17435 48238 17437 48244
rect 17437 48238 17489 48244
rect 17489 48238 17491 48244
rect 17435 48226 17491 48238
rect 17435 48188 17437 48226
rect 17437 48188 17489 48226
rect 17489 48188 17491 48226
rect 18523 48686 18525 48724
rect 18525 48686 18577 48724
rect 18577 48686 18579 48724
rect 18523 48674 18579 48686
rect 18523 48668 18525 48674
rect 18525 48668 18577 48674
rect 18577 48668 18579 48674
rect 18523 48622 18525 48644
rect 18525 48622 18577 48644
rect 18577 48622 18579 48644
rect 18523 48610 18579 48622
rect 18523 48588 18525 48610
rect 18525 48588 18577 48610
rect 18577 48588 18579 48610
rect 18523 48558 18525 48564
rect 18525 48558 18577 48564
rect 18577 48558 18579 48564
rect 18523 48546 18579 48558
rect 18523 48508 18525 48546
rect 18525 48508 18577 48546
rect 18577 48508 18579 48546
rect 18523 48482 18579 48484
rect 18523 48430 18525 48482
rect 18525 48430 18577 48482
rect 18577 48430 18579 48482
rect 18523 48428 18579 48430
rect 18523 48366 18525 48404
rect 18525 48366 18577 48404
rect 18577 48366 18579 48404
rect 18523 48354 18579 48366
rect 18523 48348 18525 48354
rect 18525 48348 18577 48354
rect 18577 48348 18579 48354
rect 18523 48302 18525 48324
rect 18525 48302 18577 48324
rect 18577 48302 18579 48324
rect 18523 48290 18579 48302
rect 18523 48268 18525 48290
rect 18525 48268 18577 48290
rect 18577 48268 18579 48290
rect 18523 48238 18525 48244
rect 18525 48238 18577 48244
rect 18577 48238 18579 48244
rect 18523 48226 18579 48238
rect 18523 48188 18525 48226
rect 18525 48188 18577 48226
rect 18577 48188 18579 48226
rect 19611 48686 19613 48724
rect 19613 48686 19665 48724
rect 19665 48686 19667 48724
rect 19611 48674 19667 48686
rect 19611 48668 19613 48674
rect 19613 48668 19665 48674
rect 19665 48668 19667 48674
rect 19611 48622 19613 48644
rect 19613 48622 19665 48644
rect 19665 48622 19667 48644
rect 19611 48610 19667 48622
rect 19611 48588 19613 48610
rect 19613 48588 19665 48610
rect 19665 48588 19667 48610
rect 19611 48558 19613 48564
rect 19613 48558 19665 48564
rect 19665 48558 19667 48564
rect 19611 48546 19667 48558
rect 19611 48508 19613 48546
rect 19613 48508 19665 48546
rect 19665 48508 19667 48546
rect 19611 48482 19667 48484
rect 19611 48430 19613 48482
rect 19613 48430 19665 48482
rect 19665 48430 19667 48482
rect 19611 48428 19667 48430
rect 19611 48366 19613 48404
rect 19613 48366 19665 48404
rect 19665 48366 19667 48404
rect 19611 48354 19667 48366
rect 19611 48348 19613 48354
rect 19613 48348 19665 48354
rect 19665 48348 19667 48354
rect 19611 48302 19613 48324
rect 19613 48302 19665 48324
rect 19665 48302 19667 48324
rect 19611 48290 19667 48302
rect 19611 48268 19613 48290
rect 19613 48268 19665 48290
rect 19665 48268 19667 48290
rect 19611 48238 19613 48244
rect 19613 48238 19665 48244
rect 19665 48238 19667 48244
rect 19611 48226 19667 48238
rect 19611 48188 19613 48226
rect 19613 48188 19665 48226
rect 19665 48188 19667 48226
rect 20699 48686 20701 48724
rect 20701 48686 20753 48724
rect 20753 48686 20755 48724
rect 20699 48674 20755 48686
rect 20699 48668 20701 48674
rect 20701 48668 20753 48674
rect 20753 48668 20755 48674
rect 20699 48622 20701 48644
rect 20701 48622 20753 48644
rect 20753 48622 20755 48644
rect 20699 48610 20755 48622
rect 20699 48588 20701 48610
rect 20701 48588 20753 48610
rect 20753 48588 20755 48610
rect 20699 48558 20701 48564
rect 20701 48558 20753 48564
rect 20753 48558 20755 48564
rect 20699 48546 20755 48558
rect 20699 48508 20701 48546
rect 20701 48508 20753 48546
rect 20753 48508 20755 48546
rect 20699 48482 20755 48484
rect 20699 48430 20701 48482
rect 20701 48430 20753 48482
rect 20753 48430 20755 48482
rect 20699 48428 20755 48430
rect 20699 48366 20701 48404
rect 20701 48366 20753 48404
rect 20753 48366 20755 48404
rect 20699 48354 20755 48366
rect 20699 48348 20701 48354
rect 20701 48348 20753 48354
rect 20753 48348 20755 48354
rect 20699 48302 20701 48324
rect 20701 48302 20753 48324
rect 20753 48302 20755 48324
rect 20699 48290 20755 48302
rect 20699 48268 20701 48290
rect 20701 48268 20753 48290
rect 20753 48268 20755 48290
rect 20699 48238 20701 48244
rect 20701 48238 20753 48244
rect 20753 48238 20755 48244
rect 20699 48226 20755 48238
rect 20699 48188 20701 48226
rect 20701 48188 20753 48226
rect 20753 48188 20755 48226
rect 21787 48686 21789 48724
rect 21789 48686 21841 48724
rect 21841 48686 21843 48724
rect 21787 48674 21843 48686
rect 21787 48668 21789 48674
rect 21789 48668 21841 48674
rect 21841 48668 21843 48674
rect 21787 48622 21789 48644
rect 21789 48622 21841 48644
rect 21841 48622 21843 48644
rect 21787 48610 21843 48622
rect 21787 48588 21789 48610
rect 21789 48588 21841 48610
rect 21841 48588 21843 48610
rect 21787 48558 21789 48564
rect 21789 48558 21841 48564
rect 21841 48558 21843 48564
rect 21787 48546 21843 48558
rect 21787 48508 21789 48546
rect 21789 48508 21841 48546
rect 21841 48508 21843 48546
rect 21787 48482 21843 48484
rect 21787 48430 21789 48482
rect 21789 48430 21841 48482
rect 21841 48430 21843 48482
rect 21787 48428 21843 48430
rect 21787 48366 21789 48404
rect 21789 48366 21841 48404
rect 21841 48366 21843 48404
rect 21787 48354 21843 48366
rect 21787 48348 21789 48354
rect 21789 48348 21841 48354
rect 21841 48348 21843 48354
rect 21787 48302 21789 48324
rect 21789 48302 21841 48324
rect 21841 48302 21843 48324
rect 21787 48290 21843 48302
rect 21787 48268 21789 48290
rect 21789 48268 21841 48290
rect 21841 48268 21843 48290
rect 21787 48238 21789 48244
rect 21789 48238 21841 48244
rect 21841 48238 21843 48244
rect 21787 48226 21843 48238
rect 21787 48188 21789 48226
rect 21789 48188 21841 48226
rect 21841 48188 21843 48226
rect 22875 48686 22877 48724
rect 22877 48686 22929 48724
rect 22929 48686 22931 48724
rect 22875 48674 22931 48686
rect 22875 48668 22877 48674
rect 22877 48668 22929 48674
rect 22929 48668 22931 48674
rect 22875 48622 22877 48644
rect 22877 48622 22929 48644
rect 22929 48622 22931 48644
rect 22875 48610 22931 48622
rect 22875 48588 22877 48610
rect 22877 48588 22929 48610
rect 22929 48588 22931 48610
rect 22875 48558 22877 48564
rect 22877 48558 22929 48564
rect 22929 48558 22931 48564
rect 22875 48546 22931 48558
rect 22875 48508 22877 48546
rect 22877 48508 22929 48546
rect 22929 48508 22931 48546
rect 22875 48482 22931 48484
rect 22875 48430 22877 48482
rect 22877 48430 22929 48482
rect 22929 48430 22931 48482
rect 22875 48428 22931 48430
rect 22875 48366 22877 48404
rect 22877 48366 22929 48404
rect 22929 48366 22931 48404
rect 22875 48354 22931 48366
rect 22875 48348 22877 48354
rect 22877 48348 22929 48354
rect 22929 48348 22931 48354
rect 22875 48302 22877 48324
rect 22877 48302 22929 48324
rect 22929 48302 22931 48324
rect 22875 48290 22931 48302
rect 22875 48268 22877 48290
rect 22877 48268 22929 48290
rect 22929 48268 22931 48290
rect 22875 48238 22877 48244
rect 22877 48238 22929 48244
rect 22929 48238 22931 48244
rect 22875 48226 22931 48238
rect 22875 48188 22877 48226
rect 22877 48188 22929 48226
rect 22929 48188 22931 48226
rect 23963 48686 23965 48724
rect 23965 48686 24017 48724
rect 24017 48686 24019 48724
rect 23963 48674 24019 48686
rect 23963 48668 23965 48674
rect 23965 48668 24017 48674
rect 24017 48668 24019 48674
rect 23963 48622 23965 48644
rect 23965 48622 24017 48644
rect 24017 48622 24019 48644
rect 23963 48610 24019 48622
rect 23963 48588 23965 48610
rect 23965 48588 24017 48610
rect 24017 48588 24019 48610
rect 23963 48558 23965 48564
rect 23965 48558 24017 48564
rect 24017 48558 24019 48564
rect 23963 48546 24019 48558
rect 23963 48508 23965 48546
rect 23965 48508 24017 48546
rect 24017 48508 24019 48546
rect 23963 48482 24019 48484
rect 23963 48430 23965 48482
rect 23965 48430 24017 48482
rect 24017 48430 24019 48482
rect 23963 48428 24019 48430
rect 23963 48366 23965 48404
rect 23965 48366 24017 48404
rect 24017 48366 24019 48404
rect 23963 48354 24019 48366
rect 23963 48348 23965 48354
rect 23965 48348 24017 48354
rect 24017 48348 24019 48354
rect 23963 48302 23965 48324
rect 23965 48302 24017 48324
rect 24017 48302 24019 48324
rect 23963 48290 24019 48302
rect 23963 48268 23965 48290
rect 23965 48268 24017 48290
rect 24017 48268 24019 48290
rect 23963 48238 23965 48244
rect 23965 48238 24017 48244
rect 24017 48238 24019 48244
rect 23963 48226 24019 48238
rect 23963 48188 23965 48226
rect 23965 48188 24017 48226
rect 24017 48188 24019 48226
rect 29403 48686 29405 48724
rect 29405 48686 29457 48724
rect 29457 48686 29459 48724
rect 29403 48674 29459 48686
rect 29403 48668 29405 48674
rect 29405 48668 29457 48674
rect 29457 48668 29459 48674
rect 29403 48622 29405 48644
rect 29405 48622 29457 48644
rect 29457 48622 29459 48644
rect 29403 48610 29459 48622
rect 29403 48588 29405 48610
rect 29405 48588 29457 48610
rect 29457 48588 29459 48610
rect 29403 48558 29405 48564
rect 29405 48558 29457 48564
rect 29457 48558 29459 48564
rect 29403 48546 29459 48558
rect 29403 48508 29405 48546
rect 29405 48508 29457 48546
rect 29457 48508 29459 48546
rect 29403 48482 29459 48484
rect 29403 48430 29405 48482
rect 29405 48430 29457 48482
rect 29457 48430 29459 48482
rect 29403 48428 29459 48430
rect 29403 48366 29405 48404
rect 29405 48366 29457 48404
rect 29457 48366 29459 48404
rect 29403 48354 29459 48366
rect 29403 48348 29405 48354
rect 29405 48348 29457 48354
rect 29457 48348 29459 48354
rect 29403 48302 29405 48324
rect 29405 48302 29457 48324
rect 29457 48302 29459 48324
rect 29403 48290 29459 48302
rect 29403 48268 29405 48290
rect 29405 48268 29457 48290
rect 29457 48268 29459 48290
rect 29403 48238 29405 48244
rect 29405 48238 29457 48244
rect 29457 48238 29459 48244
rect 29403 48226 29459 48238
rect 29403 48188 29405 48226
rect 29405 48188 29457 48226
rect 29457 48188 29459 48226
rect 30491 48686 30493 48724
rect 30493 48686 30545 48724
rect 30545 48686 30547 48724
rect 30491 48674 30547 48686
rect 30491 48668 30493 48674
rect 30493 48668 30545 48674
rect 30545 48668 30547 48674
rect 30491 48622 30493 48644
rect 30493 48622 30545 48644
rect 30545 48622 30547 48644
rect 30491 48610 30547 48622
rect 30491 48588 30493 48610
rect 30493 48588 30545 48610
rect 30545 48588 30547 48610
rect 30491 48558 30493 48564
rect 30493 48558 30545 48564
rect 30545 48558 30547 48564
rect 30491 48546 30547 48558
rect 30491 48508 30493 48546
rect 30493 48508 30545 48546
rect 30545 48508 30547 48546
rect 30491 48482 30547 48484
rect 30491 48430 30493 48482
rect 30493 48430 30545 48482
rect 30545 48430 30547 48482
rect 30491 48428 30547 48430
rect 30491 48366 30493 48404
rect 30493 48366 30545 48404
rect 30545 48366 30547 48404
rect 30491 48354 30547 48366
rect 30491 48348 30493 48354
rect 30493 48348 30545 48354
rect 30545 48348 30547 48354
rect 30491 48302 30493 48324
rect 30493 48302 30545 48324
rect 30545 48302 30547 48324
rect 30491 48290 30547 48302
rect 30491 48268 30493 48290
rect 30493 48268 30545 48290
rect 30545 48268 30547 48290
rect 30491 48238 30493 48244
rect 30493 48238 30545 48244
rect 30545 48238 30547 48244
rect 30491 48226 30547 48238
rect 30491 48188 30493 48226
rect 30493 48188 30545 48226
rect 30545 48188 30547 48226
rect 31579 48686 31581 48724
rect 31581 48686 31633 48724
rect 31633 48686 31635 48724
rect 31579 48674 31635 48686
rect 31579 48668 31581 48674
rect 31581 48668 31633 48674
rect 31633 48668 31635 48674
rect 31579 48622 31581 48644
rect 31581 48622 31633 48644
rect 31633 48622 31635 48644
rect 31579 48610 31635 48622
rect 31579 48588 31581 48610
rect 31581 48588 31633 48610
rect 31633 48588 31635 48610
rect 31579 48558 31581 48564
rect 31581 48558 31633 48564
rect 31633 48558 31635 48564
rect 31579 48546 31635 48558
rect 31579 48508 31581 48546
rect 31581 48508 31633 48546
rect 31633 48508 31635 48546
rect 31579 48482 31635 48484
rect 31579 48430 31581 48482
rect 31581 48430 31633 48482
rect 31633 48430 31635 48482
rect 31579 48428 31635 48430
rect 31579 48366 31581 48404
rect 31581 48366 31633 48404
rect 31633 48366 31635 48404
rect 31579 48354 31635 48366
rect 31579 48348 31581 48354
rect 31581 48348 31633 48354
rect 31633 48348 31635 48354
rect 31579 48302 31581 48324
rect 31581 48302 31633 48324
rect 31633 48302 31635 48324
rect 31579 48290 31635 48302
rect 31579 48268 31581 48290
rect 31581 48268 31633 48290
rect 31633 48268 31635 48290
rect 31579 48238 31581 48244
rect 31581 48238 31633 48244
rect 31633 48238 31635 48244
rect 31579 48226 31635 48238
rect 31579 48188 31581 48226
rect 31581 48188 31633 48226
rect 31633 48188 31635 48226
rect 10216 47638 10512 47640
rect 17980 46683 17982 46721
rect 17982 46683 18034 46721
rect 18034 46683 18036 46721
rect 17980 46671 18036 46683
rect 17980 46665 17982 46671
rect 17982 46665 18034 46671
rect 18034 46665 18036 46671
rect 17980 46619 17982 46641
rect 17982 46619 18034 46641
rect 18034 46619 18036 46641
rect 17980 46607 18036 46619
rect 17980 46585 17982 46607
rect 17982 46585 18034 46607
rect 18034 46585 18036 46607
rect 17980 46555 17982 46561
rect 17982 46555 18034 46561
rect 18034 46555 18036 46561
rect 17980 46543 18036 46555
rect 17980 46505 17982 46543
rect 17982 46505 18034 46543
rect 18034 46505 18036 46543
rect 17980 46479 18036 46481
rect 17980 46427 17982 46479
rect 17982 46427 18034 46479
rect 18034 46427 18036 46479
rect 17980 46425 18036 46427
rect 17980 46363 17982 46401
rect 17982 46363 18034 46401
rect 18034 46363 18036 46401
rect 17980 46351 18036 46363
rect 17980 46345 17982 46351
rect 17982 46345 18034 46351
rect 18034 46345 18036 46351
rect -5891 39858 -5755 46234
rect 17980 46299 17982 46321
rect 17982 46299 18034 46321
rect 18034 46299 18036 46321
rect 17980 46287 18036 46299
rect 17980 46265 17982 46287
rect 17982 46265 18034 46287
rect 18034 46265 18036 46287
rect 17980 46235 17982 46241
rect 17982 46235 18034 46241
rect 18034 46235 18036 46241
rect 17980 46223 18036 46235
rect 17980 46185 17982 46223
rect 17982 46185 18034 46223
rect 18034 46185 18036 46223
rect 19068 46683 19070 46721
rect 19070 46683 19122 46721
rect 19122 46683 19124 46721
rect 19068 46671 19124 46683
rect 19068 46665 19070 46671
rect 19070 46665 19122 46671
rect 19122 46665 19124 46671
rect 19068 46619 19070 46641
rect 19070 46619 19122 46641
rect 19122 46619 19124 46641
rect 19068 46607 19124 46619
rect 19068 46585 19070 46607
rect 19070 46585 19122 46607
rect 19122 46585 19124 46607
rect 19068 46555 19070 46561
rect 19070 46555 19122 46561
rect 19122 46555 19124 46561
rect 19068 46543 19124 46555
rect 19068 46505 19070 46543
rect 19070 46505 19122 46543
rect 19122 46505 19124 46543
rect 19068 46479 19124 46481
rect 19068 46427 19070 46479
rect 19070 46427 19122 46479
rect 19122 46427 19124 46479
rect 19068 46425 19124 46427
rect 19068 46363 19070 46401
rect 19070 46363 19122 46401
rect 19122 46363 19124 46401
rect 19068 46351 19124 46363
rect 19068 46345 19070 46351
rect 19070 46345 19122 46351
rect 19122 46345 19124 46351
rect 19068 46299 19070 46321
rect 19070 46299 19122 46321
rect 19122 46299 19124 46321
rect 19068 46287 19124 46299
rect 19068 46265 19070 46287
rect 19070 46265 19122 46287
rect 19122 46265 19124 46287
rect 19068 46235 19070 46241
rect 19070 46235 19122 46241
rect 19122 46235 19124 46241
rect 19068 46223 19124 46235
rect 19068 46185 19070 46223
rect 19070 46185 19122 46223
rect 19122 46185 19124 46223
rect 20156 46683 20158 46721
rect 20158 46683 20210 46721
rect 20210 46683 20212 46721
rect 20156 46671 20212 46683
rect 20156 46665 20158 46671
rect 20158 46665 20210 46671
rect 20210 46665 20212 46671
rect 20156 46619 20158 46641
rect 20158 46619 20210 46641
rect 20210 46619 20212 46641
rect 20156 46607 20212 46619
rect 20156 46585 20158 46607
rect 20158 46585 20210 46607
rect 20210 46585 20212 46607
rect 20156 46555 20158 46561
rect 20158 46555 20210 46561
rect 20210 46555 20212 46561
rect 20156 46543 20212 46555
rect 20156 46505 20158 46543
rect 20158 46505 20210 46543
rect 20210 46505 20212 46543
rect 20156 46479 20212 46481
rect 20156 46427 20158 46479
rect 20158 46427 20210 46479
rect 20210 46427 20212 46479
rect 20156 46425 20212 46427
rect 20156 46363 20158 46401
rect 20158 46363 20210 46401
rect 20210 46363 20212 46401
rect 20156 46351 20212 46363
rect 20156 46345 20158 46351
rect 20158 46345 20210 46351
rect 20210 46345 20212 46351
rect 20156 46299 20158 46321
rect 20158 46299 20210 46321
rect 20210 46299 20212 46321
rect 20156 46287 20212 46299
rect 20156 46265 20158 46287
rect 20158 46265 20210 46287
rect 20210 46265 20212 46287
rect 20156 46235 20158 46241
rect 20158 46235 20210 46241
rect 20210 46235 20212 46241
rect 20156 46223 20212 46235
rect 20156 46185 20158 46223
rect 20158 46185 20210 46223
rect 20210 46185 20212 46223
rect 21244 46683 21246 46721
rect 21246 46683 21298 46721
rect 21298 46683 21300 46721
rect 21244 46671 21300 46683
rect 21244 46665 21246 46671
rect 21246 46665 21298 46671
rect 21298 46665 21300 46671
rect 21244 46619 21246 46641
rect 21246 46619 21298 46641
rect 21298 46619 21300 46641
rect 21244 46607 21300 46619
rect 21244 46585 21246 46607
rect 21246 46585 21298 46607
rect 21298 46585 21300 46607
rect 21244 46555 21246 46561
rect 21246 46555 21298 46561
rect 21298 46555 21300 46561
rect 21244 46543 21300 46555
rect 21244 46505 21246 46543
rect 21246 46505 21298 46543
rect 21298 46505 21300 46543
rect 21244 46479 21300 46481
rect 21244 46427 21246 46479
rect 21246 46427 21298 46479
rect 21298 46427 21300 46479
rect 21244 46425 21300 46427
rect 21244 46363 21246 46401
rect 21246 46363 21298 46401
rect 21298 46363 21300 46401
rect 21244 46351 21300 46363
rect 21244 46345 21246 46351
rect 21246 46345 21298 46351
rect 21298 46345 21300 46351
rect 21244 46299 21246 46321
rect 21246 46299 21298 46321
rect 21298 46299 21300 46321
rect 21244 46287 21300 46299
rect 21244 46265 21246 46287
rect 21246 46265 21298 46287
rect 21298 46265 21300 46287
rect 21244 46235 21246 46241
rect 21246 46235 21298 46241
rect 21298 46235 21300 46241
rect 21244 46223 21300 46235
rect 21244 46185 21246 46223
rect 21246 46185 21298 46223
rect 21298 46185 21300 46223
rect 22332 46683 22334 46721
rect 22334 46683 22386 46721
rect 22386 46683 22388 46721
rect 22332 46671 22388 46683
rect 22332 46665 22334 46671
rect 22334 46665 22386 46671
rect 22386 46665 22388 46671
rect 22332 46619 22334 46641
rect 22334 46619 22386 46641
rect 22386 46619 22388 46641
rect 22332 46607 22388 46619
rect 22332 46585 22334 46607
rect 22334 46585 22386 46607
rect 22386 46585 22388 46607
rect 22332 46555 22334 46561
rect 22334 46555 22386 46561
rect 22386 46555 22388 46561
rect 22332 46543 22388 46555
rect 22332 46505 22334 46543
rect 22334 46505 22386 46543
rect 22386 46505 22388 46543
rect 22332 46479 22388 46481
rect 22332 46427 22334 46479
rect 22334 46427 22386 46479
rect 22386 46427 22388 46479
rect 22332 46425 22388 46427
rect 22332 46363 22334 46401
rect 22334 46363 22386 46401
rect 22386 46363 22388 46401
rect 22332 46351 22388 46363
rect 22332 46345 22334 46351
rect 22334 46345 22386 46351
rect 22386 46345 22388 46351
rect 22332 46299 22334 46321
rect 22334 46299 22386 46321
rect 22386 46299 22388 46321
rect 22332 46287 22388 46299
rect 22332 46265 22334 46287
rect 22334 46265 22386 46287
rect 22386 46265 22388 46287
rect 22332 46235 22334 46241
rect 22334 46235 22386 46241
rect 22386 46235 22388 46241
rect 22332 46223 22388 46235
rect 22332 46185 22334 46223
rect 22334 46185 22386 46223
rect 22386 46185 22388 46223
rect 24508 46683 24510 46721
rect 24510 46683 24562 46721
rect 24562 46683 24564 46721
rect 24508 46671 24564 46683
rect 24508 46665 24510 46671
rect 24510 46665 24562 46671
rect 24562 46665 24564 46671
rect 24508 46619 24510 46641
rect 24510 46619 24562 46641
rect 24562 46619 24564 46641
rect 24508 46607 24564 46619
rect 24508 46585 24510 46607
rect 24510 46585 24562 46607
rect 24562 46585 24564 46607
rect 24508 46555 24510 46561
rect 24510 46555 24562 46561
rect 24562 46555 24564 46561
rect 24508 46543 24564 46555
rect 24508 46505 24510 46543
rect 24510 46505 24562 46543
rect 24562 46505 24564 46543
rect 24508 46479 24564 46481
rect 24508 46427 24510 46479
rect 24510 46427 24562 46479
rect 24562 46427 24564 46479
rect 24508 46425 24564 46427
rect 24508 46363 24510 46401
rect 24510 46363 24562 46401
rect 24562 46363 24564 46401
rect 24508 46351 24564 46363
rect 24508 46345 24510 46351
rect 24510 46345 24562 46351
rect 24562 46345 24564 46351
rect 24508 46299 24510 46321
rect 24510 46299 24562 46321
rect 24562 46299 24564 46321
rect 24508 46287 24564 46299
rect 24508 46265 24510 46287
rect 24510 46265 24562 46287
rect 24562 46265 24564 46287
rect 24508 46235 24510 46241
rect 24510 46235 24562 46241
rect 24562 46235 24564 46241
rect 24508 46223 24564 46235
rect 24508 46185 24510 46223
rect 24510 46185 24562 46223
rect 24562 46185 24564 46223
rect 25596 46683 25598 46721
rect 25598 46683 25650 46721
rect 25650 46683 25652 46721
rect 25596 46671 25652 46683
rect 25596 46665 25598 46671
rect 25598 46665 25650 46671
rect 25650 46665 25652 46671
rect 25596 46619 25598 46641
rect 25598 46619 25650 46641
rect 25650 46619 25652 46641
rect 25596 46607 25652 46619
rect 25596 46585 25598 46607
rect 25598 46585 25650 46607
rect 25650 46585 25652 46607
rect 25596 46555 25598 46561
rect 25598 46555 25650 46561
rect 25650 46555 25652 46561
rect 25596 46543 25652 46555
rect 25596 46505 25598 46543
rect 25598 46505 25650 46543
rect 25650 46505 25652 46543
rect 25596 46479 25652 46481
rect 25596 46427 25598 46479
rect 25598 46427 25650 46479
rect 25650 46427 25652 46479
rect 25596 46425 25652 46427
rect 25596 46363 25598 46401
rect 25598 46363 25650 46401
rect 25650 46363 25652 46401
rect 25596 46351 25652 46363
rect 25596 46345 25598 46351
rect 25598 46345 25650 46351
rect 25650 46345 25652 46351
rect 25596 46299 25598 46321
rect 25598 46299 25650 46321
rect 25650 46299 25652 46321
rect 25596 46287 25652 46299
rect 25596 46265 25598 46287
rect 25598 46265 25650 46287
rect 25650 46265 25652 46287
rect 25596 46235 25598 46241
rect 25598 46235 25650 46241
rect 25650 46235 25652 46241
rect 25596 46223 25652 46235
rect 25596 46185 25598 46223
rect 25598 46185 25650 46223
rect 25650 46185 25652 46223
rect 26684 46683 26686 46721
rect 26686 46683 26738 46721
rect 26738 46683 26740 46721
rect 26684 46671 26740 46683
rect 26684 46665 26686 46671
rect 26686 46665 26738 46671
rect 26738 46665 26740 46671
rect 26684 46619 26686 46641
rect 26686 46619 26738 46641
rect 26738 46619 26740 46641
rect 26684 46607 26740 46619
rect 26684 46585 26686 46607
rect 26686 46585 26738 46607
rect 26738 46585 26740 46607
rect 26684 46555 26686 46561
rect 26686 46555 26738 46561
rect 26738 46555 26740 46561
rect 26684 46543 26740 46555
rect 26684 46505 26686 46543
rect 26686 46505 26738 46543
rect 26738 46505 26740 46543
rect 26684 46479 26740 46481
rect 26684 46427 26686 46479
rect 26686 46427 26738 46479
rect 26738 46427 26740 46479
rect 26684 46425 26740 46427
rect 26684 46363 26686 46401
rect 26686 46363 26738 46401
rect 26738 46363 26740 46401
rect 26684 46351 26740 46363
rect 26684 46345 26686 46351
rect 26686 46345 26738 46351
rect 26738 46345 26740 46351
rect 26684 46299 26686 46321
rect 26686 46299 26738 46321
rect 26738 46299 26740 46321
rect 26684 46287 26740 46299
rect 26684 46265 26686 46287
rect 26686 46265 26738 46287
rect 26738 46265 26740 46287
rect 26684 46235 26686 46241
rect 26686 46235 26738 46241
rect 26738 46235 26740 46241
rect 26684 46223 26740 46235
rect 26684 46185 26686 46223
rect 26686 46185 26738 46223
rect 26738 46185 26740 46223
rect 27772 46683 27774 46721
rect 27774 46683 27826 46721
rect 27826 46683 27828 46721
rect 27772 46671 27828 46683
rect 27772 46665 27774 46671
rect 27774 46665 27826 46671
rect 27826 46665 27828 46671
rect 27772 46619 27774 46641
rect 27774 46619 27826 46641
rect 27826 46619 27828 46641
rect 27772 46607 27828 46619
rect 27772 46585 27774 46607
rect 27774 46585 27826 46607
rect 27826 46585 27828 46607
rect 27772 46555 27774 46561
rect 27774 46555 27826 46561
rect 27826 46555 27828 46561
rect 27772 46543 27828 46555
rect 27772 46505 27774 46543
rect 27774 46505 27826 46543
rect 27826 46505 27828 46543
rect 27772 46479 27828 46481
rect 27772 46427 27774 46479
rect 27774 46427 27826 46479
rect 27826 46427 27828 46479
rect 27772 46425 27828 46427
rect 27772 46363 27774 46401
rect 27774 46363 27826 46401
rect 27826 46363 27828 46401
rect 27772 46351 27828 46363
rect 27772 46345 27774 46351
rect 27774 46345 27826 46351
rect 27826 46345 27828 46351
rect 27772 46299 27774 46321
rect 27774 46299 27826 46321
rect 27826 46299 27828 46321
rect 27772 46287 27828 46299
rect 27772 46265 27774 46287
rect 27774 46265 27826 46287
rect 27826 46265 27828 46287
rect 27772 46235 27774 46241
rect 27774 46235 27826 46241
rect 27826 46235 27828 46241
rect 27772 46223 27828 46235
rect 27772 46185 27774 46223
rect 27774 46185 27826 46223
rect 27826 46185 27828 46223
rect 28860 46683 28862 46721
rect 28862 46683 28914 46721
rect 28914 46683 28916 46721
rect 28860 46671 28916 46683
rect 28860 46665 28862 46671
rect 28862 46665 28914 46671
rect 28914 46665 28916 46671
rect 28860 46619 28862 46641
rect 28862 46619 28914 46641
rect 28914 46619 28916 46641
rect 28860 46607 28916 46619
rect 28860 46585 28862 46607
rect 28862 46585 28914 46607
rect 28914 46585 28916 46607
rect 28860 46555 28862 46561
rect 28862 46555 28914 46561
rect 28914 46555 28916 46561
rect 28860 46543 28916 46555
rect 28860 46505 28862 46543
rect 28862 46505 28914 46543
rect 28914 46505 28916 46543
rect 28860 46479 28916 46481
rect 28860 46427 28862 46479
rect 28862 46427 28914 46479
rect 28914 46427 28916 46479
rect 28860 46425 28916 46427
rect 28860 46363 28862 46401
rect 28862 46363 28914 46401
rect 28914 46363 28916 46401
rect 28860 46351 28916 46363
rect 28860 46345 28862 46351
rect 28862 46345 28914 46351
rect 28914 46345 28916 46351
rect 28860 46299 28862 46321
rect 28862 46299 28914 46321
rect 28914 46299 28916 46321
rect 28860 46287 28916 46299
rect 28860 46265 28862 46287
rect 28862 46265 28914 46287
rect 28914 46265 28916 46287
rect 28860 46235 28862 46241
rect 28862 46235 28914 46241
rect 28914 46235 28916 46241
rect 28860 46223 28916 46235
rect 28860 46185 28862 46223
rect 28862 46185 28914 46223
rect 28914 46185 28916 46223
rect 29948 46683 29950 46721
rect 29950 46683 30002 46721
rect 30002 46683 30004 46721
rect 29948 46671 30004 46683
rect 29948 46665 29950 46671
rect 29950 46665 30002 46671
rect 30002 46665 30004 46671
rect 29948 46619 29950 46641
rect 29950 46619 30002 46641
rect 30002 46619 30004 46641
rect 29948 46607 30004 46619
rect 29948 46585 29950 46607
rect 29950 46585 30002 46607
rect 30002 46585 30004 46607
rect 29948 46555 29950 46561
rect 29950 46555 30002 46561
rect 30002 46555 30004 46561
rect 29948 46543 30004 46555
rect 29948 46505 29950 46543
rect 29950 46505 30002 46543
rect 30002 46505 30004 46543
rect 29948 46479 30004 46481
rect 29948 46427 29950 46479
rect 29950 46427 30002 46479
rect 30002 46427 30004 46479
rect 29948 46425 30004 46427
rect 29948 46363 29950 46401
rect 29950 46363 30002 46401
rect 30002 46363 30004 46401
rect 29948 46351 30004 46363
rect 29948 46345 29950 46351
rect 29950 46345 30002 46351
rect 30002 46345 30004 46351
rect 29948 46299 29950 46321
rect 29950 46299 30002 46321
rect 30002 46299 30004 46321
rect 29948 46287 30004 46299
rect 29948 46265 29950 46287
rect 29950 46265 30002 46287
rect 30002 46265 30004 46287
rect 29948 46235 29950 46241
rect 29950 46235 30002 46241
rect 30002 46235 30004 46241
rect 29948 46223 30004 46235
rect 29948 46185 29950 46223
rect 29950 46185 30002 46223
rect 30002 46185 30004 46223
rect 31036 46683 31038 46721
rect 31038 46683 31090 46721
rect 31090 46683 31092 46721
rect 31036 46671 31092 46683
rect 31036 46665 31038 46671
rect 31038 46665 31090 46671
rect 31090 46665 31092 46671
rect 31036 46619 31038 46641
rect 31038 46619 31090 46641
rect 31090 46619 31092 46641
rect 31036 46607 31092 46619
rect 31036 46585 31038 46607
rect 31038 46585 31090 46607
rect 31090 46585 31092 46607
rect 31036 46555 31038 46561
rect 31038 46555 31090 46561
rect 31090 46555 31092 46561
rect 31036 46543 31092 46555
rect 31036 46505 31038 46543
rect 31038 46505 31090 46543
rect 31090 46505 31092 46543
rect 31036 46479 31092 46481
rect 31036 46427 31038 46479
rect 31038 46427 31090 46479
rect 31090 46427 31092 46479
rect 31036 46425 31092 46427
rect 31036 46363 31038 46401
rect 31038 46363 31090 46401
rect 31090 46363 31092 46401
rect 31036 46351 31092 46363
rect 31036 46345 31038 46351
rect 31038 46345 31090 46351
rect 31090 46345 31092 46351
rect 31036 46299 31038 46321
rect 31038 46299 31090 46321
rect 31090 46299 31092 46321
rect 31036 46287 31092 46299
rect 31036 46265 31038 46287
rect 31038 46265 31090 46287
rect 31090 46265 31092 46287
rect 40593 46315 40649 46371
rect 31036 46235 31038 46241
rect 31038 46235 31090 46241
rect 31090 46235 31092 46241
rect 31036 46223 31092 46235
rect 31036 46185 31038 46223
rect 31038 46185 31090 46223
rect 31090 46185 31092 46223
rect 383 44333 519 45829
rect 364 39871 374 41367
rect 374 39871 490 41367
rect 490 39871 500 41367
rect 10217 39889 10513 46105
rect 18249 45742 18305 45744
rect 18249 45690 18251 45742
rect 18251 45690 18303 45742
rect 18303 45690 18305 45742
rect 18249 45688 18305 45690
rect 18795 45742 18851 45744
rect 18795 45690 18797 45742
rect 18797 45690 18849 45742
rect 18849 45690 18851 45742
rect 18795 45688 18851 45690
rect 19341 45733 19397 45735
rect 19341 45681 19343 45733
rect 19343 45681 19395 45733
rect 19395 45681 19397 45733
rect 19341 45679 19397 45681
rect 19886 45732 19942 45734
rect 19886 45680 19888 45732
rect 19888 45680 19940 45732
rect 19940 45680 19942 45732
rect 19886 45678 19942 45680
rect 21517 45720 21573 45722
rect 21517 45668 21519 45720
rect 21519 45668 21571 45720
rect 21571 45668 21573 45720
rect 21517 45666 21573 45668
rect 22060 45717 22116 45719
rect 22060 45665 22062 45717
rect 22062 45665 22114 45717
rect 22114 45665 22116 45717
rect 22060 45663 22116 45665
rect 22602 45716 22658 45718
rect 22602 45664 22604 45716
rect 22604 45664 22656 45716
rect 22656 45664 22658 45716
rect 22602 45662 22658 45664
rect 23149 45721 23205 45723
rect 23149 45669 23151 45721
rect 23151 45669 23203 45721
rect 23203 45669 23205 45721
rect 23149 45667 23205 45669
rect 25867 45732 25923 45734
rect 25867 45680 25869 45732
rect 25869 45680 25921 45732
rect 25921 45680 25923 45732
rect 25867 45678 25923 45680
rect 26410 45736 26466 45738
rect 26410 45684 26412 45736
rect 26412 45684 26464 45736
rect 26464 45684 26466 45736
rect 26410 45682 26466 45684
rect 26952 45730 27008 45732
rect 26952 45678 26954 45730
rect 26954 45678 27006 45730
rect 27006 45678 27008 45730
rect 26952 45676 27008 45678
rect 27509 45721 27565 45723
rect 27509 45669 27511 45721
rect 27511 45669 27563 45721
rect 27563 45669 27565 45721
rect 27509 45667 27565 45669
rect 29133 45732 29189 45734
rect 29133 45680 29135 45732
rect 29135 45680 29187 45732
rect 29187 45680 29189 45732
rect 29133 45678 29189 45680
rect 29677 45725 29733 45727
rect 29677 45673 29679 45725
rect 29679 45673 29731 45725
rect 29731 45673 29733 45725
rect 29677 45671 29733 45673
rect 30227 45729 30283 45731
rect 30227 45677 30229 45729
rect 30229 45677 30281 45729
rect 30281 45677 30283 45729
rect 30227 45675 30283 45677
rect 30760 45729 30816 45731
rect 30760 45677 30762 45729
rect 30762 45677 30814 45729
rect 30814 45677 30816 45729
rect 30760 45675 30816 45677
rect 39561 44885 39617 44887
rect 39561 44833 39563 44885
rect 39563 44833 39615 44885
rect 39615 44833 39617 44885
rect 39561 44831 39617 44833
rect 41150 45759 41206 45815
rect 40992 44931 41048 44987
rect 39561 44695 39617 44697
rect 39561 44643 39563 44695
rect 39563 44643 39615 44695
rect 39615 44643 39617 44695
rect 39561 44641 39617 44643
rect 39561 43735 39617 43737
rect 39561 43683 39563 43735
rect 39563 43683 39615 43735
rect 39615 43683 39617 43735
rect 39561 43681 39617 43683
rect 44762 45066 44818 45068
rect 44842 45066 44898 45068
rect 44922 45066 44978 45068
rect 45002 45066 45058 45068
rect 45082 45066 45138 45068
rect 45162 45066 45218 45068
rect 45242 45066 45298 45068
rect 44762 45014 44780 45066
rect 44780 45014 44818 45066
rect 44842 45014 44844 45066
rect 44844 45014 44896 45066
rect 44896 45014 44898 45066
rect 44922 45014 44960 45066
rect 44960 45014 44972 45066
rect 44972 45014 44978 45066
rect 45002 45014 45024 45066
rect 45024 45014 45036 45066
rect 45036 45014 45058 45066
rect 45082 45014 45088 45066
rect 45088 45014 45100 45066
rect 45100 45014 45138 45066
rect 45162 45014 45164 45066
rect 45164 45014 45216 45066
rect 45216 45014 45218 45066
rect 45242 45014 45280 45066
rect 45280 45014 45298 45066
rect 44762 45012 44818 45014
rect 44842 45012 44898 45014
rect 44922 45012 44978 45014
rect 45002 45012 45058 45014
rect 45082 45012 45138 45014
rect 45162 45012 45218 45014
rect 45242 45012 45298 45014
rect 40892 44547 40948 44603
rect 40992 43781 41048 43837
rect 39561 43545 39617 43547
rect 39561 43493 39563 43545
rect 39563 43493 39615 43545
rect 39615 43493 39617 43545
rect 39561 43491 39617 43493
rect 46304 44911 46520 44929
rect 46304 44731 46322 44911
rect 46322 44731 46502 44911
rect 46502 44731 46520 44911
rect 46304 44713 46520 44731
rect 41547 44520 41603 44522
rect 41627 44520 41683 44522
rect 41707 44520 41763 44522
rect 41787 44520 41843 44522
rect 41547 44468 41593 44520
rect 41593 44468 41603 44520
rect 41627 44468 41657 44520
rect 41657 44468 41669 44520
rect 41669 44468 41683 44520
rect 41707 44468 41721 44520
rect 41721 44468 41733 44520
rect 41733 44468 41763 44520
rect 41787 44468 41797 44520
rect 41797 44468 41843 44520
rect 41547 44466 41603 44468
rect 41627 44466 41683 44468
rect 41707 44466 41763 44468
rect 41787 44466 41843 44468
rect 44801 43915 44857 43917
rect 44881 43915 44937 43917
rect 44961 43915 45017 43917
rect 45041 43915 45097 43917
rect 45121 43915 45177 43917
rect 45201 43915 45257 43917
rect 44801 43863 44831 43915
rect 44831 43863 44843 43915
rect 44843 43863 44857 43915
rect 44881 43863 44895 43915
rect 44895 43863 44907 43915
rect 44907 43863 44937 43915
rect 44961 43863 44971 43915
rect 44971 43863 45017 43915
rect 45041 43863 45087 43915
rect 45087 43863 45097 43915
rect 45121 43863 45151 43915
rect 45151 43863 45163 43915
rect 45163 43863 45177 43915
rect 45201 43863 45215 43915
rect 45215 43863 45227 43915
rect 45227 43863 45257 43915
rect 44801 43861 44857 43863
rect 44881 43861 44937 43863
rect 44961 43861 45017 43863
rect 45041 43861 45097 43863
rect 45121 43861 45177 43863
rect 45201 43861 45257 43863
rect 46292 43760 46508 43778
rect 46292 43580 46310 43760
rect 46310 43580 46490 43760
rect 46490 43580 46508 43760
rect 46292 43562 46508 43580
rect 40892 43397 40948 43453
rect 41545 43370 41601 43372
rect 41625 43370 41681 43372
rect 41705 43370 41761 43372
rect 41785 43370 41841 43372
rect 41545 43318 41591 43370
rect 41591 43318 41601 43370
rect 41625 43318 41655 43370
rect 41655 43318 41667 43370
rect 41667 43318 41681 43370
rect 41705 43318 41719 43370
rect 41719 43318 41731 43370
rect 41731 43318 41761 43370
rect 41785 43318 41795 43370
rect 41795 43318 41841 43370
rect 41545 43316 41601 43318
rect 41625 43316 41681 43318
rect 41705 43316 41761 43318
rect 41785 43316 41841 43318
rect 40593 42625 40649 42681
rect 39561 41195 39617 41197
rect 39561 41143 39563 41195
rect 39563 41143 39615 41195
rect 39615 41143 39617 41195
rect 39561 41141 39617 41143
rect 41150 42069 41206 42125
rect 40992 41241 41048 41297
rect 39561 41005 39617 41007
rect 39561 40953 39563 41005
rect 39563 40953 39615 41005
rect 39615 40953 39617 41005
rect 39561 40951 39617 40953
rect 39561 39925 39617 39927
rect 39561 39873 39563 39925
rect 39563 39873 39615 39925
rect 39615 39873 39617 39925
rect 39561 39871 39617 39873
rect 44791 41373 44847 41375
rect 44871 41373 44927 41375
rect 44951 41373 45007 41375
rect 45031 41373 45087 41375
rect 45111 41373 45167 41375
rect 45191 41373 45247 41375
rect 44791 41321 44821 41373
rect 44821 41321 44833 41373
rect 44833 41321 44847 41373
rect 44871 41321 44885 41373
rect 44885 41321 44897 41373
rect 44897 41321 44927 41373
rect 44951 41321 44961 41373
rect 44961 41321 45007 41373
rect 45031 41321 45077 41373
rect 45077 41321 45087 41373
rect 45111 41321 45141 41373
rect 45141 41321 45153 41373
rect 45153 41321 45167 41373
rect 45191 41321 45205 41373
rect 45205 41321 45217 41373
rect 45217 41321 45247 41373
rect 44791 41319 44847 41321
rect 44871 41319 44927 41321
rect 44951 41319 45007 41321
rect 45031 41319 45087 41321
rect 45111 41319 45167 41321
rect 45191 41319 45247 41321
rect 40892 40857 40948 40913
rect 40992 39971 41048 40027
rect -27062 39681 -27060 39727
rect -27060 39681 -27008 39727
rect -27008 39681 -27006 39727
rect -27062 39671 -27006 39681
rect -5664 39688 -5662 39824
rect -5662 39688 -170 39824
rect -170 39688 -168 39824
rect 39561 39735 39617 39737
rect 39561 39683 39563 39735
rect 39563 39683 39615 39735
rect 39615 39683 39617 39735
rect 39561 39681 39617 39683
rect 46150 41228 46366 41246
rect 46150 41048 46168 41228
rect 46168 41048 46348 41228
rect 46348 41048 46366 41228
rect 46150 41030 46366 41048
rect 41463 40829 41519 40831
rect 41543 40829 41599 40831
rect 41623 40829 41679 40831
rect 41703 40829 41759 40831
rect 41463 40777 41509 40829
rect 41509 40777 41519 40829
rect 41543 40777 41573 40829
rect 41573 40777 41585 40829
rect 41585 40777 41599 40829
rect 41623 40777 41637 40829
rect 41637 40777 41649 40829
rect 41649 40777 41679 40829
rect 41703 40777 41713 40829
rect 41713 40777 41759 40829
rect 41463 40775 41519 40777
rect 41543 40775 41599 40777
rect 41623 40775 41679 40777
rect 41703 40775 41759 40777
rect 44791 40103 44847 40105
rect 44871 40103 44927 40105
rect 44951 40103 45007 40105
rect 45031 40103 45087 40105
rect 45111 40103 45167 40105
rect 45191 40103 45247 40105
rect 44791 40051 44821 40103
rect 44821 40051 44833 40103
rect 44833 40051 44847 40103
rect 44871 40051 44885 40103
rect 44885 40051 44897 40103
rect 44897 40051 44927 40103
rect 44951 40051 44961 40103
rect 44961 40051 45007 40103
rect 45031 40051 45077 40103
rect 45077 40051 45087 40103
rect 45111 40051 45141 40103
rect 45141 40051 45153 40103
rect 45153 40051 45167 40103
rect 45191 40051 45205 40103
rect 45205 40051 45217 40103
rect 45217 40051 45247 40103
rect 44791 40049 44847 40051
rect 44871 40049 44927 40051
rect 44951 40049 45007 40051
rect 45031 40049 45087 40051
rect 45111 40049 45167 40051
rect 45191 40049 45247 40051
rect 46121 39938 46337 39956
rect 46121 39758 46139 39938
rect 46139 39758 46319 39938
rect 46319 39758 46337 39938
rect 46121 39740 46337 39758
rect -27062 39617 -27060 39647
rect -27060 39617 -27008 39647
rect -27008 39617 -27006 39647
rect -27062 39605 -27006 39617
rect -27062 39591 -27060 39605
rect -27060 39591 -27008 39605
rect -27008 39591 -27006 39605
rect 40892 39587 40948 39643
rect -27062 39553 -27060 39567
rect -27060 39553 -27008 39567
rect -27008 39553 -27006 39567
rect -27062 39541 -27006 39553
rect -27062 39511 -27060 39541
rect -27060 39511 -27008 39541
rect -27008 39511 -27006 39541
rect 41461 39560 41517 39562
rect 41541 39560 41597 39562
rect 41621 39560 41677 39562
rect 41701 39560 41757 39562
rect -18873 39468 -18871 39498
rect -18871 39468 -18819 39498
rect -18819 39468 -18817 39498
rect -18873 39456 -18817 39468
rect -18873 39442 -18871 39456
rect -18871 39442 -18819 39456
rect -18819 39442 -18817 39456
rect 41461 39508 41507 39560
rect 41507 39508 41517 39560
rect 41541 39508 41571 39560
rect 41571 39508 41583 39560
rect 41583 39508 41597 39560
rect 41621 39508 41635 39560
rect 41635 39508 41647 39560
rect 41647 39508 41677 39560
rect 41701 39508 41711 39560
rect 41711 39508 41757 39560
rect 41461 39506 41517 39508
rect 41541 39506 41597 39508
rect 41621 39506 41677 39508
rect 41701 39506 41757 39508
rect -18873 39404 -18871 39418
rect -18871 39404 -18819 39418
rect -18819 39404 -18817 39418
rect -18873 39392 -18817 39404
rect -18873 39362 -18871 39392
rect -18871 39362 -18819 39392
rect -18819 39362 -18817 39392
rect -18873 39328 -18817 39338
rect -18873 39282 -18871 39328
rect -18871 39282 -18819 39328
rect -18819 39282 -18817 39328
rect -18873 39212 -18871 39258
rect -18871 39212 -18819 39258
rect -18819 39212 -18817 39258
rect -18873 39202 -18817 39212
rect -31808 39098 -31806 39144
rect -31806 39098 -31754 39144
rect -31754 39098 -31752 39144
rect -31808 39088 -31752 39098
rect -31808 39034 -31806 39064
rect -31806 39034 -31754 39064
rect -31754 39034 -31752 39064
rect -31808 39022 -31752 39034
rect -31808 39008 -31806 39022
rect -31806 39008 -31754 39022
rect -31754 39008 -31752 39022
rect -31808 38970 -31806 38984
rect -31806 38970 -31754 38984
rect -31754 38970 -31752 38984
rect -31808 38958 -31752 38970
rect -31808 38928 -31806 38958
rect -31806 38928 -31754 38958
rect -31754 38928 -31752 38958
rect -31808 38894 -31752 38904
rect -31808 38848 -31806 38894
rect -31806 38848 -31754 38894
rect -31754 38848 -31752 38894
rect -27068 39066 -27066 39104
rect -27066 39066 -27014 39104
rect -27014 39066 -27012 39104
rect -27068 39054 -27012 39066
rect -27068 39048 -27066 39054
rect -27066 39048 -27014 39054
rect -27014 39048 -27012 39054
rect -27068 39002 -27066 39024
rect -27066 39002 -27014 39024
rect -27014 39002 -27012 39024
rect -27068 38990 -27012 39002
rect -27068 38968 -27066 38990
rect -27066 38968 -27014 38990
rect -27014 38968 -27012 38990
rect -27068 38938 -27066 38944
rect -27066 38938 -27014 38944
rect -27014 38938 -27012 38944
rect -27068 38926 -27012 38938
rect -27068 38888 -27066 38926
rect -27066 38888 -27014 38926
rect -27014 38888 -27012 38926
rect -27068 38862 -27012 38864
rect -27068 38810 -27066 38862
rect -27066 38810 -27014 38862
rect -27014 38810 -27012 38862
rect -27068 38808 -27012 38810
rect -27068 38746 -27066 38784
rect -27066 38746 -27014 38784
rect -27014 38746 -27012 38784
rect -27068 38734 -27012 38746
rect -27068 38728 -27066 38734
rect -27066 38728 -27014 38734
rect -27014 38728 -27012 38734
rect -27068 38682 -27066 38704
rect -27066 38682 -27014 38704
rect -27014 38682 -27012 38704
rect -27068 38670 -27012 38682
rect -27068 38648 -27066 38670
rect -27066 38648 -27014 38670
rect -27014 38648 -27012 38670
rect -31807 38595 -31751 38605
rect -31807 38549 -31805 38595
rect -31805 38549 -31753 38595
rect -31753 38549 -31751 38595
rect -31807 38479 -31805 38525
rect -31805 38479 -31753 38525
rect -31753 38479 -31751 38525
rect -31807 38469 -31751 38479
rect -31807 38415 -31805 38445
rect -31805 38415 -31753 38445
rect -31753 38415 -31751 38445
rect -31807 38403 -31751 38415
rect -31807 38389 -31805 38403
rect -31805 38389 -31753 38403
rect -31753 38389 -31751 38403
rect -27068 38618 -27066 38624
rect -27066 38618 -27014 38624
rect -27014 38618 -27012 38624
rect -27068 38606 -27012 38618
rect -27068 38568 -27066 38606
rect -27066 38568 -27014 38606
rect -27014 38568 -27012 38606
rect -27068 38542 -27012 38544
rect -27068 38490 -27066 38542
rect -27066 38490 -27014 38542
rect -27014 38490 -27012 38542
rect -27068 38488 -27012 38490
rect -31807 38351 -31805 38365
rect -31805 38351 -31753 38365
rect -31753 38351 -31751 38365
rect -31807 38339 -31751 38351
rect -31807 38309 -31805 38339
rect -31805 38309 -31753 38339
rect -31753 38309 -31751 38339
rect -29610 38407 -29554 38409
rect -29530 38407 -29474 38409
rect -29450 38407 -29394 38409
rect -29370 38407 -29314 38409
rect -29290 38407 -29234 38409
rect -29210 38407 -29154 38409
rect -29610 38355 -29600 38407
rect -29600 38355 -29554 38407
rect -29530 38355 -29484 38407
rect -29484 38355 -29474 38407
rect -29450 38355 -29420 38407
rect -29420 38355 -29408 38407
rect -29408 38355 -29394 38407
rect -29370 38355 -29356 38407
rect -29356 38355 -29344 38407
rect -29344 38355 -29314 38407
rect -29290 38355 -29280 38407
rect -29280 38355 -29234 38407
rect -29210 38355 -29164 38407
rect -29164 38355 -29154 38407
rect -29610 38353 -29554 38355
rect -29530 38353 -29474 38355
rect -29450 38353 -29394 38355
rect -29370 38353 -29314 38355
rect -29290 38353 -29234 38355
rect -29210 38353 -29154 38355
rect -27068 38426 -27066 38464
rect -27066 38426 -27014 38464
rect -27014 38426 -27012 38464
rect -27068 38414 -27012 38426
rect -27068 38408 -27066 38414
rect -27066 38408 -27014 38414
rect -27014 38408 -27012 38414
rect -31807 38275 -31751 38285
rect -31807 38229 -31805 38275
rect -31805 38229 -31753 38275
rect -31753 38229 -31751 38275
rect -27068 38362 -27066 38384
rect -27066 38362 -27014 38384
rect -27014 38362 -27012 38384
rect -27068 38350 -27012 38362
rect -27068 38328 -27066 38350
rect -27066 38328 -27014 38350
rect -27014 38328 -27012 38350
rect -31807 38159 -31805 38205
rect -31805 38159 -31753 38205
rect -31753 38159 -31751 38205
rect -31807 38149 -31751 38159
rect -27068 38298 -27066 38304
rect -27066 38298 -27014 38304
rect -27014 38298 -27012 38304
rect -27068 38286 -27012 38298
rect -27068 38248 -27066 38286
rect -27066 38248 -27014 38286
rect -27014 38248 -27012 38286
rect -18873 39148 -18871 39178
rect -18871 39148 -18819 39178
rect -18819 39148 -18817 39178
rect -18873 39136 -18817 39148
rect -18873 39122 -18871 39136
rect -18871 39122 -18819 39136
rect -18819 39122 -18817 39136
rect -18873 39084 -18871 39098
rect -18871 39084 -18819 39098
rect -18819 39084 -18817 39098
rect -18873 39072 -18817 39084
rect -18873 39042 -18871 39072
rect -18871 39042 -18819 39072
rect -18819 39042 -18817 39072
rect -18873 39008 -18817 39018
rect -18873 38962 -18871 39008
rect -18871 38962 -18819 39008
rect -18819 38962 -18817 39008
rect -18873 38892 -18871 38938
rect -18871 38892 -18819 38938
rect -18819 38892 -18817 38938
rect -18873 38882 -18817 38892
rect -18873 38828 -18871 38858
rect -18871 38828 -18819 38858
rect -18819 38828 -18817 38858
rect -18873 38816 -18817 38828
rect -18873 38802 -18871 38816
rect -18871 38802 -18819 38816
rect -18819 38802 -18817 38816
rect 1477 38818 1533 38874
rect 2526 38851 2582 38869
rect 2526 38813 2528 38851
rect 2528 38813 2580 38851
rect 2580 38813 2582 38851
rect -18873 38764 -18871 38778
rect -18871 38764 -18819 38778
rect -18819 38764 -18817 38778
rect -18873 38752 -18817 38764
rect -18873 38722 -18871 38752
rect -18871 38722 -18819 38752
rect -18819 38722 -18817 38752
rect -18873 38688 -18817 38698
rect -18873 38642 -18871 38688
rect -18871 38642 -18819 38688
rect -18819 38642 -18817 38688
rect 2526 38787 2582 38789
rect 2526 38735 2528 38787
rect 2528 38735 2580 38787
rect 2580 38735 2582 38787
rect 2526 38733 2582 38735
rect 2526 38671 2528 38709
rect 2528 38671 2580 38709
rect 2580 38671 2582 38709
rect 2526 38653 2582 38671
rect -18873 38572 -18871 38618
rect -18871 38572 -18819 38618
rect -18819 38572 -18817 38618
rect -18873 38562 -18817 38572
rect -18873 38508 -18871 38538
rect -18871 38508 -18819 38538
rect -18819 38508 -18817 38538
rect -18873 38496 -18817 38508
rect -18873 38482 -18871 38496
rect -18871 38482 -18819 38496
rect -18819 38482 -18817 38496
rect -18873 38444 -18871 38458
rect -18871 38444 -18819 38458
rect -18819 38444 -18817 38458
rect -18873 38432 -18817 38444
rect -18873 38402 -18871 38432
rect -18871 38402 -18819 38432
rect -18819 38402 -18817 38432
rect -18873 38368 -18817 38378
rect -18873 38322 -18871 38368
rect -18871 38322 -18819 38368
rect -18819 38322 -18817 38368
rect -18873 38252 -18871 38298
rect -18871 38252 -18819 38298
rect -18819 38252 -18817 38298
rect -18873 38242 -18817 38252
rect -35508 37540 -35292 37558
rect -35508 37360 -35490 37540
rect -35490 37360 -35310 37540
rect -35310 37360 -35292 37540
rect -35508 37342 -35292 37360
rect -18873 38188 -18871 38218
rect -18871 38188 -18819 38218
rect -18819 38188 -18817 38218
rect -18873 38176 -18817 38188
rect -18873 38162 -18871 38176
rect -18871 38162 -18819 38176
rect -18819 38162 -18817 38176
rect -18873 38124 -18871 38138
rect -18871 38124 -18819 38138
rect -18819 38124 -18817 38138
rect -18873 38112 -18817 38124
rect -18873 38082 -18871 38112
rect -18871 38082 -18819 38112
rect -18819 38082 -18817 38112
rect 2536 38394 2592 38396
rect 2536 38342 2538 38394
rect 2538 38342 2590 38394
rect 2590 38342 2592 38394
rect 2536 38340 2592 38342
rect 2536 38278 2538 38316
rect 2538 38278 2590 38316
rect 2590 38278 2592 38316
rect 2536 38266 2592 38278
rect 2536 38260 2538 38266
rect 2538 38260 2590 38266
rect 2590 38260 2592 38266
rect 2536 38214 2538 38236
rect 2538 38214 2590 38236
rect 2590 38214 2592 38236
rect 2536 38202 2592 38214
rect 2536 38180 2538 38202
rect 2538 38180 2590 38202
rect 2590 38180 2592 38202
rect 2536 38150 2538 38156
rect 2538 38150 2590 38156
rect 2590 38150 2592 38156
rect 2536 38138 2592 38150
rect 2536 38100 2538 38138
rect 2538 38100 2590 38138
rect 2590 38100 2592 38138
rect -18873 38048 -18817 38058
rect -18873 38002 -18871 38048
rect -18871 38002 -18819 38048
rect -18819 38002 -18817 38048
rect 2000 38009 2056 38065
rect 2536 38074 2592 38076
rect 2536 38022 2538 38074
rect 2538 38022 2590 38074
rect 2590 38022 2592 38074
rect 2536 38020 2592 38022
rect -18873 37932 -18871 37978
rect -18871 37932 -18819 37978
rect -18819 37932 -18817 37978
rect -18873 37922 -18817 37932
rect -18873 37868 -18871 37898
rect -18871 37868 -18819 37898
rect -18819 37868 -18817 37898
rect -18873 37856 -18817 37868
rect -18873 37842 -18871 37856
rect -18871 37842 -18819 37856
rect -18819 37842 -18817 37856
rect -18873 37804 -18871 37818
rect -18871 37804 -18819 37818
rect -18819 37804 -18817 37818
rect -18873 37792 -18817 37804
rect -18873 37762 -18871 37792
rect -18871 37762 -18819 37792
rect -18819 37762 -18817 37792
rect -18873 37728 -18817 37738
rect -18873 37682 -18871 37728
rect -18871 37682 -18819 37728
rect -18819 37682 -18817 37728
rect -18873 37612 -18871 37658
rect -18871 37612 -18819 37658
rect -18819 37612 -18817 37658
rect -18873 37602 -18817 37612
rect -18873 37548 -18871 37578
rect -18871 37548 -18819 37578
rect -18819 37548 -18817 37578
rect -18873 37536 -18817 37548
rect -18873 37522 -18871 37536
rect -18871 37522 -18819 37536
rect -18819 37522 -18817 37536
rect -18873 37484 -18871 37498
rect -18871 37484 -18819 37498
rect -18819 37484 -18817 37498
rect -18873 37472 -18817 37484
rect -18873 37442 -18871 37472
rect -18871 37442 -18819 37472
rect -18819 37442 -18817 37472
rect -29626 37317 -29570 37319
rect -29546 37317 -29490 37319
rect -29466 37317 -29410 37319
rect -29386 37317 -29330 37319
rect -29306 37317 -29250 37319
rect -29226 37317 -29170 37319
rect -29626 37265 -29596 37317
rect -29596 37265 -29584 37317
rect -29584 37265 -29570 37317
rect -29546 37265 -29532 37317
rect -29532 37265 -29520 37317
rect -29520 37265 -29490 37317
rect -29466 37265 -29456 37317
rect -29456 37265 -29410 37317
rect -29386 37265 -29340 37317
rect -29340 37265 -29330 37317
rect -29306 37265 -29276 37317
rect -29276 37265 -29264 37317
rect -29264 37265 -29250 37317
rect -29226 37265 -29212 37317
rect -29212 37265 -29200 37317
rect -29200 37265 -29170 37317
rect -29626 37263 -29570 37265
rect -29546 37263 -29490 37265
rect -29466 37263 -29410 37265
rect -29386 37263 -29330 37265
rect -29306 37263 -29250 37265
rect -29226 37263 -29170 37265
rect -27065 37299 -27063 37337
rect -27063 37299 -27011 37337
rect -27011 37299 -27009 37337
rect -27065 37287 -27009 37299
rect -27065 37281 -27063 37287
rect -27063 37281 -27011 37287
rect -27011 37281 -27009 37287
rect -27065 37235 -27063 37257
rect -27063 37235 -27011 37257
rect -27011 37235 -27009 37257
rect -27065 37223 -27009 37235
rect -27065 37201 -27063 37223
rect -27063 37201 -27011 37223
rect -27011 37201 -27009 37223
rect -27065 37171 -27063 37177
rect -27063 37171 -27011 37177
rect -27011 37171 -27009 37177
rect -27065 37159 -27009 37171
rect -27065 37121 -27063 37159
rect -27063 37121 -27011 37159
rect -27011 37121 -27009 37159
rect -27065 37095 -27009 37097
rect -27065 37043 -27063 37095
rect -27063 37043 -27011 37095
rect -27011 37043 -27009 37095
rect -27065 37041 -27009 37043
rect -27065 36979 -27063 37017
rect -27063 36979 -27011 37017
rect -27011 36979 -27009 37017
rect -27065 36967 -27009 36979
rect -27065 36961 -27063 36967
rect -27063 36961 -27011 36967
rect -27011 36961 -27009 36967
rect -27065 36915 -27063 36937
rect -27063 36915 -27011 36937
rect -27011 36915 -27009 36937
rect -27065 36903 -27009 36915
rect -27065 36881 -27063 36903
rect -27063 36881 -27011 36903
rect -27011 36881 -27009 36903
rect -27065 36851 -27063 36857
rect -27063 36851 -27011 36857
rect -27011 36851 -27009 36857
rect -27065 36839 -27009 36851
rect -27065 36801 -27063 36839
rect -27063 36801 -27011 36839
rect -27011 36801 -27009 36839
rect -27065 36775 -27009 36777
rect -27065 36723 -27063 36775
rect -27063 36723 -27011 36775
rect -27011 36723 -27009 36775
rect -27065 36721 -27009 36723
rect -27065 36659 -27063 36697
rect -27063 36659 -27011 36697
rect -27011 36659 -27009 36697
rect -27065 36647 -27009 36659
rect -27065 36641 -27063 36647
rect -27063 36641 -27011 36647
rect -27011 36641 -27009 36647
rect -27065 36595 -27063 36617
rect -27063 36595 -27011 36617
rect -27011 36595 -27009 36617
rect -27065 36583 -27009 36595
rect -27065 36561 -27063 36583
rect -27063 36561 -27011 36583
rect -27011 36561 -27009 36583
rect -27065 36531 -27063 36537
rect -27063 36531 -27011 36537
rect -27011 36531 -27009 36537
rect -27065 36519 -27009 36531
rect -27065 36481 -27063 36519
rect -27063 36481 -27011 36519
rect -27011 36481 -27009 36519
rect -18873 37408 -18817 37418
rect -18873 37362 -18871 37408
rect -18871 37362 -18819 37408
rect -18819 37362 -18817 37408
rect -18873 37292 -18871 37338
rect -18871 37292 -18819 37338
rect -18819 37292 -18817 37338
rect -18873 37282 -18817 37292
rect -18873 37228 -18871 37258
rect -18871 37228 -18819 37258
rect -18819 37228 -18817 37258
rect -18873 37216 -18817 37228
rect -18873 37202 -18871 37216
rect -18871 37202 -18819 37216
rect -18819 37202 -18817 37216
rect -18873 37164 -18871 37178
rect -18871 37164 -18819 37178
rect -18819 37164 -18817 37178
rect -18873 37152 -18817 37164
rect -18873 37122 -18871 37152
rect -18871 37122 -18819 37152
rect -18819 37122 -18817 37152
rect -18873 37088 -18817 37098
rect -18873 37042 -18871 37088
rect -18871 37042 -18819 37088
rect -18819 37042 -18817 37088
rect 1477 37069 1533 37125
rect 2172 37093 2174 37131
rect 2174 37093 2226 37131
rect 2226 37093 2228 37131
rect 2172 37081 2228 37093
rect 2172 37075 2174 37081
rect 2174 37075 2226 37081
rect 2226 37075 2228 37081
rect -18873 36972 -18871 37018
rect -18871 36972 -18819 37018
rect -18819 36972 -18817 37018
rect -18873 36962 -18817 36972
rect -18873 36908 -18871 36938
rect -18871 36908 -18819 36938
rect -18819 36908 -18817 36938
rect -18873 36896 -18817 36908
rect -18873 36882 -18871 36896
rect -18871 36882 -18819 36896
rect -18819 36882 -18817 36896
rect 2172 37029 2174 37051
rect 2174 37029 2226 37051
rect 2226 37029 2228 37051
rect 2172 37017 2228 37029
rect 2172 36995 2174 37017
rect 2174 36995 2226 37017
rect 2226 36995 2228 37017
rect 2172 36965 2174 36971
rect 2174 36965 2226 36971
rect 2226 36965 2228 36971
rect 2172 36953 2228 36965
rect 2172 36915 2174 36953
rect 2174 36915 2226 36953
rect 2226 36915 2228 36953
rect -18873 36844 -18871 36858
rect -18871 36844 -18819 36858
rect -18819 36844 -18817 36858
rect -18873 36832 -18817 36844
rect -18873 36802 -18871 36832
rect -18871 36802 -18819 36832
rect -18819 36802 -18817 36832
rect -18873 36768 -18817 36778
rect -18873 36722 -18871 36768
rect -18871 36722 -18819 36768
rect -18819 36722 -18817 36768
rect -18873 36652 -18871 36698
rect -18871 36652 -18819 36698
rect -18819 36652 -18817 36698
rect -18873 36642 -18817 36652
rect -18873 36588 -18871 36618
rect -18871 36588 -18819 36618
rect -18819 36588 -18817 36618
rect -18873 36576 -18817 36588
rect -18873 36562 -18871 36576
rect -18871 36562 -18819 36576
rect -18819 36562 -18817 36576
rect -18873 36524 -18871 36538
rect -18871 36524 -18819 36538
rect -18819 36524 -18817 36538
rect -18873 36512 -18817 36524
rect -18873 36482 -18871 36512
rect -18871 36482 -18819 36512
rect -18819 36482 -18817 36512
rect -18873 36448 -18817 36458
rect -18873 36402 -18871 36448
rect -18871 36402 -18819 36448
rect -18819 36402 -18817 36448
rect -18873 36332 -18871 36378
rect -18871 36332 -18819 36378
rect -18819 36332 -18817 36378
rect -18873 36322 -18817 36332
rect 2173 36645 2229 36647
rect 2173 36593 2175 36645
rect 2175 36593 2227 36645
rect 2227 36593 2229 36645
rect 2173 36591 2229 36593
rect 2173 36529 2175 36567
rect 2175 36529 2227 36567
rect 2227 36529 2229 36567
rect 2173 36517 2229 36529
rect 2173 36511 2175 36517
rect 2175 36511 2227 36517
rect 2227 36511 2229 36517
rect 2173 36465 2175 36487
rect 2175 36465 2227 36487
rect 2227 36465 2229 36487
rect 2173 36453 2229 36465
rect 2173 36431 2175 36453
rect 2175 36431 2227 36453
rect 2227 36431 2229 36453
rect 2173 36401 2175 36407
rect 2175 36401 2227 36407
rect 2227 36401 2229 36407
rect 2173 36389 2229 36401
rect 2173 36351 2175 36389
rect 2175 36351 2227 36389
rect 2227 36351 2229 36389
rect -18873 36268 -18871 36298
rect -18871 36268 -18819 36298
rect -18819 36268 -18817 36298
rect -18873 36256 -18817 36268
rect -18873 36242 -18871 36256
rect -18871 36242 -18819 36256
rect -18819 36242 -18817 36256
rect 2000 36259 2056 36315
rect 2173 36325 2229 36327
rect 2173 36273 2175 36325
rect 2175 36273 2227 36325
rect 2227 36273 2229 36325
rect 2173 36271 2229 36273
rect -27065 36090 -27063 36120
rect -27063 36090 -27011 36120
rect -27011 36090 -27009 36120
rect -27065 36078 -27009 36090
rect -27065 36064 -27063 36078
rect -27063 36064 -27011 36078
rect -27011 36064 -27009 36078
rect -18873 36204 -18871 36218
rect -18871 36204 -18819 36218
rect -18819 36204 -18817 36218
rect -18873 36192 -18817 36204
rect -18873 36162 -18871 36192
rect -18871 36162 -18819 36192
rect -18819 36162 -18817 36192
rect -27065 36026 -27063 36040
rect -27063 36026 -27011 36040
rect -27011 36026 -27009 36040
rect -27065 36014 -27009 36026
rect -27065 35984 -27063 36014
rect -27063 35984 -27011 36014
rect -27011 35984 -27009 36014
rect 2952 36085 3008 36087
rect 3032 36085 3088 36087
rect 3112 36085 3168 36087
rect 3192 36085 3248 36087
rect 3272 36085 3328 36087
rect 2952 36033 2954 36085
rect 2954 36033 3006 36085
rect 3006 36033 3008 36085
rect 3032 36033 3070 36085
rect 3070 36033 3082 36085
rect 3082 36033 3088 36085
rect 3112 36033 3134 36085
rect 3134 36033 3146 36085
rect 3146 36033 3168 36085
rect 3192 36033 3198 36085
rect 3198 36033 3210 36085
rect 3210 36033 3248 36085
rect 3272 36033 3274 36085
rect 3274 36033 3326 36085
rect 3326 36033 3328 36085
rect 2952 36031 3008 36033
rect 3032 36031 3088 36033
rect 3112 36031 3168 36033
rect 3192 36031 3248 36033
rect 3272 36031 3328 36033
rect 3588 36088 3644 36090
rect 3668 36088 3724 36090
rect 3748 36088 3804 36090
rect 3588 36036 3606 36088
rect 3606 36036 3644 36088
rect 3668 36036 3670 36088
rect 3670 36036 3722 36088
rect 3722 36036 3724 36088
rect 3748 36036 3786 36088
rect 3786 36036 3804 36088
rect 3588 36034 3644 36036
rect 3668 36034 3724 36036
rect 3748 36034 3804 36036
rect -27065 35950 -27009 35960
rect -27065 35904 -27063 35950
rect -27063 35904 -27011 35950
rect -27011 35904 -27009 35950
rect -27065 35834 -27063 35880
rect -27063 35834 -27011 35880
rect -27011 35834 -27009 35880
rect -27065 35824 -27009 35834
rect 6349 36537 6405 36593
rect 5055 36087 5111 36089
rect 5135 36087 5191 36089
rect 5215 36087 5271 36089
rect 5295 36087 5351 36089
rect 5055 36035 5081 36087
rect 5081 36035 5111 36087
rect 5135 36035 5145 36087
rect 5145 36035 5191 36087
rect 5215 36035 5261 36087
rect 5261 36035 5271 36087
rect 5295 36035 5325 36087
rect 5325 36035 5351 36087
rect 5055 36033 5111 36035
rect 5135 36033 5191 36035
rect 5215 36033 5271 36035
rect 5295 36033 5351 36035
rect 5579 36088 5635 36090
rect 5659 36088 5715 36090
rect 5739 36088 5795 36090
rect 5579 36036 5597 36088
rect 5597 36036 5635 36088
rect 5659 36036 5661 36088
rect 5661 36036 5713 36088
rect 5713 36036 5715 36088
rect 5739 36036 5777 36088
rect 5777 36036 5795 36088
rect 5579 36034 5635 36036
rect 5659 36034 5715 36036
rect 5739 36034 5795 36036
rect 6349 36193 6405 36249
rect 6938 36080 6994 36082
rect 7018 36080 7074 36082
rect 7098 36080 7154 36082
rect 6938 36028 6956 36080
rect 6956 36028 6994 36080
rect 7018 36028 7020 36080
rect 7020 36028 7072 36080
rect 7072 36028 7074 36080
rect 7098 36028 7136 36080
rect 7136 36028 7154 36080
rect 6938 36026 6994 36028
rect 7018 36026 7074 36028
rect 7098 36026 7154 36028
rect 7384 36087 7440 36089
rect 7464 36087 7520 36089
rect 7544 36087 7600 36089
rect 7624 36087 7680 36089
rect 7384 36035 7410 36087
rect 7410 36035 7440 36087
rect 7464 36035 7474 36087
rect 7474 36035 7520 36087
rect 7544 36035 7590 36087
rect 7590 36035 7600 36087
rect 7624 36035 7654 36087
rect 7654 36035 7680 36087
rect 7384 36033 7440 36035
rect 7464 36033 7520 36035
rect 7544 36033 7600 36035
rect 7624 36033 7680 36035
rect 8946 36086 9002 36088
rect 9026 36086 9082 36088
rect 9106 36086 9162 36088
rect 9186 36086 9242 36088
rect 9266 36086 9322 36088
rect 8946 36034 8948 36086
rect 8948 36034 9000 36086
rect 9000 36034 9002 36086
rect 9026 36034 9064 36086
rect 9064 36034 9076 36086
rect 9076 36034 9082 36086
rect 9106 36034 9128 36086
rect 9128 36034 9140 36086
rect 9140 36034 9162 36086
rect 9186 36034 9192 36086
rect 9192 36034 9204 36086
rect 9204 36034 9242 36086
rect 9266 36034 9268 36086
rect 9268 36034 9320 36086
rect 9320 36034 9322 36086
rect 8946 36032 9002 36034
rect 9026 36032 9082 36034
rect 9106 36032 9162 36034
rect 9186 36032 9242 36034
rect 9266 36032 9322 36034
rect 9580 36083 9636 36085
rect 9660 36083 9716 36085
rect 9740 36083 9796 36085
rect 9580 36031 9598 36083
rect 9598 36031 9636 36083
rect 9660 36031 9662 36083
rect 9662 36031 9714 36083
rect 9714 36031 9716 36083
rect 9740 36031 9778 36083
rect 9778 36031 9796 36083
rect 9580 36029 9636 36031
rect 9660 36029 9716 36031
rect 9740 36029 9796 36031
rect -27065 35770 -27063 35800
rect -27063 35770 -27011 35800
rect -27011 35770 -27009 35800
rect -27065 35758 -27009 35770
rect -27065 35744 -27063 35758
rect -27063 35744 -27011 35758
rect -27011 35744 -27009 35758
rect -27065 35706 -27063 35720
rect -27063 35706 -27011 35720
rect -27011 35706 -27009 35720
rect -27065 35694 -27009 35706
rect -27065 35664 -27063 35694
rect -27063 35664 -27011 35694
rect -27011 35664 -27009 35694
rect -27065 35630 -27009 35640
rect -27065 35584 -27063 35630
rect -27063 35584 -27011 35630
rect -27011 35584 -27009 35630
rect -27065 35514 -27063 35560
rect -27063 35514 -27011 35560
rect -27011 35514 -27009 35560
rect -27065 35504 -27009 35514
rect -27065 35450 -27063 35480
rect -27063 35450 -27011 35480
rect -27011 35450 -27009 35480
rect -27065 35438 -27009 35450
rect -27065 35424 -27063 35438
rect -27063 35424 -27011 35438
rect -27011 35424 -27009 35438
rect -27065 35386 -27063 35400
rect -27063 35386 -27011 35400
rect -27011 35386 -27009 35400
rect -27065 35374 -27009 35386
rect -27065 35344 -27063 35374
rect -27063 35344 -27011 35374
rect -27011 35344 -27009 35374
rect -27065 35310 -27009 35320
rect -27065 35264 -27063 35310
rect -27063 35264 -27011 35310
rect -27011 35264 -27009 35310
rect -27065 35194 -27063 35240
rect -27063 35194 -27011 35240
rect -27011 35194 -27009 35240
rect -27065 35184 -27009 35194
rect -27065 35130 -27063 35160
rect -27063 35130 -27011 35160
rect -27011 35130 -27009 35160
rect -27065 35118 -27009 35130
rect -27065 35104 -27063 35118
rect -27063 35104 -27011 35118
rect -27011 35104 -27009 35118
rect -27065 35066 -27063 35080
rect -27063 35066 -27011 35080
rect -27011 35066 -27009 35080
rect -27065 35054 -27009 35066
rect -27065 35024 -27063 35054
rect -27063 35024 -27011 35054
rect -27011 35024 -27009 35054
rect -27068 34664 -27012 34682
rect -27068 34626 -27066 34664
rect -27066 34626 -27014 34664
rect -27014 34626 -27012 34664
rect -9365 34670 -9309 34672
rect -9365 34618 -9363 34670
rect -9363 34618 -9311 34670
rect -9311 34618 -9309 34670
rect -9365 34616 -9309 34618
rect -27068 34600 -27012 34602
rect -27068 34548 -27066 34600
rect -27066 34548 -27014 34600
rect -27014 34548 -27012 34600
rect -27068 34546 -27012 34548
rect -27068 34484 -27066 34522
rect -27066 34484 -27014 34522
rect -27014 34484 -27012 34522
rect -27068 34472 -27012 34484
rect -27068 34466 -27066 34472
rect -27066 34466 -27014 34472
rect -27014 34466 -27012 34472
rect -27068 34420 -27066 34442
rect -27066 34420 -27014 34442
rect -27014 34420 -27012 34442
rect -27068 34408 -27012 34420
rect -27068 34386 -27066 34408
rect -27066 34386 -27014 34408
rect -27014 34386 -27012 34408
rect -27068 34356 -27066 34362
rect -27066 34356 -27014 34362
rect -27014 34356 -27012 34362
rect -27068 34344 -27012 34356
rect -27068 34306 -27066 34344
rect -27066 34306 -27014 34344
rect -27014 34306 -27012 34344
rect -27068 34280 -27012 34282
rect -27068 34228 -27066 34280
rect -27066 34228 -27014 34280
rect -27014 34228 -27012 34280
rect -27068 34226 -27012 34228
rect -27068 34164 -27066 34202
rect -27066 34164 -27014 34202
rect -27014 34164 -27012 34202
rect -27068 34152 -27012 34164
rect -27068 34146 -27066 34152
rect -27066 34146 -27014 34152
rect -27014 34146 -27012 34152
rect 5936 34135 5992 34191
rect -27068 34100 -27066 34122
rect -27066 34100 -27014 34122
rect -27014 34100 -27012 34122
rect -27068 34088 -27012 34100
rect -27068 34066 -27066 34088
rect -27066 34066 -27014 34088
rect -27014 34066 -27012 34088
rect -27068 34036 -27066 34042
rect -27066 34036 -27014 34042
rect -27014 34036 -27012 34042
rect -27068 34024 -27012 34036
rect -27068 33986 -27066 34024
rect -27066 33986 -27014 34024
rect -27014 33986 -27012 34024
rect -27068 33960 -27012 33962
rect -27068 33908 -27066 33960
rect -27066 33908 -27014 33960
rect -27014 33908 -27012 33960
rect -27068 33906 -27012 33908
rect -27068 33844 -27066 33882
rect -27066 33844 -27014 33882
rect -27014 33844 -27012 33882
rect -27068 33832 -27012 33844
rect -27068 33826 -27066 33832
rect -27066 33826 -27014 33832
rect -27014 33826 -27012 33832
rect -27068 33780 -27066 33802
rect -27066 33780 -27014 33802
rect -27014 33780 -27012 33802
rect -27068 33768 -27012 33780
rect -27068 33746 -27066 33768
rect -27066 33746 -27014 33768
rect -27014 33746 -27012 33768
rect 6742 33790 6798 33846
rect -27068 33716 -27066 33722
rect -27066 33716 -27014 33722
rect -27014 33716 -27012 33722
rect -27068 33704 -27012 33716
rect -27068 33666 -27066 33704
rect -27066 33666 -27014 33704
rect -27014 33666 -27012 33704
rect -27068 33640 -27012 33642
rect -27068 33588 -27066 33640
rect -27066 33588 -27014 33640
rect -27014 33588 -27012 33640
rect -27068 33586 -27012 33588
rect -27068 33524 -27066 33562
rect -27066 33524 -27014 33562
rect -27014 33524 -27012 33562
rect -27068 33506 -27012 33524
rect -21514 33491 -21458 33547
rect -6944 33173 -6888 33175
rect -6944 33121 -6942 33173
rect -6942 33121 -6890 33173
rect -6890 33121 -6888 33173
rect -6944 33119 -6888 33121
rect -27073 32830 -27071 32860
rect -27071 32830 -27019 32860
rect -27019 32830 -27017 32860
rect -27073 32818 -27017 32830
rect -27073 32804 -27071 32818
rect -27071 32804 -27019 32818
rect -27019 32804 -27017 32818
rect -27073 32766 -27071 32780
rect -27071 32766 -27019 32780
rect -27019 32766 -27017 32780
rect -27073 32754 -27017 32766
rect -27073 32724 -27071 32754
rect -27071 32724 -27019 32754
rect -27019 32724 -27017 32754
rect -27073 32690 -27017 32700
rect -27073 32644 -27071 32690
rect -27071 32644 -27019 32690
rect -27019 32644 -27017 32690
rect -27073 32574 -27071 32620
rect -27071 32574 -27019 32620
rect -27019 32574 -27017 32620
rect -27073 32564 -27017 32574
rect -27073 32510 -27071 32540
rect -27071 32510 -27019 32540
rect -27019 32510 -27017 32540
rect -27073 32498 -27017 32510
rect -27073 32484 -27071 32498
rect -27071 32484 -27019 32498
rect -27019 32484 -27017 32498
rect -27073 32446 -27071 32460
rect -27071 32446 -27019 32460
rect -27019 32446 -27017 32460
rect -27073 32434 -27017 32446
rect -27073 32404 -27071 32434
rect -27071 32404 -27019 32434
rect -27019 32404 -27017 32434
rect 5321 32285 5377 32341
rect 7368 32292 7424 32348
rect 7969 31751 8025 31807
rect 4358 30426 4414 30428
rect 4358 30374 4360 30426
rect 4360 30374 4412 30426
rect 4412 30374 4414 30426
rect 4358 30372 4414 30374
rect 8332 30431 8388 30433
rect 8332 30379 8334 30431
rect 8334 30379 8386 30431
rect 8386 30379 8388 30431
rect 8332 30377 8388 30379
rect 3330 30245 3386 30301
rect -12689 29746 -12633 29748
rect -12689 29694 -12687 29746
rect -12687 29694 -12635 29746
rect -12635 29694 -12633 29746
rect -12689 29692 -12633 29694
rect 1917 29692 1973 29748
rect 16725 29692 16781 29748
rect -13465 29323 -13409 29325
rect -13465 29271 -13463 29323
rect -13463 29271 -13411 29323
rect -13411 29271 -13409 29323
rect -13465 29269 -13409 29271
rect 1917 29269 1973 29325
rect 17416 29269 17472 29325
rect -38151 26588 -38095 26590
rect -38071 26588 -38015 26590
rect -37991 26588 -37935 26590
rect -37911 26588 -37855 26590
rect -37831 26588 -37775 26590
rect -37751 26588 -37695 26590
rect -37671 26588 -37615 26590
rect -37591 26588 -37535 26590
rect -37511 26588 -37455 26590
rect -37431 26588 -37375 26590
rect -37351 26588 -37295 26590
rect -37271 26588 -37215 26590
rect -37191 26588 -37135 26590
rect -37111 26588 -37055 26590
rect -37031 26588 -36975 26590
rect -36951 26588 -36895 26590
rect -36871 26588 -36815 26590
rect -36791 26588 -36735 26590
rect -36711 26588 -36655 26590
rect -36631 26588 -36575 26590
rect -36551 26588 -36495 26590
rect -36471 26588 -36415 26590
rect -36391 26588 -36335 26590
rect -36311 26588 -36255 26590
rect -36231 26588 -36175 26590
rect -36151 26588 -36095 26590
rect -36071 26588 -36015 26590
rect -35991 26588 -35935 26590
rect -35911 26588 -35855 26590
rect -35831 26588 -35775 26590
rect -35751 26588 -35695 26590
rect -35671 26588 -35615 26590
rect -35591 26588 -35535 26590
rect -35511 26588 -35455 26590
rect -35431 26588 -35375 26590
rect -35351 26588 -35295 26590
rect -35271 26588 -35215 26590
rect -35191 26588 -35135 26590
rect -35111 26588 -35055 26590
rect -35031 26588 -34975 26590
rect -34951 26588 -34895 26590
rect -38151 26536 -38129 26588
rect -38129 26536 -38117 26588
rect -38117 26536 -38095 26588
rect -38071 26536 -38065 26588
rect -38065 26536 -38053 26588
rect -38053 26536 -38015 26588
rect -37991 26536 -37989 26588
rect -37989 26536 -37937 26588
rect -37937 26536 -37935 26588
rect -37911 26536 -37873 26588
rect -37873 26536 -37861 26588
rect -37861 26536 -37855 26588
rect -37831 26536 -37809 26588
rect -37809 26536 -37797 26588
rect -37797 26536 -37775 26588
rect -37751 26536 -37745 26588
rect -37745 26536 -37733 26588
rect -37733 26536 -37695 26588
rect -37671 26536 -37669 26588
rect -37669 26536 -37617 26588
rect -37617 26536 -37615 26588
rect -37591 26536 -37553 26588
rect -37553 26536 -37541 26588
rect -37541 26536 -37535 26588
rect -37511 26536 -37489 26588
rect -37489 26536 -37477 26588
rect -37477 26536 -37455 26588
rect -37431 26536 -37425 26588
rect -37425 26536 -37413 26588
rect -37413 26536 -37375 26588
rect -37351 26536 -37349 26588
rect -37349 26536 -37297 26588
rect -37297 26536 -37295 26588
rect -37271 26536 -37233 26588
rect -37233 26536 -37221 26588
rect -37221 26536 -37215 26588
rect -37191 26536 -37169 26588
rect -37169 26536 -37157 26588
rect -37157 26536 -37135 26588
rect -37111 26536 -37105 26588
rect -37105 26536 -37093 26588
rect -37093 26536 -37055 26588
rect -37031 26536 -37029 26588
rect -37029 26536 -36977 26588
rect -36977 26536 -36975 26588
rect -36951 26536 -36913 26588
rect -36913 26536 -36901 26588
rect -36901 26536 -36895 26588
rect -36871 26536 -36849 26588
rect -36849 26536 -36837 26588
rect -36837 26536 -36815 26588
rect -36791 26536 -36785 26588
rect -36785 26536 -36773 26588
rect -36773 26536 -36735 26588
rect -36711 26536 -36709 26588
rect -36709 26536 -36657 26588
rect -36657 26536 -36655 26588
rect -36631 26536 -36593 26588
rect -36593 26536 -36581 26588
rect -36581 26536 -36575 26588
rect -36551 26536 -36529 26588
rect -36529 26536 -36517 26588
rect -36517 26536 -36495 26588
rect -36471 26536 -36465 26588
rect -36465 26536 -36453 26588
rect -36453 26536 -36415 26588
rect -36391 26536 -36389 26588
rect -36389 26536 -36337 26588
rect -36337 26536 -36335 26588
rect -36311 26536 -36273 26588
rect -36273 26536 -36261 26588
rect -36261 26536 -36255 26588
rect -36231 26536 -36209 26588
rect -36209 26536 -36197 26588
rect -36197 26536 -36175 26588
rect -36151 26536 -36145 26588
rect -36145 26536 -36133 26588
rect -36133 26536 -36095 26588
rect -36071 26536 -36069 26588
rect -36069 26536 -36017 26588
rect -36017 26536 -36015 26588
rect -35991 26536 -35953 26588
rect -35953 26536 -35941 26588
rect -35941 26536 -35935 26588
rect -35911 26536 -35889 26588
rect -35889 26536 -35877 26588
rect -35877 26536 -35855 26588
rect -35831 26536 -35825 26588
rect -35825 26536 -35813 26588
rect -35813 26536 -35775 26588
rect -35751 26536 -35749 26588
rect -35749 26536 -35697 26588
rect -35697 26536 -35695 26588
rect -35671 26536 -35633 26588
rect -35633 26536 -35621 26588
rect -35621 26536 -35615 26588
rect -35591 26536 -35569 26588
rect -35569 26536 -35557 26588
rect -35557 26536 -35535 26588
rect -35511 26536 -35505 26588
rect -35505 26536 -35493 26588
rect -35493 26536 -35455 26588
rect -35431 26536 -35429 26588
rect -35429 26536 -35377 26588
rect -35377 26536 -35375 26588
rect -35351 26536 -35313 26588
rect -35313 26536 -35301 26588
rect -35301 26536 -35295 26588
rect -35271 26536 -35249 26588
rect -35249 26536 -35237 26588
rect -35237 26536 -35215 26588
rect -35191 26536 -35185 26588
rect -35185 26536 -35173 26588
rect -35173 26536 -35135 26588
rect -35111 26536 -35109 26588
rect -35109 26536 -35057 26588
rect -35057 26536 -35055 26588
rect -35031 26536 -34993 26588
rect -34993 26536 -34981 26588
rect -34981 26536 -34975 26588
rect -34951 26536 -34929 26588
rect -34929 26536 -34917 26588
rect -34917 26536 -34895 26588
rect -38151 26534 -38095 26536
rect -38071 26534 -38015 26536
rect -37991 26534 -37935 26536
rect -37911 26534 -37855 26536
rect -37831 26534 -37775 26536
rect -37751 26534 -37695 26536
rect -37671 26534 -37615 26536
rect -37591 26534 -37535 26536
rect -37511 26534 -37455 26536
rect -37431 26534 -37375 26536
rect -37351 26534 -37295 26536
rect -37271 26534 -37215 26536
rect -37191 26534 -37135 26536
rect -37111 26534 -37055 26536
rect -37031 26534 -36975 26536
rect -36951 26534 -36895 26536
rect -36871 26534 -36815 26536
rect -36791 26534 -36735 26536
rect -36711 26534 -36655 26536
rect -36631 26534 -36575 26536
rect -36551 26534 -36495 26536
rect -36471 26534 -36415 26536
rect -36391 26534 -36335 26536
rect -36311 26534 -36255 26536
rect -36231 26534 -36175 26536
rect -36151 26534 -36095 26536
rect -36071 26534 -36015 26536
rect -35991 26534 -35935 26536
rect -35911 26534 -35855 26536
rect -35831 26534 -35775 26536
rect -35751 26534 -35695 26536
rect -35671 26534 -35615 26536
rect -35591 26534 -35535 26536
rect -35511 26534 -35455 26536
rect -35431 26534 -35375 26536
rect -35351 26534 -35295 26536
rect -35271 26534 -35215 26536
rect -35191 26534 -35135 26536
rect -35111 26534 -35055 26536
rect -35031 26534 -34975 26536
rect -34951 26534 -34895 26536
rect 4705 28748 4761 28804
rect 7964 28840 8020 28842
rect 7964 28788 7966 28840
rect 7966 28788 8018 28840
rect 8018 28788 8020 28840
rect 7964 28786 8020 28788
rect -15691 28037 -15689 28059
rect -15689 28037 -15637 28059
rect -15637 28037 -15635 28059
rect -15691 28025 -15635 28037
rect -15691 28003 -15689 28025
rect -15689 28003 -15637 28025
rect -15637 28003 -15635 28025
rect -15691 27973 -15689 27979
rect -15689 27973 -15637 27979
rect -15637 27973 -15635 27979
rect -15691 27961 -15635 27973
rect -15691 27923 -15689 27961
rect -15689 27923 -15637 27961
rect -15637 27923 -15635 27961
rect -15691 27897 -15635 27899
rect -15691 27845 -15689 27897
rect -15689 27845 -15637 27897
rect -15637 27845 -15635 27897
rect -15691 27843 -15635 27845
rect -15691 27781 -15689 27819
rect -15689 27781 -15637 27819
rect -15637 27781 -15635 27819
rect -15691 27769 -15635 27781
rect -15691 27763 -15689 27769
rect -15689 27763 -15637 27769
rect -15637 27763 -15635 27769
rect -15691 27717 -15689 27739
rect -15689 27717 -15637 27739
rect -15637 27717 -15635 27739
rect -15691 27705 -15635 27717
rect -15691 27683 -15689 27705
rect -15689 27683 -15637 27705
rect -15637 27683 -15635 27705
rect -17599 27552 -17543 27608
rect -17599 26323 -17543 26379
rect -15709 26252 -15653 26270
rect -15709 26214 -15707 26252
rect -15707 26214 -15655 26252
rect -15655 26214 -15653 26252
rect -15709 26188 -15653 26190
rect -15709 26136 -15707 26188
rect -15707 26136 -15655 26188
rect -15655 26136 -15653 26188
rect -15709 26134 -15653 26136
rect -15709 26072 -15707 26110
rect -15707 26072 -15655 26110
rect -15655 26072 -15653 26110
rect -15709 26054 -15653 26072
rect -12381 28059 -12325 28061
rect -12381 28007 -12379 28059
rect -12379 28007 -12327 28059
rect -12327 28007 -12325 28059
rect -12381 28005 -12325 28007
rect -12381 27943 -12379 27981
rect -12379 27943 -12327 27981
rect -12327 27943 -12325 27981
rect -12381 27931 -12325 27943
rect -12381 27925 -12379 27931
rect -12379 27925 -12327 27931
rect -12327 27925 -12325 27931
rect -12381 27879 -12379 27901
rect -12379 27879 -12327 27901
rect -12327 27879 -12325 27901
rect -12381 27867 -12325 27879
rect -12381 27845 -12379 27867
rect -12379 27845 -12327 27867
rect -12327 27845 -12325 27867
rect -12381 27815 -12379 27821
rect -12379 27815 -12327 27821
rect -12327 27815 -12325 27821
rect -12381 27803 -12325 27815
rect -12381 27765 -12379 27803
rect -12379 27765 -12327 27803
rect -12327 27765 -12325 27803
rect -12381 27739 -12325 27741
rect -12381 27687 -12379 27739
rect -12379 27687 -12327 27739
rect -12327 27687 -12325 27739
rect -12381 27685 -12325 27687
rect -12374 27402 -12318 27420
rect -12374 27364 -12372 27402
rect -12372 27364 -12320 27402
rect -12320 27364 -12318 27402
rect -12374 27338 -12318 27340
rect -12374 27286 -12372 27338
rect -12372 27286 -12320 27338
rect -12320 27286 -12318 27338
rect -12374 27284 -12318 27286
rect -12374 27222 -12372 27260
rect -12372 27222 -12320 27260
rect -12320 27222 -12318 27260
rect -12374 27204 -12318 27222
rect -12377 26457 -12321 26459
rect -12377 26405 -12375 26457
rect -12375 26405 -12323 26457
rect -12323 26405 -12321 26457
rect -12377 26403 -12321 26405
rect -12377 26341 -12375 26379
rect -12375 26341 -12323 26379
rect -12323 26341 -12321 26379
rect -12377 26329 -12321 26341
rect -12377 26323 -12375 26329
rect -12375 26323 -12323 26329
rect -12323 26323 -12321 26329
rect -12377 26277 -12375 26299
rect -12375 26277 -12323 26299
rect -12323 26277 -12321 26299
rect -12377 26265 -12321 26277
rect -12377 26243 -12375 26265
rect -12375 26243 -12323 26265
rect -12323 26243 -12321 26265
rect -12377 26213 -12375 26219
rect -12375 26213 -12323 26219
rect -12323 26213 -12321 26219
rect -12377 26201 -12321 26213
rect -12377 26163 -12375 26201
rect -12375 26163 -12323 26201
rect -12323 26163 -12321 26201
rect -12377 26137 -12321 26139
rect -12377 26085 -12375 26137
rect -12375 26085 -12323 26137
rect -12323 26085 -12321 26137
rect -12377 26083 -12321 26085
rect -12381 25803 -12325 25821
rect -12381 25765 -12379 25803
rect -12379 25765 -12327 25803
rect -12327 25765 -12325 25803
rect -12381 25739 -12325 25741
rect -12381 25687 -12379 25739
rect -12379 25687 -12327 25739
rect -12327 25687 -12325 25739
rect -12381 25685 -12325 25687
rect -25437 25450 -25381 25476
rect -25437 25420 -25435 25450
rect -25435 25420 -25383 25450
rect -25383 25420 -25381 25450
rect -25437 25386 -25381 25396
rect -25437 25340 -25435 25386
rect -25435 25340 -25383 25386
rect -25383 25340 -25381 25386
rect -25437 25270 -25435 25316
rect -25435 25270 -25383 25316
rect -25383 25270 -25381 25316
rect -25437 25260 -25381 25270
rect -25437 25206 -25435 25236
rect -25435 25206 -25383 25236
rect -25383 25206 -25381 25236
rect -25437 25180 -25381 25206
rect -40583 25143 -40367 25161
rect -40583 24963 -40565 25143
rect -40565 24963 -40385 25143
rect -40385 24963 -40367 25143
rect -40583 24945 -40367 24963
rect -38145 23580 -38089 23582
rect -38065 23580 -38009 23582
rect -37985 23580 -37929 23582
rect -37905 23580 -37849 23582
rect -37825 23580 -37769 23582
rect -37745 23580 -37689 23582
rect -37665 23580 -37609 23582
rect -37585 23580 -37529 23582
rect -37505 23580 -37449 23582
rect -37425 23580 -37369 23582
rect -37345 23580 -37289 23582
rect -37265 23580 -37209 23582
rect -37185 23580 -37129 23582
rect -37105 23580 -37049 23582
rect -37025 23580 -36969 23582
rect -36945 23580 -36889 23582
rect -36865 23580 -36809 23582
rect -36785 23580 -36729 23582
rect -36705 23580 -36649 23582
rect -36625 23580 -36569 23582
rect -36545 23580 -36489 23582
rect -36465 23580 -36409 23582
rect -36385 23580 -36329 23582
rect -36305 23580 -36249 23582
rect -36225 23580 -36169 23582
rect -36145 23580 -36089 23582
rect -36065 23580 -36009 23582
rect -35985 23580 -35929 23582
rect -35905 23580 -35849 23582
rect -35825 23580 -35769 23582
rect -35745 23580 -35689 23582
rect -35665 23580 -35609 23582
rect -35585 23580 -35529 23582
rect -35505 23580 -35449 23582
rect -35425 23580 -35369 23582
rect -35345 23580 -35289 23582
rect -35265 23580 -35209 23582
rect -35185 23580 -35129 23582
rect -35105 23580 -35049 23582
rect -35025 23580 -34969 23582
rect -34945 23580 -34889 23582
rect -38145 23528 -38123 23580
rect -38123 23528 -38111 23580
rect -38111 23528 -38089 23580
rect -38065 23528 -38059 23580
rect -38059 23528 -38047 23580
rect -38047 23528 -38009 23580
rect -37985 23528 -37983 23580
rect -37983 23528 -37931 23580
rect -37931 23528 -37929 23580
rect -37905 23528 -37867 23580
rect -37867 23528 -37855 23580
rect -37855 23528 -37849 23580
rect -37825 23528 -37803 23580
rect -37803 23528 -37791 23580
rect -37791 23528 -37769 23580
rect -37745 23528 -37739 23580
rect -37739 23528 -37727 23580
rect -37727 23528 -37689 23580
rect -37665 23528 -37663 23580
rect -37663 23528 -37611 23580
rect -37611 23528 -37609 23580
rect -37585 23528 -37547 23580
rect -37547 23528 -37535 23580
rect -37535 23528 -37529 23580
rect -37505 23528 -37483 23580
rect -37483 23528 -37471 23580
rect -37471 23528 -37449 23580
rect -37425 23528 -37419 23580
rect -37419 23528 -37407 23580
rect -37407 23528 -37369 23580
rect -37345 23528 -37343 23580
rect -37343 23528 -37291 23580
rect -37291 23528 -37289 23580
rect -37265 23528 -37227 23580
rect -37227 23528 -37215 23580
rect -37215 23528 -37209 23580
rect -37185 23528 -37163 23580
rect -37163 23528 -37151 23580
rect -37151 23528 -37129 23580
rect -37105 23528 -37099 23580
rect -37099 23528 -37087 23580
rect -37087 23528 -37049 23580
rect -37025 23528 -37023 23580
rect -37023 23528 -36971 23580
rect -36971 23528 -36969 23580
rect -36945 23528 -36907 23580
rect -36907 23528 -36895 23580
rect -36895 23528 -36889 23580
rect -36865 23528 -36843 23580
rect -36843 23528 -36831 23580
rect -36831 23528 -36809 23580
rect -36785 23528 -36779 23580
rect -36779 23528 -36767 23580
rect -36767 23528 -36729 23580
rect -36705 23528 -36703 23580
rect -36703 23528 -36651 23580
rect -36651 23528 -36649 23580
rect -36625 23528 -36587 23580
rect -36587 23528 -36575 23580
rect -36575 23528 -36569 23580
rect -36545 23528 -36523 23580
rect -36523 23528 -36511 23580
rect -36511 23528 -36489 23580
rect -36465 23528 -36459 23580
rect -36459 23528 -36447 23580
rect -36447 23528 -36409 23580
rect -36385 23528 -36383 23580
rect -36383 23528 -36331 23580
rect -36331 23528 -36329 23580
rect -36305 23528 -36267 23580
rect -36267 23528 -36255 23580
rect -36255 23528 -36249 23580
rect -36225 23528 -36203 23580
rect -36203 23528 -36191 23580
rect -36191 23528 -36169 23580
rect -36145 23528 -36139 23580
rect -36139 23528 -36127 23580
rect -36127 23528 -36089 23580
rect -36065 23528 -36063 23580
rect -36063 23528 -36011 23580
rect -36011 23528 -36009 23580
rect -35985 23528 -35947 23580
rect -35947 23528 -35935 23580
rect -35935 23528 -35929 23580
rect -35905 23528 -35883 23580
rect -35883 23528 -35871 23580
rect -35871 23528 -35849 23580
rect -35825 23528 -35819 23580
rect -35819 23528 -35807 23580
rect -35807 23528 -35769 23580
rect -35745 23528 -35743 23580
rect -35743 23528 -35691 23580
rect -35691 23528 -35689 23580
rect -35665 23528 -35627 23580
rect -35627 23528 -35615 23580
rect -35615 23528 -35609 23580
rect -35585 23528 -35563 23580
rect -35563 23528 -35551 23580
rect -35551 23528 -35529 23580
rect -35505 23528 -35499 23580
rect -35499 23528 -35487 23580
rect -35487 23528 -35449 23580
rect -35425 23528 -35423 23580
rect -35423 23528 -35371 23580
rect -35371 23528 -35369 23580
rect -35345 23528 -35307 23580
rect -35307 23528 -35295 23580
rect -35295 23528 -35289 23580
rect -35265 23528 -35243 23580
rect -35243 23528 -35231 23580
rect -35231 23528 -35209 23580
rect -35185 23528 -35179 23580
rect -35179 23528 -35167 23580
rect -35167 23528 -35129 23580
rect -35105 23528 -35103 23580
rect -35103 23528 -35051 23580
rect -35051 23528 -35049 23580
rect -35025 23528 -34987 23580
rect -34987 23528 -34975 23580
rect -34975 23528 -34969 23580
rect -34945 23528 -34923 23580
rect -34923 23528 -34911 23580
rect -34911 23528 -34889 23580
rect -38145 23526 -38089 23528
rect -38065 23526 -38009 23528
rect -37985 23526 -37929 23528
rect -37905 23526 -37849 23528
rect -37825 23526 -37769 23528
rect -37745 23526 -37689 23528
rect -37665 23526 -37609 23528
rect -37585 23526 -37529 23528
rect -37505 23526 -37449 23528
rect -37425 23526 -37369 23528
rect -37345 23526 -37289 23528
rect -37265 23526 -37209 23528
rect -37185 23526 -37129 23528
rect -37105 23526 -37049 23528
rect -37025 23526 -36969 23528
rect -36945 23526 -36889 23528
rect -36865 23526 -36809 23528
rect -36785 23526 -36729 23528
rect -36705 23526 -36649 23528
rect -36625 23526 -36569 23528
rect -36545 23526 -36489 23528
rect -36465 23526 -36409 23528
rect -36385 23526 -36329 23528
rect -36305 23526 -36249 23528
rect -36225 23526 -36169 23528
rect -36145 23526 -36089 23528
rect -36065 23526 -36009 23528
rect -35985 23526 -35929 23528
rect -35905 23526 -35849 23528
rect -35825 23526 -35769 23528
rect -35745 23526 -35689 23528
rect -35665 23526 -35609 23528
rect -35585 23526 -35529 23528
rect -35505 23526 -35449 23528
rect -35425 23526 -35369 23528
rect -35345 23526 -35289 23528
rect -35265 23526 -35209 23528
rect -35185 23526 -35129 23528
rect -35105 23526 -35049 23528
rect -35025 23526 -34969 23528
rect -34945 23526 -34889 23528
rect -38143 19052 -38087 19054
rect -38063 19052 -38007 19054
rect -37983 19052 -37927 19054
rect -37903 19052 -37847 19054
rect -37823 19052 -37767 19054
rect -37743 19052 -37687 19054
rect -37663 19052 -37607 19054
rect -37583 19052 -37527 19054
rect -37503 19052 -37447 19054
rect -37423 19052 -37367 19054
rect -37343 19052 -37287 19054
rect -37263 19052 -37207 19054
rect -37183 19052 -37127 19054
rect -37103 19052 -37047 19054
rect -37023 19052 -36967 19054
rect -36943 19052 -36887 19054
rect -36863 19052 -36807 19054
rect -36783 19052 -36727 19054
rect -36703 19052 -36647 19054
rect -36623 19052 -36567 19054
rect -36543 19052 -36487 19054
rect -36463 19052 -36407 19054
rect -36383 19052 -36327 19054
rect -36303 19052 -36247 19054
rect -36223 19052 -36167 19054
rect -36143 19052 -36087 19054
rect -36063 19052 -36007 19054
rect -35983 19052 -35927 19054
rect -35903 19052 -35847 19054
rect -35823 19052 -35767 19054
rect -35743 19052 -35687 19054
rect -35663 19052 -35607 19054
rect -35583 19052 -35527 19054
rect -35503 19052 -35447 19054
rect -35423 19052 -35367 19054
rect -35343 19052 -35287 19054
rect -35263 19052 -35207 19054
rect -35183 19052 -35127 19054
rect -35103 19052 -35047 19054
rect -35023 19052 -34967 19054
rect -34943 19052 -34887 19054
rect -38143 19000 -38141 19052
rect -38141 19000 -38089 19052
rect -38089 19000 -38087 19052
rect -38063 19000 -38025 19052
rect -38025 19000 -38013 19052
rect -38013 19000 -38007 19052
rect -37983 19000 -37961 19052
rect -37961 19000 -37949 19052
rect -37949 19000 -37927 19052
rect -37903 19000 -37897 19052
rect -37897 19000 -37885 19052
rect -37885 19000 -37847 19052
rect -37823 19000 -37821 19052
rect -37821 19000 -37769 19052
rect -37769 19000 -37767 19052
rect -37743 19000 -37705 19052
rect -37705 19000 -37693 19052
rect -37693 19000 -37687 19052
rect -37663 19000 -37641 19052
rect -37641 19000 -37629 19052
rect -37629 19000 -37607 19052
rect -37583 19000 -37577 19052
rect -37577 19000 -37565 19052
rect -37565 19000 -37527 19052
rect -37503 19000 -37501 19052
rect -37501 19000 -37449 19052
rect -37449 19000 -37447 19052
rect -37423 19000 -37385 19052
rect -37385 19000 -37373 19052
rect -37373 19000 -37367 19052
rect -37343 19000 -37321 19052
rect -37321 19000 -37309 19052
rect -37309 19000 -37287 19052
rect -37263 19000 -37257 19052
rect -37257 19000 -37245 19052
rect -37245 19000 -37207 19052
rect -37183 19000 -37181 19052
rect -37181 19000 -37129 19052
rect -37129 19000 -37127 19052
rect -37103 19000 -37065 19052
rect -37065 19000 -37053 19052
rect -37053 19000 -37047 19052
rect -37023 19000 -37001 19052
rect -37001 19000 -36989 19052
rect -36989 19000 -36967 19052
rect -36943 19000 -36937 19052
rect -36937 19000 -36925 19052
rect -36925 19000 -36887 19052
rect -36863 19000 -36861 19052
rect -36861 19000 -36809 19052
rect -36809 19000 -36807 19052
rect -36783 19000 -36745 19052
rect -36745 19000 -36733 19052
rect -36733 19000 -36727 19052
rect -36703 19000 -36681 19052
rect -36681 19000 -36669 19052
rect -36669 19000 -36647 19052
rect -36623 19000 -36617 19052
rect -36617 19000 -36605 19052
rect -36605 19000 -36567 19052
rect -36543 19000 -36541 19052
rect -36541 19000 -36489 19052
rect -36489 19000 -36487 19052
rect -36463 19000 -36425 19052
rect -36425 19000 -36413 19052
rect -36413 19000 -36407 19052
rect -36383 19000 -36361 19052
rect -36361 19000 -36349 19052
rect -36349 19000 -36327 19052
rect -36303 19000 -36297 19052
rect -36297 19000 -36285 19052
rect -36285 19000 -36247 19052
rect -36223 19000 -36221 19052
rect -36221 19000 -36169 19052
rect -36169 19000 -36167 19052
rect -36143 19000 -36105 19052
rect -36105 19000 -36093 19052
rect -36093 19000 -36087 19052
rect -36063 19000 -36041 19052
rect -36041 19000 -36029 19052
rect -36029 19000 -36007 19052
rect -35983 19000 -35977 19052
rect -35977 19000 -35965 19052
rect -35965 19000 -35927 19052
rect -35903 19000 -35901 19052
rect -35901 19000 -35849 19052
rect -35849 19000 -35847 19052
rect -35823 19000 -35785 19052
rect -35785 19000 -35773 19052
rect -35773 19000 -35767 19052
rect -35743 19000 -35721 19052
rect -35721 19000 -35709 19052
rect -35709 19000 -35687 19052
rect -35663 19000 -35657 19052
rect -35657 19000 -35645 19052
rect -35645 19000 -35607 19052
rect -35583 19000 -35581 19052
rect -35581 19000 -35529 19052
rect -35529 19000 -35527 19052
rect -35503 19000 -35465 19052
rect -35465 19000 -35453 19052
rect -35453 19000 -35447 19052
rect -35423 19000 -35401 19052
rect -35401 19000 -35389 19052
rect -35389 19000 -35367 19052
rect -35343 19000 -35337 19052
rect -35337 19000 -35325 19052
rect -35325 19000 -35287 19052
rect -35263 19000 -35261 19052
rect -35261 19000 -35209 19052
rect -35209 19000 -35207 19052
rect -35183 19000 -35145 19052
rect -35145 19000 -35133 19052
rect -35133 19000 -35127 19052
rect -35103 19000 -35081 19052
rect -35081 19000 -35069 19052
rect -35069 19000 -35047 19052
rect -35023 19000 -35017 19052
rect -35017 19000 -35005 19052
rect -35005 19000 -34967 19052
rect -34943 19000 -34941 19052
rect -34941 19000 -34889 19052
rect -34889 19000 -34887 19052
rect -38143 18998 -38087 19000
rect -38063 18998 -38007 19000
rect -37983 18998 -37927 19000
rect -37903 18998 -37847 19000
rect -37823 18998 -37767 19000
rect -37743 18998 -37687 19000
rect -37663 18998 -37607 19000
rect -37583 18998 -37527 19000
rect -37503 18998 -37447 19000
rect -37423 18998 -37367 19000
rect -37343 18998 -37287 19000
rect -37263 18998 -37207 19000
rect -37183 18998 -37127 19000
rect -37103 18998 -37047 19000
rect -37023 18998 -36967 19000
rect -36943 18998 -36887 19000
rect -36863 18998 -36807 19000
rect -36783 18998 -36727 19000
rect -36703 18998 -36647 19000
rect -36623 18998 -36567 19000
rect -36543 18998 -36487 19000
rect -36463 18998 -36407 19000
rect -36383 18998 -36327 19000
rect -36303 18998 -36247 19000
rect -36223 18998 -36167 19000
rect -36143 18998 -36087 19000
rect -36063 18998 -36007 19000
rect -35983 18998 -35927 19000
rect -35903 18998 -35847 19000
rect -35823 18998 -35767 19000
rect -35743 18998 -35687 19000
rect -35663 18998 -35607 19000
rect -35583 18998 -35527 19000
rect -35503 18998 -35447 19000
rect -35423 18998 -35367 19000
rect -35343 18998 -35287 19000
rect -35263 18998 -35207 19000
rect -35183 18998 -35127 19000
rect -35103 18998 -35047 19000
rect -35023 18998 -34967 19000
rect -34943 18998 -34887 19000
rect -40586 17602 -40370 17620
rect -40586 17422 -40568 17602
rect -40568 17422 -40388 17602
rect -40388 17422 -40370 17602
rect -40586 17404 -40370 17422
rect -38141 16057 -38085 16059
rect -38061 16057 -38005 16059
rect -37981 16057 -37925 16059
rect -37901 16057 -37845 16059
rect -37821 16057 -37765 16059
rect -37741 16057 -37685 16059
rect -37661 16057 -37605 16059
rect -37581 16057 -37525 16059
rect -37501 16057 -37445 16059
rect -37421 16057 -37365 16059
rect -37341 16057 -37285 16059
rect -37261 16057 -37205 16059
rect -37181 16057 -37125 16059
rect -37101 16057 -37045 16059
rect -37021 16057 -36965 16059
rect -36941 16057 -36885 16059
rect -36861 16057 -36805 16059
rect -36781 16057 -36725 16059
rect -36701 16057 -36645 16059
rect -36621 16057 -36565 16059
rect -36541 16057 -36485 16059
rect -36461 16057 -36405 16059
rect -36381 16057 -36325 16059
rect -36301 16057 -36245 16059
rect -36221 16057 -36165 16059
rect -36141 16057 -36085 16059
rect -36061 16057 -36005 16059
rect -35981 16057 -35925 16059
rect -35901 16057 -35845 16059
rect -35821 16057 -35765 16059
rect -35741 16057 -35685 16059
rect -35661 16057 -35605 16059
rect -35581 16057 -35525 16059
rect -35501 16057 -35445 16059
rect -35421 16057 -35365 16059
rect -35341 16057 -35285 16059
rect -35261 16057 -35205 16059
rect -35181 16057 -35125 16059
rect -35101 16057 -35045 16059
rect -35021 16057 -34965 16059
rect -34941 16057 -34885 16059
rect -38141 16005 -38119 16057
rect -38119 16005 -38107 16057
rect -38107 16005 -38085 16057
rect -38061 16005 -38055 16057
rect -38055 16005 -38043 16057
rect -38043 16005 -38005 16057
rect -37981 16005 -37979 16057
rect -37979 16005 -37927 16057
rect -37927 16005 -37925 16057
rect -37901 16005 -37863 16057
rect -37863 16005 -37851 16057
rect -37851 16005 -37845 16057
rect -37821 16005 -37799 16057
rect -37799 16005 -37787 16057
rect -37787 16005 -37765 16057
rect -37741 16005 -37735 16057
rect -37735 16005 -37723 16057
rect -37723 16005 -37685 16057
rect -37661 16005 -37659 16057
rect -37659 16005 -37607 16057
rect -37607 16005 -37605 16057
rect -37581 16005 -37543 16057
rect -37543 16005 -37531 16057
rect -37531 16005 -37525 16057
rect -37501 16005 -37479 16057
rect -37479 16005 -37467 16057
rect -37467 16005 -37445 16057
rect -37421 16005 -37415 16057
rect -37415 16005 -37403 16057
rect -37403 16005 -37365 16057
rect -37341 16005 -37339 16057
rect -37339 16005 -37287 16057
rect -37287 16005 -37285 16057
rect -37261 16005 -37223 16057
rect -37223 16005 -37211 16057
rect -37211 16005 -37205 16057
rect -37181 16005 -37159 16057
rect -37159 16005 -37147 16057
rect -37147 16005 -37125 16057
rect -37101 16005 -37095 16057
rect -37095 16005 -37083 16057
rect -37083 16005 -37045 16057
rect -37021 16005 -37019 16057
rect -37019 16005 -36967 16057
rect -36967 16005 -36965 16057
rect -36941 16005 -36903 16057
rect -36903 16005 -36891 16057
rect -36891 16005 -36885 16057
rect -36861 16005 -36839 16057
rect -36839 16005 -36827 16057
rect -36827 16005 -36805 16057
rect -36781 16005 -36775 16057
rect -36775 16005 -36763 16057
rect -36763 16005 -36725 16057
rect -36701 16005 -36699 16057
rect -36699 16005 -36647 16057
rect -36647 16005 -36645 16057
rect -36621 16005 -36583 16057
rect -36583 16005 -36571 16057
rect -36571 16005 -36565 16057
rect -36541 16005 -36519 16057
rect -36519 16005 -36507 16057
rect -36507 16005 -36485 16057
rect -36461 16005 -36455 16057
rect -36455 16005 -36443 16057
rect -36443 16005 -36405 16057
rect -36381 16005 -36379 16057
rect -36379 16005 -36327 16057
rect -36327 16005 -36325 16057
rect -36301 16005 -36263 16057
rect -36263 16005 -36251 16057
rect -36251 16005 -36245 16057
rect -36221 16005 -36199 16057
rect -36199 16005 -36187 16057
rect -36187 16005 -36165 16057
rect -36141 16005 -36135 16057
rect -36135 16005 -36123 16057
rect -36123 16005 -36085 16057
rect -36061 16005 -36059 16057
rect -36059 16005 -36007 16057
rect -36007 16005 -36005 16057
rect -35981 16005 -35943 16057
rect -35943 16005 -35931 16057
rect -35931 16005 -35925 16057
rect -35901 16005 -35879 16057
rect -35879 16005 -35867 16057
rect -35867 16005 -35845 16057
rect -35821 16005 -35815 16057
rect -35815 16005 -35803 16057
rect -35803 16005 -35765 16057
rect -35741 16005 -35739 16057
rect -35739 16005 -35687 16057
rect -35687 16005 -35685 16057
rect -35661 16005 -35623 16057
rect -35623 16005 -35611 16057
rect -35611 16005 -35605 16057
rect -35581 16005 -35559 16057
rect -35559 16005 -35547 16057
rect -35547 16005 -35525 16057
rect -35501 16005 -35495 16057
rect -35495 16005 -35483 16057
rect -35483 16005 -35445 16057
rect -35421 16005 -35419 16057
rect -35419 16005 -35367 16057
rect -35367 16005 -35365 16057
rect -35341 16005 -35303 16057
rect -35303 16005 -35291 16057
rect -35291 16005 -35285 16057
rect -35261 16005 -35239 16057
rect -35239 16005 -35227 16057
rect -35227 16005 -35205 16057
rect -35181 16005 -35175 16057
rect -35175 16005 -35163 16057
rect -35163 16005 -35125 16057
rect -35101 16005 -35099 16057
rect -35099 16005 -35047 16057
rect -35047 16005 -35045 16057
rect -35021 16005 -34983 16057
rect -34983 16005 -34971 16057
rect -34971 16005 -34965 16057
rect -34941 16005 -34919 16057
rect -34919 16005 -34907 16057
rect -34907 16005 -34885 16057
rect -38141 16003 -38085 16005
rect -38061 16003 -38005 16005
rect -37981 16003 -37925 16005
rect -37901 16003 -37845 16005
rect -37821 16003 -37765 16005
rect -37741 16003 -37685 16005
rect -37661 16003 -37605 16005
rect -37581 16003 -37525 16005
rect -37501 16003 -37445 16005
rect -37421 16003 -37365 16005
rect -37341 16003 -37285 16005
rect -37261 16003 -37205 16005
rect -37181 16003 -37125 16005
rect -37101 16003 -37045 16005
rect -37021 16003 -36965 16005
rect -36941 16003 -36885 16005
rect -36861 16003 -36805 16005
rect -36781 16003 -36725 16005
rect -36701 16003 -36645 16005
rect -36621 16003 -36565 16005
rect -36541 16003 -36485 16005
rect -36461 16003 -36405 16005
rect -36381 16003 -36325 16005
rect -36301 16003 -36245 16005
rect -36221 16003 -36165 16005
rect -36141 16003 -36085 16005
rect -36061 16003 -36005 16005
rect -35981 16003 -35925 16005
rect -35901 16003 -35845 16005
rect -35821 16003 -35765 16005
rect -35741 16003 -35685 16005
rect -35661 16003 -35605 16005
rect -35581 16003 -35525 16005
rect -35501 16003 -35445 16005
rect -35421 16003 -35365 16005
rect -35341 16003 -35285 16005
rect -35261 16003 -35205 16005
rect -35181 16003 -35125 16005
rect -35101 16003 -35045 16005
rect -35021 16003 -34965 16005
rect -34941 16003 -34885 16005
rect -25437 24919 -25381 24937
rect -25437 24881 -25435 24919
rect -25435 24881 -25383 24919
rect -25383 24881 -25381 24919
rect -25437 24855 -25381 24857
rect -25437 24803 -25435 24855
rect -25435 24803 -25383 24855
rect -25383 24803 -25381 24855
rect -25437 24801 -25381 24803
rect -25437 24739 -25435 24777
rect -25435 24739 -25383 24777
rect -25383 24739 -25381 24777
rect -25437 24721 -25381 24739
rect -15708 25418 -15652 25420
rect -15708 25366 -15706 25418
rect -15706 25366 -15654 25418
rect -15654 25366 -15652 25418
rect -15708 25364 -15652 25366
rect -15708 25302 -15706 25340
rect -15706 25302 -15654 25340
rect -15654 25302 -15652 25340
rect -15708 25290 -15652 25302
rect -15708 25284 -15706 25290
rect -15706 25284 -15654 25290
rect -15654 25284 -15652 25290
rect -15708 25238 -15706 25260
rect -15706 25238 -15654 25260
rect -15654 25238 -15652 25260
rect -15708 25226 -15652 25238
rect -15708 25204 -15706 25226
rect -15706 25204 -15654 25226
rect -15654 25204 -15652 25226
rect -15708 25174 -15706 25180
rect -15706 25174 -15654 25180
rect -15654 25174 -15652 25180
rect -15708 25162 -15652 25174
rect -15708 25124 -15706 25162
rect -15706 25124 -15654 25162
rect -15654 25124 -15652 25162
rect -15708 25098 -15652 25100
rect -15708 25046 -15706 25098
rect -15706 25046 -15654 25098
rect -15654 25046 -15652 25098
rect -15708 25044 -15652 25046
rect -17599 24910 -17543 24966
rect -13985 25604 -13929 25660
rect -12381 25623 -12379 25661
rect -12379 25623 -12327 25661
rect -12327 25623 -12325 25661
rect -12381 25605 -12325 25623
rect -14406 24812 -14350 24868
rect -17599 23681 -17543 23737
rect -15720 23611 -15664 23629
rect -15720 23573 -15718 23611
rect -15718 23573 -15666 23611
rect -15666 23573 -15664 23611
rect -15720 23547 -15664 23549
rect -15720 23495 -15718 23547
rect -15718 23495 -15666 23547
rect -15666 23495 -15664 23547
rect -15720 23493 -15664 23495
rect -15720 23431 -15718 23469
rect -15718 23431 -15666 23469
rect -15666 23431 -15664 23469
rect -15720 23413 -15664 23431
rect -12389 24655 -12387 24693
rect -12387 24655 -12335 24693
rect -12335 24655 -12333 24693
rect -12389 24643 -12333 24655
rect -12389 24637 -12387 24643
rect -12387 24637 -12335 24643
rect -12335 24637 -12333 24643
rect -12389 24591 -12387 24613
rect -12387 24591 -12335 24613
rect -12335 24591 -12333 24613
rect -12389 24579 -12333 24591
rect -12389 24557 -12387 24579
rect -12387 24557 -12335 24579
rect -12335 24557 -12333 24579
rect -12389 24527 -12387 24533
rect -12387 24527 -12335 24533
rect -12335 24527 -12333 24533
rect -12389 24515 -12333 24527
rect -12389 24477 -12387 24515
rect -12387 24477 -12335 24515
rect -12335 24477 -12333 24515
rect -12385 24211 -12329 24229
rect -12385 24173 -12383 24211
rect -12383 24173 -12331 24211
rect -12331 24173 -12329 24211
rect -12385 24147 -12329 24149
rect -12385 24095 -12383 24147
rect -12383 24095 -12331 24147
rect -12331 24095 -12329 24147
rect -12385 24093 -12329 24095
rect -12385 24031 -12383 24069
rect -12383 24031 -12331 24069
rect -12331 24031 -12329 24069
rect -12385 24013 -12329 24031
rect -12382 23253 -12326 23255
rect -12382 23201 -12380 23253
rect -12380 23201 -12328 23253
rect -12328 23201 -12326 23253
rect -12382 23199 -12326 23201
rect -12382 23137 -12380 23175
rect -12380 23137 -12328 23175
rect -12328 23137 -12326 23175
rect -12382 23125 -12326 23137
rect -12382 23119 -12380 23125
rect -12380 23119 -12328 23125
rect -12328 23119 -12326 23125
rect -12382 23073 -12380 23095
rect -12380 23073 -12328 23095
rect -12328 23073 -12326 23095
rect -12382 23061 -12326 23073
rect -12382 23039 -12380 23061
rect -12380 23039 -12328 23061
rect -12328 23039 -12326 23061
rect -12382 23009 -12380 23015
rect -12380 23009 -12328 23015
rect -12328 23009 -12326 23015
rect -12382 22997 -12326 23009
rect -12382 22959 -12380 22997
rect -12380 22959 -12328 22997
rect -12328 22959 -12326 22997
rect -12382 22933 -12326 22935
rect -12382 22881 -12380 22933
rect -12380 22881 -12328 22933
rect -12328 22881 -12326 22933
rect -12382 22879 -12326 22881
rect -12385 22601 -12329 22619
rect -12385 22563 -12383 22601
rect -12383 22563 -12331 22601
rect -12331 22563 -12329 22601
rect -12385 22537 -12329 22539
rect -12385 22485 -12383 22537
rect -12383 22485 -12331 22537
rect -12331 22485 -12329 22537
rect -12385 22483 -12329 22485
rect -12385 22421 -12383 22459
rect -12383 22421 -12331 22459
rect -12331 22421 -12329 22459
rect -12385 22403 -12329 22421
rect -25448 17844 -25446 17882
rect -25446 17844 -25394 17882
rect -25394 17844 -25392 17882
rect -25448 17832 -25392 17844
rect -25448 17826 -25446 17832
rect -25446 17826 -25394 17832
rect -25394 17826 -25392 17832
rect -25448 17780 -25446 17802
rect -25446 17780 -25394 17802
rect -25394 17780 -25392 17802
rect -25448 17768 -25392 17780
rect -25448 17746 -25446 17768
rect -25446 17746 -25394 17768
rect -25394 17746 -25392 17768
rect -25448 17716 -25446 17722
rect -25446 17716 -25394 17722
rect -25394 17716 -25392 17722
rect -25448 17704 -25392 17716
rect -25448 17666 -25446 17704
rect -25446 17666 -25394 17704
rect -25394 17666 -25392 17704
rect -25442 17376 -25386 17394
rect -25442 17338 -25440 17376
rect -25440 17338 -25388 17376
rect -25388 17338 -25386 17376
rect -25442 17312 -25386 17314
rect -25442 17260 -25440 17312
rect -25440 17260 -25388 17312
rect -25388 17260 -25386 17312
rect -25442 17258 -25386 17260
rect -25442 17196 -25440 17234
rect -25440 17196 -25388 17234
rect -25388 17196 -25386 17234
rect -25442 17178 -25386 17196
rect -24166 16189 -24110 16245
rect -27916 15381 -27860 15437
rect -25509 14371 -25507 14409
rect -25507 14371 -25455 14409
rect -25455 14371 -25453 14409
rect -25509 14359 -25453 14371
rect -25509 14353 -25507 14359
rect -25507 14353 -25455 14359
rect -25455 14353 -25453 14359
rect -25509 14307 -25507 14329
rect -25507 14307 -25455 14329
rect -25455 14307 -25453 14329
rect -25509 14295 -25453 14307
rect -25509 14273 -25507 14295
rect -25507 14273 -25455 14295
rect -25455 14273 -25453 14295
rect -25509 14243 -25507 14249
rect -25507 14243 -25455 14249
rect -25455 14243 -25453 14249
rect -25509 14231 -25453 14243
rect -25509 14193 -25507 14231
rect -25507 14193 -25455 14231
rect -25455 14193 -25453 14231
rect -25510 13897 -25454 13915
rect -25510 13859 -25508 13897
rect -25508 13859 -25456 13897
rect -25456 13859 -25454 13897
rect -25510 13833 -25454 13835
rect -25510 13781 -25508 13833
rect -25508 13781 -25456 13833
rect -25456 13781 -25454 13833
rect -25510 13779 -25454 13781
rect -25510 13717 -25508 13755
rect -25508 13717 -25456 13755
rect -25456 13717 -25454 13755
rect -25510 13699 -25454 13717
rect -18219 14067 -18163 14069
rect -18219 14015 -18217 14067
rect -18217 14015 -18165 14067
rect -18165 14015 -18163 14067
rect -18219 14013 -18163 14015
rect 4332 28535 4388 28591
rect 8342 28532 8398 28588
rect -5275 27472 -5219 27528
rect -3914 26795 -3858 26851
rect 19875 25949 19931 26005
rect 19877 25538 19933 25594
rect 5721 24576 5777 24578
rect 5721 24524 5723 24576
rect 5723 24524 5775 24576
rect 5775 24524 5777 24576
rect 5721 24522 5777 24524
rect 7072 24532 7128 24588
rect 5721 24460 5723 24498
rect 5723 24460 5775 24498
rect 5775 24460 5777 24498
rect 5721 24448 5777 24460
rect 5721 24442 5723 24448
rect 5723 24442 5775 24448
rect 5775 24442 5777 24448
rect 5721 24396 5723 24418
rect 5723 24396 5775 24418
rect 5775 24396 5777 24418
rect 5721 24384 5777 24396
rect 5721 24362 5723 24384
rect 5723 24362 5775 24384
rect 5775 24362 5777 24384
rect 5721 24332 5723 24338
rect 5723 24332 5775 24338
rect 5775 24332 5777 24338
rect 5721 24320 5777 24332
rect 5721 24282 5723 24320
rect 5723 24282 5775 24320
rect 5775 24282 5777 24320
rect 5721 24256 5777 24258
rect 5721 24204 5723 24256
rect 5723 24204 5775 24256
rect 5775 24204 5777 24256
rect 5721 24202 5777 24204
rect 42895 24145 42951 24147
rect 42975 24145 43031 24147
rect 43055 24145 43111 24147
rect 43135 24145 43191 24147
rect 43215 24145 43271 24147
rect 43295 24145 43351 24147
rect 43375 24145 43431 24147
rect 43455 24145 43511 24147
rect 43535 24145 43591 24147
rect 43615 24145 43671 24147
rect 43695 24145 43751 24147
rect 43775 24145 43831 24147
rect 43855 24145 43911 24147
rect 43935 24145 43991 24147
rect 44015 24145 44071 24147
rect 44095 24145 44151 24147
rect 44175 24145 44231 24147
rect 44255 24145 44311 24147
rect 44335 24145 44391 24147
rect 44415 24145 44471 24147
rect 44495 24145 44551 24147
rect 44575 24145 44631 24147
rect 44655 24145 44711 24147
rect 44735 24145 44791 24147
rect 44815 24145 44871 24147
rect 44895 24145 44951 24147
rect 44975 24145 45031 24147
rect 45055 24145 45111 24147
rect 45135 24145 45191 24147
rect 45215 24145 45271 24147
rect 45295 24145 45351 24147
rect 45375 24145 45431 24147
rect 45455 24145 45511 24147
rect 45535 24145 45591 24147
rect 45615 24145 45671 24147
rect 45695 24145 45751 24147
rect 45775 24145 45831 24147
rect 45855 24145 45911 24147
rect 45935 24145 45991 24147
rect 46015 24145 46071 24147
rect 46095 24145 46151 24147
rect 42895 24093 42917 24145
rect 42917 24093 42929 24145
rect 42929 24093 42951 24145
rect 42975 24093 42981 24145
rect 42981 24093 42993 24145
rect 42993 24093 43031 24145
rect 43055 24093 43057 24145
rect 43057 24093 43109 24145
rect 43109 24093 43111 24145
rect 43135 24093 43173 24145
rect 43173 24093 43185 24145
rect 43185 24093 43191 24145
rect 43215 24093 43237 24145
rect 43237 24093 43249 24145
rect 43249 24093 43271 24145
rect 43295 24093 43301 24145
rect 43301 24093 43313 24145
rect 43313 24093 43351 24145
rect 43375 24093 43377 24145
rect 43377 24093 43429 24145
rect 43429 24093 43431 24145
rect 43455 24093 43493 24145
rect 43493 24093 43505 24145
rect 43505 24093 43511 24145
rect 43535 24093 43557 24145
rect 43557 24093 43569 24145
rect 43569 24093 43591 24145
rect 43615 24093 43621 24145
rect 43621 24093 43633 24145
rect 43633 24093 43671 24145
rect 43695 24093 43697 24145
rect 43697 24093 43749 24145
rect 43749 24093 43751 24145
rect 43775 24093 43813 24145
rect 43813 24093 43825 24145
rect 43825 24093 43831 24145
rect 43855 24093 43877 24145
rect 43877 24093 43889 24145
rect 43889 24093 43911 24145
rect 43935 24093 43941 24145
rect 43941 24093 43953 24145
rect 43953 24093 43991 24145
rect 44015 24093 44017 24145
rect 44017 24093 44069 24145
rect 44069 24093 44071 24145
rect 44095 24093 44133 24145
rect 44133 24093 44145 24145
rect 44145 24093 44151 24145
rect 44175 24093 44197 24145
rect 44197 24093 44209 24145
rect 44209 24093 44231 24145
rect 44255 24093 44261 24145
rect 44261 24093 44273 24145
rect 44273 24093 44311 24145
rect 44335 24093 44337 24145
rect 44337 24093 44389 24145
rect 44389 24093 44391 24145
rect 44415 24093 44453 24145
rect 44453 24093 44465 24145
rect 44465 24093 44471 24145
rect 44495 24093 44517 24145
rect 44517 24093 44529 24145
rect 44529 24093 44551 24145
rect 44575 24093 44581 24145
rect 44581 24093 44593 24145
rect 44593 24093 44631 24145
rect 44655 24093 44657 24145
rect 44657 24093 44709 24145
rect 44709 24093 44711 24145
rect 44735 24093 44773 24145
rect 44773 24093 44785 24145
rect 44785 24093 44791 24145
rect 44815 24093 44837 24145
rect 44837 24093 44849 24145
rect 44849 24093 44871 24145
rect 44895 24093 44901 24145
rect 44901 24093 44913 24145
rect 44913 24093 44951 24145
rect 44975 24093 44977 24145
rect 44977 24093 45029 24145
rect 45029 24093 45031 24145
rect 45055 24093 45093 24145
rect 45093 24093 45105 24145
rect 45105 24093 45111 24145
rect 45135 24093 45157 24145
rect 45157 24093 45169 24145
rect 45169 24093 45191 24145
rect 45215 24093 45221 24145
rect 45221 24093 45233 24145
rect 45233 24093 45271 24145
rect 45295 24093 45297 24145
rect 45297 24093 45349 24145
rect 45349 24093 45351 24145
rect 45375 24093 45413 24145
rect 45413 24093 45425 24145
rect 45425 24093 45431 24145
rect 45455 24093 45477 24145
rect 45477 24093 45489 24145
rect 45489 24093 45511 24145
rect 45535 24093 45541 24145
rect 45541 24093 45553 24145
rect 45553 24093 45591 24145
rect 45615 24093 45617 24145
rect 45617 24093 45669 24145
rect 45669 24093 45671 24145
rect 45695 24093 45733 24145
rect 45733 24093 45745 24145
rect 45745 24093 45751 24145
rect 45775 24093 45797 24145
rect 45797 24093 45809 24145
rect 45809 24093 45831 24145
rect 45855 24093 45861 24145
rect 45861 24093 45873 24145
rect 45873 24093 45911 24145
rect 45935 24093 45937 24145
rect 45937 24093 45989 24145
rect 45989 24093 45991 24145
rect 46015 24093 46053 24145
rect 46053 24093 46065 24145
rect 46065 24093 46071 24145
rect 46095 24093 46117 24145
rect 46117 24093 46129 24145
rect 46129 24093 46151 24145
rect 42895 24091 42951 24093
rect 42975 24091 43031 24093
rect 43055 24091 43111 24093
rect 43135 24091 43191 24093
rect 43215 24091 43271 24093
rect 43295 24091 43351 24093
rect 43375 24091 43431 24093
rect 43455 24091 43511 24093
rect 43535 24091 43591 24093
rect 43615 24091 43671 24093
rect 43695 24091 43751 24093
rect 43775 24091 43831 24093
rect 43855 24091 43911 24093
rect 43935 24091 43991 24093
rect 44015 24091 44071 24093
rect 44095 24091 44151 24093
rect 44175 24091 44231 24093
rect 44255 24091 44311 24093
rect 44335 24091 44391 24093
rect 44415 24091 44471 24093
rect 44495 24091 44551 24093
rect 44575 24091 44631 24093
rect 44655 24091 44711 24093
rect 44735 24091 44791 24093
rect 44815 24091 44871 24093
rect 44895 24091 44951 24093
rect 44975 24091 45031 24093
rect 45055 24091 45111 24093
rect 45135 24091 45191 24093
rect 45215 24091 45271 24093
rect 45295 24091 45351 24093
rect 45375 24091 45431 24093
rect 45455 24091 45511 24093
rect 45535 24091 45591 24093
rect 45615 24091 45671 24093
rect 45695 24091 45751 24093
rect 45775 24091 45831 24093
rect 45855 24091 45911 24093
rect 45935 24091 45991 24093
rect 46015 24091 46071 24093
rect 46095 24091 46151 24093
rect 36070 23958 36126 24014
rect 35156 23860 35212 23862
rect 35156 23808 35158 23860
rect 35158 23808 35210 23860
rect 35210 23808 35212 23860
rect 35156 23806 35212 23808
rect 7095 23592 7151 23648
rect 39355 23693 39411 23711
rect 39355 23655 39357 23693
rect 39357 23655 39409 23693
rect 39409 23655 39411 23693
rect 37827 23557 37829 23579
rect 37829 23557 37881 23579
rect 37881 23557 37883 23579
rect 37827 23545 37883 23557
rect 37827 23523 37829 23545
rect 37829 23523 37881 23545
rect 37881 23523 37883 23545
rect 39355 23629 39411 23631
rect 39355 23577 39357 23629
rect 39357 23577 39409 23629
rect 39409 23577 39411 23629
rect 39355 23575 39411 23577
rect 39355 23513 39357 23551
rect 39357 23513 39409 23551
rect 39409 23513 39411 23551
rect 39355 23495 39411 23513
rect 8797 23327 8853 23329
rect 8877 23327 8933 23329
rect 8797 23275 8807 23327
rect 8807 23275 8853 23327
rect 8877 23275 8923 23327
rect 8923 23275 8933 23327
rect 8797 23273 8853 23275
rect 8877 23273 8933 23275
rect 37834 23140 37836 23178
rect 37836 23140 37888 23178
rect 37888 23140 37890 23178
rect 37834 23128 37890 23140
rect 37834 23122 37836 23128
rect 37836 23122 37888 23128
rect 37888 23122 37890 23128
rect 2554 23057 2610 23059
rect 2554 23005 2556 23057
rect 2556 23005 2608 23057
rect 2608 23005 2610 23057
rect 2554 23003 2610 23005
rect 10206 23057 10262 23059
rect 10206 23005 10208 23057
rect 10208 23005 10260 23057
rect 10260 23005 10262 23057
rect 10206 23003 10262 23005
rect 37834 23076 37836 23098
rect 37836 23076 37888 23098
rect 37888 23076 37890 23098
rect 37834 23064 37890 23076
rect 37834 23042 37836 23064
rect 37836 23042 37888 23064
rect 37888 23042 37890 23064
rect 37834 23012 37836 23018
rect 37836 23012 37888 23018
rect 37888 23012 37890 23018
rect 37834 23000 37890 23012
rect 37834 22962 37836 23000
rect 37836 22962 37888 23000
rect 37888 22962 37890 23000
rect 39350 23146 39352 23184
rect 39352 23146 39404 23184
rect 39404 23146 39406 23184
rect 39350 23134 39406 23146
rect 39350 23128 39352 23134
rect 39352 23128 39404 23134
rect 39404 23128 39406 23134
rect 39350 23082 39352 23104
rect 39352 23082 39404 23104
rect 39404 23082 39406 23104
rect 39350 23070 39406 23082
rect 39350 23048 39352 23070
rect 39352 23048 39404 23070
rect 39404 23048 39406 23070
rect 39350 23018 39352 23024
rect 39352 23018 39404 23024
rect 39404 23018 39406 23024
rect 39350 23006 39406 23018
rect 39350 22968 39352 23006
rect 39352 22968 39404 23006
rect 39404 22968 39406 23006
rect 35122 22632 35258 22768
rect 35782 22725 35838 22727
rect 35862 22725 35918 22727
rect 35942 22725 35998 22727
rect 35782 22673 35820 22725
rect 35820 22673 35832 22725
rect 35832 22673 35838 22725
rect 35862 22673 35884 22725
rect 35884 22673 35896 22725
rect 35896 22673 35918 22725
rect 35942 22673 35948 22725
rect 35948 22673 35960 22725
rect 35960 22673 35998 22725
rect 35782 22671 35838 22673
rect 35862 22671 35918 22673
rect 35942 22671 35998 22673
rect 47566 22706 47782 22724
rect 47566 22526 47584 22706
rect 47584 22526 47764 22706
rect 47764 22526 47782 22706
rect 47566 22508 47782 22526
rect 39355 22367 39411 22385
rect 39355 22329 39357 22367
rect 39357 22329 39409 22367
rect 39409 22329 39411 22367
rect 37833 22221 37835 22243
rect 37835 22221 37887 22243
rect 37887 22221 37889 22243
rect 37833 22209 37889 22221
rect 37833 22187 37835 22209
rect 37835 22187 37887 22209
rect 37887 22187 37889 22209
rect 39355 22303 39411 22305
rect 39355 22251 39357 22303
rect 39357 22251 39409 22303
rect 39409 22251 39411 22303
rect 39355 22249 39411 22251
rect 39355 22187 39357 22225
rect 39357 22187 39409 22225
rect 39409 22187 39411 22225
rect 39355 22169 39411 22187
rect -967 21565 -911 21621
rect 6311 21565 6367 21621
rect 37828 21760 37830 21790
rect 37830 21760 37882 21790
rect 37882 21760 37884 21790
rect 37828 21748 37884 21760
rect 37828 21734 37830 21748
rect 37830 21734 37882 21748
rect 37882 21734 37884 21748
rect 37828 21696 37830 21710
rect 37830 21696 37882 21710
rect 37882 21696 37884 21710
rect 37828 21684 37884 21696
rect 37828 21654 37830 21684
rect 37830 21654 37882 21684
rect 37882 21654 37884 21684
rect 39356 21780 39358 21818
rect 39358 21780 39410 21818
rect 39410 21780 39412 21818
rect 39356 21768 39412 21780
rect 39356 21762 39358 21768
rect 39358 21762 39410 21768
rect 39410 21762 39412 21768
rect 39356 21716 39358 21738
rect 39358 21716 39410 21738
rect 39410 21716 39412 21738
rect 39356 21704 39412 21716
rect 39356 21682 39358 21704
rect 39358 21682 39410 21704
rect 39410 21682 39412 21704
rect 39356 21652 39358 21658
rect 39358 21652 39410 21658
rect 39410 21652 39412 21658
rect 39356 21640 39412 21652
rect 39356 21602 39358 21640
rect 39358 21602 39410 21640
rect 39410 21602 39412 21640
rect 35156 21579 35212 21581
rect 35156 21527 35158 21579
rect 35158 21527 35210 21579
rect 35210 21527 35212 21579
rect 35156 21525 35212 21527
rect 35481 21319 35537 21375
rect 42893 21149 42949 21151
rect 42973 21149 43029 21151
rect 43053 21149 43109 21151
rect 43133 21149 43189 21151
rect 43213 21149 43269 21151
rect 43293 21149 43349 21151
rect 43373 21149 43429 21151
rect 43453 21149 43509 21151
rect 43533 21149 43589 21151
rect 43613 21149 43669 21151
rect 43693 21149 43749 21151
rect 43773 21149 43829 21151
rect 43853 21149 43909 21151
rect 43933 21149 43989 21151
rect 44013 21149 44069 21151
rect 44093 21149 44149 21151
rect 44173 21149 44229 21151
rect 44253 21149 44309 21151
rect 44333 21149 44389 21151
rect 44413 21149 44469 21151
rect 44493 21149 44549 21151
rect 44573 21149 44629 21151
rect 44653 21149 44709 21151
rect 44733 21149 44789 21151
rect 44813 21149 44869 21151
rect 44893 21149 44949 21151
rect 44973 21149 45029 21151
rect 45053 21149 45109 21151
rect 45133 21149 45189 21151
rect 45213 21149 45269 21151
rect 45293 21149 45349 21151
rect 45373 21149 45429 21151
rect 45453 21149 45509 21151
rect 45533 21149 45589 21151
rect 45613 21149 45669 21151
rect 45693 21149 45749 21151
rect 45773 21149 45829 21151
rect 45853 21149 45909 21151
rect 45933 21149 45989 21151
rect 46013 21149 46069 21151
rect 46093 21149 46149 21151
rect 42893 21097 42915 21149
rect 42915 21097 42927 21149
rect 42927 21097 42949 21149
rect 42973 21097 42979 21149
rect 42979 21097 42991 21149
rect 42991 21097 43029 21149
rect 43053 21097 43055 21149
rect 43055 21097 43107 21149
rect 43107 21097 43109 21149
rect 43133 21097 43171 21149
rect 43171 21097 43183 21149
rect 43183 21097 43189 21149
rect 43213 21097 43235 21149
rect 43235 21097 43247 21149
rect 43247 21097 43269 21149
rect 43293 21097 43299 21149
rect 43299 21097 43311 21149
rect 43311 21097 43349 21149
rect 43373 21097 43375 21149
rect 43375 21097 43427 21149
rect 43427 21097 43429 21149
rect 43453 21097 43491 21149
rect 43491 21097 43503 21149
rect 43503 21097 43509 21149
rect 43533 21097 43555 21149
rect 43555 21097 43567 21149
rect 43567 21097 43589 21149
rect 43613 21097 43619 21149
rect 43619 21097 43631 21149
rect 43631 21097 43669 21149
rect 43693 21097 43695 21149
rect 43695 21097 43747 21149
rect 43747 21097 43749 21149
rect 43773 21097 43811 21149
rect 43811 21097 43823 21149
rect 43823 21097 43829 21149
rect 43853 21097 43875 21149
rect 43875 21097 43887 21149
rect 43887 21097 43909 21149
rect 43933 21097 43939 21149
rect 43939 21097 43951 21149
rect 43951 21097 43989 21149
rect 44013 21097 44015 21149
rect 44015 21097 44067 21149
rect 44067 21097 44069 21149
rect 44093 21097 44131 21149
rect 44131 21097 44143 21149
rect 44143 21097 44149 21149
rect 44173 21097 44195 21149
rect 44195 21097 44207 21149
rect 44207 21097 44229 21149
rect 44253 21097 44259 21149
rect 44259 21097 44271 21149
rect 44271 21097 44309 21149
rect 44333 21097 44335 21149
rect 44335 21097 44387 21149
rect 44387 21097 44389 21149
rect 44413 21097 44451 21149
rect 44451 21097 44463 21149
rect 44463 21097 44469 21149
rect 44493 21097 44515 21149
rect 44515 21097 44527 21149
rect 44527 21097 44549 21149
rect 44573 21097 44579 21149
rect 44579 21097 44591 21149
rect 44591 21097 44629 21149
rect 44653 21097 44655 21149
rect 44655 21097 44707 21149
rect 44707 21097 44709 21149
rect 44733 21097 44771 21149
rect 44771 21097 44783 21149
rect 44783 21097 44789 21149
rect 44813 21097 44835 21149
rect 44835 21097 44847 21149
rect 44847 21097 44869 21149
rect 44893 21097 44899 21149
rect 44899 21097 44911 21149
rect 44911 21097 44949 21149
rect 44973 21097 44975 21149
rect 44975 21097 45027 21149
rect 45027 21097 45029 21149
rect 45053 21097 45091 21149
rect 45091 21097 45103 21149
rect 45103 21097 45109 21149
rect 45133 21097 45155 21149
rect 45155 21097 45167 21149
rect 45167 21097 45189 21149
rect 45213 21097 45219 21149
rect 45219 21097 45231 21149
rect 45231 21097 45269 21149
rect 45293 21097 45295 21149
rect 45295 21097 45347 21149
rect 45347 21097 45349 21149
rect 45373 21097 45411 21149
rect 45411 21097 45423 21149
rect 45423 21097 45429 21149
rect 45453 21097 45475 21149
rect 45475 21097 45487 21149
rect 45487 21097 45509 21149
rect 45533 21097 45539 21149
rect 45539 21097 45551 21149
rect 45551 21097 45589 21149
rect 45613 21097 45615 21149
rect 45615 21097 45667 21149
rect 45667 21097 45669 21149
rect 45693 21097 45731 21149
rect 45731 21097 45743 21149
rect 45743 21097 45749 21149
rect 45773 21097 45795 21149
rect 45795 21097 45807 21149
rect 45807 21097 45829 21149
rect 45853 21097 45859 21149
rect 45859 21097 45871 21149
rect 45871 21097 45909 21149
rect 45933 21097 45935 21149
rect 45935 21097 45987 21149
rect 45987 21097 45989 21149
rect 46013 21097 46051 21149
rect 46051 21097 46063 21149
rect 46063 21097 46069 21149
rect 46093 21097 46115 21149
rect 46115 21097 46127 21149
rect 46127 21097 46149 21149
rect 42893 21095 42949 21097
rect 42973 21095 43029 21097
rect 43053 21095 43109 21097
rect 43133 21095 43189 21097
rect 43213 21095 43269 21097
rect 43293 21095 43349 21097
rect 43373 21095 43429 21097
rect 43453 21095 43509 21097
rect 43533 21095 43589 21097
rect 43613 21095 43669 21097
rect 43693 21095 43749 21097
rect 43773 21095 43829 21097
rect 43853 21095 43909 21097
rect 43933 21095 43989 21097
rect 44013 21095 44069 21097
rect 44093 21095 44149 21097
rect 44173 21095 44229 21097
rect 44253 21095 44309 21097
rect 44333 21095 44389 21097
rect 44413 21095 44469 21097
rect 44493 21095 44549 21097
rect 44573 21095 44629 21097
rect 44653 21095 44709 21097
rect 44733 21095 44789 21097
rect 44813 21095 44869 21097
rect 44893 21095 44949 21097
rect 44973 21095 45029 21097
rect 45053 21095 45109 21097
rect 45133 21095 45189 21097
rect 45213 21095 45269 21097
rect 45293 21095 45349 21097
rect 45373 21095 45429 21097
rect 45453 21095 45509 21097
rect 45533 21095 45589 21097
rect 45613 21095 45669 21097
rect 45693 21095 45749 21097
rect 45773 21095 45829 21097
rect 45853 21095 45909 21097
rect 45933 21095 45989 21097
rect 46013 21095 46069 21097
rect 46093 21095 46149 21097
rect 14692 21021 14748 21023
rect 14692 20969 14694 21021
rect 14694 20969 14746 21021
rect 14746 20969 14748 21021
rect 14692 20967 14748 20969
rect 6314 20897 6370 20953
rect -967 20655 -911 20711
rect -14148 15310 -14092 15366
rect -13060 14135 -13004 14137
rect -13060 14083 -13058 14135
rect -13058 14083 -13006 14135
rect -13006 14083 -13004 14135
rect -13060 14081 -13004 14083
rect 55 19453 111 19509
rect -752 19152 -696 19208
rect 14691 19267 14747 19323
rect 4877 19158 5173 19168
rect 3065 19100 3121 19102
rect 3065 19048 3067 19100
rect 3067 19048 3119 19100
rect 3119 19048 3121 19100
rect 3065 19046 3121 19048
rect 4877 19042 5173 19158
rect 4877 19032 5173 19042
rect 7089 19100 7145 19102
rect 7089 19048 7091 19100
rect 7091 19048 7143 19100
rect 7143 19048 7145 19100
rect 7089 19046 7145 19048
rect 8985 19100 9041 19102
rect 8985 19048 8987 19100
rect 8987 19048 9039 19100
rect 9039 19048 9041 19100
rect 8985 19046 9041 19048
rect 10236 19052 10292 19054
rect 10236 19000 10238 19052
rect 10238 19000 10290 19052
rect 10290 19000 10292 19052
rect 10236 18998 10292 19000
rect 23693 19376 23749 19378
rect 23693 19324 23695 19376
rect 23695 19324 23747 19376
rect 23747 19324 23749 19376
rect 23693 19322 23749 19324
rect 20975 19002 21031 19058
rect 5711 18850 5767 18906
rect 7710 18850 7766 18906
rect 4903 18591 4959 18647
rect 6901 18591 6957 18647
rect 8284 18712 8340 18714
rect 8284 18660 8286 18712
rect 8286 18660 8338 18712
rect 8338 18660 8340 18712
rect 8284 18658 8340 18660
rect 13578 18682 13634 18684
rect 13578 18630 13580 18682
rect 13580 18630 13632 18682
rect 13632 18630 13634 18682
rect 13578 18628 13634 18630
rect 3711 18252 3767 18308
rect 9710 18252 9766 18308
rect 2902 17971 2958 18027
rect 8903 17971 8959 18027
rect 237 17766 293 17768
rect 237 17714 239 17766
rect 239 17714 291 17766
rect 291 17714 293 17766
rect 237 17712 293 17714
rect -817 17519 -761 17521
rect -817 17467 -815 17519
rect -815 17467 -763 17519
rect -763 17467 -761 17519
rect -817 17465 -761 17467
rect 14693 17482 14749 17538
rect 23693 17546 23749 17548
rect 23693 17494 23695 17546
rect 23695 17494 23747 17546
rect 23747 17494 23749 17546
rect 23693 17492 23749 17494
rect 4299 17283 4355 17285
rect 4299 17231 4301 17283
rect 4301 17231 4353 17283
rect 4353 17231 4355 17283
rect 4299 17229 4355 17231
rect 6231 17283 6287 17285
rect 6231 17231 6233 17283
rect 6233 17231 6285 17283
rect 6285 17231 6287 17283
rect 6231 17229 6287 17231
rect -10412 17097 -10356 17153
rect 13607 17023 13663 17079
rect -10411 16228 -10355 16284
rect 267 16274 11123 16410
rect -5782 15702 -5726 15704
rect -5782 15650 -5780 15702
rect -5780 15650 -5728 15702
rect -5728 15650 -5726 15702
rect -5782 15648 -5726 15650
rect -3004 15394 -2948 15450
rect -4895 14379 -4893 14409
rect -4893 14379 -4841 14409
rect -4841 14379 -4839 14409
rect -4895 14367 -4839 14379
rect -4895 14353 -4893 14367
rect -4893 14353 -4841 14367
rect -4841 14353 -4839 14367
rect -4895 14315 -4893 14329
rect -4893 14315 -4841 14329
rect -4841 14315 -4839 14329
rect -4895 14303 -4839 14315
rect -4895 14273 -4893 14303
rect -4893 14273 -4841 14303
rect -4841 14273 -4839 14303
rect -4903 13922 -4901 13960
rect -4901 13922 -4849 13960
rect -4849 13922 -4847 13960
rect -4903 13910 -4847 13922
rect -4903 13904 -4901 13910
rect -4901 13904 -4849 13910
rect -4849 13904 -4847 13910
rect -4903 13858 -4901 13880
rect -4901 13858 -4849 13880
rect -4849 13858 -4847 13880
rect -4903 13846 -4847 13858
rect -4903 13824 -4901 13846
rect -4901 13824 -4849 13846
rect -4849 13824 -4847 13846
rect -4903 13794 -4901 13800
rect -4901 13794 -4849 13800
rect -4849 13794 -4847 13800
rect -4903 13782 -4847 13794
rect -4903 13744 -4901 13782
rect -4901 13744 -4849 13782
rect -4849 13744 -4847 13782
rect -6158 10821 -6102 10823
rect -6078 10821 -6022 10823
rect -5998 10821 -5942 10823
rect -6158 10769 -6140 10821
rect -6140 10769 -6102 10821
rect -6078 10769 -6076 10821
rect -6076 10769 -6024 10821
rect -6024 10769 -6022 10821
rect -5998 10769 -5960 10821
rect -5960 10769 -5942 10821
rect -6158 10767 -6102 10769
rect -6078 10767 -6022 10769
rect -5998 10767 -5942 10769
rect -10966 10163 -10910 10219
rect -5702 10820 -5646 10822
rect -5622 10820 -5566 10822
rect -5542 10820 -5486 10822
rect -5462 10820 -5406 10822
rect -5702 10768 -5676 10820
rect -5676 10768 -5646 10820
rect -5622 10768 -5612 10820
rect -5612 10768 -5566 10820
rect -5542 10768 -5496 10820
rect -5496 10768 -5486 10820
rect -5462 10768 -5432 10820
rect -5432 10768 -5406 10820
rect -5702 10766 -5646 10768
rect -5622 10766 -5566 10768
rect -5542 10766 -5486 10768
rect -5462 10766 -5406 10768
rect -6152 10144 -6096 10200
rect -6156 9578 -6100 9580
rect -6076 9578 -6020 9580
rect -5996 9578 -5940 9580
rect -6156 9526 -6138 9578
rect -6138 9526 -6100 9578
rect -6076 9526 -6074 9578
rect -6074 9526 -6022 9578
rect -6022 9526 -6020 9578
rect -5996 9526 -5958 9578
rect -5958 9526 -5940 9578
rect -6156 9524 -6100 9526
rect -6076 9524 -6020 9526
rect -5996 9524 -5940 9526
rect -3131 14928 -3129 14966
rect -3129 14928 -3077 14966
rect -3077 14928 -3075 14966
rect -3131 14916 -3075 14928
rect -3131 14910 -3129 14916
rect -3129 14910 -3077 14916
rect -3077 14910 -3075 14916
rect -3131 14864 -3129 14886
rect -3129 14864 -3077 14886
rect -3077 14864 -3075 14886
rect -3131 14852 -3075 14864
rect -3131 14830 -3129 14852
rect -3129 14830 -3077 14852
rect -3077 14830 -3075 14852
rect -3131 14800 -3129 14806
rect -3129 14800 -3077 14806
rect -3077 14800 -3075 14806
rect -3131 14788 -3075 14800
rect -3131 14750 -3129 14788
rect -3129 14750 -3077 14788
rect -3077 14750 -3075 14788
rect -3019 14584 -2963 14640
rect -2594 13077 -2538 13133
rect -1795 13115 -1739 13117
rect -1795 13063 -1793 13115
rect -1793 13063 -1741 13115
rect -1741 13063 -1739 13115
rect -1795 13061 -1739 13063
rect -1795 12999 -1793 13037
rect -1793 12999 -1741 13037
rect -1741 12999 -1739 13037
rect -1795 12987 -1739 12999
rect -1795 12981 -1793 12987
rect -1793 12981 -1741 12987
rect -1741 12981 -1739 12987
rect -1795 12935 -1793 12957
rect -1793 12935 -1741 12957
rect -1741 12935 -1739 12957
rect -1795 12923 -1739 12935
rect -1795 12901 -1793 12923
rect -1793 12901 -1741 12923
rect -1741 12901 -1739 12923
rect -1795 12871 -1793 12877
rect -1793 12871 -1741 12877
rect -1741 12871 -1739 12877
rect -1795 12859 -1739 12871
rect -1795 12821 -1793 12859
rect -1793 12821 -1741 12859
rect -1741 12821 -1739 12859
rect -1795 12795 -1739 12797
rect -1795 12743 -1793 12795
rect -1793 12743 -1741 12795
rect -1741 12743 -1739 12795
rect -1795 12741 -1739 12743
rect -5357 10144 -5301 10200
rect -4785 10173 -4729 10229
rect -4444 10173 -4388 10229
rect -5702 9578 -5646 9580
rect -5622 9578 -5566 9580
rect -5542 9578 -5486 9580
rect -5462 9578 -5406 9580
rect -5702 9526 -5656 9578
rect -5656 9526 -5646 9578
rect -5622 9526 -5592 9578
rect -5592 9526 -5580 9578
rect -5580 9526 -5566 9578
rect -5542 9526 -5528 9578
rect -5528 9526 -5516 9578
rect -5516 9526 -5486 9578
rect -5462 9526 -5452 9578
rect -5452 9526 -5406 9578
rect -5702 9524 -5646 9526
rect -5622 9524 -5566 9526
rect -5542 9524 -5486 9526
rect -5462 9524 -5406 9526
rect -16745 7547 -16689 7603
rect -7211 7213 -6755 7231
rect -7211 7033 -7201 7213
rect -7201 7033 -6765 7213
rect -6765 7033 -6755 7213
rect -7211 7015 -6755 7033
rect -25512 6608 -25510 6646
rect -25510 6608 -25458 6646
rect -25458 6608 -25456 6646
rect -25512 6596 -25456 6608
rect -25512 6590 -25510 6596
rect -25510 6590 -25458 6596
rect -25458 6590 -25456 6596
rect -25512 6544 -25510 6566
rect -25510 6544 -25458 6566
rect -25458 6544 -25456 6566
rect -25512 6532 -25456 6544
rect -25512 6510 -25510 6532
rect -25510 6510 -25458 6532
rect -25458 6510 -25456 6532
rect -25512 6480 -25510 6486
rect -25510 6480 -25458 6486
rect -25458 6480 -25456 6486
rect -25512 6468 -25456 6480
rect -25512 6430 -25510 6468
rect -25510 6430 -25458 6468
rect -25458 6430 -25456 6468
rect -18247 6297 -18191 6299
rect -18247 6245 -18245 6297
rect -18245 6245 -18193 6297
rect -18193 6245 -18191 6297
rect -18247 6243 -18191 6245
rect -13071 6307 -13015 6309
rect -13071 6255 -13069 6307
rect -13069 6255 -13017 6307
rect -13017 6255 -13015 6307
rect -13071 6253 -13015 6255
rect -4905 6665 -4849 6691
rect -4905 6635 -4903 6665
rect -4903 6635 -4851 6665
rect -4851 6635 -4849 6665
rect -4905 6601 -4849 6611
rect -4905 6555 -4903 6601
rect -4903 6555 -4851 6601
rect -4851 6555 -4849 6601
rect -4905 6485 -4903 6531
rect -4903 6485 -4851 6531
rect -4851 6485 -4849 6531
rect -4905 6475 -4849 6485
rect -4905 6421 -4903 6451
rect -4903 6421 -4851 6451
rect -4851 6421 -4849 6451
rect -4905 6395 -4849 6421
rect -25513 6121 -25511 6159
rect -25511 6121 -25459 6159
rect -25459 6121 -25457 6159
rect -25513 6109 -25457 6121
rect -25513 6103 -25511 6109
rect -25511 6103 -25459 6109
rect -25459 6103 -25457 6109
rect -25513 6057 -25511 6079
rect -25511 6057 -25459 6079
rect -25459 6057 -25457 6079
rect -25513 6045 -25457 6057
rect -25513 6023 -25511 6045
rect -25511 6023 -25459 6045
rect -25459 6023 -25457 6045
rect -25513 5993 -25511 5999
rect -25511 5993 -25459 5999
rect -25459 5993 -25457 5999
rect -25513 5981 -25457 5993
rect -25513 5943 -25511 5981
rect -25511 5943 -25459 5981
rect -25459 5943 -25457 5981
rect -4902 6094 -4900 6124
rect -4900 6094 -4848 6124
rect -4848 6094 -4846 6124
rect -4902 6082 -4846 6094
rect -4902 6068 -4900 6082
rect -4900 6068 -4848 6082
rect -4848 6068 -4846 6082
rect -4902 6030 -4900 6044
rect -4900 6030 -4848 6044
rect -4848 6030 -4846 6044
rect -4902 6018 -4846 6030
rect -4902 5988 -4900 6018
rect -4900 5988 -4848 6018
rect -4848 5988 -4846 6018
rect -1494 12403 -1438 12405
rect -1494 12351 -1492 12403
rect -1492 12351 -1440 12403
rect -1440 12351 -1438 12403
rect -1494 12349 -1438 12351
rect -2881 12268 -2825 12324
rect -1922 11475 -1866 11531
rect -1754 11520 -1698 11522
rect -1754 11468 -1752 11520
rect -1752 11468 -1700 11520
rect -1700 11468 -1698 11520
rect -1754 11466 -1698 11468
rect -1754 11404 -1752 11442
rect -1752 11404 -1700 11442
rect -1700 11404 -1698 11442
rect -1754 11392 -1698 11404
rect -1754 11386 -1752 11392
rect -1752 11386 -1700 11392
rect -1700 11386 -1698 11392
rect -1754 11340 -1752 11362
rect -1752 11340 -1700 11362
rect -1700 11340 -1698 11362
rect -1754 11328 -1698 11340
rect -1754 11306 -1752 11328
rect -1752 11306 -1700 11328
rect -1700 11306 -1698 11328
rect -1754 11276 -1752 11282
rect -1752 11276 -1700 11282
rect -1700 11276 -1698 11282
rect -1754 11264 -1698 11276
rect -1754 11226 -1752 11264
rect -1752 11226 -1700 11264
rect -1700 11226 -1698 11264
rect -1754 11200 -1698 11202
rect -1754 11148 -1752 11200
rect -1752 11148 -1700 11200
rect -1700 11148 -1698 11200
rect -1754 11146 -1698 11148
rect -2208 10669 -2152 10725
rect -1494 10777 -1438 10779
rect -1494 10725 -1492 10777
rect -1492 10725 -1440 10777
rect -1440 10725 -1438 10777
rect -1494 10723 -1438 10725
rect -1922 9877 -1866 9933
rect -1755 9917 -1699 9919
rect -1755 9865 -1753 9917
rect -1753 9865 -1701 9917
rect -1701 9865 -1699 9917
rect -1755 9863 -1699 9865
rect -1755 9801 -1753 9839
rect -1753 9801 -1701 9839
rect -1701 9801 -1699 9839
rect -1755 9789 -1699 9801
rect -1755 9783 -1753 9789
rect -1753 9783 -1701 9789
rect -1701 9783 -1699 9789
rect -1755 9737 -1753 9759
rect -1753 9737 -1701 9759
rect -1701 9737 -1699 9759
rect -1755 9725 -1699 9737
rect -1755 9703 -1753 9725
rect -1753 9703 -1701 9725
rect -1701 9703 -1699 9725
rect -1755 9673 -1753 9679
rect -1753 9673 -1701 9679
rect -1701 9673 -1699 9679
rect -1755 9661 -1699 9673
rect -1755 9623 -1753 9661
rect -1753 9623 -1701 9661
rect -1701 9623 -1699 9661
rect -1755 9597 -1699 9599
rect -1755 9545 -1753 9597
rect -1753 9545 -1701 9597
rect -1701 9545 -1699 9597
rect -1755 9543 -1699 9545
rect -2208 9069 -2152 9125
rect -1494 9119 -1438 9121
rect -1494 9067 -1492 9119
rect -1492 9067 -1440 9119
rect -1440 9067 -1438 9119
rect -1494 9065 -1438 9067
rect -2594 8275 -2538 8331
rect -1752 8316 -1696 8318
rect -1752 8264 -1750 8316
rect -1750 8264 -1698 8316
rect -1698 8264 -1696 8316
rect -1752 8262 -1696 8264
rect -1752 8200 -1750 8238
rect -1750 8200 -1698 8238
rect -1698 8200 -1696 8238
rect -1752 8188 -1696 8200
rect -1752 8182 -1750 8188
rect -1750 8182 -1698 8188
rect -1698 8182 -1696 8188
rect -1752 8136 -1750 8158
rect -1750 8136 -1698 8158
rect -1698 8136 -1696 8158
rect -1752 8124 -1696 8136
rect -1752 8102 -1750 8124
rect -1750 8102 -1698 8124
rect -1698 8102 -1696 8124
rect -1752 8072 -1750 8078
rect -1750 8072 -1698 8078
rect -1698 8072 -1696 8078
rect -1752 8060 -1696 8072
rect -1752 8022 -1750 8060
rect -1750 8022 -1698 8060
rect -1698 8022 -1696 8060
rect -1752 7996 -1696 7998
rect -1752 7944 -1750 7996
rect -1750 7944 -1698 7996
rect -1698 7944 -1696 7996
rect -1752 7942 -1696 7944
rect -2881 7467 -2825 7523
rect -1494 7580 -1438 7582
rect -1494 7528 -1492 7580
rect -1492 7528 -1440 7580
rect -1440 7528 -1438 7580
rect -1494 7526 -1438 7528
rect -1494 7186 -1492 7224
rect -1492 7186 -1440 7224
rect -1440 7186 -1438 7224
rect -1494 7174 -1438 7186
rect -1494 7168 -1492 7174
rect -1492 7168 -1440 7174
rect -1440 7168 -1438 7174
rect -1494 7122 -1492 7144
rect -1492 7122 -1440 7144
rect -1440 7122 -1438 7144
rect -1494 7110 -1438 7122
rect -1494 7088 -1492 7110
rect -1492 7088 -1440 7110
rect -1440 7088 -1438 7110
rect -1494 7058 -1492 7064
rect -1492 7058 -1440 7064
rect -1440 7058 -1438 7064
rect -1494 7046 -1438 7058
rect -1494 7008 -1492 7046
rect -1492 7008 -1440 7046
rect -1440 7008 -1438 7046
rect -1494 6445 -1438 6447
rect -1494 6393 -1492 6445
rect -1492 6393 -1440 6445
rect -1440 6393 -1438 6445
rect -1494 6391 -1438 6393
rect -3046 5982 -2990 6038
rect -3180 5506 -3178 5544
rect -3178 5506 -3126 5544
rect -3126 5506 -3124 5544
rect -3180 5494 -3124 5506
rect -3180 5488 -3178 5494
rect -3178 5488 -3126 5494
rect -3126 5488 -3124 5494
rect -3180 5442 -3178 5464
rect -3178 5442 -3126 5464
rect -3126 5442 -3124 5464
rect -3180 5430 -3124 5442
rect -3180 5408 -3178 5430
rect -3178 5408 -3126 5430
rect -3126 5408 -3124 5430
rect -3180 5378 -3178 5384
rect -3178 5378 -3126 5384
rect -3126 5378 -3124 5384
rect -3180 5366 -3124 5378
rect -3180 5328 -3178 5366
rect -3178 5328 -3126 5366
rect -3126 5328 -3124 5366
rect -3024 5173 -2968 5229
rect -10762 4987 -10706 5043
rect 39 16160 175 16162
rect 39 10668 49 16160
rect 49 10668 165 16160
rect 165 10668 175 16160
rect 39 10666 175 10668
rect 11251 16163 11387 16173
rect 11251 14447 11261 16163
rect 11261 14447 11377 16163
rect 11377 14447 11387 16163
rect 11251 14437 11387 14447
rect 23690 15782 23746 15784
rect 23690 15730 23692 15782
rect 23692 15730 23744 15782
rect 23744 15730 23746 15782
rect 23690 15728 23746 15730
rect 14690 15651 14746 15707
rect 20932 15490 20988 15492
rect 20932 15438 20934 15490
rect 20934 15438 20986 15490
rect 20986 15438 20988 15490
rect 20932 15436 20988 15438
rect 14694 15222 14750 15224
rect 14694 15170 14696 15222
rect 14696 15170 14748 15222
rect 14748 15170 14750 15222
rect 14694 15168 14750 15170
rect 11292 13884 11348 13940
rect 11292 13804 11348 13860
rect 11292 13724 11348 13780
rect 11292 13644 11348 13700
rect 11292 13564 11348 13620
rect 11292 13484 11348 13540
rect 11292 13404 11348 13460
rect 11292 13324 11348 13380
rect 11292 13244 11348 13300
rect 11292 13164 11348 13220
rect 11292 13084 11348 13140
rect 11292 13004 11348 13060
rect 14689 13959 14745 13961
rect 14689 13907 14691 13959
rect 14691 13907 14743 13959
rect 14743 13907 14745 13959
rect 14689 13905 14745 13907
rect 23690 13991 23746 13993
rect 23690 13939 23692 13991
rect 23692 13939 23744 13991
rect 23744 13939 23746 13991
rect 23690 13937 23746 13939
rect 13640 13468 13696 13524
rect 11252 12100 11388 12110
rect 11252 11344 11262 12100
rect 11262 11344 11378 12100
rect 11378 11344 11388 12100
rect 11252 11334 11388 11344
rect 14706 12174 14762 12176
rect 14706 12122 14708 12174
rect 14708 12122 14760 12174
rect 14760 12122 14762 12174
rect 14706 12120 14762 12122
rect 23695 12184 23751 12186
rect 23695 12132 23697 12184
rect 23697 12132 23749 12184
rect 23749 12132 23751 12184
rect 23695 12130 23751 12132
rect 20989 11846 21045 11902
rect 13703 11616 13759 11672
rect 6502 10378 11198 10514
rect 14695 10377 14751 10379
rect 14695 10325 14697 10377
rect 14697 10325 14749 10377
rect 14749 10325 14751 10377
rect 14695 10323 14751 10325
rect 23695 10374 23751 10376
rect 23695 10322 23697 10374
rect 23697 10322 23749 10374
rect 23749 10322 23751 10374
rect 23695 10320 23751 10322
rect 35493 8471 35549 8527
rect 36070 9094 36126 9150
rect 36635 8409 36691 8465
rect 35028 8277 35084 8279
rect 35028 8225 35030 8277
rect 35030 8225 35082 8277
rect 35082 8225 35084 8277
rect 35028 8223 35084 8225
rect 38582 8023 38638 8033
rect 38582 7977 38584 8023
rect 38584 7977 38636 8023
rect 38636 7977 38638 8023
rect 38582 7907 38584 7953
rect 38584 7907 38636 7953
rect 38636 7907 38638 7953
rect 38582 7897 38638 7907
rect 40112 8065 40114 8095
rect 40114 8065 40166 8095
rect 40166 8065 40168 8095
rect 40112 8053 40168 8065
rect 40112 8039 40114 8053
rect 40114 8039 40166 8053
rect 40166 8039 40168 8053
rect 40112 8001 40114 8015
rect 40114 8001 40166 8015
rect 40166 8001 40168 8015
rect 40112 7989 40168 8001
rect 40112 7959 40114 7989
rect 40114 7959 40166 7989
rect 40166 7959 40168 7989
rect 36308 7873 36364 7875
rect 36388 7873 36444 7875
rect 36468 7873 36524 7875
rect 36308 7821 36326 7873
rect 36326 7821 36364 7873
rect 36388 7821 36390 7873
rect 36390 7821 36442 7873
rect 36442 7821 36444 7873
rect 36468 7821 36506 7873
rect 36506 7821 36524 7873
rect 36308 7819 36364 7821
rect 36388 7819 36444 7821
rect 36468 7819 36524 7821
rect 38580 7507 38582 7537
rect 38582 7507 38634 7537
rect 38634 7507 38636 7537
rect 38580 7495 38636 7507
rect 38580 7481 38582 7495
rect 38582 7481 38634 7495
rect 38634 7481 38636 7495
rect 38580 7443 38582 7457
rect 38582 7443 38634 7457
rect 38634 7443 38636 7457
rect 38580 7431 38636 7443
rect 38580 7401 38582 7431
rect 38582 7401 38634 7431
rect 38634 7401 38636 7431
rect 40099 7520 40101 7550
rect 40101 7520 40153 7550
rect 40153 7520 40155 7550
rect 40099 7508 40155 7520
rect 40099 7494 40101 7508
rect 40101 7494 40153 7508
rect 40153 7494 40155 7508
rect 40099 7456 40101 7470
rect 40101 7456 40153 7470
rect 40153 7456 40155 7470
rect 40099 7444 40155 7456
rect 40099 7414 40101 7444
rect 40101 7414 40153 7444
rect 40153 7414 40155 7444
rect 36378 7332 36434 7334
rect 36458 7332 36514 7334
rect 36378 7280 36388 7332
rect 36388 7280 36434 7332
rect 36458 7280 36504 7332
rect 36504 7280 36514 7332
rect 36378 7278 36434 7280
rect 36458 7278 36514 7280
rect 35032 7217 35088 7219
rect 35032 7165 35034 7217
rect 35034 7165 35086 7217
rect 35086 7165 35088 7217
rect 35032 7163 35088 7165
rect 42634 7213 42690 7215
rect 42714 7213 42770 7215
rect 42794 7213 42850 7215
rect 42874 7213 42930 7215
rect 42954 7213 43010 7215
rect 43034 7213 43090 7215
rect 43114 7213 43170 7215
rect 43194 7213 43250 7215
rect 43274 7213 43330 7215
rect 43354 7213 43410 7215
rect 43434 7213 43490 7215
rect 43514 7213 43570 7215
rect 43594 7213 43650 7215
rect 43674 7213 43730 7215
rect 43754 7213 43810 7215
rect 43834 7213 43890 7215
rect 43914 7213 43970 7215
rect 43994 7213 44050 7215
rect 44074 7213 44130 7215
rect 44154 7213 44210 7215
rect 44234 7213 44290 7215
rect 44314 7213 44370 7215
rect 44394 7213 44450 7215
rect 44474 7213 44530 7215
rect 44554 7213 44610 7215
rect 44634 7213 44690 7215
rect 44714 7213 44770 7215
rect 44794 7213 44850 7215
rect 44874 7213 44930 7215
rect 44954 7213 45010 7215
rect 45034 7213 45090 7215
rect 45114 7213 45170 7215
rect 45194 7213 45250 7215
rect 45274 7213 45330 7215
rect 45354 7213 45410 7215
rect 45434 7213 45490 7215
rect 45514 7213 45570 7215
rect 45594 7213 45650 7215
rect 45674 7213 45730 7215
rect 45754 7213 45810 7215
rect 45834 7213 45890 7215
rect 42634 7161 42656 7213
rect 42656 7161 42668 7213
rect 42668 7161 42690 7213
rect 42714 7161 42720 7213
rect 42720 7161 42732 7213
rect 42732 7161 42770 7213
rect 42794 7161 42796 7213
rect 42796 7161 42848 7213
rect 42848 7161 42850 7213
rect 42874 7161 42912 7213
rect 42912 7161 42924 7213
rect 42924 7161 42930 7213
rect 42954 7161 42976 7213
rect 42976 7161 42988 7213
rect 42988 7161 43010 7213
rect 43034 7161 43040 7213
rect 43040 7161 43052 7213
rect 43052 7161 43090 7213
rect 43114 7161 43116 7213
rect 43116 7161 43168 7213
rect 43168 7161 43170 7213
rect 43194 7161 43232 7213
rect 43232 7161 43244 7213
rect 43244 7161 43250 7213
rect 43274 7161 43296 7213
rect 43296 7161 43308 7213
rect 43308 7161 43330 7213
rect 43354 7161 43360 7213
rect 43360 7161 43372 7213
rect 43372 7161 43410 7213
rect 43434 7161 43436 7213
rect 43436 7161 43488 7213
rect 43488 7161 43490 7213
rect 43514 7161 43552 7213
rect 43552 7161 43564 7213
rect 43564 7161 43570 7213
rect 43594 7161 43616 7213
rect 43616 7161 43628 7213
rect 43628 7161 43650 7213
rect 43674 7161 43680 7213
rect 43680 7161 43692 7213
rect 43692 7161 43730 7213
rect 43754 7161 43756 7213
rect 43756 7161 43808 7213
rect 43808 7161 43810 7213
rect 43834 7161 43872 7213
rect 43872 7161 43884 7213
rect 43884 7161 43890 7213
rect 43914 7161 43936 7213
rect 43936 7161 43948 7213
rect 43948 7161 43970 7213
rect 43994 7161 44000 7213
rect 44000 7161 44012 7213
rect 44012 7161 44050 7213
rect 44074 7161 44076 7213
rect 44076 7161 44128 7213
rect 44128 7161 44130 7213
rect 44154 7161 44192 7213
rect 44192 7161 44204 7213
rect 44204 7161 44210 7213
rect 44234 7161 44256 7213
rect 44256 7161 44268 7213
rect 44268 7161 44290 7213
rect 44314 7161 44320 7213
rect 44320 7161 44332 7213
rect 44332 7161 44370 7213
rect 44394 7161 44396 7213
rect 44396 7161 44448 7213
rect 44448 7161 44450 7213
rect 44474 7161 44512 7213
rect 44512 7161 44524 7213
rect 44524 7161 44530 7213
rect 44554 7161 44576 7213
rect 44576 7161 44588 7213
rect 44588 7161 44610 7213
rect 44634 7161 44640 7213
rect 44640 7161 44652 7213
rect 44652 7161 44690 7213
rect 44714 7161 44716 7213
rect 44716 7161 44768 7213
rect 44768 7161 44770 7213
rect 44794 7161 44832 7213
rect 44832 7161 44844 7213
rect 44844 7161 44850 7213
rect 44874 7161 44896 7213
rect 44896 7161 44908 7213
rect 44908 7161 44930 7213
rect 44954 7161 44960 7213
rect 44960 7161 44972 7213
rect 44972 7161 45010 7213
rect 45034 7161 45036 7213
rect 45036 7161 45088 7213
rect 45088 7161 45090 7213
rect 45114 7161 45152 7213
rect 45152 7161 45164 7213
rect 45164 7161 45170 7213
rect 45194 7161 45216 7213
rect 45216 7161 45228 7213
rect 45228 7161 45250 7213
rect 45274 7161 45280 7213
rect 45280 7161 45292 7213
rect 45292 7161 45330 7213
rect 45354 7161 45356 7213
rect 45356 7161 45408 7213
rect 45408 7161 45410 7213
rect 45434 7161 45472 7213
rect 45472 7161 45484 7213
rect 45484 7161 45490 7213
rect 45514 7161 45536 7213
rect 45536 7161 45548 7213
rect 45548 7161 45570 7213
rect 45594 7161 45600 7213
rect 45600 7161 45612 7213
rect 45612 7161 45650 7213
rect 45674 7161 45676 7213
rect 45676 7161 45728 7213
rect 45728 7161 45730 7213
rect 45754 7161 45792 7213
rect 45792 7161 45804 7213
rect 45804 7161 45810 7213
rect 45834 7161 45856 7213
rect 45856 7161 45868 7213
rect 45868 7161 45890 7213
rect 42634 7159 42690 7161
rect 42714 7159 42770 7161
rect 42794 7159 42850 7161
rect 42874 7159 42930 7161
rect 42954 7159 43010 7161
rect 43034 7159 43090 7161
rect 43114 7159 43170 7161
rect 43194 7159 43250 7161
rect 43274 7159 43330 7161
rect 43354 7159 43410 7161
rect 43434 7159 43490 7161
rect 43514 7159 43570 7161
rect 43594 7159 43650 7161
rect 43674 7159 43730 7161
rect 43754 7159 43810 7161
rect 43834 7159 43890 7161
rect 43914 7159 43970 7161
rect 43994 7159 44050 7161
rect 44074 7159 44130 7161
rect 44154 7159 44210 7161
rect 44234 7159 44290 7161
rect 44314 7159 44370 7161
rect 44394 7159 44450 7161
rect 44474 7159 44530 7161
rect 44554 7159 44610 7161
rect 44634 7159 44690 7161
rect 44714 7159 44770 7161
rect 44794 7159 44850 7161
rect 44874 7159 44930 7161
rect 44954 7159 45010 7161
rect 45034 7159 45090 7161
rect 45114 7159 45170 7161
rect 45194 7159 45250 7161
rect 45274 7159 45330 7161
rect 45354 7159 45410 7161
rect 45434 7159 45490 7161
rect 45514 7159 45570 7161
rect 45594 7159 45650 7161
rect 45674 7159 45730 7161
rect 45754 7159 45810 7161
rect 45834 7159 45890 7161
rect 35031 6948 35087 6950
rect 35031 6896 35033 6948
rect 35033 6896 35085 6948
rect 35085 6896 35087 6948
rect 35031 6894 35087 6896
rect 36366 6784 36422 6786
rect 36366 6732 36368 6784
rect 36368 6732 36420 6784
rect 36420 6732 36422 6784
rect 36366 6730 36422 6732
rect 38582 6650 38584 6672
rect 38584 6650 38636 6672
rect 38636 6650 38638 6672
rect 38582 6638 38638 6650
rect 38582 6616 38584 6638
rect 38584 6616 38636 6638
rect 38636 6616 38638 6638
rect 40104 6729 40106 6759
rect 40106 6729 40158 6759
rect 40158 6729 40160 6759
rect 40104 6717 40160 6729
rect 40104 6703 40106 6717
rect 40106 6703 40158 6717
rect 40158 6703 40160 6717
rect 40104 6665 40106 6679
rect 40106 6665 40158 6679
rect 40158 6665 40160 6679
rect 40104 6653 40160 6665
rect 40104 6623 40106 6653
rect 40106 6623 40158 6653
rect 40158 6623 40160 6653
rect 36991 6243 37047 6245
rect 36991 6191 36993 6243
rect 36993 6191 37045 6243
rect 37045 6191 37047 6243
rect 36991 6189 37047 6191
rect 38575 6176 38577 6206
rect 38577 6176 38629 6206
rect 38629 6176 38631 6206
rect 38575 6164 38631 6176
rect 38575 6150 38577 6164
rect 38577 6150 38629 6164
rect 38629 6150 38631 6164
rect 38575 6112 38577 6126
rect 38577 6112 38629 6126
rect 38629 6112 38631 6126
rect 38575 6100 38631 6112
rect 38575 6070 38577 6100
rect 38577 6070 38629 6100
rect 38629 6070 38631 6100
rect 40104 6173 40106 6203
rect 40106 6173 40158 6203
rect 40158 6173 40160 6203
rect 40104 6161 40160 6173
rect 40104 6147 40106 6161
rect 40106 6147 40158 6161
rect 40158 6147 40160 6161
rect 40104 6109 40106 6123
rect 40106 6109 40158 6123
rect 40158 6109 40160 6123
rect 40104 6097 40160 6109
rect 40104 6067 40106 6097
rect 40106 6067 40158 6097
rect 40158 6067 40160 6097
rect 35031 5879 35087 5881
rect 35031 5827 35033 5879
rect 35033 5827 35085 5879
rect 35085 5827 35087 5879
rect 35031 5825 35087 5827
rect 35991 5701 36047 5703
rect 36071 5701 36127 5703
rect 35991 5649 36001 5701
rect 36001 5649 36047 5701
rect 36071 5649 36117 5701
rect 36117 5649 36127 5701
rect 35991 5647 36047 5649
rect 36071 5647 36127 5649
rect 47483 5772 47699 5790
rect 47483 5592 47501 5772
rect 47501 5592 47681 5772
rect 47681 5592 47699 5772
rect 47483 5574 47699 5592
rect 35028 5556 35084 5558
rect 35028 5504 35030 5556
rect 35030 5504 35082 5556
rect 35082 5504 35084 5556
rect 35028 5502 35084 5504
rect 38583 5260 38585 5282
rect 38585 5260 38637 5282
rect 38637 5260 38639 5282
rect 38583 5248 38639 5260
rect 38583 5226 38585 5248
rect 38585 5226 38637 5248
rect 38637 5226 38639 5248
rect 40121 5349 40123 5379
rect 40123 5349 40175 5379
rect 40175 5349 40177 5379
rect 40121 5337 40177 5349
rect 40121 5323 40123 5337
rect 40123 5323 40175 5337
rect 40175 5323 40177 5337
rect 40121 5285 40123 5299
rect 40123 5285 40175 5299
rect 40175 5285 40177 5299
rect 40121 5273 40177 5285
rect 40121 5243 40123 5273
rect 40123 5243 40175 5273
rect 40175 5243 40177 5273
rect 36516 5153 36572 5155
rect 36596 5153 36652 5155
rect 36676 5153 36732 5155
rect 36516 5101 36534 5153
rect 36534 5101 36572 5153
rect 36596 5101 36598 5153
rect 36598 5101 36650 5153
rect 36650 5101 36652 5153
rect 36676 5101 36714 5153
rect 36714 5101 36732 5153
rect 36516 5099 36572 5101
rect 36596 5099 36652 5101
rect 36676 5099 36732 5101
rect 38574 4823 38576 4853
rect 38576 4823 38628 4853
rect 38628 4823 38630 4853
rect 38574 4811 38630 4823
rect 38574 4797 38576 4811
rect 38576 4797 38628 4811
rect 38628 4797 38630 4811
rect 38574 4759 38576 4773
rect 38576 4759 38628 4773
rect 38628 4759 38630 4773
rect 38574 4747 38630 4759
rect 38574 4717 38576 4747
rect 38576 4717 38628 4747
rect 38628 4717 38630 4747
rect 40104 4801 40106 4831
rect 40106 4801 40158 4831
rect 40158 4801 40160 4831
rect 40104 4789 40160 4801
rect 40104 4775 40106 4789
rect 40106 4775 40158 4789
rect 40158 4775 40160 4789
rect 40104 4737 40106 4751
rect 40106 4737 40158 4751
rect 40158 4737 40160 4751
rect 40104 4725 40160 4737
rect 40104 4695 40106 4725
rect 40106 4695 40158 4725
rect 40158 4695 40160 4725
rect 36368 4610 36424 4612
rect 36448 4610 36504 4612
rect 36368 4558 36378 4610
rect 36378 4558 36424 4610
rect 36448 4558 36494 4610
rect 36494 4558 36504 4610
rect 36368 4556 36424 4558
rect 36448 4556 36504 4558
rect 35039 4486 35095 4488
rect 35039 4434 35041 4486
rect 35041 4434 35093 4486
rect 35093 4434 35095 4486
rect 35039 4432 35095 4434
rect 35028 4181 35084 4183
rect 35028 4129 35030 4181
rect 35030 4129 35082 4181
rect 35082 4129 35084 4181
rect 35028 4127 35084 4129
rect 42611 4214 42667 4216
rect 42691 4214 42747 4216
rect 42771 4214 42827 4216
rect 42851 4214 42907 4216
rect 42931 4214 42987 4216
rect 43011 4214 43067 4216
rect 43091 4214 43147 4216
rect 43171 4214 43227 4216
rect 43251 4214 43307 4216
rect 43331 4214 43387 4216
rect 43411 4214 43467 4216
rect 43491 4214 43547 4216
rect 43571 4214 43627 4216
rect 43651 4214 43707 4216
rect 43731 4214 43787 4216
rect 43811 4214 43867 4216
rect 43891 4214 43947 4216
rect 43971 4214 44027 4216
rect 44051 4214 44107 4216
rect 44131 4214 44187 4216
rect 44211 4214 44267 4216
rect 44291 4214 44347 4216
rect 44371 4214 44427 4216
rect 44451 4214 44507 4216
rect 44531 4214 44587 4216
rect 44611 4214 44667 4216
rect 44691 4214 44747 4216
rect 44771 4214 44827 4216
rect 44851 4214 44907 4216
rect 44931 4214 44987 4216
rect 45011 4214 45067 4216
rect 45091 4214 45147 4216
rect 45171 4214 45227 4216
rect 45251 4214 45307 4216
rect 45331 4214 45387 4216
rect 45411 4214 45467 4216
rect 45491 4214 45547 4216
rect 45571 4214 45627 4216
rect 45651 4214 45707 4216
rect 45731 4214 45787 4216
rect 45811 4214 45867 4216
rect 45891 4214 45947 4216
rect 42611 4162 42621 4214
rect 42621 4162 42667 4214
rect 42691 4162 42737 4214
rect 42737 4162 42747 4214
rect 42771 4162 42801 4214
rect 42801 4162 42813 4214
rect 42813 4162 42827 4214
rect 42851 4162 42865 4214
rect 42865 4162 42877 4214
rect 42877 4162 42907 4214
rect 42931 4162 42941 4214
rect 42941 4162 42987 4214
rect 43011 4162 43057 4214
rect 43057 4162 43067 4214
rect 43091 4162 43121 4214
rect 43121 4162 43133 4214
rect 43133 4162 43147 4214
rect 43171 4162 43185 4214
rect 43185 4162 43197 4214
rect 43197 4162 43227 4214
rect 43251 4162 43261 4214
rect 43261 4162 43307 4214
rect 43331 4162 43377 4214
rect 43377 4162 43387 4214
rect 43411 4162 43441 4214
rect 43441 4162 43453 4214
rect 43453 4162 43467 4214
rect 43491 4162 43505 4214
rect 43505 4162 43517 4214
rect 43517 4162 43547 4214
rect 43571 4162 43581 4214
rect 43581 4162 43627 4214
rect 43651 4162 43697 4214
rect 43697 4162 43707 4214
rect 43731 4162 43761 4214
rect 43761 4162 43773 4214
rect 43773 4162 43787 4214
rect 43811 4162 43825 4214
rect 43825 4162 43837 4214
rect 43837 4162 43867 4214
rect 43891 4162 43901 4214
rect 43901 4162 43947 4214
rect 43971 4162 44017 4214
rect 44017 4162 44027 4214
rect 44051 4162 44081 4214
rect 44081 4162 44093 4214
rect 44093 4162 44107 4214
rect 44131 4162 44145 4214
rect 44145 4162 44157 4214
rect 44157 4162 44187 4214
rect 44211 4162 44221 4214
rect 44221 4162 44267 4214
rect 44291 4162 44337 4214
rect 44337 4162 44347 4214
rect 44371 4162 44401 4214
rect 44401 4162 44413 4214
rect 44413 4162 44427 4214
rect 44451 4162 44465 4214
rect 44465 4162 44477 4214
rect 44477 4162 44507 4214
rect 44531 4162 44541 4214
rect 44541 4162 44587 4214
rect 44611 4162 44657 4214
rect 44657 4162 44667 4214
rect 44691 4162 44721 4214
rect 44721 4162 44733 4214
rect 44733 4162 44747 4214
rect 44771 4162 44785 4214
rect 44785 4162 44797 4214
rect 44797 4162 44827 4214
rect 44851 4162 44861 4214
rect 44861 4162 44907 4214
rect 44931 4162 44977 4214
rect 44977 4162 44987 4214
rect 45011 4162 45041 4214
rect 45041 4162 45053 4214
rect 45053 4162 45067 4214
rect 45091 4162 45105 4214
rect 45105 4162 45117 4214
rect 45117 4162 45147 4214
rect 45171 4162 45181 4214
rect 45181 4162 45227 4214
rect 45251 4162 45297 4214
rect 45297 4162 45307 4214
rect 45331 4162 45361 4214
rect 45361 4162 45373 4214
rect 45373 4162 45387 4214
rect 45411 4162 45425 4214
rect 45425 4162 45437 4214
rect 45437 4162 45467 4214
rect 45491 4162 45501 4214
rect 45501 4162 45547 4214
rect 45571 4162 45617 4214
rect 45617 4162 45627 4214
rect 45651 4162 45681 4214
rect 45681 4162 45693 4214
rect 45693 4162 45707 4214
rect 45731 4162 45745 4214
rect 45745 4162 45757 4214
rect 45757 4162 45787 4214
rect 45811 4162 45821 4214
rect 45821 4162 45867 4214
rect 45891 4162 45937 4214
rect 45937 4162 45947 4214
rect 42611 4160 42667 4162
rect 42691 4160 42747 4162
rect 42771 4160 42827 4162
rect 42851 4160 42907 4162
rect 42931 4160 42987 4162
rect 43011 4160 43067 4162
rect 43091 4160 43147 4162
rect 43171 4160 43227 4162
rect 43251 4160 43307 4162
rect 43331 4160 43387 4162
rect 43411 4160 43467 4162
rect 43491 4160 43547 4162
rect 43571 4160 43627 4162
rect 43651 4160 43707 4162
rect 43731 4160 43787 4162
rect 43811 4160 43867 4162
rect 43891 4160 43947 4162
rect 43971 4160 44027 4162
rect 44051 4160 44107 4162
rect 44131 4160 44187 4162
rect 44211 4160 44267 4162
rect 44291 4160 44347 4162
rect 44371 4160 44427 4162
rect 44451 4160 44507 4162
rect 44531 4160 44587 4162
rect 44611 4160 44667 4162
rect 44691 4160 44747 4162
rect 44771 4160 44827 4162
rect 44851 4160 44907 4162
rect 44931 4160 44987 4162
rect 45011 4160 45067 4162
rect 45091 4160 45147 4162
rect 45171 4160 45227 4162
rect 45251 4160 45307 4162
rect 45331 4160 45387 4162
rect 45411 4160 45467 4162
rect 45491 4160 45547 4162
rect 45571 4160 45627 4162
rect 45651 4160 45707 4162
rect 45731 4160 45787 4162
rect 45811 4160 45867 4162
rect 45891 4160 45947 4162
rect 36992 4067 37048 4069
rect 36992 4015 36994 4067
rect 36994 4015 37046 4067
rect 37046 4015 37048 4067
rect 36992 4013 37048 4015
rect 40111 3970 40113 4000
rect 40113 3970 40165 4000
rect 40165 3970 40167 4000
rect 40111 3958 40167 3970
rect 40111 3944 40113 3958
rect 40113 3944 40165 3958
rect 40165 3944 40167 3958
rect 38583 3915 38639 3925
rect 38583 3869 38585 3915
rect 38585 3869 38637 3915
rect 38637 3869 38639 3915
rect 38583 3799 38585 3845
rect 38585 3799 38637 3845
rect 38637 3799 38639 3845
rect 38583 3789 38639 3799
rect 40111 3906 40113 3920
rect 40113 3906 40165 3920
rect 40165 3906 40167 3920
rect 40111 3894 40167 3906
rect 40111 3864 40113 3894
rect 40113 3864 40165 3894
rect 40165 3864 40167 3894
rect 36394 3521 36450 3523
rect 36394 3469 36416 3521
rect 36416 3469 36428 3521
rect 36428 3469 36450 3521
rect 36394 3467 36450 3469
rect 38577 3423 38579 3453
rect 38579 3423 38631 3453
rect 38631 3423 38633 3453
rect 38577 3411 38633 3423
rect 38577 3397 38579 3411
rect 38579 3397 38631 3411
rect 38631 3397 38633 3411
rect 38577 3359 38579 3373
rect 38579 3359 38631 3373
rect 38631 3359 38633 3373
rect 38577 3347 38633 3359
rect 38577 3317 38579 3347
rect 38579 3317 38631 3347
rect 38631 3317 38633 3347
rect 40101 3417 40103 3447
rect 40103 3417 40155 3447
rect 40155 3417 40157 3447
rect 40101 3405 40157 3417
rect 40101 3391 40103 3405
rect 40103 3391 40155 3405
rect 40155 3391 40157 3405
rect 40101 3353 40103 3367
rect 40103 3353 40155 3367
rect 40155 3353 40157 3367
rect 40101 3341 40157 3353
rect 40101 3311 40103 3341
rect 40103 3311 40155 3341
rect 40155 3311 40157 3341
rect 35035 3116 35091 3118
rect 35035 3064 35037 3116
rect 35037 3064 35089 3116
rect 35089 3064 35091 3116
rect 35035 3062 35091 3064
rect 35493 1531 35549 1587
rect 36070 2154 36126 2210
rect 36635 1469 36691 1525
rect 35028 1337 35084 1339
rect 35028 1285 35030 1337
rect 35030 1285 35082 1337
rect 35082 1285 35084 1337
rect 35028 1283 35084 1285
rect 38582 1083 38638 1093
rect 38582 1037 38584 1083
rect 38584 1037 38636 1083
rect 38636 1037 38638 1083
rect 38582 967 38584 1013
rect 38584 967 38636 1013
rect 38636 967 38638 1013
rect 38582 957 38638 967
rect 40112 1125 40114 1155
rect 40114 1125 40166 1155
rect 40166 1125 40168 1155
rect 40112 1113 40168 1125
rect 40112 1099 40114 1113
rect 40114 1099 40166 1113
rect 40166 1099 40168 1113
rect 40112 1061 40114 1075
rect 40114 1061 40166 1075
rect 40166 1061 40168 1075
rect 40112 1049 40168 1061
rect 40112 1019 40114 1049
rect 40114 1019 40166 1049
rect 40166 1019 40168 1049
rect 36308 933 36364 935
rect 36388 933 36444 935
rect 36468 933 36524 935
rect 36308 881 36326 933
rect 36326 881 36364 933
rect 36388 881 36390 933
rect 36390 881 36442 933
rect 36442 881 36444 933
rect 36468 881 36506 933
rect 36506 881 36524 933
rect 36308 879 36364 881
rect 36388 879 36444 881
rect 36468 879 36524 881
rect 38580 567 38582 597
rect 38582 567 38634 597
rect 38634 567 38636 597
rect 38580 555 38636 567
rect 38580 541 38582 555
rect 38582 541 38634 555
rect 38634 541 38636 555
rect 38580 503 38582 517
rect 38582 503 38634 517
rect 38634 503 38636 517
rect 38580 491 38636 503
rect 38580 461 38582 491
rect 38582 461 38634 491
rect 38634 461 38636 491
rect 40099 580 40101 610
rect 40101 580 40153 610
rect 40153 580 40155 610
rect 40099 568 40155 580
rect 40099 554 40101 568
rect 40101 554 40153 568
rect 40153 554 40155 568
rect 40099 516 40101 530
rect 40101 516 40153 530
rect 40153 516 40155 530
rect 40099 504 40155 516
rect 40099 474 40101 504
rect 40101 474 40153 504
rect 40153 474 40155 504
rect 36378 392 36434 394
rect 36458 392 36514 394
rect 36378 340 36388 392
rect 36388 340 36434 392
rect 36458 340 36504 392
rect 36504 340 36514 392
rect 36378 338 36434 340
rect 36458 338 36514 340
rect 326 207 21102 217
rect 326 91 352 207
rect 352 91 21076 207
rect 21076 91 21102 207
rect 326 81 21102 91
rect 35032 277 35088 279
rect 35032 225 35034 277
rect 35034 225 35086 277
rect 35086 225 35088 277
rect 35032 223 35088 225
rect 42636 280 42692 282
rect 42716 280 42772 282
rect 42796 280 42852 282
rect 42876 280 42932 282
rect 42956 280 43012 282
rect 43036 280 43092 282
rect 43116 280 43172 282
rect 43196 280 43252 282
rect 43276 280 43332 282
rect 43356 280 43412 282
rect 43436 280 43492 282
rect 43516 280 43572 282
rect 43596 280 43652 282
rect 43676 280 43732 282
rect 43756 280 43812 282
rect 43836 280 43892 282
rect 43916 280 43972 282
rect 43996 280 44052 282
rect 44076 280 44132 282
rect 44156 280 44212 282
rect 44236 280 44292 282
rect 44316 280 44372 282
rect 44396 280 44452 282
rect 44476 280 44532 282
rect 44556 280 44612 282
rect 44636 280 44692 282
rect 44716 280 44772 282
rect 44796 280 44852 282
rect 44876 280 44932 282
rect 44956 280 45012 282
rect 45036 280 45092 282
rect 45116 280 45172 282
rect 45196 280 45252 282
rect 45276 280 45332 282
rect 45356 280 45412 282
rect 45436 280 45492 282
rect 45516 280 45572 282
rect 45596 280 45652 282
rect 45676 280 45732 282
rect 45756 280 45812 282
rect 45836 280 45892 282
rect 42636 228 42658 280
rect 42658 228 42670 280
rect 42670 228 42692 280
rect 42716 228 42722 280
rect 42722 228 42734 280
rect 42734 228 42772 280
rect 42796 228 42798 280
rect 42798 228 42850 280
rect 42850 228 42852 280
rect 42876 228 42914 280
rect 42914 228 42926 280
rect 42926 228 42932 280
rect 42956 228 42978 280
rect 42978 228 42990 280
rect 42990 228 43012 280
rect 43036 228 43042 280
rect 43042 228 43054 280
rect 43054 228 43092 280
rect 43116 228 43118 280
rect 43118 228 43170 280
rect 43170 228 43172 280
rect 43196 228 43234 280
rect 43234 228 43246 280
rect 43246 228 43252 280
rect 43276 228 43298 280
rect 43298 228 43310 280
rect 43310 228 43332 280
rect 43356 228 43362 280
rect 43362 228 43374 280
rect 43374 228 43412 280
rect 43436 228 43438 280
rect 43438 228 43490 280
rect 43490 228 43492 280
rect 43516 228 43554 280
rect 43554 228 43566 280
rect 43566 228 43572 280
rect 43596 228 43618 280
rect 43618 228 43630 280
rect 43630 228 43652 280
rect 43676 228 43682 280
rect 43682 228 43694 280
rect 43694 228 43732 280
rect 43756 228 43758 280
rect 43758 228 43810 280
rect 43810 228 43812 280
rect 43836 228 43874 280
rect 43874 228 43886 280
rect 43886 228 43892 280
rect 43916 228 43938 280
rect 43938 228 43950 280
rect 43950 228 43972 280
rect 43996 228 44002 280
rect 44002 228 44014 280
rect 44014 228 44052 280
rect 44076 228 44078 280
rect 44078 228 44130 280
rect 44130 228 44132 280
rect 44156 228 44194 280
rect 44194 228 44206 280
rect 44206 228 44212 280
rect 44236 228 44258 280
rect 44258 228 44270 280
rect 44270 228 44292 280
rect 44316 228 44322 280
rect 44322 228 44334 280
rect 44334 228 44372 280
rect 44396 228 44398 280
rect 44398 228 44450 280
rect 44450 228 44452 280
rect 44476 228 44514 280
rect 44514 228 44526 280
rect 44526 228 44532 280
rect 44556 228 44578 280
rect 44578 228 44590 280
rect 44590 228 44612 280
rect 44636 228 44642 280
rect 44642 228 44654 280
rect 44654 228 44692 280
rect 44716 228 44718 280
rect 44718 228 44770 280
rect 44770 228 44772 280
rect 44796 228 44834 280
rect 44834 228 44846 280
rect 44846 228 44852 280
rect 44876 228 44898 280
rect 44898 228 44910 280
rect 44910 228 44932 280
rect 44956 228 44962 280
rect 44962 228 44974 280
rect 44974 228 45012 280
rect 45036 228 45038 280
rect 45038 228 45090 280
rect 45090 228 45092 280
rect 45116 228 45154 280
rect 45154 228 45166 280
rect 45166 228 45172 280
rect 45196 228 45218 280
rect 45218 228 45230 280
rect 45230 228 45252 280
rect 45276 228 45282 280
rect 45282 228 45294 280
rect 45294 228 45332 280
rect 45356 228 45358 280
rect 45358 228 45410 280
rect 45410 228 45412 280
rect 45436 228 45474 280
rect 45474 228 45486 280
rect 45486 228 45492 280
rect 45516 228 45538 280
rect 45538 228 45550 280
rect 45550 228 45572 280
rect 45596 228 45602 280
rect 45602 228 45614 280
rect 45614 228 45652 280
rect 45676 228 45678 280
rect 45678 228 45730 280
rect 45730 228 45732 280
rect 45756 228 45794 280
rect 45794 228 45806 280
rect 45806 228 45812 280
rect 45836 228 45858 280
rect 45858 228 45870 280
rect 45870 228 45892 280
rect 42636 226 42692 228
rect 42716 226 42772 228
rect 42796 226 42852 228
rect 42876 226 42932 228
rect 42956 226 43012 228
rect 43036 226 43092 228
rect 43116 226 43172 228
rect 43196 226 43252 228
rect 43276 226 43332 228
rect 43356 226 43412 228
rect 43436 226 43492 228
rect 43516 226 43572 228
rect 43596 226 43652 228
rect 43676 226 43732 228
rect 43756 226 43812 228
rect 43836 226 43892 228
rect 43916 226 43972 228
rect 43996 226 44052 228
rect 44076 226 44132 228
rect 44156 226 44212 228
rect 44236 226 44292 228
rect 44316 226 44372 228
rect 44396 226 44452 228
rect 44476 226 44532 228
rect 44556 226 44612 228
rect 44636 226 44692 228
rect 44716 226 44772 228
rect 44796 226 44852 228
rect 44876 226 44932 228
rect 44956 226 45012 228
rect 45036 226 45092 228
rect 45116 226 45172 228
rect 45196 226 45252 228
rect 45276 226 45332 228
rect 45356 226 45412 228
rect 45436 226 45492 228
rect 45516 226 45572 228
rect 45596 226 45652 228
rect 45676 226 45732 228
rect 45756 226 45812 228
rect 45836 226 45892 228
rect 35031 8 35087 10
rect 35031 -44 35033 8
rect 35033 -44 35085 8
rect 35085 -44 35087 8
rect 35031 -46 35087 -44
rect 36366 -156 36422 -154
rect 36366 -208 36368 -156
rect 36368 -208 36420 -156
rect 36420 -208 36422 -156
rect 36366 -210 36422 -208
rect 38582 -290 38584 -268
rect 38584 -290 38636 -268
rect 38636 -290 38638 -268
rect 38582 -302 38638 -290
rect 38582 -324 38584 -302
rect 38584 -324 38636 -302
rect 38636 -324 38638 -302
rect 40104 -211 40106 -181
rect 40106 -211 40158 -181
rect 40158 -211 40160 -181
rect 40104 -223 40160 -211
rect 40104 -237 40106 -223
rect 40106 -237 40158 -223
rect 40158 -237 40160 -223
rect 40104 -275 40106 -261
rect 40106 -275 40158 -261
rect 40158 -275 40160 -261
rect 40104 -287 40160 -275
rect 40104 -317 40106 -287
rect 40106 -317 40158 -287
rect 40158 -317 40160 -287
rect 36991 -697 37047 -695
rect 36991 -749 36993 -697
rect 36993 -749 37045 -697
rect 37045 -749 37047 -697
rect 36991 -751 37047 -749
rect 38575 -764 38577 -734
rect 38577 -764 38629 -734
rect 38629 -764 38631 -734
rect 38575 -776 38631 -764
rect 38575 -790 38577 -776
rect 38577 -790 38629 -776
rect 38629 -790 38631 -776
rect 38575 -828 38577 -814
rect 38577 -828 38629 -814
rect 38629 -828 38631 -814
rect 38575 -840 38631 -828
rect 38575 -870 38577 -840
rect 38577 -870 38629 -840
rect 38629 -870 38631 -840
rect 40104 -767 40106 -737
rect 40106 -767 40158 -737
rect 40158 -767 40160 -737
rect 40104 -779 40160 -767
rect 40104 -793 40106 -779
rect 40106 -793 40158 -779
rect 40158 -793 40160 -779
rect 40104 -831 40106 -817
rect 40106 -831 40158 -817
rect 40158 -831 40160 -817
rect 40104 -843 40160 -831
rect 40104 -873 40106 -843
rect 40106 -873 40158 -843
rect 40158 -873 40160 -843
rect 35031 -1061 35087 -1059
rect 35031 -1113 35033 -1061
rect 35033 -1113 35085 -1061
rect 35085 -1113 35087 -1061
rect 35031 -1115 35087 -1113
rect 35991 -1239 36047 -1237
rect 36071 -1239 36127 -1237
rect 35991 -1291 36001 -1239
rect 36001 -1291 36047 -1239
rect 36071 -1291 36117 -1239
rect 36117 -1291 36127 -1239
rect 35991 -1293 36047 -1291
rect 36071 -1293 36127 -1291
rect 47499 -1168 47715 -1150
rect 47499 -1348 47517 -1168
rect 47517 -1348 47697 -1168
rect 47697 -1348 47715 -1168
rect 47499 -1366 47715 -1348
rect 35028 -1384 35084 -1382
rect 35028 -1436 35030 -1384
rect 35030 -1436 35082 -1384
rect 35082 -1436 35084 -1384
rect 35028 -1438 35084 -1436
rect 38583 -1680 38585 -1658
rect 38585 -1680 38637 -1658
rect 38637 -1680 38639 -1658
rect 38583 -1692 38639 -1680
rect 38583 -1714 38585 -1692
rect 38585 -1714 38637 -1692
rect 38637 -1714 38639 -1692
rect 40121 -1591 40123 -1561
rect 40123 -1591 40175 -1561
rect 40175 -1591 40177 -1561
rect 40121 -1603 40177 -1591
rect 40121 -1617 40123 -1603
rect 40123 -1617 40175 -1603
rect 40175 -1617 40177 -1603
rect 40121 -1655 40123 -1641
rect 40123 -1655 40175 -1641
rect 40175 -1655 40177 -1641
rect 40121 -1667 40177 -1655
rect 40121 -1697 40123 -1667
rect 40123 -1697 40175 -1667
rect 40175 -1697 40177 -1667
rect 36516 -1787 36572 -1785
rect 36596 -1787 36652 -1785
rect 36676 -1787 36732 -1785
rect 36516 -1839 36534 -1787
rect 36534 -1839 36572 -1787
rect 36596 -1839 36598 -1787
rect 36598 -1839 36650 -1787
rect 36650 -1839 36652 -1787
rect 36676 -1839 36714 -1787
rect 36714 -1839 36732 -1787
rect 36516 -1841 36572 -1839
rect 36596 -1841 36652 -1839
rect 36676 -1841 36732 -1839
rect 38574 -2117 38576 -2087
rect 38576 -2117 38628 -2087
rect 38628 -2117 38630 -2087
rect 38574 -2129 38630 -2117
rect 38574 -2143 38576 -2129
rect 38576 -2143 38628 -2129
rect 38628 -2143 38630 -2129
rect 38574 -2181 38576 -2167
rect 38576 -2181 38628 -2167
rect 38628 -2181 38630 -2167
rect 38574 -2193 38630 -2181
rect 38574 -2223 38576 -2193
rect 38576 -2223 38628 -2193
rect 38628 -2223 38630 -2193
rect 40104 -2139 40106 -2109
rect 40106 -2139 40158 -2109
rect 40158 -2139 40160 -2109
rect 40104 -2151 40160 -2139
rect 40104 -2165 40106 -2151
rect 40106 -2165 40158 -2151
rect 40158 -2165 40160 -2151
rect 40104 -2203 40106 -2189
rect 40106 -2203 40158 -2189
rect 40158 -2203 40160 -2189
rect 40104 -2215 40160 -2203
rect 40104 -2245 40106 -2215
rect 40106 -2245 40158 -2215
rect 40158 -2245 40160 -2215
rect 36368 -2330 36424 -2328
rect 36448 -2330 36504 -2328
rect 36368 -2382 36378 -2330
rect 36378 -2382 36424 -2330
rect 36448 -2382 36494 -2330
rect 36494 -2382 36504 -2330
rect 36368 -2384 36424 -2382
rect 36448 -2384 36504 -2382
rect 35039 -2454 35095 -2452
rect 35039 -2506 35041 -2454
rect 35041 -2506 35093 -2454
rect 35093 -2506 35095 -2454
rect 35039 -2508 35095 -2506
rect 35028 -2759 35084 -2757
rect 35028 -2811 35030 -2759
rect 35030 -2811 35082 -2759
rect 35082 -2811 35084 -2759
rect 35028 -2813 35084 -2811
rect 42592 -2726 42648 -2724
rect 42672 -2726 42728 -2724
rect 42752 -2726 42808 -2724
rect 42832 -2726 42888 -2724
rect 42912 -2726 42968 -2724
rect 42992 -2726 43048 -2724
rect 43072 -2726 43128 -2724
rect 43152 -2726 43208 -2724
rect 43232 -2726 43288 -2724
rect 43312 -2726 43368 -2724
rect 43392 -2726 43448 -2724
rect 43472 -2726 43528 -2724
rect 43552 -2726 43608 -2724
rect 43632 -2726 43688 -2724
rect 43712 -2726 43768 -2724
rect 43792 -2726 43848 -2724
rect 43872 -2726 43928 -2724
rect 43952 -2726 44008 -2724
rect 44032 -2726 44088 -2724
rect 44112 -2726 44168 -2724
rect 44192 -2726 44248 -2724
rect 44272 -2726 44328 -2724
rect 44352 -2726 44408 -2724
rect 44432 -2726 44488 -2724
rect 44512 -2726 44568 -2724
rect 44592 -2726 44648 -2724
rect 44672 -2726 44728 -2724
rect 44752 -2726 44808 -2724
rect 44832 -2726 44888 -2724
rect 44912 -2726 44968 -2724
rect 44992 -2726 45048 -2724
rect 45072 -2726 45128 -2724
rect 45152 -2726 45208 -2724
rect 45232 -2726 45288 -2724
rect 45312 -2726 45368 -2724
rect 45392 -2726 45448 -2724
rect 45472 -2726 45528 -2724
rect 45552 -2726 45608 -2724
rect 45632 -2726 45688 -2724
rect 45712 -2726 45768 -2724
rect 45792 -2726 45848 -2724
rect 45872 -2726 45928 -2724
rect 42592 -2778 42602 -2726
rect 42602 -2778 42648 -2726
rect 42672 -2778 42718 -2726
rect 42718 -2778 42728 -2726
rect 42752 -2778 42782 -2726
rect 42782 -2778 42794 -2726
rect 42794 -2778 42808 -2726
rect 42832 -2778 42846 -2726
rect 42846 -2778 42858 -2726
rect 42858 -2778 42888 -2726
rect 42912 -2778 42922 -2726
rect 42922 -2778 42968 -2726
rect 42992 -2778 43038 -2726
rect 43038 -2778 43048 -2726
rect 43072 -2778 43102 -2726
rect 43102 -2778 43114 -2726
rect 43114 -2778 43128 -2726
rect 43152 -2778 43166 -2726
rect 43166 -2778 43178 -2726
rect 43178 -2778 43208 -2726
rect 43232 -2778 43242 -2726
rect 43242 -2778 43288 -2726
rect 43312 -2778 43358 -2726
rect 43358 -2778 43368 -2726
rect 43392 -2778 43422 -2726
rect 43422 -2778 43434 -2726
rect 43434 -2778 43448 -2726
rect 43472 -2778 43486 -2726
rect 43486 -2778 43498 -2726
rect 43498 -2778 43528 -2726
rect 43552 -2778 43562 -2726
rect 43562 -2778 43608 -2726
rect 43632 -2778 43678 -2726
rect 43678 -2778 43688 -2726
rect 43712 -2778 43742 -2726
rect 43742 -2778 43754 -2726
rect 43754 -2778 43768 -2726
rect 43792 -2778 43806 -2726
rect 43806 -2778 43818 -2726
rect 43818 -2778 43848 -2726
rect 43872 -2778 43882 -2726
rect 43882 -2778 43928 -2726
rect 43952 -2778 43998 -2726
rect 43998 -2778 44008 -2726
rect 44032 -2778 44062 -2726
rect 44062 -2778 44074 -2726
rect 44074 -2778 44088 -2726
rect 44112 -2778 44126 -2726
rect 44126 -2778 44138 -2726
rect 44138 -2778 44168 -2726
rect 44192 -2778 44202 -2726
rect 44202 -2778 44248 -2726
rect 44272 -2778 44318 -2726
rect 44318 -2778 44328 -2726
rect 44352 -2778 44382 -2726
rect 44382 -2778 44394 -2726
rect 44394 -2778 44408 -2726
rect 44432 -2778 44446 -2726
rect 44446 -2778 44458 -2726
rect 44458 -2778 44488 -2726
rect 44512 -2778 44522 -2726
rect 44522 -2778 44568 -2726
rect 44592 -2778 44638 -2726
rect 44638 -2778 44648 -2726
rect 44672 -2778 44702 -2726
rect 44702 -2778 44714 -2726
rect 44714 -2778 44728 -2726
rect 44752 -2778 44766 -2726
rect 44766 -2778 44778 -2726
rect 44778 -2778 44808 -2726
rect 44832 -2778 44842 -2726
rect 44842 -2778 44888 -2726
rect 44912 -2778 44958 -2726
rect 44958 -2778 44968 -2726
rect 44992 -2778 45022 -2726
rect 45022 -2778 45034 -2726
rect 45034 -2778 45048 -2726
rect 45072 -2778 45086 -2726
rect 45086 -2778 45098 -2726
rect 45098 -2778 45128 -2726
rect 45152 -2778 45162 -2726
rect 45162 -2778 45208 -2726
rect 45232 -2778 45278 -2726
rect 45278 -2778 45288 -2726
rect 45312 -2778 45342 -2726
rect 45342 -2778 45354 -2726
rect 45354 -2778 45368 -2726
rect 45392 -2778 45406 -2726
rect 45406 -2778 45418 -2726
rect 45418 -2778 45448 -2726
rect 45472 -2778 45482 -2726
rect 45482 -2778 45528 -2726
rect 45552 -2778 45598 -2726
rect 45598 -2778 45608 -2726
rect 45632 -2778 45662 -2726
rect 45662 -2778 45674 -2726
rect 45674 -2778 45688 -2726
rect 45712 -2778 45726 -2726
rect 45726 -2778 45738 -2726
rect 45738 -2778 45768 -2726
rect 45792 -2778 45802 -2726
rect 45802 -2778 45848 -2726
rect 45872 -2778 45918 -2726
rect 45918 -2778 45928 -2726
rect 42592 -2780 42648 -2778
rect 42672 -2780 42728 -2778
rect 42752 -2780 42808 -2778
rect 42832 -2780 42888 -2778
rect 42912 -2780 42968 -2778
rect 42992 -2780 43048 -2778
rect 43072 -2780 43128 -2778
rect 43152 -2780 43208 -2778
rect 43232 -2780 43288 -2778
rect 43312 -2780 43368 -2778
rect 43392 -2780 43448 -2778
rect 43472 -2780 43528 -2778
rect 43552 -2780 43608 -2778
rect 43632 -2780 43688 -2778
rect 43712 -2780 43768 -2778
rect 43792 -2780 43848 -2778
rect 43872 -2780 43928 -2778
rect 43952 -2780 44008 -2778
rect 44032 -2780 44088 -2778
rect 44112 -2780 44168 -2778
rect 44192 -2780 44248 -2778
rect 44272 -2780 44328 -2778
rect 44352 -2780 44408 -2778
rect 44432 -2780 44488 -2778
rect 44512 -2780 44568 -2778
rect 44592 -2780 44648 -2778
rect 44672 -2780 44728 -2778
rect 44752 -2780 44808 -2778
rect 44832 -2780 44888 -2778
rect 44912 -2780 44968 -2778
rect 44992 -2780 45048 -2778
rect 45072 -2780 45128 -2778
rect 45152 -2780 45208 -2778
rect 45232 -2780 45288 -2778
rect 45312 -2780 45368 -2778
rect 45392 -2780 45448 -2778
rect 45472 -2780 45528 -2778
rect 45552 -2780 45608 -2778
rect 45632 -2780 45688 -2778
rect 45712 -2780 45768 -2778
rect 45792 -2780 45848 -2778
rect 45872 -2780 45928 -2778
rect 36992 -2873 37048 -2871
rect 36992 -2925 36994 -2873
rect 36994 -2925 37046 -2873
rect 37046 -2925 37048 -2873
rect 36992 -2927 37048 -2925
rect 40111 -2970 40113 -2940
rect 40113 -2970 40165 -2940
rect 40165 -2970 40167 -2940
rect 40111 -2982 40167 -2970
rect 40111 -2996 40113 -2982
rect 40113 -2996 40165 -2982
rect 40165 -2996 40167 -2982
rect 38583 -3025 38639 -3015
rect 38583 -3071 38585 -3025
rect 38585 -3071 38637 -3025
rect 38637 -3071 38639 -3025
rect 38583 -3141 38585 -3095
rect 38585 -3141 38637 -3095
rect 38637 -3141 38639 -3095
rect 38583 -3151 38639 -3141
rect 40111 -3034 40113 -3020
rect 40113 -3034 40165 -3020
rect 40165 -3034 40167 -3020
rect 40111 -3046 40167 -3034
rect 40111 -3076 40113 -3046
rect 40113 -3076 40165 -3046
rect 40165 -3076 40167 -3046
rect 36394 -3419 36450 -3417
rect 36394 -3471 36416 -3419
rect 36416 -3471 36428 -3419
rect 36428 -3471 36450 -3419
rect 36394 -3473 36450 -3471
rect 38577 -3517 38579 -3487
rect 38579 -3517 38631 -3487
rect 38631 -3517 38633 -3487
rect 38577 -3529 38633 -3517
rect 38577 -3543 38579 -3529
rect 38579 -3543 38631 -3529
rect 38631 -3543 38633 -3529
rect 38577 -3581 38579 -3567
rect 38579 -3581 38631 -3567
rect 38631 -3581 38633 -3567
rect 38577 -3593 38633 -3581
rect 38577 -3623 38579 -3593
rect 38579 -3623 38631 -3593
rect 38631 -3623 38633 -3593
rect 40101 -3523 40103 -3493
rect 40103 -3523 40155 -3493
rect 40155 -3523 40157 -3493
rect 40101 -3535 40157 -3523
rect 40101 -3549 40103 -3535
rect 40103 -3549 40155 -3535
rect 40155 -3549 40157 -3535
rect 40101 -3587 40103 -3573
rect 40103 -3587 40155 -3573
rect 40155 -3587 40157 -3573
rect 40101 -3599 40157 -3587
rect 40101 -3629 40103 -3599
rect 40103 -3629 40155 -3599
rect 40155 -3629 40157 -3599
rect 35035 -3824 35091 -3822
rect 35035 -3876 35037 -3824
rect 35037 -3876 35089 -3824
rect 35089 -3876 35091 -3824
rect 35035 -3878 35091 -3876
rect -3577 -6850 -3521 -6848
rect -3577 -6902 -3575 -6850
rect -3575 -6902 -3523 -6850
rect -3523 -6902 -3521 -6850
rect -3577 -6904 -3521 -6902
rect -3577 -6966 -3575 -6928
rect -3575 -6966 -3523 -6928
rect -3523 -6966 -3521 -6928
rect -3577 -6978 -3521 -6966
rect -3577 -6984 -3575 -6978
rect -3575 -6984 -3523 -6978
rect -3523 -6984 -3521 -6978
rect -3577 -7030 -3575 -7008
rect -3575 -7030 -3523 -7008
rect -3523 -7030 -3521 -7008
rect -3577 -7042 -3521 -7030
rect -3577 -7064 -3575 -7042
rect -3575 -7064 -3523 -7042
rect -3523 -7064 -3521 -7042
rect -3577 -7094 -3575 -7088
rect -3575 -7094 -3523 -7088
rect -3523 -7094 -3521 -7088
rect -3577 -7106 -3521 -7094
rect -3577 -7144 -3575 -7106
rect -3575 -7144 -3523 -7106
rect -3523 -7144 -3521 -7106
rect -3577 -7170 -3521 -7168
rect -3577 -7222 -3575 -7170
rect -3575 -7222 -3523 -7170
rect -3523 -7222 -3521 -7170
rect -3577 -7224 -3521 -7222
rect -3577 -7286 -3575 -7248
rect -3575 -7286 -3523 -7248
rect -3523 -7286 -3521 -7248
rect -3577 -7298 -3521 -7286
rect -3577 -7304 -3575 -7298
rect -3575 -7304 -3523 -7298
rect -3523 -7304 -3521 -7298
rect -3577 -7350 -3575 -7328
rect -3575 -7350 -3523 -7328
rect -3523 -7350 -3521 -7328
rect -3577 -7362 -3521 -7350
rect -3577 -7384 -3575 -7362
rect -3575 -7384 -3523 -7362
rect -3523 -7384 -3521 -7362
rect -3577 -7414 -3575 -7408
rect -3575 -7414 -3523 -7408
rect -3523 -7414 -3521 -7408
rect -3577 -7426 -3521 -7414
rect -3577 -7464 -3575 -7426
rect -3575 -7464 -3523 -7426
rect -3523 -7464 -3521 -7426
rect -3577 -7490 -3521 -7488
rect -3577 -7542 -3575 -7490
rect -3575 -7542 -3523 -7490
rect -3523 -7542 -3521 -7490
rect -3577 -7544 -3521 -7542
rect -3577 -7606 -3575 -7568
rect -3575 -7606 -3523 -7568
rect -3523 -7606 -3521 -7568
rect -3577 -7618 -3521 -7606
rect -3577 -7624 -3575 -7618
rect -3575 -7624 -3523 -7618
rect -3523 -7624 -3521 -7618
rect -3577 -7670 -3575 -7648
rect -3575 -7670 -3523 -7648
rect -3523 -7670 -3521 -7648
rect -3577 -7682 -3521 -7670
rect -3577 -7704 -3575 -7682
rect -3575 -7704 -3523 -7682
rect -3523 -7704 -3521 -7682
rect -3577 -7734 -3575 -7728
rect -3575 -7734 -3523 -7728
rect -3523 -7734 -3521 -7728
rect -3577 -7746 -3521 -7734
rect -3577 -7784 -3575 -7746
rect -3575 -7784 -3523 -7746
rect -3523 -7784 -3521 -7746
rect -3577 -7810 -3521 -7808
rect -3577 -7862 -3575 -7810
rect -3575 -7862 -3523 -7810
rect -3523 -7862 -3521 -7810
rect -3577 -7864 -3521 -7862
rect -3577 -7926 -3575 -7888
rect -3575 -7926 -3523 -7888
rect -3523 -7926 -3521 -7888
rect -3577 -7938 -3521 -7926
rect -3577 -7944 -3575 -7938
rect -3575 -7944 -3523 -7938
rect -3523 -7944 -3521 -7938
rect -3577 -7990 -3575 -7968
rect -3575 -7990 -3523 -7968
rect -3523 -7990 -3521 -7968
rect -3577 -8002 -3521 -7990
rect -3577 -8024 -3575 -8002
rect -3575 -8024 -3523 -8002
rect -3523 -8024 -3521 -8002
rect -3577 -8054 -3575 -8048
rect -3575 -8054 -3523 -8048
rect -3523 -8054 -3521 -8048
rect -3577 -8066 -3521 -8054
rect -3577 -8104 -3575 -8066
rect -3575 -8104 -3523 -8066
rect -3523 -8104 -3521 -8066
rect -3577 -8130 -3521 -8128
rect -3577 -8182 -3575 -8130
rect -3575 -8182 -3523 -8130
rect -3523 -8182 -3521 -8130
rect -3577 -8184 -3521 -8182
rect -3577 -8246 -3575 -8208
rect -3575 -8246 -3523 -8208
rect -3523 -8246 -3521 -8208
rect -3577 -8258 -3521 -8246
rect -3577 -8264 -3575 -8258
rect -3575 -8264 -3523 -8258
rect -3523 -8264 -3521 -8258
rect -3577 -8310 -3575 -8288
rect -3575 -8310 -3523 -8288
rect -3523 -8310 -3521 -8288
rect -3577 -8322 -3521 -8310
rect -3577 -8344 -3575 -8322
rect -3575 -8344 -3523 -8322
rect -3523 -8344 -3521 -8322
rect -3577 -8374 -3575 -8368
rect -3575 -8374 -3523 -8368
rect -3523 -8374 -3521 -8368
rect -3577 -8386 -3521 -8374
rect -3577 -8424 -3575 -8386
rect -3575 -8424 -3523 -8386
rect -3523 -8424 -3521 -8386
rect -3577 -8450 -3521 -8448
rect -3577 -8502 -3575 -8450
rect -3575 -8502 -3523 -8450
rect -3523 -8502 -3521 -8450
rect -3577 -8504 -3521 -8502
rect -3577 -8566 -3575 -8528
rect -3575 -8566 -3523 -8528
rect -3523 -8566 -3521 -8528
rect -3577 -8578 -3521 -8566
rect -3577 -8584 -3575 -8578
rect -3575 -8584 -3523 -8578
rect -3523 -8584 -3521 -8578
rect -3577 -8630 -3575 -8608
rect -3575 -8630 -3523 -8608
rect -3523 -8630 -3521 -8608
rect -3577 -8642 -3521 -8630
rect -3577 -8664 -3575 -8642
rect -3575 -8664 -3523 -8642
rect -3523 -8664 -3521 -8642
rect -3577 -8694 -3575 -8688
rect -3575 -8694 -3523 -8688
rect -3523 -8694 -3521 -8688
rect -3577 -8706 -3521 -8694
rect -3577 -8744 -3575 -8706
rect -3575 -8744 -3523 -8706
rect -3523 -8744 -3521 -8706
rect -3577 -8770 -3521 -8768
rect -3577 -8822 -3575 -8770
rect -3575 -8822 -3523 -8770
rect -3523 -8822 -3521 -8770
rect -3577 -8824 -3521 -8822
rect -3577 -8886 -3575 -8848
rect -3575 -8886 -3523 -8848
rect -3523 -8886 -3521 -8848
rect -3577 -8898 -3521 -8886
rect -3577 -8904 -3575 -8898
rect -3575 -8904 -3523 -8898
rect -3523 -8904 -3521 -8898
rect -3577 -8950 -3575 -8928
rect -3575 -8950 -3523 -8928
rect -3523 -8950 -3521 -8928
rect -3577 -8962 -3521 -8950
rect -3577 -8984 -3575 -8962
rect -3575 -8984 -3523 -8962
rect -3523 -8984 -3521 -8962
rect -3577 -9014 -3575 -9008
rect -3575 -9014 -3523 -9008
rect -3523 -9014 -3521 -9008
rect -3577 -9026 -3521 -9014
rect -3577 -9064 -3575 -9026
rect -3575 -9064 -3523 -9026
rect -3523 -9064 -3521 -9026
rect -3577 -9090 -3521 -9088
rect -3577 -9142 -3575 -9090
rect -3575 -9142 -3523 -9090
rect -3523 -9142 -3521 -9090
rect -3577 -9144 -3521 -9142
rect -3577 -9206 -3575 -9168
rect -3575 -9206 -3523 -9168
rect -3523 -9206 -3521 -9168
rect -3577 -9218 -3521 -9206
rect -3577 -9224 -3575 -9218
rect -3575 -9224 -3523 -9218
rect -3523 -9224 -3521 -9218
rect -3577 -9270 -3575 -9248
rect -3575 -9270 -3523 -9248
rect -3523 -9270 -3521 -9248
rect -3577 -9282 -3521 -9270
rect -3577 -9304 -3575 -9282
rect -3575 -9304 -3523 -9282
rect -3523 -9304 -3521 -9282
rect -3577 -9334 -3575 -9328
rect -3575 -9334 -3523 -9328
rect -3523 -9334 -3521 -9328
rect -3577 -9346 -3521 -9334
rect -3577 -9384 -3575 -9346
rect -3575 -9384 -3523 -9346
rect -3523 -9384 -3521 -9346
rect -3577 -9410 -3521 -9408
rect -3577 -9462 -3575 -9410
rect -3575 -9462 -3523 -9410
rect -3523 -9462 -3521 -9410
rect -3577 -9464 -3521 -9462
rect -3577 -9526 -3575 -9488
rect -3575 -9526 -3523 -9488
rect -3523 -9526 -3521 -9488
rect -3577 -9538 -3521 -9526
rect -3577 -9544 -3575 -9538
rect -3575 -9544 -3523 -9538
rect -3523 -9544 -3521 -9538
rect -3577 -9590 -3575 -9568
rect -3575 -9590 -3523 -9568
rect -3523 -9590 -3521 -9568
rect -3577 -9602 -3521 -9590
rect -3577 -9624 -3575 -9602
rect -3575 -9624 -3523 -9602
rect -3523 -9624 -3521 -9602
rect -3577 -9654 -3575 -9648
rect -3575 -9654 -3523 -9648
rect -3523 -9654 -3521 -9648
rect -3577 -9666 -3521 -9654
rect -3577 -9704 -3575 -9666
rect -3575 -9704 -3523 -9666
rect -3523 -9704 -3521 -9666
rect -3577 -9730 -3521 -9728
rect -3577 -9782 -3575 -9730
rect -3575 -9782 -3523 -9730
rect -3523 -9782 -3521 -9730
rect -3577 -9784 -3521 -9782
rect -3577 -9846 -3575 -9808
rect -3575 -9846 -3523 -9808
rect -3523 -9846 -3521 -9808
rect -3577 -9858 -3521 -9846
rect -3577 -9864 -3575 -9858
rect -3575 -9864 -3523 -9858
rect -3523 -9864 -3521 -9858
rect -3577 -9910 -3575 -9888
rect -3575 -9910 -3523 -9888
rect -3523 -9910 -3521 -9888
rect -3577 -9922 -3521 -9910
rect -3577 -9944 -3575 -9922
rect -3575 -9944 -3523 -9922
rect -3523 -9944 -3521 -9922
rect -3577 -9974 -3575 -9968
rect -3575 -9974 -3523 -9968
rect -3523 -9974 -3521 -9968
rect -3577 -9986 -3521 -9974
rect -3577 -10024 -3575 -9986
rect -3575 -10024 -3523 -9986
rect -3523 -10024 -3521 -9986
rect -3577 -10050 -3521 -10048
rect -3577 -10102 -3575 -10050
rect -3575 -10102 -3523 -10050
rect -3523 -10102 -3521 -10050
rect -3577 -10104 -3521 -10102
rect -571 -6857 -515 -6855
rect -571 -6909 -569 -6857
rect -569 -6909 -517 -6857
rect -517 -6909 -515 -6857
rect -571 -6911 -515 -6909
rect -571 -6973 -569 -6935
rect -569 -6973 -517 -6935
rect -517 -6973 -515 -6935
rect -571 -6985 -515 -6973
rect -571 -6991 -569 -6985
rect -569 -6991 -517 -6985
rect -517 -6991 -515 -6985
rect -571 -7037 -569 -7015
rect -569 -7037 -517 -7015
rect -517 -7037 -515 -7015
rect -571 -7049 -515 -7037
rect -571 -7071 -569 -7049
rect -569 -7071 -517 -7049
rect -517 -7071 -515 -7049
rect -571 -7101 -569 -7095
rect -569 -7101 -517 -7095
rect -517 -7101 -515 -7095
rect -571 -7113 -515 -7101
rect -571 -7151 -569 -7113
rect -569 -7151 -517 -7113
rect -517 -7151 -515 -7113
rect -571 -7177 -515 -7175
rect -571 -7229 -569 -7177
rect -569 -7229 -517 -7177
rect -517 -7229 -515 -7177
rect -571 -7231 -515 -7229
rect -571 -7293 -569 -7255
rect -569 -7293 -517 -7255
rect -517 -7293 -515 -7255
rect -571 -7305 -515 -7293
rect -571 -7311 -569 -7305
rect -569 -7311 -517 -7305
rect -517 -7311 -515 -7305
rect -571 -7357 -569 -7335
rect -569 -7357 -517 -7335
rect -517 -7357 -515 -7335
rect -571 -7369 -515 -7357
rect -571 -7391 -569 -7369
rect -569 -7391 -517 -7369
rect -517 -7391 -515 -7369
rect -571 -7421 -569 -7415
rect -569 -7421 -517 -7415
rect -517 -7421 -515 -7415
rect -571 -7433 -515 -7421
rect -571 -7471 -569 -7433
rect -569 -7471 -517 -7433
rect -517 -7471 -515 -7433
rect -571 -7497 -515 -7495
rect -571 -7549 -569 -7497
rect -569 -7549 -517 -7497
rect -517 -7549 -515 -7497
rect -571 -7551 -515 -7549
rect -571 -7613 -569 -7575
rect -569 -7613 -517 -7575
rect -517 -7613 -515 -7575
rect -571 -7625 -515 -7613
rect -571 -7631 -569 -7625
rect -569 -7631 -517 -7625
rect -517 -7631 -515 -7625
rect -571 -7677 -569 -7655
rect -569 -7677 -517 -7655
rect -517 -7677 -515 -7655
rect -571 -7689 -515 -7677
rect -571 -7711 -569 -7689
rect -569 -7711 -517 -7689
rect -517 -7711 -515 -7689
rect -571 -7741 -569 -7735
rect -569 -7741 -517 -7735
rect -517 -7741 -515 -7735
rect -571 -7753 -515 -7741
rect -571 -7791 -569 -7753
rect -569 -7791 -517 -7753
rect -517 -7791 -515 -7753
rect -571 -7817 -515 -7815
rect -571 -7869 -569 -7817
rect -569 -7869 -517 -7817
rect -517 -7869 -515 -7817
rect -571 -7871 -515 -7869
rect -571 -7933 -569 -7895
rect -569 -7933 -517 -7895
rect -517 -7933 -515 -7895
rect -571 -7945 -515 -7933
rect -571 -7951 -569 -7945
rect -569 -7951 -517 -7945
rect -517 -7951 -515 -7945
rect -571 -7997 -569 -7975
rect -569 -7997 -517 -7975
rect -517 -7997 -515 -7975
rect -571 -8009 -515 -7997
rect -571 -8031 -569 -8009
rect -569 -8031 -517 -8009
rect -517 -8031 -515 -8009
rect -571 -8061 -569 -8055
rect -569 -8061 -517 -8055
rect -517 -8061 -515 -8055
rect -571 -8073 -515 -8061
rect -571 -8111 -569 -8073
rect -569 -8111 -517 -8073
rect -517 -8111 -515 -8073
rect -571 -8137 -515 -8135
rect -571 -8189 -569 -8137
rect -569 -8189 -517 -8137
rect -517 -8189 -515 -8137
rect -571 -8191 -515 -8189
rect -571 -8253 -569 -8215
rect -569 -8253 -517 -8215
rect -517 -8253 -515 -8215
rect -571 -8265 -515 -8253
rect -571 -8271 -569 -8265
rect -569 -8271 -517 -8265
rect -517 -8271 -515 -8265
rect -571 -8317 -569 -8295
rect -569 -8317 -517 -8295
rect -517 -8317 -515 -8295
rect -571 -8329 -515 -8317
rect -571 -8351 -569 -8329
rect -569 -8351 -517 -8329
rect -517 -8351 -515 -8329
rect -571 -8381 -569 -8375
rect -569 -8381 -517 -8375
rect -517 -8381 -515 -8375
rect -571 -8393 -515 -8381
rect -571 -8431 -569 -8393
rect -569 -8431 -517 -8393
rect -517 -8431 -515 -8393
rect -571 -8457 -515 -8455
rect -571 -8509 -569 -8457
rect -569 -8509 -517 -8457
rect -517 -8509 -515 -8457
rect -571 -8511 -515 -8509
rect -571 -8573 -569 -8535
rect -569 -8573 -517 -8535
rect -517 -8573 -515 -8535
rect -571 -8585 -515 -8573
rect -571 -8591 -569 -8585
rect -569 -8591 -517 -8585
rect -517 -8591 -515 -8585
rect -571 -8637 -569 -8615
rect -569 -8637 -517 -8615
rect -517 -8637 -515 -8615
rect -571 -8649 -515 -8637
rect -571 -8671 -569 -8649
rect -569 -8671 -517 -8649
rect -517 -8671 -515 -8649
rect -571 -8701 -569 -8695
rect -569 -8701 -517 -8695
rect -517 -8701 -515 -8695
rect -571 -8713 -515 -8701
rect -571 -8751 -569 -8713
rect -569 -8751 -517 -8713
rect -517 -8751 -515 -8713
rect -571 -8777 -515 -8775
rect -571 -8829 -569 -8777
rect -569 -8829 -517 -8777
rect -517 -8829 -515 -8777
rect -571 -8831 -515 -8829
rect -571 -8893 -569 -8855
rect -569 -8893 -517 -8855
rect -517 -8893 -515 -8855
rect -571 -8905 -515 -8893
rect -571 -8911 -569 -8905
rect -569 -8911 -517 -8905
rect -517 -8911 -515 -8905
rect -571 -8957 -569 -8935
rect -569 -8957 -517 -8935
rect -517 -8957 -515 -8935
rect -571 -8969 -515 -8957
rect -571 -8991 -569 -8969
rect -569 -8991 -517 -8969
rect -517 -8991 -515 -8969
rect -571 -9021 -569 -9015
rect -569 -9021 -517 -9015
rect -517 -9021 -515 -9015
rect -571 -9033 -515 -9021
rect -571 -9071 -569 -9033
rect -569 -9071 -517 -9033
rect -517 -9071 -515 -9033
rect -571 -9097 -515 -9095
rect -571 -9149 -569 -9097
rect -569 -9149 -517 -9097
rect -517 -9149 -515 -9097
rect -571 -9151 -515 -9149
rect -571 -9213 -569 -9175
rect -569 -9213 -517 -9175
rect -517 -9213 -515 -9175
rect -571 -9225 -515 -9213
rect -571 -9231 -569 -9225
rect -569 -9231 -517 -9225
rect -517 -9231 -515 -9225
rect -571 -9277 -569 -9255
rect -569 -9277 -517 -9255
rect -517 -9277 -515 -9255
rect -571 -9289 -515 -9277
rect -571 -9311 -569 -9289
rect -569 -9311 -517 -9289
rect -517 -9311 -515 -9289
rect -571 -9341 -569 -9335
rect -569 -9341 -517 -9335
rect -517 -9341 -515 -9335
rect -571 -9353 -515 -9341
rect -571 -9391 -569 -9353
rect -569 -9391 -517 -9353
rect -517 -9391 -515 -9353
rect -571 -9417 -515 -9415
rect -571 -9469 -569 -9417
rect -569 -9469 -517 -9417
rect -517 -9469 -515 -9417
rect -571 -9471 -515 -9469
rect -571 -9533 -569 -9495
rect -569 -9533 -517 -9495
rect -517 -9533 -515 -9495
rect -571 -9545 -515 -9533
rect -571 -9551 -569 -9545
rect -569 -9551 -517 -9545
rect -517 -9551 -515 -9545
rect -571 -9597 -569 -9575
rect -569 -9597 -517 -9575
rect -517 -9597 -515 -9575
rect -571 -9609 -515 -9597
rect -571 -9631 -569 -9609
rect -569 -9631 -517 -9609
rect -517 -9631 -515 -9609
rect -571 -9661 -569 -9655
rect -569 -9661 -517 -9655
rect -517 -9661 -515 -9655
rect -571 -9673 -515 -9661
rect -571 -9711 -569 -9673
rect -569 -9711 -517 -9673
rect -517 -9711 -515 -9673
rect -571 -9737 -515 -9735
rect -571 -9789 -569 -9737
rect -569 -9789 -517 -9737
rect -517 -9789 -515 -9737
rect -571 -9791 -515 -9789
rect -571 -9853 -569 -9815
rect -569 -9853 -517 -9815
rect -517 -9853 -515 -9815
rect -571 -9865 -515 -9853
rect -571 -9871 -569 -9865
rect -569 -9871 -517 -9865
rect -517 -9871 -515 -9865
rect -571 -9917 -569 -9895
rect -569 -9917 -517 -9895
rect -517 -9917 -515 -9895
rect -571 -9929 -515 -9917
rect -571 -9951 -569 -9929
rect -569 -9951 -517 -9929
rect -517 -9951 -515 -9929
rect -571 -9981 -569 -9975
rect -569 -9981 -517 -9975
rect -517 -9981 -515 -9975
rect -571 -9993 -515 -9981
rect -571 -10031 -569 -9993
rect -569 -10031 -517 -9993
rect -517 -10031 -515 -9993
rect -571 -10057 -515 -10055
rect -571 -10109 -569 -10057
rect -569 -10109 -517 -10057
rect -517 -10109 -515 -10057
rect -571 -10111 -515 -10109
rect -2169 -12110 -1953 -12092
rect -2169 -12290 -2151 -12110
rect -2151 -12290 -1971 -12110
rect -1971 -12290 -1953 -12110
rect -2169 -12308 -1953 -12290
<< metal3 >>
rect -17013 85607 -16777 90441
rect -17013 85371 -15174 85607
rect -15410 78145 -15174 85371
rect 10990 85579 11226 90441
rect 22915 85752 23151 90441
rect 10990 85343 12843 85579
rect 22915 85516 24892 85752
rect -15420 78130 -15164 78145
rect -15420 77914 -15400 78130
rect -15184 77914 -15164 78130
rect 12607 78116 12843 85343
rect 24656 78117 24892 85516
rect -15420 77899 -15164 77914
rect 12596 78101 12852 78116
rect 12596 77885 12616 78101
rect 12832 77885 12852 78101
rect 12596 77870 12852 77885
rect 24646 78102 24902 78117
rect 24646 77886 24666 78102
rect 24882 77886 24902 78102
rect 24646 77871 24902 77886
rect 14134 76743 14282 76750
rect -16859 76692 -16738 76728
rect -16859 76628 -16831 76692
rect -16767 76628 -16738 76692
rect -16859 76612 -16738 76628
rect -16859 76548 -16831 76612
rect -16767 76548 -16738 76612
rect -16859 76532 -16738 76548
rect -16859 76468 -16831 76532
rect -16767 76468 -16738 76532
rect -16859 76452 -16738 76468
rect -16859 76388 -16831 76452
rect -16767 76388 -16738 76452
rect -16859 76372 -16738 76388
rect -16859 76308 -16831 76372
rect -16767 76308 -16738 76372
rect -16859 76292 -16738 76308
rect -16859 76228 -16831 76292
rect -16767 76228 -16738 76292
rect -16859 76212 -16738 76228
rect -16859 76148 -16831 76212
rect -16767 76148 -16738 76212
rect -16859 76132 -16738 76148
rect -16859 76068 -16831 76132
rect -16767 76068 -16738 76132
rect -16859 76052 -16738 76068
rect -16859 75988 -16831 76052
rect -16767 75988 -16738 76052
rect -16859 75972 -16738 75988
rect -16859 75908 -16831 75972
rect -16767 75908 -16738 75972
rect -16859 75892 -16738 75908
rect -16859 75828 -16831 75892
rect -16767 75828 -16738 75892
rect -16859 75812 -16738 75828
rect -16859 75748 -16831 75812
rect -16767 75748 -16738 75812
rect -16859 75732 -16738 75748
rect -16859 75668 -16831 75732
rect -16767 75668 -16738 75732
rect -16859 75652 -16738 75668
rect -16859 75588 -16831 75652
rect -16767 75588 -16738 75652
rect -16859 75572 -16738 75588
rect -16859 75508 -16831 75572
rect -16767 75508 -16738 75572
rect -16859 75492 -16738 75508
rect -16859 75428 -16831 75492
rect -16767 75428 -16738 75492
rect -16859 75412 -16738 75428
rect -16859 75348 -16831 75412
rect -16767 75348 -16738 75412
rect -16859 75332 -16738 75348
rect -16859 75268 -16831 75332
rect -16767 75268 -16738 75332
rect -16859 75252 -16738 75268
rect -16859 75188 -16831 75252
rect -16767 75188 -16738 75252
rect -16859 75172 -16738 75188
rect -16859 75108 -16831 75172
rect -16767 75108 -16738 75172
rect -16859 75092 -16738 75108
rect -16859 75028 -16831 75092
rect -16767 75028 -16738 75092
rect -16859 75012 -16738 75028
rect -16859 74948 -16831 75012
rect -16767 74948 -16738 75012
rect -16859 74932 -16738 74948
rect -16859 74868 -16831 74932
rect -16767 74868 -16738 74932
rect -16859 74852 -16738 74868
rect -16859 74788 -16831 74852
rect -16767 74788 -16738 74852
rect -16859 74772 -16738 74788
rect -16859 74708 -16831 74772
rect -16767 74708 -16738 74772
rect -16859 74692 -16738 74708
rect -16859 74628 -16831 74692
rect -16767 74628 -16738 74692
rect -16859 74612 -16738 74628
rect -16859 74548 -16831 74612
rect -16767 74548 -16738 74612
rect -16859 74532 -16738 74548
rect -16859 74468 -16831 74532
rect -16767 74468 -16738 74532
rect -16859 74452 -16738 74468
rect -16859 74388 -16831 74452
rect -16767 74388 -16738 74452
rect -16859 74372 -16738 74388
rect -16859 74308 -16831 74372
rect -16767 74308 -16738 74372
rect -16859 74292 -16738 74308
rect -16859 74228 -16831 74292
rect -16767 74228 -16738 74292
rect -16859 74212 -16738 74228
rect -16859 74148 -16831 74212
rect -16767 74148 -16738 74212
rect -16859 74132 -16738 74148
rect -16859 74068 -16831 74132
rect -16767 74068 -16738 74132
rect -16859 74052 -16738 74068
rect -16859 73988 -16831 74052
rect -16767 73988 -16738 74052
rect -16859 73972 -16738 73988
rect -16859 73908 -16831 73972
rect -16767 73908 -16738 73972
rect -16859 73892 -16738 73908
rect -16859 73828 -16831 73892
rect -16767 73828 -16738 73892
rect -16859 73812 -16738 73828
rect -16859 73748 -16831 73812
rect -16767 73748 -16738 73812
rect -16859 73732 -16738 73748
rect -16859 73668 -16831 73732
rect -16767 73668 -16738 73732
rect -16859 73652 -16738 73668
rect -16859 73588 -16831 73652
rect -16767 73588 -16738 73652
rect -16859 73572 -16738 73588
rect -16859 73508 -16831 73572
rect -16767 73508 -16738 73572
rect -16859 73492 -16738 73508
rect -16859 73428 -16831 73492
rect -16767 73428 -16738 73492
rect -16859 73393 -16738 73428
rect -13858 76698 -13737 76734
rect -13858 76634 -13830 76698
rect -13766 76634 -13737 76698
rect -13858 76618 -13737 76634
rect -13858 76554 -13830 76618
rect -13766 76554 -13737 76618
rect -13858 76538 -13737 76554
rect -13858 76474 -13830 76538
rect -13766 76474 -13737 76538
rect -13858 76458 -13737 76474
rect -13858 76394 -13830 76458
rect -13766 76394 -13737 76458
rect -13858 76378 -13737 76394
rect -13858 76314 -13830 76378
rect -13766 76314 -13737 76378
rect -13858 76298 -13737 76314
rect -13858 76234 -13830 76298
rect -13766 76234 -13737 76298
rect -13858 76218 -13737 76234
rect -13858 76154 -13830 76218
rect -13766 76154 -13737 76218
rect -13858 76138 -13737 76154
rect -13858 76074 -13830 76138
rect -13766 76074 -13737 76138
rect -13858 76058 -13737 76074
rect -13858 75994 -13830 76058
rect -13766 75994 -13737 76058
rect -13858 75978 -13737 75994
rect -13858 75914 -13830 75978
rect -13766 75914 -13737 75978
rect -13858 75898 -13737 75914
rect -13858 75834 -13830 75898
rect -13766 75834 -13737 75898
rect -13858 75818 -13737 75834
rect -13858 75754 -13830 75818
rect -13766 75754 -13737 75818
rect -13858 75738 -13737 75754
rect -13858 75674 -13830 75738
rect -13766 75674 -13737 75738
rect -13858 75658 -13737 75674
rect -13858 75594 -13830 75658
rect -13766 75594 -13737 75658
rect -13858 75578 -13737 75594
rect -13858 75514 -13830 75578
rect -13766 75514 -13737 75578
rect -13858 75498 -13737 75514
rect -13858 75434 -13830 75498
rect -13766 75434 -13737 75498
rect -13858 75418 -13737 75434
rect -13858 75354 -13830 75418
rect -13766 75354 -13737 75418
rect -13858 75338 -13737 75354
rect -13858 75274 -13830 75338
rect -13766 75274 -13737 75338
rect -13858 75258 -13737 75274
rect -13858 75194 -13830 75258
rect -13766 75194 -13737 75258
rect -13858 75178 -13737 75194
rect -13858 75114 -13830 75178
rect -13766 75114 -13737 75178
rect -13858 75098 -13737 75114
rect -13858 75034 -13830 75098
rect -13766 75034 -13737 75098
rect -13858 75018 -13737 75034
rect -13858 74954 -13830 75018
rect -13766 74954 -13737 75018
rect -13858 74938 -13737 74954
rect -13858 74874 -13830 74938
rect -13766 74874 -13737 74938
rect -13858 74858 -13737 74874
rect -13858 74794 -13830 74858
rect -13766 74794 -13737 74858
rect -13858 74778 -13737 74794
rect -13858 74714 -13830 74778
rect -13766 74714 -13737 74778
rect -13858 74698 -13737 74714
rect -13858 74634 -13830 74698
rect -13766 74634 -13737 74698
rect -13858 74618 -13737 74634
rect -13858 74554 -13830 74618
rect -13766 74554 -13737 74618
rect -13858 74538 -13737 74554
rect -13858 74474 -13830 74538
rect -13766 74474 -13737 74538
rect -13858 74458 -13737 74474
rect -13858 74394 -13830 74458
rect -13766 74394 -13737 74458
rect -13858 74378 -13737 74394
rect -13858 74314 -13830 74378
rect -13766 74314 -13737 74378
rect -13858 74298 -13737 74314
rect -13858 74234 -13830 74298
rect -13766 74234 -13737 74298
rect -13858 74218 -13737 74234
rect -13858 74154 -13830 74218
rect -13766 74154 -13737 74218
rect -13858 74138 -13737 74154
rect -13858 74074 -13830 74138
rect -13766 74074 -13737 74138
rect -13858 74058 -13737 74074
rect -13858 73994 -13830 74058
rect -13766 73994 -13737 74058
rect -13858 73978 -13737 73994
rect -13858 73914 -13830 73978
rect -13766 73914 -13737 73978
rect -13858 73898 -13737 73914
rect -13858 73834 -13830 73898
rect -13766 73834 -13737 73898
rect -13858 73818 -13737 73834
rect -13858 73754 -13830 73818
rect -13766 73754 -13737 73818
rect -13858 73738 -13737 73754
rect -13858 73674 -13830 73738
rect -13766 73674 -13737 73738
rect -13858 73658 -13737 73674
rect -13858 73594 -13830 73658
rect -13766 73594 -13737 73658
rect -13858 73578 -13737 73594
rect -13858 73514 -13830 73578
rect -13766 73514 -13737 73578
rect -13858 73498 -13737 73514
rect -13858 73434 -13830 73498
rect -13766 73434 -13737 73498
rect -13858 73399 -13737 73434
rect 11133 76730 11281 76737
rect 11133 76694 11179 76730
rect 11235 76694 11281 76730
rect 11133 76630 11175 76694
rect 11239 76630 11281 76694
rect 11133 76614 11179 76630
rect 11235 76614 11281 76630
rect 11133 76550 11175 76614
rect 11239 76550 11281 76614
rect 11133 76534 11179 76550
rect 11235 76534 11281 76550
rect 11133 76470 11175 76534
rect 11239 76470 11281 76534
rect 11133 76454 11179 76470
rect 11235 76454 11281 76470
rect 11133 76390 11175 76454
rect 11239 76390 11281 76454
rect 11133 76374 11179 76390
rect 11235 76374 11281 76390
rect 11133 76310 11175 76374
rect 11239 76310 11281 76374
rect 11133 76294 11179 76310
rect 11235 76294 11281 76310
rect 11133 76230 11175 76294
rect 11239 76230 11281 76294
rect 11133 76214 11179 76230
rect 11235 76214 11281 76230
rect 11133 76150 11175 76214
rect 11239 76150 11281 76214
rect 11133 76134 11179 76150
rect 11235 76134 11281 76150
rect 11133 76070 11175 76134
rect 11239 76070 11281 76134
rect 11133 76054 11179 76070
rect 11235 76054 11281 76070
rect 11133 75990 11175 76054
rect 11239 75990 11281 76054
rect 11133 75974 11179 75990
rect 11235 75974 11281 75990
rect 11133 75910 11175 75974
rect 11239 75910 11281 75974
rect 11133 75894 11179 75910
rect 11235 75894 11281 75910
rect 11133 75830 11175 75894
rect 11239 75830 11281 75894
rect 11133 75814 11179 75830
rect 11235 75814 11281 75830
rect 11133 75750 11175 75814
rect 11239 75750 11281 75814
rect 11133 75734 11179 75750
rect 11235 75734 11281 75750
rect 11133 75670 11175 75734
rect 11239 75670 11281 75734
rect 11133 75654 11179 75670
rect 11235 75654 11281 75670
rect 11133 75590 11175 75654
rect 11239 75590 11281 75654
rect 11133 75574 11179 75590
rect 11235 75574 11281 75590
rect 11133 75510 11175 75574
rect 11239 75510 11281 75574
rect 11133 75494 11179 75510
rect 11235 75494 11281 75510
rect 11133 75430 11175 75494
rect 11239 75430 11281 75494
rect 11133 75414 11179 75430
rect 11235 75414 11281 75430
rect 11133 75350 11175 75414
rect 11239 75350 11281 75414
rect 11133 75334 11179 75350
rect 11235 75334 11281 75350
rect 11133 75270 11175 75334
rect 11239 75270 11281 75334
rect 11133 75254 11179 75270
rect 11235 75254 11281 75270
rect 11133 75190 11175 75254
rect 11239 75190 11281 75254
rect 11133 75174 11179 75190
rect 11235 75174 11281 75190
rect 11133 75110 11175 75174
rect 11239 75110 11281 75174
rect 11133 75094 11179 75110
rect 11235 75094 11281 75110
rect 11133 75030 11175 75094
rect 11239 75030 11281 75094
rect 11133 75014 11179 75030
rect 11235 75014 11281 75030
rect 11133 74950 11175 75014
rect 11239 74950 11281 75014
rect 11133 74934 11179 74950
rect 11235 74934 11281 74950
rect 11133 74870 11175 74934
rect 11239 74870 11281 74934
rect 11133 74854 11179 74870
rect 11235 74854 11281 74870
rect 11133 74790 11175 74854
rect 11239 74790 11281 74854
rect 11133 74774 11179 74790
rect 11235 74774 11281 74790
rect 11133 74710 11175 74774
rect 11239 74710 11281 74774
rect 11133 74694 11179 74710
rect 11235 74694 11281 74710
rect 11133 74630 11175 74694
rect 11239 74630 11281 74694
rect 11133 74614 11179 74630
rect 11235 74614 11281 74630
rect 11133 74550 11175 74614
rect 11239 74550 11281 74614
rect 11133 74534 11179 74550
rect 11235 74534 11281 74550
rect 11133 74470 11175 74534
rect 11239 74470 11281 74534
rect 11133 74454 11179 74470
rect 11235 74454 11281 74470
rect 11133 74390 11175 74454
rect 11239 74390 11281 74454
rect 11133 74374 11179 74390
rect 11235 74374 11281 74390
rect 11133 74310 11175 74374
rect 11239 74310 11281 74374
rect 11133 74294 11179 74310
rect 11235 74294 11281 74310
rect 11133 74230 11175 74294
rect 11239 74230 11281 74294
rect 11133 74214 11179 74230
rect 11235 74214 11281 74230
rect 11133 74150 11175 74214
rect 11239 74150 11281 74214
rect 11133 74134 11179 74150
rect 11235 74134 11281 74150
rect 11133 74070 11175 74134
rect 11239 74070 11281 74134
rect 11133 74054 11179 74070
rect 11235 74054 11281 74070
rect 11133 73990 11175 74054
rect 11239 73990 11281 74054
rect 11133 73974 11179 73990
rect 11235 73974 11281 73990
rect 11133 73910 11175 73974
rect 11239 73910 11281 73974
rect 11133 73894 11179 73910
rect 11235 73894 11281 73910
rect 11133 73830 11175 73894
rect 11239 73830 11281 73894
rect 11133 73814 11179 73830
rect 11235 73814 11281 73830
rect 11133 73750 11175 73814
rect 11239 73750 11281 73814
rect 11133 73734 11179 73750
rect 11235 73734 11281 73750
rect 11133 73670 11175 73734
rect 11239 73670 11281 73734
rect 11133 73654 11179 73670
rect 11235 73654 11281 73670
rect 11133 73590 11175 73654
rect 11239 73590 11281 73654
rect 11133 73574 11179 73590
rect 11235 73574 11281 73590
rect 11133 73510 11175 73574
rect 11239 73510 11281 73574
rect 11133 73494 11179 73510
rect 11235 73494 11281 73510
rect 11133 73430 11175 73494
rect 11239 73430 11281 73494
rect 11133 73394 11179 73430
rect 11235 73394 11281 73430
rect 14134 76707 14180 76743
rect 14236 76707 14282 76743
rect 14134 76643 14176 76707
rect 14240 76643 14282 76707
rect 14134 76627 14180 76643
rect 14236 76627 14282 76643
rect 14134 76563 14176 76627
rect 14240 76563 14282 76627
rect 14134 76547 14180 76563
rect 14236 76547 14282 76563
rect 14134 76483 14176 76547
rect 14240 76483 14282 76547
rect 14134 76467 14180 76483
rect 14236 76467 14282 76483
rect 14134 76403 14176 76467
rect 14240 76403 14282 76467
rect 14134 76387 14180 76403
rect 14236 76387 14282 76403
rect 14134 76323 14176 76387
rect 14240 76323 14282 76387
rect 14134 76307 14180 76323
rect 14236 76307 14282 76323
rect 14134 76243 14176 76307
rect 14240 76243 14282 76307
rect 14134 76227 14180 76243
rect 14236 76227 14282 76243
rect 14134 76163 14176 76227
rect 14240 76163 14282 76227
rect 14134 76147 14180 76163
rect 14236 76147 14282 76163
rect 14134 76083 14176 76147
rect 14240 76083 14282 76147
rect 14134 76067 14180 76083
rect 14236 76067 14282 76083
rect 14134 76003 14176 76067
rect 14240 76003 14282 76067
rect 14134 75987 14180 76003
rect 14236 75987 14282 76003
rect 14134 75923 14176 75987
rect 14240 75923 14282 75987
rect 14134 75907 14180 75923
rect 14236 75907 14282 75923
rect 14134 75843 14176 75907
rect 14240 75843 14282 75907
rect 14134 75827 14180 75843
rect 14236 75827 14282 75843
rect 14134 75763 14176 75827
rect 14240 75763 14282 75827
rect 14134 75747 14180 75763
rect 14236 75747 14282 75763
rect 14134 75683 14176 75747
rect 14240 75683 14282 75747
rect 14134 75667 14180 75683
rect 14236 75667 14282 75683
rect 14134 75603 14176 75667
rect 14240 75603 14282 75667
rect 14134 75587 14180 75603
rect 14236 75587 14282 75603
rect 14134 75523 14176 75587
rect 14240 75523 14282 75587
rect 14134 75507 14180 75523
rect 14236 75507 14282 75523
rect 14134 75443 14176 75507
rect 14240 75443 14282 75507
rect 14134 75427 14180 75443
rect 14236 75427 14282 75443
rect 14134 75363 14176 75427
rect 14240 75363 14282 75427
rect 14134 75347 14180 75363
rect 14236 75347 14282 75363
rect 14134 75283 14176 75347
rect 14240 75283 14282 75347
rect 14134 75267 14180 75283
rect 14236 75267 14282 75283
rect 14134 75203 14176 75267
rect 14240 75203 14282 75267
rect 14134 75187 14180 75203
rect 14236 75187 14282 75203
rect 14134 75123 14176 75187
rect 14240 75123 14282 75187
rect 14134 75107 14180 75123
rect 14236 75107 14282 75123
rect 14134 75043 14176 75107
rect 14240 75043 14282 75107
rect 14134 75027 14180 75043
rect 14236 75027 14282 75043
rect 14134 74963 14176 75027
rect 14240 74963 14282 75027
rect 14134 74947 14180 74963
rect 14236 74947 14282 74963
rect 14134 74883 14176 74947
rect 14240 74883 14282 74947
rect 14134 74867 14180 74883
rect 14236 74867 14282 74883
rect 14134 74803 14176 74867
rect 14240 74803 14282 74867
rect 14134 74787 14180 74803
rect 14236 74787 14282 74803
rect 14134 74723 14176 74787
rect 14240 74723 14282 74787
rect 14134 74707 14180 74723
rect 14236 74707 14282 74723
rect 14134 74643 14176 74707
rect 14240 74643 14282 74707
rect 14134 74627 14180 74643
rect 14236 74627 14282 74643
rect 14134 74563 14176 74627
rect 14240 74563 14282 74627
rect 14134 74547 14180 74563
rect 14236 74547 14282 74563
rect 14134 74483 14176 74547
rect 14240 74483 14282 74547
rect 14134 74467 14180 74483
rect 14236 74467 14282 74483
rect 14134 74403 14176 74467
rect 14240 74403 14282 74467
rect 14134 74387 14180 74403
rect 14236 74387 14282 74403
rect 14134 74323 14176 74387
rect 14240 74323 14282 74387
rect 14134 74307 14180 74323
rect 14236 74307 14282 74323
rect 14134 74243 14176 74307
rect 14240 74243 14282 74307
rect 14134 74227 14180 74243
rect 14236 74227 14282 74243
rect 14134 74163 14176 74227
rect 14240 74163 14282 74227
rect 14134 74147 14180 74163
rect 14236 74147 14282 74163
rect 14134 74083 14176 74147
rect 14240 74083 14282 74147
rect 14134 74067 14180 74083
rect 14236 74067 14282 74083
rect 14134 74003 14176 74067
rect 14240 74003 14282 74067
rect 14134 73987 14180 74003
rect 14236 73987 14282 74003
rect 14134 73923 14176 73987
rect 14240 73923 14282 73987
rect 14134 73907 14180 73923
rect 14236 73907 14282 73923
rect 14134 73843 14176 73907
rect 14240 73843 14282 73907
rect 14134 73827 14180 73843
rect 14236 73827 14282 73843
rect 14134 73763 14176 73827
rect 14240 73763 14282 73827
rect 14134 73747 14180 73763
rect 14236 73747 14282 73763
rect 14134 73683 14176 73747
rect 14240 73683 14282 73747
rect 14134 73667 14180 73683
rect 14236 73667 14282 73683
rect 14134 73603 14176 73667
rect 14240 73603 14282 73667
rect 14134 73587 14180 73603
rect 14236 73587 14282 73603
rect 14134 73523 14176 73587
rect 14240 73523 14282 73587
rect 14134 73507 14180 73523
rect 14236 73507 14282 73523
rect 14134 73443 14176 73507
rect 14240 73443 14282 73507
rect 14134 73407 14180 73443
rect 14236 73407 14282 73443
rect 14134 73400 14282 73407
rect 57721 75975 62907 76211
rect 11133 73387 11281 73394
rect -16697 71802 -16560 71832
rect -16697 71738 -16664 71802
rect -16600 71738 -16560 71802
rect -16697 71706 -16560 71738
rect -15509 71798 -15392 71820
rect -15509 71734 -15486 71798
rect -15422 71734 -15392 71798
rect -15509 71709 -15392 71734
rect -15292 71805 -15176 71835
rect -15292 71741 -15269 71805
rect -15205 71741 -15176 71805
rect -15292 71714 -15176 71741
rect -14161 71802 -14041 71826
rect -14161 71738 -14135 71802
rect -14071 71738 -14041 71802
rect -14161 71709 -14041 71738
rect -16577 70298 -16469 70319
rect -16577 70234 -16554 70298
rect -16490 70234 -16469 70298
rect -16577 70206 -16469 70234
rect -15464 70284 -15355 70304
rect -15464 70220 -15440 70284
rect -15376 70220 -15355 70284
rect -15464 70197 -15355 70220
rect -15249 70285 -15140 70310
rect -15249 70221 -15227 70285
rect -15163 70221 -15140 70285
rect -15249 70197 -15140 70221
rect -14091 70285 -13954 70311
rect -14091 70221 -14063 70285
rect -13999 70221 -13954 70285
rect -14091 70197 -13954 70221
rect 57721 69420 57957 75975
rect 36555 69334 57957 69420
rect 36555 69270 36631 69334
rect 36695 69270 57957 69334
rect 36555 69184 57957 69270
rect -13963 68741 62907 68813
rect -16718 68703 -16634 68708
rect -13963 68703 36066 68741
rect -16718 68699 36066 68703
rect -16718 68643 -16704 68699
rect -16648 68677 36066 68699
rect 36130 68677 62907 68741
rect -16648 68643 62907 68677
rect -16718 68639 62907 68643
rect -16718 68634 -16634 68639
rect -13963 68577 62907 68639
rect -15432 68492 -15348 68520
rect -15432 68428 -15422 68492
rect -15358 68428 -15348 68492
rect -15432 68412 -15348 68428
rect -15432 68348 -15422 68412
rect -15358 68348 -15348 68412
rect -15432 68332 -15348 68348
rect -15432 68268 -15422 68332
rect -15358 68268 -15348 68332
rect -15973 68255 -15880 68266
rect -15973 68191 -15959 68255
rect -15895 68191 -15880 68255
rect -15973 68175 -15880 68191
rect -15973 68111 -15959 68175
rect -15895 68111 -15880 68175
rect -15432 68252 -15348 68268
rect -15432 68188 -15422 68252
rect -15358 68188 -15348 68252
rect -15432 68161 -15348 68188
rect -14889 68258 -14796 68269
rect -14889 68194 -14875 68258
rect -14811 68194 -14796 68258
rect -14889 68178 -14796 68194
rect -15973 68100 -15880 68111
rect -14889 68114 -14875 68178
rect -14811 68114 -14796 68178
rect -14889 68103 -14796 68114
rect -13966 68081 58032 68169
rect -14209 68073 -14125 68078
rect -13966 68073 35477 68081
rect -14209 68069 35477 68073
rect -14209 68013 -14195 68069
rect -14139 68017 35477 68069
rect 35541 68017 58032 68081
rect -14139 68013 58032 68017
rect -14209 68009 58032 68013
rect -14209 68004 -14125 68009
rect -13966 67933 58032 68009
rect -16605 67613 -16482 67643
rect -16605 67549 -16577 67613
rect -16513 67549 -16482 67613
rect -16605 67518 -16482 67549
rect -15449 67607 -15330 67633
rect -15449 67543 -15422 67607
rect -15358 67543 -15330 67607
rect -15449 67513 -15330 67543
rect -14328 67618 -14211 67641
rect -14328 67554 -14304 67618
rect -14240 67554 -14211 67618
rect -14328 67526 -14211 67554
rect -13106 66705 -13096 66769
rect -13032 66705 -8073 66769
rect -8009 66705 -7999 66769
rect -12325 66382 -12315 66446
rect -12251 66382 -7266 66446
rect -7202 66382 -7192 66446
rect -11313 65949 -11305 66013
rect -11241 65949 -2673 66013
rect -2609 65949 -2599 66013
rect -10544 65696 -10536 65760
rect -10472 65696 -1866 65760
rect -1802 65696 -1792 65760
rect -8083 65265 -8073 65329
rect -8009 65265 -7999 65329
rect -2683 65265 -2673 65329
rect -2609 65265 -2599 65329
rect -7276 65012 -7266 65076
rect -7202 65012 -7192 65076
rect -1876 65012 -1866 65076
rect -1802 65012 -1792 65076
rect 17420 64728 17506 64748
rect 17420 64664 17431 64728
rect 17495 64664 17506 64728
rect 17420 64648 17506 64664
rect 17420 64584 17431 64648
rect 17495 64584 17506 64648
rect 17420 64568 17506 64584
rect 17420 64504 17431 64568
rect 17495 64504 17506 64568
rect 17420 64488 17506 64504
rect 17420 64424 17431 64488
rect 17495 64424 17506 64488
rect 17420 64408 17506 64424
rect 17420 64344 17431 64408
rect 17495 64344 17506 64408
rect 17420 64328 17506 64344
rect 17420 64264 17431 64328
rect 17495 64264 17506 64328
rect 17420 64248 17506 64264
rect 17420 64184 17431 64248
rect 17495 64184 17506 64248
rect 17420 64164 17506 64184
rect 23948 64728 24034 64748
rect 23948 64664 23959 64728
rect 24023 64664 24034 64728
rect 23948 64648 24034 64664
rect 23948 64584 23959 64648
rect 24023 64584 24034 64648
rect 23948 64568 24034 64584
rect 23948 64504 23959 64568
rect 24023 64504 24034 64568
rect 23948 64488 24034 64504
rect 23948 64424 23959 64488
rect 24023 64424 24034 64488
rect 23948 64408 24034 64424
rect 23948 64344 23959 64408
rect 24023 64344 24034 64408
rect 23948 64328 24034 64344
rect 23948 64264 23959 64328
rect 24023 64264 24034 64328
rect 23948 64248 24034 64264
rect 23948 64184 23959 64248
rect 24023 64184 24034 64248
rect 23948 64164 24034 64184
rect 31564 64728 31650 64748
rect 31564 64664 31575 64728
rect 31639 64664 31650 64728
rect 31564 64648 31650 64664
rect 31564 64584 31575 64648
rect 31639 64584 31650 64648
rect 31564 64568 31650 64584
rect 31564 64504 31575 64568
rect 31639 64504 31650 64568
rect 31564 64488 31650 64504
rect 31564 64424 31575 64488
rect 31639 64424 31650 64488
rect 31564 64408 31650 64424
rect 31564 64344 31575 64408
rect 31639 64344 31650 64408
rect 31564 64328 31650 64344
rect 31564 64264 31575 64328
rect 31639 64264 31650 64328
rect 31564 64248 31650 64264
rect 31564 64184 31575 64248
rect 31639 64184 31650 64248
rect 31564 64164 31650 64184
rect -11081 63533 -10727 63557
rect -11081 63229 -11056 63533
rect -10752 63402 -10727 63533
rect -9894 63402 -9432 63407
rect -10752 63338 -10187 63402
rect -10123 63338 -10113 63402
rect -9894 63338 -9855 63402
rect -9791 63338 -9775 63402
rect -9711 63338 -9695 63402
rect -9631 63338 -9615 63402
rect -9551 63338 -9535 63402
rect -9471 63338 -9432 63402
rect -10752 63229 -10727 63338
rect -9894 63333 -9432 63338
rect -8083 63404 -7621 63409
rect -8083 63340 -8044 63404
rect -7980 63340 -7964 63404
rect -7900 63340 -7884 63404
rect -7820 63340 -7804 63404
rect -7740 63340 -7724 63404
rect -7660 63340 -7621 63404
rect -8083 63335 -7621 63340
rect -6288 63400 -5826 63405
rect -6288 63336 -6249 63400
rect -6185 63336 -6169 63400
rect -6105 63336 -6089 63400
rect -6025 63336 -6009 63400
rect -5945 63336 -5929 63400
rect -5865 63336 -5826 63400
rect -6288 63331 -5826 63336
rect -4489 63398 -4027 63403
rect -4489 63334 -4450 63398
rect -4386 63334 -4370 63398
rect -4306 63334 -4290 63398
rect -4226 63334 -4210 63398
rect -4146 63334 -4130 63398
rect -4066 63334 -4027 63398
rect -4489 63329 -4027 63334
rect -2698 63402 -2236 63407
rect -2698 63338 -2659 63402
rect -2595 63338 -2579 63402
rect -2515 63338 -2499 63402
rect -2435 63338 -2419 63402
rect -2355 63338 -2339 63402
rect -2275 63338 -2236 63402
rect -2698 63333 -2236 63338
rect -896 63398 -434 63403
rect -896 63334 -857 63398
rect -793 63334 -777 63398
rect -713 63334 -697 63398
rect -633 63334 -617 63398
rect -553 63334 -537 63398
rect -473 63334 -434 63398
rect -896 63329 -434 63334
rect -11081 63205 -10727 63229
rect 747 63224 1297 63237
rect -6949 63198 -6689 63211
rect -6949 62974 -6931 63198
rect -6707 62974 -6689 63198
rect 747 63000 790 63224
rect 1254 63000 1297 63224
rect 747 62987 1297 63000
rect -6949 62961 -6689 62974
rect 17965 62725 18051 62745
rect 17965 62661 17976 62725
rect 18040 62661 18051 62725
rect 17965 62645 18051 62661
rect 17965 62581 17976 62645
rect 18040 62581 18051 62645
rect 17965 62565 18051 62581
rect 17965 62501 17976 62565
rect 18040 62501 18051 62565
rect 17965 62485 18051 62501
rect 17965 62421 17976 62485
rect 18040 62421 18051 62485
rect 17965 62405 18051 62421
rect 17965 62341 17976 62405
rect 18040 62341 18051 62405
rect 17965 62325 18051 62341
rect 17965 62261 17976 62325
rect 18040 62261 18051 62325
rect 17965 62245 18051 62261
rect 17965 62181 17976 62245
rect 18040 62181 18051 62245
rect 17965 62161 18051 62181
rect 19053 62725 19139 62745
rect 19053 62661 19064 62725
rect 19128 62661 19139 62725
rect 19053 62645 19139 62661
rect 19053 62581 19064 62645
rect 19128 62581 19139 62645
rect 19053 62565 19139 62581
rect 19053 62501 19064 62565
rect 19128 62501 19139 62565
rect 19053 62485 19139 62501
rect 19053 62421 19064 62485
rect 19128 62421 19139 62485
rect 19053 62405 19139 62421
rect 19053 62341 19064 62405
rect 19128 62341 19139 62405
rect 19053 62325 19139 62341
rect 19053 62261 19064 62325
rect 19128 62261 19139 62325
rect 19053 62245 19139 62261
rect 19053 62181 19064 62245
rect 19128 62181 19139 62245
rect 19053 62161 19139 62181
rect 21229 62725 21315 62745
rect 21229 62661 21240 62725
rect 21304 62661 21315 62725
rect 21229 62645 21315 62661
rect 21229 62581 21240 62645
rect 21304 62581 21315 62645
rect 21229 62565 21315 62581
rect 21229 62501 21240 62565
rect 21304 62501 21315 62565
rect 21229 62485 21315 62501
rect 21229 62421 21240 62485
rect 21304 62421 21315 62485
rect 21229 62405 21315 62421
rect 21229 62341 21240 62405
rect 21304 62341 21315 62405
rect 21229 62325 21315 62341
rect 21229 62261 21240 62325
rect 21304 62261 21315 62325
rect 21229 62245 21315 62261
rect 21229 62181 21240 62245
rect 21304 62181 21315 62245
rect 21229 62161 21315 62181
rect 22317 62725 22403 62745
rect 22317 62661 22328 62725
rect 22392 62661 22403 62725
rect 22317 62645 22403 62661
rect 22317 62581 22328 62645
rect 22392 62581 22403 62645
rect 22317 62565 22403 62581
rect 22317 62501 22328 62565
rect 22392 62501 22403 62565
rect 22317 62485 22403 62501
rect 22317 62421 22328 62485
rect 22392 62421 22403 62485
rect 22317 62405 22403 62421
rect 22317 62341 22328 62405
rect 22392 62341 22403 62405
rect 22317 62325 22403 62341
rect 22317 62261 22328 62325
rect 22392 62261 22403 62325
rect 22317 62245 22403 62261
rect 22317 62181 22328 62245
rect 22392 62181 22403 62245
rect 22317 62161 22403 62181
rect 23405 62725 23491 62745
rect 23405 62661 23416 62725
rect 23480 62661 23491 62725
rect 23405 62645 23491 62661
rect 23405 62581 23416 62645
rect 23480 62581 23491 62645
rect 23405 62565 23491 62581
rect 23405 62501 23416 62565
rect 23480 62501 23491 62565
rect 23405 62485 23491 62501
rect 23405 62421 23416 62485
rect 23480 62421 23491 62485
rect 23405 62405 23491 62421
rect 23405 62341 23416 62405
rect 23480 62341 23491 62405
rect 23405 62325 23491 62341
rect 23405 62261 23416 62325
rect 23480 62261 23491 62325
rect 23405 62245 23491 62261
rect 23405 62181 23416 62245
rect 23480 62181 23491 62245
rect 23405 62161 23491 62181
rect 24493 62725 24579 62745
rect 24493 62661 24504 62725
rect 24568 62661 24579 62725
rect 24493 62645 24579 62661
rect 24493 62581 24504 62645
rect 24568 62581 24579 62645
rect 24493 62565 24579 62581
rect 24493 62501 24504 62565
rect 24568 62501 24579 62565
rect 24493 62485 24579 62501
rect 24493 62421 24504 62485
rect 24568 62421 24579 62485
rect 24493 62405 24579 62421
rect 24493 62341 24504 62405
rect 24568 62341 24579 62405
rect 24493 62325 24579 62341
rect 24493 62261 24504 62325
rect 24568 62261 24579 62325
rect 24493 62245 24579 62261
rect 24493 62181 24504 62245
rect 24568 62181 24579 62245
rect 24493 62161 24579 62181
rect 25581 62725 25667 62745
rect 25581 62661 25592 62725
rect 25656 62661 25667 62725
rect 25581 62645 25667 62661
rect 25581 62581 25592 62645
rect 25656 62581 25667 62645
rect 25581 62565 25667 62581
rect 25581 62501 25592 62565
rect 25656 62501 25667 62565
rect 25581 62485 25667 62501
rect 25581 62421 25592 62485
rect 25656 62421 25667 62485
rect 25581 62405 25667 62421
rect 25581 62341 25592 62405
rect 25656 62341 25667 62405
rect 25581 62325 25667 62341
rect 25581 62261 25592 62325
rect 25656 62261 25667 62325
rect 25581 62245 25667 62261
rect 25581 62181 25592 62245
rect 25656 62181 25667 62245
rect 25581 62161 25667 62181
rect 26669 62725 26755 62745
rect 26669 62661 26680 62725
rect 26744 62661 26755 62725
rect 26669 62645 26755 62661
rect 26669 62581 26680 62645
rect 26744 62581 26755 62645
rect 26669 62565 26755 62581
rect 26669 62501 26680 62565
rect 26744 62501 26755 62565
rect 26669 62485 26755 62501
rect 26669 62421 26680 62485
rect 26744 62421 26755 62485
rect 26669 62405 26755 62421
rect 26669 62341 26680 62405
rect 26744 62341 26755 62405
rect 26669 62325 26755 62341
rect 26669 62261 26680 62325
rect 26744 62261 26755 62325
rect 26669 62245 26755 62261
rect 26669 62181 26680 62245
rect 26744 62181 26755 62245
rect 26669 62161 26755 62181
rect 28845 62725 28931 62745
rect 28845 62661 28856 62725
rect 28920 62661 28931 62725
rect 28845 62645 28931 62661
rect 28845 62581 28856 62645
rect 28920 62581 28931 62645
rect 28845 62565 28931 62581
rect 28845 62501 28856 62565
rect 28920 62501 28931 62565
rect 28845 62485 28931 62501
rect 28845 62421 28856 62485
rect 28920 62421 28931 62485
rect 28845 62405 28931 62421
rect 28845 62341 28856 62405
rect 28920 62341 28931 62405
rect 28845 62325 28931 62341
rect 28845 62261 28856 62325
rect 28920 62261 28931 62325
rect 28845 62245 28931 62261
rect 28845 62181 28856 62245
rect 28920 62181 28931 62245
rect 28845 62161 28931 62181
rect 29933 62725 30019 62745
rect 29933 62661 29944 62725
rect 30008 62661 30019 62725
rect 29933 62645 30019 62661
rect 29933 62581 29944 62645
rect 30008 62581 30019 62645
rect 29933 62565 30019 62581
rect 29933 62501 29944 62565
rect 30008 62501 30019 62565
rect 29933 62485 30019 62501
rect 29933 62421 29944 62485
rect 30008 62421 30019 62485
rect 29933 62405 30019 62421
rect 29933 62341 29944 62405
rect 30008 62341 30019 62405
rect 29933 62325 30019 62341
rect 29933 62261 29944 62325
rect 30008 62261 30019 62325
rect 29933 62245 30019 62261
rect 29933 62181 29944 62245
rect 30008 62181 30019 62245
rect 29933 62161 30019 62181
rect 31021 62725 31107 62745
rect 31021 62661 31032 62725
rect 31096 62661 31107 62725
rect 31021 62645 31107 62661
rect 31021 62581 31032 62645
rect 31096 62581 31107 62645
rect 31021 62565 31107 62581
rect 31021 62501 31032 62565
rect 31096 62501 31107 62565
rect 31021 62485 31107 62501
rect 31021 62421 31032 62485
rect 31096 62421 31107 62485
rect 31021 62405 31107 62421
rect 31021 62341 31032 62405
rect 31096 62341 31107 62405
rect 31021 62325 31107 62341
rect 31021 62261 31032 62325
rect 31096 62261 31107 62325
rect 31021 62245 31107 62261
rect 31021 62181 31032 62245
rect 31096 62181 31107 62245
rect 31021 62161 31107 62181
rect 57796 61375 58032 67933
rect 57796 61139 62907 61375
rect 337 60806 529 60832
rect -8583 54595 -8471 54619
rect -8583 54531 -8557 54595
rect -8493 54531 -8471 54595
rect -8583 54507 -8471 54531
rect -6889 54596 -6772 54625
rect -6889 54532 -6866 54596
rect -6802 54532 -6772 54596
rect -6889 54508 -6772 54532
rect -5179 54595 -5082 54614
rect -5179 54531 -5161 54595
rect -5097 54531 -5082 54595
rect -5179 54511 -5082 54531
rect -3385 54595 -3280 54622
rect -3385 54531 -3365 54595
rect -3301 54531 -3280 54595
rect -3385 54512 -3280 54531
rect -1556 54595 -1453 54615
rect -1556 54531 -1536 54595
rect -1472 54531 -1453 54595
rect -1556 54511 -1453 54531
rect -9714 54403 -9452 54408
rect -9714 54339 -9695 54403
rect -9631 54339 -9615 54403
rect -9551 54339 -9535 54403
rect -9471 54339 -9452 54403
rect -9714 54334 -9452 54339
rect -7919 54402 -7657 54407
rect -7919 54338 -7900 54402
rect -7836 54338 -7820 54402
rect -7756 54338 -7740 54402
rect -7676 54338 -7657 54402
rect -7919 54333 -7657 54338
rect -6119 54404 -5857 54409
rect -6119 54340 -6100 54404
rect -6036 54340 -6020 54404
rect -5956 54340 -5940 54404
rect -5876 54340 -5857 54404
rect -6119 54335 -5857 54340
rect -4321 54403 -4059 54408
rect -4321 54339 -4302 54403
rect -4238 54339 -4222 54403
rect -4158 54339 -4142 54403
rect -4078 54339 -4059 54403
rect -4321 54334 -4059 54339
rect -2523 54404 -2261 54409
rect -2523 54340 -2504 54404
rect -2440 54340 -2424 54404
rect -2360 54340 -2344 54404
rect -2280 54340 -2261 54404
rect -2523 54335 -2261 54340
rect -720 54403 -458 54408
rect -720 54339 -701 54403
rect -637 54339 -621 54403
rect -557 54339 -541 54403
rect -477 54339 -458 54403
rect -720 54334 -458 54339
rect 156 54404 258 54424
rect 156 54340 176 54404
rect 240 54340 258 54404
rect 156 54319 258 54340
rect -7275 54019 -7265 54083
rect -7201 54019 -7191 54083
rect -1875 54019 -1865 54083
rect -1801 54019 -1791 54083
rect -8083 53766 -8073 53830
rect -8009 53766 -7999 53830
rect -2683 53766 -2673 53830
rect -2609 53766 -2599 53830
rect -10546 53338 -10536 53402
rect -10472 53338 -1865 53402
rect -1801 53338 -1791 53402
rect -11315 53082 -11305 53146
rect -11241 53082 -2673 53146
rect -2609 53082 -2599 53146
rect 337 53142 361 60806
rect 505 53142 529 60806
rect 337 53116 529 53142
rect 10167 60818 10561 60841
rect -12325 52649 -12315 52713
rect -12251 52649 -7265 52713
rect -7201 52649 -7191 52713
rect -13106 52326 -13096 52390
rect -13032 52326 -8073 52390
rect -8009 52326 -7999 52390
rect -8864 51243 -8760 51254
rect -8864 51179 -8844 51243
rect -8780 51179 -8760 51243
rect -8864 51163 -8760 51179
rect -8864 51099 -8844 51163
rect -8780 51099 -8760 51163
rect -7742 51247 -7634 51272
rect -7742 51183 -7722 51247
rect -7658 51183 -7634 51247
rect -7742 51162 -7634 51183
rect -8864 51083 -8760 51099
rect -8864 51019 -8844 51083
rect -8780 51019 -8760 51083
rect -8864 51009 -8760 51019
rect -5698 51046 -3878 51071
rect -5698 50902 -5660 51046
rect -3916 50902 -3878 51046
rect -5698 50878 -3878 50902
rect -3372 51057 -2526 51079
rect -3372 50913 -3341 51057
rect -2557 50913 -2526 51057
rect -3372 50891 -2526 50913
rect -1665 51047 -755 51069
rect -1665 50903 -1642 51047
rect -778 50903 -755 51047
rect -1665 50881 -755 50903
rect -8884 50776 -8770 50796
rect -8884 50712 -8859 50776
rect -8795 50712 -8770 50776
rect -88 50771 131 50779
rect -88 50735 -47 50771
rect 89 50735 131 50771
rect -8884 50696 -8770 50712
rect -8884 50632 -8859 50696
rect -8795 50632 -8770 50696
rect -8884 50617 -8770 50632
rect -19102 50616 -8770 50617
rect -19102 50596 -8859 50616
rect -19102 50532 -19005 50596
rect -18941 50552 -8859 50596
rect -8795 50552 -8770 50616
rect -18941 50536 -8770 50552
rect -18941 50532 -8859 50536
rect -19102 50512 -8859 50532
rect -8884 50472 -8859 50512
rect -8795 50472 -8770 50536
rect -8884 50456 -8770 50472
rect -5942 50720 -5738 50725
rect -8884 50392 -8859 50456
rect -8795 50392 -8770 50456
rect -8884 50373 -8770 50392
rect -8497 50441 -8398 50461
rect -8497 50377 -8480 50441
rect -8416 50377 -8398 50441
rect -8497 50357 -8398 50377
rect -57094 50072 -28000 50155
rect -57094 50008 -8480 50072
rect -8416 50008 -8406 50072
rect -57094 49919 -28000 50008
rect -27080 49720 -26716 49725
rect -27080 49656 -27050 49720
rect -26986 49656 -26970 49720
rect -26906 49656 -26890 49720
rect -26826 49656 -26810 49720
rect -26746 49656 -26716 49720
rect -27080 49651 -26716 49656
rect -26472 49418 -26408 50008
rect -26070 49424 -25986 49429
rect -26070 49420 -7722 49424
rect -26472 49409 -26147 49418
rect -26472 49353 -26391 49409
rect -26335 49353 -26311 49409
rect -26255 49353 -26231 49409
rect -26175 49353 -26147 49409
rect -26070 49364 -26056 49420
rect -26000 49364 -7722 49420
rect -26070 49360 -7722 49364
rect -7658 49360 -7648 49424
rect -26070 49355 -25986 49360
rect -26472 49349 -26147 49353
rect -26418 49344 -26147 49349
rect -25994 49178 -25630 49183
rect -25994 49114 -25964 49178
rect -25900 49114 -25884 49178
rect -25820 49114 -25804 49178
rect -25740 49114 -25724 49178
rect -25660 49114 -25630 49178
rect -25994 49109 -25630 49114
rect -5942 47776 -5912 50720
rect -5768 47776 -5738 50720
rect -5942 47771 -5738 47776
rect -88 47791 -51 50735
rect 93 47791 131 50735
rect -88 47755 -47 47791
rect 89 47755 131 47791
rect -88 47747 131 47755
rect 10167 47634 10212 60818
rect 10516 47634 10561 60818
rect 17420 60728 17506 60748
rect 17420 60664 17431 60728
rect 17495 60664 17506 60728
rect 17420 60648 17506 60664
rect 17420 60584 17431 60648
rect 17495 60584 17506 60648
rect 17420 60568 17506 60584
rect 17420 60504 17431 60568
rect 17495 60504 17506 60568
rect 17420 60488 17506 60504
rect 17420 60424 17431 60488
rect 17495 60424 17506 60488
rect 17420 60408 17506 60424
rect 17420 60344 17431 60408
rect 17495 60344 17506 60408
rect 17420 60328 17506 60344
rect 17420 60264 17431 60328
rect 17495 60264 17506 60328
rect 17420 60248 17506 60264
rect 17420 60184 17431 60248
rect 17495 60184 17506 60248
rect 17420 60164 17506 60184
rect 18508 60728 18594 60748
rect 18508 60664 18519 60728
rect 18583 60664 18594 60728
rect 18508 60648 18594 60664
rect 18508 60584 18519 60648
rect 18583 60584 18594 60648
rect 18508 60568 18594 60584
rect 18508 60504 18519 60568
rect 18583 60504 18594 60568
rect 18508 60488 18594 60504
rect 18508 60424 18519 60488
rect 18583 60424 18594 60488
rect 18508 60408 18594 60424
rect 18508 60344 18519 60408
rect 18583 60344 18594 60408
rect 18508 60328 18594 60344
rect 18508 60264 18519 60328
rect 18583 60264 18594 60328
rect 18508 60248 18594 60264
rect 18508 60184 18519 60248
rect 18583 60184 18594 60248
rect 18508 60164 18594 60184
rect 19596 60728 19682 60748
rect 19596 60664 19607 60728
rect 19671 60664 19682 60728
rect 19596 60648 19682 60664
rect 19596 60584 19607 60648
rect 19671 60584 19682 60648
rect 19596 60568 19682 60584
rect 19596 60504 19607 60568
rect 19671 60504 19682 60568
rect 19596 60488 19682 60504
rect 19596 60424 19607 60488
rect 19671 60424 19682 60488
rect 19596 60408 19682 60424
rect 19596 60344 19607 60408
rect 19671 60344 19682 60408
rect 19596 60328 19682 60344
rect 19596 60264 19607 60328
rect 19671 60264 19682 60328
rect 19596 60248 19682 60264
rect 19596 60184 19607 60248
rect 19671 60184 19682 60248
rect 19596 60164 19682 60184
rect 20684 60728 20770 60748
rect 20684 60664 20695 60728
rect 20759 60664 20770 60728
rect 20684 60648 20770 60664
rect 20684 60584 20695 60648
rect 20759 60584 20770 60648
rect 20684 60568 20770 60584
rect 20684 60504 20695 60568
rect 20759 60504 20770 60568
rect 20684 60488 20770 60504
rect 20684 60424 20695 60488
rect 20759 60424 20770 60488
rect 20684 60408 20770 60424
rect 20684 60344 20695 60408
rect 20759 60344 20770 60408
rect 20684 60328 20770 60344
rect 20684 60264 20695 60328
rect 20759 60264 20770 60328
rect 20684 60248 20770 60264
rect 20684 60184 20695 60248
rect 20759 60184 20770 60248
rect 20684 60164 20770 60184
rect 21772 60728 21858 60748
rect 21772 60664 21783 60728
rect 21847 60664 21858 60728
rect 21772 60648 21858 60664
rect 21772 60584 21783 60648
rect 21847 60584 21858 60648
rect 21772 60568 21858 60584
rect 21772 60504 21783 60568
rect 21847 60504 21858 60568
rect 21772 60488 21858 60504
rect 21772 60424 21783 60488
rect 21847 60424 21858 60488
rect 21772 60408 21858 60424
rect 21772 60344 21783 60408
rect 21847 60344 21858 60408
rect 21772 60328 21858 60344
rect 21772 60264 21783 60328
rect 21847 60264 21858 60328
rect 21772 60248 21858 60264
rect 21772 60184 21783 60248
rect 21847 60184 21858 60248
rect 21772 60164 21858 60184
rect 22860 60728 22946 60748
rect 22860 60664 22871 60728
rect 22935 60664 22946 60728
rect 22860 60648 22946 60664
rect 22860 60584 22871 60648
rect 22935 60584 22946 60648
rect 22860 60568 22946 60584
rect 22860 60504 22871 60568
rect 22935 60504 22946 60568
rect 22860 60488 22946 60504
rect 22860 60424 22871 60488
rect 22935 60424 22946 60488
rect 22860 60408 22946 60424
rect 22860 60344 22871 60408
rect 22935 60344 22946 60408
rect 22860 60328 22946 60344
rect 22860 60264 22871 60328
rect 22935 60264 22946 60328
rect 22860 60248 22946 60264
rect 22860 60184 22871 60248
rect 22935 60184 22946 60248
rect 22860 60164 22946 60184
rect 23948 60728 24034 60748
rect 23948 60664 23959 60728
rect 24023 60664 24034 60728
rect 23948 60648 24034 60664
rect 23948 60584 23959 60648
rect 24023 60584 24034 60648
rect 23948 60568 24034 60584
rect 23948 60504 23959 60568
rect 24023 60504 24034 60568
rect 23948 60488 24034 60504
rect 23948 60424 23959 60488
rect 24023 60424 24034 60488
rect 23948 60408 24034 60424
rect 23948 60344 23959 60408
rect 24023 60344 24034 60408
rect 23948 60328 24034 60344
rect 23948 60264 23959 60328
rect 24023 60264 24034 60328
rect 23948 60248 24034 60264
rect 23948 60184 23959 60248
rect 24023 60184 24034 60248
rect 23948 60164 24034 60184
rect 25036 60728 25122 60748
rect 25036 60664 25047 60728
rect 25111 60664 25122 60728
rect 25036 60648 25122 60664
rect 25036 60584 25047 60648
rect 25111 60584 25122 60648
rect 25036 60568 25122 60584
rect 25036 60504 25047 60568
rect 25111 60504 25122 60568
rect 25036 60488 25122 60504
rect 25036 60424 25047 60488
rect 25111 60424 25122 60488
rect 25036 60408 25122 60424
rect 25036 60344 25047 60408
rect 25111 60344 25122 60408
rect 25036 60328 25122 60344
rect 25036 60264 25047 60328
rect 25111 60264 25122 60328
rect 25036 60248 25122 60264
rect 25036 60184 25047 60248
rect 25111 60184 25122 60248
rect 25036 60164 25122 60184
rect 26124 60728 26210 60748
rect 26124 60664 26135 60728
rect 26199 60664 26210 60728
rect 26124 60648 26210 60664
rect 26124 60584 26135 60648
rect 26199 60584 26210 60648
rect 26124 60568 26210 60584
rect 26124 60504 26135 60568
rect 26199 60504 26210 60568
rect 26124 60488 26210 60504
rect 26124 60424 26135 60488
rect 26199 60424 26210 60488
rect 26124 60408 26210 60424
rect 26124 60344 26135 60408
rect 26199 60344 26210 60408
rect 26124 60328 26210 60344
rect 26124 60264 26135 60328
rect 26199 60264 26210 60328
rect 26124 60248 26210 60264
rect 26124 60184 26135 60248
rect 26199 60184 26210 60248
rect 26124 60164 26210 60184
rect 27212 60728 27298 60748
rect 27212 60664 27223 60728
rect 27287 60664 27298 60728
rect 27212 60648 27298 60664
rect 27212 60584 27223 60648
rect 27287 60584 27298 60648
rect 27212 60568 27298 60584
rect 27212 60504 27223 60568
rect 27287 60504 27298 60568
rect 27212 60488 27298 60504
rect 27212 60424 27223 60488
rect 27287 60424 27298 60488
rect 27212 60408 27298 60424
rect 27212 60344 27223 60408
rect 27287 60344 27298 60408
rect 27212 60328 27298 60344
rect 27212 60264 27223 60328
rect 27287 60264 27298 60328
rect 27212 60248 27298 60264
rect 27212 60184 27223 60248
rect 27287 60184 27298 60248
rect 27212 60164 27298 60184
rect 28300 60728 28386 60748
rect 28300 60664 28311 60728
rect 28375 60664 28386 60728
rect 28300 60648 28386 60664
rect 28300 60584 28311 60648
rect 28375 60584 28386 60648
rect 28300 60568 28386 60584
rect 28300 60504 28311 60568
rect 28375 60504 28386 60568
rect 28300 60488 28386 60504
rect 28300 60424 28311 60488
rect 28375 60424 28386 60488
rect 28300 60408 28386 60424
rect 28300 60344 28311 60408
rect 28375 60344 28386 60408
rect 28300 60328 28386 60344
rect 28300 60264 28311 60328
rect 28375 60264 28386 60328
rect 28300 60248 28386 60264
rect 28300 60184 28311 60248
rect 28375 60184 28386 60248
rect 28300 60164 28386 60184
rect 29388 60728 29474 60748
rect 29388 60664 29399 60728
rect 29463 60664 29474 60728
rect 29388 60648 29474 60664
rect 29388 60584 29399 60648
rect 29463 60584 29474 60648
rect 29388 60568 29474 60584
rect 29388 60504 29399 60568
rect 29463 60504 29474 60568
rect 29388 60488 29474 60504
rect 29388 60424 29399 60488
rect 29463 60424 29474 60488
rect 29388 60408 29474 60424
rect 29388 60344 29399 60408
rect 29463 60344 29474 60408
rect 29388 60328 29474 60344
rect 29388 60264 29399 60328
rect 29463 60264 29474 60328
rect 29388 60248 29474 60264
rect 29388 60184 29399 60248
rect 29463 60184 29474 60248
rect 29388 60164 29474 60184
rect 30476 60728 30562 60748
rect 30476 60664 30487 60728
rect 30551 60664 30562 60728
rect 30476 60648 30562 60664
rect 30476 60584 30487 60648
rect 30551 60584 30562 60648
rect 30476 60568 30562 60584
rect 30476 60504 30487 60568
rect 30551 60504 30562 60568
rect 30476 60488 30562 60504
rect 30476 60424 30487 60488
rect 30551 60424 30562 60488
rect 30476 60408 30562 60424
rect 30476 60344 30487 60408
rect 30551 60344 30562 60408
rect 30476 60328 30562 60344
rect 30476 60264 30487 60328
rect 30551 60264 30562 60328
rect 30476 60248 30562 60264
rect 30476 60184 30487 60248
rect 30551 60184 30562 60248
rect 30476 60164 30562 60184
rect 31564 60728 31650 60748
rect 31564 60664 31575 60728
rect 31639 60664 31650 60728
rect 31564 60648 31650 60664
rect 31564 60584 31575 60648
rect 31639 60584 31650 60648
rect 31564 60568 31650 60584
rect 31564 60504 31575 60568
rect 31639 60504 31650 60568
rect 31564 60488 31650 60504
rect 31564 60424 31575 60488
rect 31639 60424 31650 60488
rect 31564 60408 31650 60424
rect 31564 60344 31575 60408
rect 31639 60344 31650 60408
rect 31564 60328 31650 60344
rect 31564 60264 31575 60328
rect 31639 60264 31650 60328
rect 31564 60248 31650 60264
rect 31564 60184 31575 60248
rect 31639 60184 31650 60248
rect 31564 60164 31650 60184
rect 17965 58725 18051 58745
rect 17965 58661 17976 58725
rect 18040 58661 18051 58725
rect 17965 58645 18051 58661
rect 17965 58581 17976 58645
rect 18040 58581 18051 58645
rect 17965 58565 18051 58581
rect 17965 58501 17976 58565
rect 18040 58501 18051 58565
rect 17965 58485 18051 58501
rect 17965 58421 17976 58485
rect 18040 58421 18051 58485
rect 17965 58405 18051 58421
rect 17965 58341 17976 58405
rect 18040 58341 18051 58405
rect 17965 58325 18051 58341
rect 17965 58261 17976 58325
rect 18040 58261 18051 58325
rect 17965 58245 18051 58261
rect 17965 58181 17976 58245
rect 18040 58181 18051 58245
rect 17965 58161 18051 58181
rect 19053 58725 19139 58745
rect 19053 58661 19064 58725
rect 19128 58661 19139 58725
rect 19053 58645 19139 58661
rect 19053 58581 19064 58645
rect 19128 58581 19139 58645
rect 19053 58565 19139 58581
rect 19053 58501 19064 58565
rect 19128 58501 19139 58565
rect 19053 58485 19139 58501
rect 19053 58421 19064 58485
rect 19128 58421 19139 58485
rect 19053 58405 19139 58421
rect 19053 58341 19064 58405
rect 19128 58341 19139 58405
rect 19053 58325 19139 58341
rect 19053 58261 19064 58325
rect 19128 58261 19139 58325
rect 19053 58245 19139 58261
rect 19053 58181 19064 58245
rect 19128 58181 19139 58245
rect 19053 58161 19139 58181
rect 20141 58725 20227 58745
rect 20141 58661 20152 58725
rect 20216 58661 20227 58725
rect 20141 58645 20227 58661
rect 20141 58581 20152 58645
rect 20216 58581 20227 58645
rect 20141 58565 20227 58581
rect 20141 58501 20152 58565
rect 20216 58501 20227 58565
rect 20141 58485 20227 58501
rect 20141 58421 20152 58485
rect 20216 58421 20227 58485
rect 20141 58405 20227 58421
rect 20141 58341 20152 58405
rect 20216 58341 20227 58405
rect 20141 58325 20227 58341
rect 20141 58261 20152 58325
rect 20216 58261 20227 58325
rect 20141 58245 20227 58261
rect 20141 58181 20152 58245
rect 20216 58181 20227 58245
rect 20141 58161 20227 58181
rect 21229 58725 21315 58745
rect 21229 58661 21240 58725
rect 21304 58661 21315 58725
rect 21229 58645 21315 58661
rect 21229 58581 21240 58645
rect 21304 58581 21315 58645
rect 21229 58565 21315 58581
rect 21229 58501 21240 58565
rect 21304 58501 21315 58565
rect 21229 58485 21315 58501
rect 21229 58421 21240 58485
rect 21304 58421 21315 58485
rect 21229 58405 21315 58421
rect 21229 58341 21240 58405
rect 21304 58341 21315 58405
rect 21229 58325 21315 58341
rect 21229 58261 21240 58325
rect 21304 58261 21315 58325
rect 21229 58245 21315 58261
rect 21229 58181 21240 58245
rect 21304 58181 21315 58245
rect 21229 58161 21315 58181
rect 22317 58725 22403 58745
rect 22317 58661 22328 58725
rect 22392 58661 22403 58725
rect 22317 58645 22403 58661
rect 22317 58581 22328 58645
rect 22392 58581 22403 58645
rect 22317 58565 22403 58581
rect 22317 58501 22328 58565
rect 22392 58501 22403 58565
rect 22317 58485 22403 58501
rect 22317 58421 22328 58485
rect 22392 58421 22403 58485
rect 22317 58405 22403 58421
rect 22317 58341 22328 58405
rect 22392 58341 22403 58405
rect 22317 58325 22403 58341
rect 22317 58261 22328 58325
rect 22392 58261 22403 58325
rect 22317 58245 22403 58261
rect 22317 58181 22328 58245
rect 22392 58181 22403 58245
rect 22317 58161 22403 58181
rect 23405 58725 23491 58745
rect 23405 58661 23416 58725
rect 23480 58661 23491 58725
rect 23405 58645 23491 58661
rect 23405 58581 23416 58645
rect 23480 58581 23491 58645
rect 23405 58565 23491 58581
rect 23405 58501 23416 58565
rect 23480 58501 23491 58565
rect 23405 58485 23491 58501
rect 23405 58421 23416 58485
rect 23480 58421 23491 58485
rect 23405 58405 23491 58421
rect 23405 58341 23416 58405
rect 23480 58341 23491 58405
rect 23405 58325 23491 58341
rect 23405 58261 23416 58325
rect 23480 58261 23491 58325
rect 23405 58245 23491 58261
rect 23405 58181 23416 58245
rect 23480 58181 23491 58245
rect 23405 58161 23491 58181
rect 24493 58725 24579 58745
rect 24493 58661 24504 58725
rect 24568 58661 24579 58725
rect 24493 58645 24579 58661
rect 24493 58581 24504 58645
rect 24568 58581 24579 58645
rect 24493 58565 24579 58581
rect 24493 58501 24504 58565
rect 24568 58501 24579 58565
rect 24493 58485 24579 58501
rect 24493 58421 24504 58485
rect 24568 58421 24579 58485
rect 24493 58405 24579 58421
rect 24493 58341 24504 58405
rect 24568 58341 24579 58405
rect 24493 58325 24579 58341
rect 24493 58261 24504 58325
rect 24568 58261 24579 58325
rect 24493 58245 24579 58261
rect 24493 58181 24504 58245
rect 24568 58181 24579 58245
rect 24493 58161 24579 58181
rect 25581 58725 25667 58745
rect 25581 58661 25592 58725
rect 25656 58661 25667 58725
rect 25581 58645 25667 58661
rect 25581 58581 25592 58645
rect 25656 58581 25667 58645
rect 25581 58565 25667 58581
rect 25581 58501 25592 58565
rect 25656 58501 25667 58565
rect 25581 58485 25667 58501
rect 25581 58421 25592 58485
rect 25656 58421 25667 58485
rect 25581 58405 25667 58421
rect 25581 58341 25592 58405
rect 25656 58341 25667 58405
rect 25581 58325 25667 58341
rect 25581 58261 25592 58325
rect 25656 58261 25667 58325
rect 25581 58245 25667 58261
rect 25581 58181 25592 58245
rect 25656 58181 25667 58245
rect 25581 58161 25667 58181
rect 26669 58725 26755 58745
rect 26669 58661 26680 58725
rect 26744 58661 26755 58725
rect 26669 58645 26755 58661
rect 26669 58581 26680 58645
rect 26744 58581 26755 58645
rect 26669 58565 26755 58581
rect 26669 58501 26680 58565
rect 26744 58501 26755 58565
rect 26669 58485 26755 58501
rect 26669 58421 26680 58485
rect 26744 58421 26755 58485
rect 26669 58405 26755 58421
rect 26669 58341 26680 58405
rect 26744 58341 26755 58405
rect 26669 58325 26755 58341
rect 26669 58261 26680 58325
rect 26744 58261 26755 58325
rect 26669 58245 26755 58261
rect 26669 58181 26680 58245
rect 26744 58181 26755 58245
rect 26669 58161 26755 58181
rect 27757 58725 27843 58745
rect 27757 58661 27768 58725
rect 27832 58661 27843 58725
rect 27757 58645 27843 58661
rect 27757 58581 27768 58645
rect 27832 58581 27843 58645
rect 27757 58565 27843 58581
rect 27757 58501 27768 58565
rect 27832 58501 27843 58565
rect 27757 58485 27843 58501
rect 27757 58421 27768 58485
rect 27832 58421 27843 58485
rect 27757 58405 27843 58421
rect 27757 58341 27768 58405
rect 27832 58341 27843 58405
rect 27757 58325 27843 58341
rect 27757 58261 27768 58325
rect 27832 58261 27843 58325
rect 27757 58245 27843 58261
rect 27757 58181 27768 58245
rect 27832 58181 27843 58245
rect 27757 58161 27843 58181
rect 28845 58725 28931 58745
rect 28845 58661 28856 58725
rect 28920 58661 28931 58725
rect 28845 58645 28931 58661
rect 28845 58581 28856 58645
rect 28920 58581 28931 58645
rect 28845 58565 28931 58581
rect 28845 58501 28856 58565
rect 28920 58501 28931 58565
rect 28845 58485 28931 58501
rect 28845 58421 28856 58485
rect 28920 58421 28931 58485
rect 28845 58405 28931 58421
rect 28845 58341 28856 58405
rect 28920 58341 28931 58405
rect 28845 58325 28931 58341
rect 28845 58261 28856 58325
rect 28920 58261 28931 58325
rect 28845 58245 28931 58261
rect 28845 58181 28856 58245
rect 28920 58181 28931 58245
rect 28845 58161 28931 58181
rect 29933 58725 30019 58745
rect 29933 58661 29944 58725
rect 30008 58661 30019 58725
rect 29933 58645 30019 58661
rect 29933 58581 29944 58645
rect 30008 58581 30019 58645
rect 29933 58565 30019 58581
rect 29933 58501 29944 58565
rect 30008 58501 30019 58565
rect 29933 58485 30019 58501
rect 29933 58421 29944 58485
rect 30008 58421 30019 58485
rect 29933 58405 30019 58421
rect 29933 58341 29944 58405
rect 30008 58341 30019 58405
rect 29933 58325 30019 58341
rect 29933 58261 29944 58325
rect 30008 58261 30019 58325
rect 29933 58245 30019 58261
rect 29933 58181 29944 58245
rect 30008 58181 30019 58245
rect 29933 58161 30019 58181
rect 31021 58725 31107 58745
rect 31021 58661 31032 58725
rect 31096 58661 31107 58725
rect 31021 58645 31107 58661
rect 31021 58581 31032 58645
rect 31096 58581 31107 58645
rect 31021 58565 31107 58581
rect 31021 58501 31032 58565
rect 31096 58501 31107 58565
rect 31021 58485 31107 58501
rect 31021 58421 31032 58485
rect 31096 58421 31107 58485
rect 31021 58405 31107 58421
rect 31021 58341 31032 58405
rect 31096 58341 31107 58405
rect 31021 58325 31107 58341
rect 31021 58261 31032 58325
rect 31096 58261 31107 58325
rect 31021 58245 31107 58261
rect 31021 58181 31032 58245
rect 31096 58181 31107 58245
rect 31021 58161 31107 58181
rect 17420 56728 17506 56748
rect 17420 56664 17431 56728
rect 17495 56664 17506 56728
rect 17420 56648 17506 56664
rect 17420 56584 17431 56648
rect 17495 56584 17506 56648
rect 17420 56568 17506 56584
rect 17420 56504 17431 56568
rect 17495 56504 17506 56568
rect 17420 56488 17506 56504
rect 17420 56424 17431 56488
rect 17495 56424 17506 56488
rect 17420 56408 17506 56424
rect 17420 56344 17431 56408
rect 17495 56344 17506 56408
rect 17420 56328 17506 56344
rect 17420 56264 17431 56328
rect 17495 56264 17506 56328
rect 17420 56248 17506 56264
rect 17420 56184 17431 56248
rect 17495 56184 17506 56248
rect 17420 56164 17506 56184
rect 18508 56728 18594 56748
rect 18508 56664 18519 56728
rect 18583 56664 18594 56728
rect 18508 56648 18594 56664
rect 18508 56584 18519 56648
rect 18583 56584 18594 56648
rect 18508 56568 18594 56584
rect 18508 56504 18519 56568
rect 18583 56504 18594 56568
rect 18508 56488 18594 56504
rect 18508 56424 18519 56488
rect 18583 56424 18594 56488
rect 18508 56408 18594 56424
rect 18508 56344 18519 56408
rect 18583 56344 18594 56408
rect 18508 56328 18594 56344
rect 18508 56264 18519 56328
rect 18583 56264 18594 56328
rect 18508 56248 18594 56264
rect 18508 56184 18519 56248
rect 18583 56184 18594 56248
rect 18508 56164 18594 56184
rect 19596 56728 19682 56748
rect 19596 56664 19607 56728
rect 19671 56664 19682 56728
rect 19596 56648 19682 56664
rect 19596 56584 19607 56648
rect 19671 56584 19682 56648
rect 19596 56568 19682 56584
rect 19596 56504 19607 56568
rect 19671 56504 19682 56568
rect 19596 56488 19682 56504
rect 19596 56424 19607 56488
rect 19671 56424 19682 56488
rect 19596 56408 19682 56424
rect 19596 56344 19607 56408
rect 19671 56344 19682 56408
rect 19596 56328 19682 56344
rect 19596 56264 19607 56328
rect 19671 56264 19682 56328
rect 19596 56248 19682 56264
rect 19596 56184 19607 56248
rect 19671 56184 19682 56248
rect 19596 56164 19682 56184
rect 20684 56728 20770 56748
rect 20684 56664 20695 56728
rect 20759 56664 20770 56728
rect 20684 56648 20770 56664
rect 20684 56584 20695 56648
rect 20759 56584 20770 56648
rect 20684 56568 20770 56584
rect 20684 56504 20695 56568
rect 20759 56504 20770 56568
rect 20684 56488 20770 56504
rect 20684 56424 20695 56488
rect 20759 56424 20770 56488
rect 20684 56408 20770 56424
rect 20684 56344 20695 56408
rect 20759 56344 20770 56408
rect 20684 56328 20770 56344
rect 20684 56264 20695 56328
rect 20759 56264 20770 56328
rect 20684 56248 20770 56264
rect 20684 56184 20695 56248
rect 20759 56184 20770 56248
rect 20684 56164 20770 56184
rect 21772 56728 21858 56748
rect 21772 56664 21783 56728
rect 21847 56664 21858 56728
rect 21772 56648 21858 56664
rect 21772 56584 21783 56648
rect 21847 56584 21858 56648
rect 21772 56568 21858 56584
rect 21772 56504 21783 56568
rect 21847 56504 21858 56568
rect 21772 56488 21858 56504
rect 21772 56424 21783 56488
rect 21847 56424 21858 56488
rect 21772 56408 21858 56424
rect 21772 56344 21783 56408
rect 21847 56344 21858 56408
rect 21772 56328 21858 56344
rect 21772 56264 21783 56328
rect 21847 56264 21858 56328
rect 21772 56248 21858 56264
rect 21772 56184 21783 56248
rect 21847 56184 21858 56248
rect 21772 56164 21858 56184
rect 22860 56728 22946 56748
rect 22860 56664 22871 56728
rect 22935 56664 22946 56728
rect 22860 56648 22946 56664
rect 22860 56584 22871 56648
rect 22935 56584 22946 56648
rect 22860 56568 22946 56584
rect 22860 56504 22871 56568
rect 22935 56504 22946 56568
rect 22860 56488 22946 56504
rect 22860 56424 22871 56488
rect 22935 56424 22946 56488
rect 22860 56408 22946 56424
rect 22860 56344 22871 56408
rect 22935 56344 22946 56408
rect 22860 56328 22946 56344
rect 22860 56264 22871 56328
rect 22935 56264 22946 56328
rect 22860 56248 22946 56264
rect 22860 56184 22871 56248
rect 22935 56184 22946 56248
rect 22860 56164 22946 56184
rect 23948 56728 24034 56748
rect 23948 56664 23959 56728
rect 24023 56664 24034 56728
rect 23948 56648 24034 56664
rect 23948 56584 23959 56648
rect 24023 56584 24034 56648
rect 23948 56568 24034 56584
rect 23948 56504 23959 56568
rect 24023 56504 24034 56568
rect 23948 56488 24034 56504
rect 23948 56424 23959 56488
rect 24023 56424 24034 56488
rect 23948 56408 24034 56424
rect 23948 56344 23959 56408
rect 24023 56344 24034 56408
rect 23948 56328 24034 56344
rect 23948 56264 23959 56328
rect 24023 56264 24034 56328
rect 23948 56248 24034 56264
rect 23948 56184 23959 56248
rect 24023 56184 24034 56248
rect 23948 56164 24034 56184
rect 25036 56728 25122 56748
rect 25036 56664 25047 56728
rect 25111 56664 25122 56728
rect 25036 56648 25122 56664
rect 25036 56584 25047 56648
rect 25111 56584 25122 56648
rect 25036 56568 25122 56584
rect 25036 56504 25047 56568
rect 25111 56504 25122 56568
rect 25036 56488 25122 56504
rect 25036 56424 25047 56488
rect 25111 56424 25122 56488
rect 25036 56408 25122 56424
rect 25036 56344 25047 56408
rect 25111 56344 25122 56408
rect 25036 56328 25122 56344
rect 25036 56264 25047 56328
rect 25111 56264 25122 56328
rect 25036 56248 25122 56264
rect 25036 56184 25047 56248
rect 25111 56184 25122 56248
rect 25036 56164 25122 56184
rect 26124 56728 26210 56748
rect 26124 56664 26135 56728
rect 26199 56664 26210 56728
rect 26124 56648 26210 56664
rect 26124 56584 26135 56648
rect 26199 56584 26210 56648
rect 26124 56568 26210 56584
rect 26124 56504 26135 56568
rect 26199 56504 26210 56568
rect 26124 56488 26210 56504
rect 26124 56424 26135 56488
rect 26199 56424 26210 56488
rect 26124 56408 26210 56424
rect 26124 56344 26135 56408
rect 26199 56344 26210 56408
rect 26124 56328 26210 56344
rect 26124 56264 26135 56328
rect 26199 56264 26210 56328
rect 26124 56248 26210 56264
rect 26124 56184 26135 56248
rect 26199 56184 26210 56248
rect 26124 56164 26210 56184
rect 27212 56728 27298 56748
rect 27212 56664 27223 56728
rect 27287 56664 27298 56728
rect 27212 56648 27298 56664
rect 27212 56584 27223 56648
rect 27287 56584 27298 56648
rect 27212 56568 27298 56584
rect 27212 56504 27223 56568
rect 27287 56504 27298 56568
rect 27212 56488 27298 56504
rect 27212 56424 27223 56488
rect 27287 56424 27298 56488
rect 27212 56408 27298 56424
rect 27212 56344 27223 56408
rect 27287 56344 27298 56408
rect 27212 56328 27298 56344
rect 27212 56264 27223 56328
rect 27287 56264 27298 56328
rect 27212 56248 27298 56264
rect 27212 56184 27223 56248
rect 27287 56184 27298 56248
rect 27212 56164 27298 56184
rect 28300 56728 28386 56748
rect 28300 56664 28311 56728
rect 28375 56664 28386 56728
rect 28300 56648 28386 56664
rect 28300 56584 28311 56648
rect 28375 56584 28386 56648
rect 28300 56568 28386 56584
rect 28300 56504 28311 56568
rect 28375 56504 28386 56568
rect 28300 56488 28386 56504
rect 28300 56424 28311 56488
rect 28375 56424 28386 56488
rect 28300 56408 28386 56424
rect 28300 56344 28311 56408
rect 28375 56344 28386 56408
rect 28300 56328 28386 56344
rect 28300 56264 28311 56328
rect 28375 56264 28386 56328
rect 28300 56248 28386 56264
rect 28300 56184 28311 56248
rect 28375 56184 28386 56248
rect 28300 56164 28386 56184
rect 29388 56728 29474 56748
rect 29388 56664 29399 56728
rect 29463 56664 29474 56728
rect 29388 56648 29474 56664
rect 29388 56584 29399 56648
rect 29463 56584 29474 56648
rect 29388 56568 29474 56584
rect 29388 56504 29399 56568
rect 29463 56504 29474 56568
rect 29388 56488 29474 56504
rect 29388 56424 29399 56488
rect 29463 56424 29474 56488
rect 29388 56408 29474 56424
rect 29388 56344 29399 56408
rect 29463 56344 29474 56408
rect 29388 56328 29474 56344
rect 29388 56264 29399 56328
rect 29463 56264 29474 56328
rect 29388 56248 29474 56264
rect 29388 56184 29399 56248
rect 29463 56184 29474 56248
rect 29388 56164 29474 56184
rect 30476 56728 30562 56748
rect 30476 56664 30487 56728
rect 30551 56664 30562 56728
rect 30476 56648 30562 56664
rect 30476 56584 30487 56648
rect 30551 56584 30562 56648
rect 30476 56568 30562 56584
rect 30476 56504 30487 56568
rect 30551 56504 30562 56568
rect 30476 56488 30562 56504
rect 30476 56424 30487 56488
rect 30551 56424 30562 56488
rect 30476 56408 30562 56424
rect 30476 56344 30487 56408
rect 30551 56344 30562 56408
rect 30476 56328 30562 56344
rect 30476 56264 30487 56328
rect 30551 56264 30562 56328
rect 30476 56248 30562 56264
rect 30476 56184 30487 56248
rect 30551 56184 30562 56248
rect 30476 56164 30562 56184
rect 31564 56728 31650 56748
rect 31564 56664 31575 56728
rect 31639 56664 31650 56728
rect 31564 56648 31650 56664
rect 31564 56584 31575 56648
rect 31639 56584 31650 56648
rect 31564 56568 31650 56584
rect 31564 56504 31575 56568
rect 31639 56504 31650 56568
rect 31564 56488 31650 56504
rect 31564 56424 31575 56488
rect 31639 56424 31650 56488
rect 31564 56408 31650 56424
rect 31564 56344 31575 56408
rect 31639 56344 31650 56408
rect 31564 56328 31650 56344
rect 31564 56264 31575 56328
rect 31639 56264 31650 56328
rect 31564 56248 31650 56264
rect 31564 56184 31575 56248
rect 31639 56184 31650 56248
rect 31564 56164 31650 56184
rect 52756 55101 62907 55337
rect 17965 54725 18051 54745
rect 17965 54661 17976 54725
rect 18040 54661 18051 54725
rect 17965 54645 18051 54661
rect 17965 54581 17976 54645
rect 18040 54581 18051 54645
rect 17965 54565 18051 54581
rect 17965 54501 17976 54565
rect 18040 54501 18051 54565
rect 17965 54485 18051 54501
rect 17965 54421 17976 54485
rect 18040 54421 18051 54485
rect 17965 54405 18051 54421
rect 17965 54341 17976 54405
rect 18040 54341 18051 54405
rect 17965 54325 18051 54341
rect 17965 54261 17976 54325
rect 18040 54261 18051 54325
rect 17965 54245 18051 54261
rect 17965 54181 17976 54245
rect 18040 54181 18051 54245
rect 17965 54161 18051 54181
rect 19053 54725 19139 54745
rect 19053 54661 19064 54725
rect 19128 54661 19139 54725
rect 19053 54645 19139 54661
rect 19053 54581 19064 54645
rect 19128 54581 19139 54645
rect 19053 54565 19139 54581
rect 19053 54501 19064 54565
rect 19128 54501 19139 54565
rect 19053 54485 19139 54501
rect 19053 54421 19064 54485
rect 19128 54421 19139 54485
rect 19053 54405 19139 54421
rect 19053 54341 19064 54405
rect 19128 54341 19139 54405
rect 19053 54325 19139 54341
rect 19053 54261 19064 54325
rect 19128 54261 19139 54325
rect 19053 54245 19139 54261
rect 19053 54181 19064 54245
rect 19128 54181 19139 54245
rect 19053 54161 19139 54181
rect 20141 54725 20227 54745
rect 20141 54661 20152 54725
rect 20216 54661 20227 54725
rect 20141 54645 20227 54661
rect 20141 54581 20152 54645
rect 20216 54581 20227 54645
rect 20141 54565 20227 54581
rect 20141 54501 20152 54565
rect 20216 54501 20227 54565
rect 20141 54485 20227 54501
rect 20141 54421 20152 54485
rect 20216 54421 20227 54485
rect 20141 54405 20227 54421
rect 20141 54341 20152 54405
rect 20216 54341 20227 54405
rect 20141 54325 20227 54341
rect 20141 54261 20152 54325
rect 20216 54261 20227 54325
rect 20141 54245 20227 54261
rect 20141 54181 20152 54245
rect 20216 54181 20227 54245
rect 20141 54161 20227 54181
rect 21229 54725 21315 54745
rect 21229 54661 21240 54725
rect 21304 54661 21315 54725
rect 21229 54645 21315 54661
rect 21229 54581 21240 54645
rect 21304 54581 21315 54645
rect 21229 54565 21315 54581
rect 21229 54501 21240 54565
rect 21304 54501 21315 54565
rect 21229 54485 21315 54501
rect 21229 54421 21240 54485
rect 21304 54421 21315 54485
rect 21229 54405 21315 54421
rect 21229 54341 21240 54405
rect 21304 54341 21315 54405
rect 21229 54325 21315 54341
rect 21229 54261 21240 54325
rect 21304 54261 21315 54325
rect 21229 54245 21315 54261
rect 21229 54181 21240 54245
rect 21304 54181 21315 54245
rect 21229 54161 21315 54181
rect 22317 54725 22403 54745
rect 22317 54661 22328 54725
rect 22392 54661 22403 54725
rect 22317 54645 22403 54661
rect 22317 54581 22328 54645
rect 22392 54581 22403 54645
rect 22317 54565 22403 54581
rect 22317 54501 22328 54565
rect 22392 54501 22403 54565
rect 22317 54485 22403 54501
rect 22317 54421 22328 54485
rect 22392 54421 22403 54485
rect 22317 54405 22403 54421
rect 22317 54341 22328 54405
rect 22392 54341 22403 54405
rect 22317 54325 22403 54341
rect 22317 54261 22328 54325
rect 22392 54261 22403 54325
rect 22317 54245 22403 54261
rect 22317 54181 22328 54245
rect 22392 54181 22403 54245
rect 22317 54161 22403 54181
rect 23405 54725 23491 54745
rect 23405 54661 23416 54725
rect 23480 54661 23491 54725
rect 23405 54645 23491 54661
rect 23405 54581 23416 54645
rect 23480 54581 23491 54645
rect 23405 54565 23491 54581
rect 23405 54501 23416 54565
rect 23480 54501 23491 54565
rect 23405 54485 23491 54501
rect 23405 54421 23416 54485
rect 23480 54421 23491 54485
rect 23405 54405 23491 54421
rect 23405 54341 23416 54405
rect 23480 54341 23491 54405
rect 23405 54325 23491 54341
rect 23405 54261 23416 54325
rect 23480 54261 23491 54325
rect 23405 54245 23491 54261
rect 23405 54181 23416 54245
rect 23480 54181 23491 54245
rect 23405 54161 23491 54181
rect 24493 54725 24579 54745
rect 24493 54661 24504 54725
rect 24568 54661 24579 54725
rect 24493 54645 24579 54661
rect 24493 54581 24504 54645
rect 24568 54581 24579 54645
rect 24493 54565 24579 54581
rect 24493 54501 24504 54565
rect 24568 54501 24579 54565
rect 24493 54485 24579 54501
rect 24493 54421 24504 54485
rect 24568 54421 24579 54485
rect 24493 54405 24579 54421
rect 24493 54341 24504 54405
rect 24568 54341 24579 54405
rect 24493 54325 24579 54341
rect 24493 54261 24504 54325
rect 24568 54261 24579 54325
rect 24493 54245 24579 54261
rect 24493 54181 24504 54245
rect 24568 54181 24579 54245
rect 24493 54161 24579 54181
rect 25581 54725 25667 54745
rect 25581 54661 25592 54725
rect 25656 54661 25667 54725
rect 25581 54645 25667 54661
rect 25581 54581 25592 54645
rect 25656 54581 25667 54645
rect 25581 54565 25667 54581
rect 25581 54501 25592 54565
rect 25656 54501 25667 54565
rect 25581 54485 25667 54501
rect 25581 54421 25592 54485
rect 25656 54421 25667 54485
rect 25581 54405 25667 54421
rect 25581 54341 25592 54405
rect 25656 54341 25667 54405
rect 25581 54325 25667 54341
rect 25581 54261 25592 54325
rect 25656 54261 25667 54325
rect 25581 54245 25667 54261
rect 25581 54181 25592 54245
rect 25656 54181 25667 54245
rect 25581 54161 25667 54181
rect 26669 54725 26755 54745
rect 26669 54661 26680 54725
rect 26744 54661 26755 54725
rect 26669 54645 26755 54661
rect 26669 54581 26680 54645
rect 26744 54581 26755 54645
rect 26669 54565 26755 54581
rect 26669 54501 26680 54565
rect 26744 54501 26755 54565
rect 26669 54485 26755 54501
rect 26669 54421 26680 54485
rect 26744 54421 26755 54485
rect 26669 54405 26755 54421
rect 26669 54341 26680 54405
rect 26744 54341 26755 54405
rect 26669 54325 26755 54341
rect 26669 54261 26680 54325
rect 26744 54261 26755 54325
rect 26669 54245 26755 54261
rect 26669 54181 26680 54245
rect 26744 54181 26755 54245
rect 26669 54161 26755 54181
rect 27757 54725 27843 54745
rect 27757 54661 27768 54725
rect 27832 54661 27843 54725
rect 27757 54645 27843 54661
rect 27757 54581 27768 54645
rect 27832 54581 27843 54645
rect 27757 54565 27843 54581
rect 27757 54501 27768 54565
rect 27832 54501 27843 54565
rect 27757 54485 27843 54501
rect 27757 54421 27768 54485
rect 27832 54421 27843 54485
rect 27757 54405 27843 54421
rect 27757 54341 27768 54405
rect 27832 54341 27843 54405
rect 27757 54325 27843 54341
rect 27757 54261 27768 54325
rect 27832 54261 27843 54325
rect 27757 54245 27843 54261
rect 27757 54181 27768 54245
rect 27832 54181 27843 54245
rect 27757 54161 27843 54181
rect 28845 54725 28931 54745
rect 28845 54661 28856 54725
rect 28920 54661 28931 54725
rect 28845 54645 28931 54661
rect 28845 54581 28856 54645
rect 28920 54581 28931 54645
rect 28845 54565 28931 54581
rect 28845 54501 28856 54565
rect 28920 54501 28931 54565
rect 28845 54485 28931 54501
rect 28845 54421 28856 54485
rect 28920 54421 28931 54485
rect 28845 54405 28931 54421
rect 28845 54341 28856 54405
rect 28920 54341 28931 54405
rect 28845 54325 28931 54341
rect 28845 54261 28856 54325
rect 28920 54261 28931 54325
rect 28845 54245 28931 54261
rect 28845 54181 28856 54245
rect 28920 54181 28931 54245
rect 28845 54161 28931 54181
rect 29933 54725 30019 54745
rect 29933 54661 29944 54725
rect 30008 54661 30019 54725
rect 29933 54645 30019 54661
rect 29933 54581 29944 54645
rect 30008 54581 30019 54645
rect 29933 54565 30019 54581
rect 29933 54501 29944 54565
rect 30008 54501 30019 54565
rect 29933 54485 30019 54501
rect 29933 54421 29944 54485
rect 30008 54421 30019 54485
rect 29933 54405 30019 54421
rect 29933 54341 29944 54405
rect 30008 54341 30019 54405
rect 29933 54325 30019 54341
rect 29933 54261 29944 54325
rect 30008 54261 30019 54325
rect 29933 54245 30019 54261
rect 29933 54181 29944 54245
rect 30008 54181 30019 54245
rect 29933 54161 30019 54181
rect 31021 54725 31107 54745
rect 31021 54661 31032 54725
rect 31096 54661 31107 54725
rect 31021 54645 31107 54661
rect 31021 54581 31032 54645
rect 31096 54581 31107 54645
rect 31021 54565 31107 54581
rect 31021 54501 31032 54565
rect 31096 54501 31107 54565
rect 31021 54485 31107 54501
rect 31021 54421 31032 54485
rect 31096 54421 31107 54485
rect 31021 54405 31107 54421
rect 31021 54341 31032 54405
rect 31096 54341 31107 54405
rect 31021 54325 31107 54341
rect 31021 54261 31032 54325
rect 31096 54261 31107 54325
rect 31021 54245 31107 54261
rect 31021 54181 31032 54245
rect 31096 54181 31107 54245
rect 31021 54161 31107 54181
rect 17420 52728 17506 52748
rect 17420 52664 17431 52728
rect 17495 52664 17506 52728
rect 17420 52648 17506 52664
rect 17420 52584 17431 52648
rect 17495 52584 17506 52648
rect 17420 52568 17506 52584
rect 17420 52504 17431 52568
rect 17495 52504 17506 52568
rect 17420 52488 17506 52504
rect 17420 52424 17431 52488
rect 17495 52424 17506 52488
rect 17420 52408 17506 52424
rect 17420 52344 17431 52408
rect 17495 52344 17506 52408
rect 17420 52328 17506 52344
rect 17420 52264 17431 52328
rect 17495 52264 17506 52328
rect 17420 52248 17506 52264
rect 17420 52184 17431 52248
rect 17495 52184 17506 52248
rect 17420 52164 17506 52184
rect 18508 52728 18594 52748
rect 18508 52664 18519 52728
rect 18583 52664 18594 52728
rect 18508 52648 18594 52664
rect 18508 52584 18519 52648
rect 18583 52584 18594 52648
rect 18508 52568 18594 52584
rect 18508 52504 18519 52568
rect 18583 52504 18594 52568
rect 18508 52488 18594 52504
rect 18508 52424 18519 52488
rect 18583 52424 18594 52488
rect 18508 52408 18594 52424
rect 18508 52344 18519 52408
rect 18583 52344 18594 52408
rect 18508 52328 18594 52344
rect 18508 52264 18519 52328
rect 18583 52264 18594 52328
rect 18508 52248 18594 52264
rect 18508 52184 18519 52248
rect 18583 52184 18594 52248
rect 18508 52164 18594 52184
rect 19596 52728 19682 52748
rect 19596 52664 19607 52728
rect 19671 52664 19682 52728
rect 19596 52648 19682 52664
rect 19596 52584 19607 52648
rect 19671 52584 19682 52648
rect 19596 52568 19682 52584
rect 19596 52504 19607 52568
rect 19671 52504 19682 52568
rect 19596 52488 19682 52504
rect 19596 52424 19607 52488
rect 19671 52424 19682 52488
rect 19596 52408 19682 52424
rect 19596 52344 19607 52408
rect 19671 52344 19682 52408
rect 19596 52328 19682 52344
rect 19596 52264 19607 52328
rect 19671 52264 19682 52328
rect 19596 52248 19682 52264
rect 19596 52184 19607 52248
rect 19671 52184 19682 52248
rect 19596 52164 19682 52184
rect 20684 52728 20770 52748
rect 20684 52664 20695 52728
rect 20759 52664 20770 52728
rect 20684 52648 20770 52664
rect 20684 52584 20695 52648
rect 20759 52584 20770 52648
rect 20684 52568 20770 52584
rect 20684 52504 20695 52568
rect 20759 52504 20770 52568
rect 20684 52488 20770 52504
rect 20684 52424 20695 52488
rect 20759 52424 20770 52488
rect 20684 52408 20770 52424
rect 20684 52344 20695 52408
rect 20759 52344 20770 52408
rect 20684 52328 20770 52344
rect 20684 52264 20695 52328
rect 20759 52264 20770 52328
rect 20684 52248 20770 52264
rect 20684 52184 20695 52248
rect 20759 52184 20770 52248
rect 20684 52164 20770 52184
rect 21772 52728 21858 52748
rect 21772 52664 21783 52728
rect 21847 52664 21858 52728
rect 21772 52648 21858 52664
rect 21772 52584 21783 52648
rect 21847 52584 21858 52648
rect 21772 52568 21858 52584
rect 21772 52504 21783 52568
rect 21847 52504 21858 52568
rect 21772 52488 21858 52504
rect 21772 52424 21783 52488
rect 21847 52424 21858 52488
rect 21772 52408 21858 52424
rect 21772 52344 21783 52408
rect 21847 52344 21858 52408
rect 21772 52328 21858 52344
rect 21772 52264 21783 52328
rect 21847 52264 21858 52328
rect 21772 52248 21858 52264
rect 21772 52184 21783 52248
rect 21847 52184 21858 52248
rect 21772 52164 21858 52184
rect 22860 52728 22946 52748
rect 22860 52664 22871 52728
rect 22935 52664 22946 52728
rect 22860 52648 22946 52664
rect 22860 52584 22871 52648
rect 22935 52584 22946 52648
rect 22860 52568 22946 52584
rect 22860 52504 22871 52568
rect 22935 52504 22946 52568
rect 22860 52488 22946 52504
rect 22860 52424 22871 52488
rect 22935 52424 22946 52488
rect 22860 52408 22946 52424
rect 22860 52344 22871 52408
rect 22935 52344 22946 52408
rect 22860 52328 22946 52344
rect 22860 52264 22871 52328
rect 22935 52264 22946 52328
rect 22860 52248 22946 52264
rect 22860 52184 22871 52248
rect 22935 52184 22946 52248
rect 22860 52164 22946 52184
rect 23948 52728 24034 52748
rect 23948 52664 23959 52728
rect 24023 52664 24034 52728
rect 23948 52648 24034 52664
rect 23948 52584 23959 52648
rect 24023 52584 24034 52648
rect 23948 52568 24034 52584
rect 23948 52504 23959 52568
rect 24023 52504 24034 52568
rect 23948 52488 24034 52504
rect 23948 52424 23959 52488
rect 24023 52424 24034 52488
rect 23948 52408 24034 52424
rect 23948 52344 23959 52408
rect 24023 52344 24034 52408
rect 23948 52328 24034 52344
rect 23948 52264 23959 52328
rect 24023 52264 24034 52328
rect 23948 52248 24034 52264
rect 23948 52184 23959 52248
rect 24023 52184 24034 52248
rect 23948 52164 24034 52184
rect 25036 52728 25122 52748
rect 25036 52664 25047 52728
rect 25111 52664 25122 52728
rect 25036 52648 25122 52664
rect 25036 52584 25047 52648
rect 25111 52584 25122 52648
rect 25036 52568 25122 52584
rect 25036 52504 25047 52568
rect 25111 52504 25122 52568
rect 25036 52488 25122 52504
rect 25036 52424 25047 52488
rect 25111 52424 25122 52488
rect 25036 52408 25122 52424
rect 25036 52344 25047 52408
rect 25111 52344 25122 52408
rect 25036 52328 25122 52344
rect 25036 52264 25047 52328
rect 25111 52264 25122 52328
rect 25036 52248 25122 52264
rect 25036 52184 25047 52248
rect 25111 52184 25122 52248
rect 25036 52164 25122 52184
rect 26124 52728 26210 52748
rect 26124 52664 26135 52728
rect 26199 52664 26210 52728
rect 26124 52648 26210 52664
rect 26124 52584 26135 52648
rect 26199 52584 26210 52648
rect 26124 52568 26210 52584
rect 26124 52504 26135 52568
rect 26199 52504 26210 52568
rect 26124 52488 26210 52504
rect 26124 52424 26135 52488
rect 26199 52424 26210 52488
rect 26124 52408 26210 52424
rect 26124 52344 26135 52408
rect 26199 52344 26210 52408
rect 26124 52328 26210 52344
rect 26124 52264 26135 52328
rect 26199 52264 26210 52328
rect 26124 52248 26210 52264
rect 26124 52184 26135 52248
rect 26199 52184 26210 52248
rect 26124 52164 26210 52184
rect 27212 52728 27298 52748
rect 27212 52664 27223 52728
rect 27287 52664 27298 52728
rect 27212 52648 27298 52664
rect 27212 52584 27223 52648
rect 27287 52584 27298 52648
rect 27212 52568 27298 52584
rect 27212 52504 27223 52568
rect 27287 52504 27298 52568
rect 27212 52488 27298 52504
rect 27212 52424 27223 52488
rect 27287 52424 27298 52488
rect 27212 52408 27298 52424
rect 27212 52344 27223 52408
rect 27287 52344 27298 52408
rect 27212 52328 27298 52344
rect 27212 52264 27223 52328
rect 27287 52264 27298 52328
rect 27212 52248 27298 52264
rect 27212 52184 27223 52248
rect 27287 52184 27298 52248
rect 27212 52164 27298 52184
rect 28300 52728 28386 52748
rect 28300 52664 28311 52728
rect 28375 52664 28386 52728
rect 28300 52648 28386 52664
rect 28300 52584 28311 52648
rect 28375 52584 28386 52648
rect 28300 52568 28386 52584
rect 28300 52504 28311 52568
rect 28375 52504 28386 52568
rect 28300 52488 28386 52504
rect 28300 52424 28311 52488
rect 28375 52424 28386 52488
rect 28300 52408 28386 52424
rect 28300 52344 28311 52408
rect 28375 52344 28386 52408
rect 28300 52328 28386 52344
rect 28300 52264 28311 52328
rect 28375 52264 28386 52328
rect 28300 52248 28386 52264
rect 28300 52184 28311 52248
rect 28375 52184 28386 52248
rect 28300 52164 28386 52184
rect 29388 52728 29474 52748
rect 29388 52664 29399 52728
rect 29463 52664 29474 52728
rect 29388 52648 29474 52664
rect 29388 52584 29399 52648
rect 29463 52584 29474 52648
rect 29388 52568 29474 52584
rect 29388 52504 29399 52568
rect 29463 52504 29474 52568
rect 29388 52488 29474 52504
rect 29388 52424 29399 52488
rect 29463 52424 29474 52488
rect 29388 52408 29474 52424
rect 29388 52344 29399 52408
rect 29463 52344 29474 52408
rect 29388 52328 29474 52344
rect 29388 52264 29399 52328
rect 29463 52264 29474 52328
rect 29388 52248 29474 52264
rect 29388 52184 29399 52248
rect 29463 52184 29474 52248
rect 29388 52164 29474 52184
rect 30476 52728 30562 52748
rect 30476 52664 30487 52728
rect 30551 52664 30562 52728
rect 30476 52648 30562 52664
rect 30476 52584 30487 52648
rect 30551 52584 30562 52648
rect 30476 52568 30562 52584
rect 30476 52504 30487 52568
rect 30551 52504 30562 52568
rect 30476 52488 30562 52504
rect 30476 52424 30487 52488
rect 30551 52424 30562 52488
rect 30476 52408 30562 52424
rect 30476 52344 30487 52408
rect 30551 52344 30562 52408
rect 30476 52328 30562 52344
rect 30476 52264 30487 52328
rect 30551 52264 30562 52328
rect 30476 52248 30562 52264
rect 30476 52184 30487 52248
rect 30551 52184 30562 52248
rect 30476 52164 30562 52184
rect 31564 52728 31650 52748
rect 31564 52664 31575 52728
rect 31639 52664 31650 52728
rect 31564 52648 31650 52664
rect 31564 52584 31575 52648
rect 31639 52584 31650 52648
rect 31564 52568 31650 52584
rect 31564 52504 31575 52568
rect 31639 52504 31650 52568
rect 31564 52488 31650 52504
rect 31564 52424 31575 52488
rect 31639 52424 31650 52488
rect 31564 52408 31650 52424
rect 31564 52344 31575 52408
rect 31639 52344 31650 52408
rect 31564 52328 31650 52344
rect 31564 52264 31575 52328
rect 31639 52264 31650 52328
rect 31564 52248 31650 52264
rect 31564 52184 31575 52248
rect 31639 52184 31650 52248
rect 31564 52164 31650 52184
rect 17965 50725 18051 50745
rect 17965 50661 17976 50725
rect 18040 50661 18051 50725
rect 17965 50645 18051 50661
rect 17965 50581 17976 50645
rect 18040 50581 18051 50645
rect 17965 50565 18051 50581
rect 17965 50501 17976 50565
rect 18040 50501 18051 50565
rect 17965 50485 18051 50501
rect 17965 50421 17976 50485
rect 18040 50421 18051 50485
rect 17965 50405 18051 50421
rect 17965 50341 17976 50405
rect 18040 50341 18051 50405
rect 17965 50325 18051 50341
rect 17965 50261 17976 50325
rect 18040 50261 18051 50325
rect 17965 50245 18051 50261
rect 17965 50181 17976 50245
rect 18040 50181 18051 50245
rect 17965 50161 18051 50181
rect 20141 50725 20227 50745
rect 20141 50661 20152 50725
rect 20216 50661 20227 50725
rect 20141 50645 20227 50661
rect 20141 50581 20152 50645
rect 20216 50581 20227 50645
rect 20141 50565 20227 50581
rect 20141 50501 20152 50565
rect 20216 50501 20227 50565
rect 20141 50485 20227 50501
rect 20141 50421 20152 50485
rect 20216 50421 20227 50485
rect 20141 50405 20227 50421
rect 20141 50341 20152 50405
rect 20216 50341 20227 50405
rect 20141 50325 20227 50341
rect 20141 50261 20152 50325
rect 20216 50261 20227 50325
rect 20141 50245 20227 50261
rect 20141 50181 20152 50245
rect 20216 50181 20227 50245
rect 20141 50161 20227 50181
rect 21229 50725 21315 50745
rect 21229 50661 21240 50725
rect 21304 50661 21315 50725
rect 21229 50645 21315 50661
rect 21229 50581 21240 50645
rect 21304 50581 21315 50645
rect 21229 50565 21315 50581
rect 21229 50501 21240 50565
rect 21304 50501 21315 50565
rect 21229 50485 21315 50501
rect 21229 50421 21240 50485
rect 21304 50421 21315 50485
rect 21229 50405 21315 50421
rect 21229 50341 21240 50405
rect 21304 50341 21315 50405
rect 21229 50325 21315 50341
rect 21229 50261 21240 50325
rect 21304 50261 21315 50325
rect 21229 50245 21315 50261
rect 21229 50181 21240 50245
rect 21304 50181 21315 50245
rect 21229 50161 21315 50181
rect 23405 50725 23491 50745
rect 23405 50661 23416 50725
rect 23480 50661 23491 50725
rect 23405 50645 23491 50661
rect 23405 50581 23416 50645
rect 23480 50581 23491 50645
rect 23405 50565 23491 50581
rect 23405 50501 23416 50565
rect 23480 50501 23491 50565
rect 23405 50485 23491 50501
rect 23405 50421 23416 50485
rect 23480 50421 23491 50485
rect 23405 50405 23491 50421
rect 23405 50341 23416 50405
rect 23480 50341 23491 50405
rect 23405 50325 23491 50341
rect 23405 50261 23416 50325
rect 23480 50261 23491 50325
rect 23405 50245 23491 50261
rect 23405 50181 23416 50245
rect 23480 50181 23491 50245
rect 23405 50161 23491 50181
rect 24493 50725 24579 50745
rect 24493 50661 24504 50725
rect 24568 50661 24579 50725
rect 24493 50645 24579 50661
rect 24493 50581 24504 50645
rect 24568 50581 24579 50645
rect 24493 50565 24579 50581
rect 24493 50501 24504 50565
rect 24568 50501 24579 50565
rect 24493 50485 24579 50501
rect 24493 50421 24504 50485
rect 24568 50421 24579 50485
rect 24493 50405 24579 50421
rect 24493 50341 24504 50405
rect 24568 50341 24579 50405
rect 24493 50325 24579 50341
rect 24493 50261 24504 50325
rect 24568 50261 24579 50325
rect 24493 50245 24579 50261
rect 24493 50181 24504 50245
rect 24568 50181 24579 50245
rect 24493 50161 24579 50181
rect 25581 50725 25667 50745
rect 25581 50661 25592 50725
rect 25656 50661 25667 50725
rect 25581 50645 25667 50661
rect 25581 50581 25592 50645
rect 25656 50581 25667 50645
rect 25581 50565 25667 50581
rect 25581 50501 25592 50565
rect 25656 50501 25667 50565
rect 25581 50485 25667 50501
rect 25581 50421 25592 50485
rect 25656 50421 25667 50485
rect 25581 50405 25667 50421
rect 25581 50341 25592 50405
rect 25656 50341 25667 50405
rect 25581 50325 25667 50341
rect 25581 50261 25592 50325
rect 25656 50261 25667 50325
rect 25581 50245 25667 50261
rect 25581 50181 25592 50245
rect 25656 50181 25667 50245
rect 25581 50161 25667 50181
rect 27757 50725 27843 50745
rect 27757 50661 27768 50725
rect 27832 50661 27843 50725
rect 27757 50645 27843 50661
rect 27757 50581 27768 50645
rect 27832 50581 27843 50645
rect 27757 50565 27843 50581
rect 27757 50501 27768 50565
rect 27832 50501 27843 50565
rect 27757 50485 27843 50501
rect 27757 50421 27768 50485
rect 27832 50421 27843 50485
rect 27757 50405 27843 50421
rect 27757 50341 27768 50405
rect 27832 50341 27843 50405
rect 27757 50325 27843 50341
rect 27757 50261 27768 50325
rect 27832 50261 27843 50325
rect 27757 50245 27843 50261
rect 27757 50181 27768 50245
rect 27832 50181 27843 50245
rect 27757 50161 27843 50181
rect 28845 50725 28931 50745
rect 28845 50661 28856 50725
rect 28920 50661 28931 50725
rect 28845 50645 28931 50661
rect 28845 50581 28856 50645
rect 28920 50581 28931 50645
rect 28845 50565 28931 50581
rect 28845 50501 28856 50565
rect 28920 50501 28931 50565
rect 28845 50485 28931 50501
rect 28845 50421 28856 50485
rect 28920 50421 28931 50485
rect 28845 50405 28931 50421
rect 28845 50341 28856 50405
rect 28920 50341 28931 50405
rect 28845 50325 28931 50341
rect 28845 50261 28856 50325
rect 28920 50261 28931 50325
rect 28845 50245 28931 50261
rect 28845 50181 28856 50245
rect 28920 50181 28931 50245
rect 28845 50161 28931 50181
rect 31021 50725 31107 50745
rect 31021 50661 31032 50725
rect 31096 50661 31107 50725
rect 31021 50645 31107 50661
rect 31021 50581 31032 50645
rect 31096 50581 31107 50645
rect 31021 50565 31107 50581
rect 31021 50501 31032 50565
rect 31096 50501 31107 50565
rect 31021 50485 31107 50501
rect 31021 50421 31032 50485
rect 31096 50421 31107 50485
rect 31021 50405 31107 50421
rect 31021 50341 31032 50405
rect 31096 50341 31107 50405
rect 31021 50325 31107 50341
rect 31021 50261 31032 50325
rect 31096 50261 31107 50325
rect 31021 50245 31107 50261
rect 31021 50181 31032 50245
rect 31096 50181 31107 50245
rect 31021 50161 31107 50181
rect 17420 48728 17506 48748
rect 17420 48664 17431 48728
rect 17495 48664 17506 48728
rect 17420 48648 17506 48664
rect 17420 48584 17431 48648
rect 17495 48584 17506 48648
rect 17420 48568 17506 48584
rect 17420 48504 17431 48568
rect 17495 48504 17506 48568
rect 17420 48488 17506 48504
rect 17420 48424 17431 48488
rect 17495 48424 17506 48488
rect 17420 48408 17506 48424
rect 17420 48344 17431 48408
rect 17495 48344 17506 48408
rect 17420 48328 17506 48344
rect 17420 48264 17431 48328
rect 17495 48264 17506 48328
rect 17420 48248 17506 48264
rect 17420 48184 17431 48248
rect 17495 48184 17506 48248
rect 17420 48164 17506 48184
rect 18508 48728 18594 48748
rect 18508 48664 18519 48728
rect 18583 48664 18594 48728
rect 18508 48648 18594 48664
rect 18508 48584 18519 48648
rect 18583 48584 18594 48648
rect 18508 48568 18594 48584
rect 18508 48504 18519 48568
rect 18583 48504 18594 48568
rect 18508 48488 18594 48504
rect 18508 48424 18519 48488
rect 18583 48424 18594 48488
rect 18508 48408 18594 48424
rect 18508 48344 18519 48408
rect 18583 48344 18594 48408
rect 18508 48328 18594 48344
rect 18508 48264 18519 48328
rect 18583 48264 18594 48328
rect 18508 48248 18594 48264
rect 18508 48184 18519 48248
rect 18583 48184 18594 48248
rect 18508 48164 18594 48184
rect 19596 48728 19682 48748
rect 19596 48664 19607 48728
rect 19671 48664 19682 48728
rect 19596 48648 19682 48664
rect 19596 48584 19607 48648
rect 19671 48584 19682 48648
rect 19596 48568 19682 48584
rect 19596 48504 19607 48568
rect 19671 48504 19682 48568
rect 19596 48488 19682 48504
rect 19596 48424 19607 48488
rect 19671 48424 19682 48488
rect 19596 48408 19682 48424
rect 19596 48344 19607 48408
rect 19671 48344 19682 48408
rect 19596 48328 19682 48344
rect 19596 48264 19607 48328
rect 19671 48264 19682 48328
rect 19596 48248 19682 48264
rect 19596 48184 19607 48248
rect 19671 48184 19682 48248
rect 19596 48164 19682 48184
rect 20684 48728 20770 48748
rect 20684 48664 20695 48728
rect 20759 48664 20770 48728
rect 20684 48648 20770 48664
rect 20684 48584 20695 48648
rect 20759 48584 20770 48648
rect 20684 48568 20770 48584
rect 20684 48504 20695 48568
rect 20759 48504 20770 48568
rect 20684 48488 20770 48504
rect 20684 48424 20695 48488
rect 20759 48424 20770 48488
rect 20684 48408 20770 48424
rect 20684 48344 20695 48408
rect 20759 48344 20770 48408
rect 20684 48328 20770 48344
rect 20684 48264 20695 48328
rect 20759 48264 20770 48328
rect 20684 48248 20770 48264
rect 20684 48184 20695 48248
rect 20759 48184 20770 48248
rect 20684 48164 20770 48184
rect 21772 48728 21858 48748
rect 21772 48664 21783 48728
rect 21847 48664 21858 48728
rect 21772 48648 21858 48664
rect 21772 48584 21783 48648
rect 21847 48584 21858 48648
rect 21772 48568 21858 48584
rect 21772 48504 21783 48568
rect 21847 48504 21858 48568
rect 21772 48488 21858 48504
rect 21772 48424 21783 48488
rect 21847 48424 21858 48488
rect 21772 48408 21858 48424
rect 21772 48344 21783 48408
rect 21847 48344 21858 48408
rect 21772 48328 21858 48344
rect 21772 48264 21783 48328
rect 21847 48264 21858 48328
rect 21772 48248 21858 48264
rect 21772 48184 21783 48248
rect 21847 48184 21858 48248
rect 21772 48164 21858 48184
rect 22860 48728 22946 48748
rect 22860 48664 22871 48728
rect 22935 48664 22946 48728
rect 22860 48648 22946 48664
rect 22860 48584 22871 48648
rect 22935 48584 22946 48648
rect 22860 48568 22946 48584
rect 22860 48504 22871 48568
rect 22935 48504 22946 48568
rect 22860 48488 22946 48504
rect 22860 48424 22871 48488
rect 22935 48424 22946 48488
rect 22860 48408 22946 48424
rect 22860 48344 22871 48408
rect 22935 48344 22946 48408
rect 22860 48328 22946 48344
rect 22860 48264 22871 48328
rect 22935 48264 22946 48328
rect 22860 48248 22946 48264
rect 22860 48184 22871 48248
rect 22935 48184 22946 48248
rect 22860 48164 22946 48184
rect 23948 48728 24034 48748
rect 23948 48664 23959 48728
rect 24023 48664 24034 48728
rect 23948 48648 24034 48664
rect 23948 48584 23959 48648
rect 24023 48584 24034 48648
rect 23948 48568 24034 48584
rect 23948 48504 23959 48568
rect 24023 48504 24034 48568
rect 23948 48488 24034 48504
rect 23948 48424 23959 48488
rect 24023 48424 24034 48488
rect 23948 48408 24034 48424
rect 23948 48344 23959 48408
rect 24023 48344 24034 48408
rect 23948 48328 24034 48344
rect 23948 48264 23959 48328
rect 24023 48264 24034 48328
rect 23948 48248 24034 48264
rect 23948 48184 23959 48248
rect 24023 48184 24034 48248
rect 23948 48164 24034 48184
rect 29388 48728 29474 48748
rect 29388 48664 29399 48728
rect 29463 48664 29474 48728
rect 29388 48648 29474 48664
rect 29388 48584 29399 48648
rect 29463 48584 29474 48648
rect 29388 48568 29474 48584
rect 29388 48504 29399 48568
rect 29463 48504 29474 48568
rect 29388 48488 29474 48504
rect 29388 48424 29399 48488
rect 29463 48424 29474 48488
rect 29388 48408 29474 48424
rect 29388 48344 29399 48408
rect 29463 48344 29474 48408
rect 29388 48328 29474 48344
rect 29388 48264 29399 48328
rect 29463 48264 29474 48328
rect 29388 48248 29474 48264
rect 29388 48184 29399 48248
rect 29463 48184 29474 48248
rect 29388 48164 29474 48184
rect 30476 48728 30562 48748
rect 30476 48664 30487 48728
rect 30551 48664 30562 48728
rect 30476 48648 30562 48664
rect 30476 48584 30487 48648
rect 30551 48584 30562 48648
rect 30476 48568 30562 48584
rect 30476 48504 30487 48568
rect 30551 48504 30562 48568
rect 30476 48488 30562 48504
rect 30476 48424 30487 48488
rect 30551 48424 30562 48488
rect 30476 48408 30562 48424
rect 30476 48344 30487 48408
rect 30551 48344 30562 48408
rect 30476 48328 30562 48344
rect 30476 48264 30487 48328
rect 30551 48264 30562 48328
rect 30476 48248 30562 48264
rect 30476 48184 30487 48248
rect 30551 48184 30562 48248
rect 30476 48164 30562 48184
rect 31564 48728 31650 48748
rect 31564 48664 31575 48728
rect 31639 48664 31650 48728
rect 31564 48648 31650 48664
rect 31564 48584 31575 48648
rect 31639 48584 31650 48648
rect 31564 48568 31650 48584
rect 31564 48504 31575 48568
rect 31639 48504 31650 48568
rect 31564 48488 31650 48504
rect 31564 48424 31575 48488
rect 31639 48424 31650 48488
rect 31564 48408 31650 48424
rect 31564 48344 31575 48408
rect 31639 48344 31650 48408
rect 31564 48328 31650 48344
rect 31564 48264 31575 48328
rect 31639 48264 31650 48328
rect 31564 48248 31650 48264
rect 31564 48184 31575 48248
rect 31639 48184 31650 48248
rect 31564 48164 31650 48184
rect 10167 47612 10561 47634
rect -23498 47192 -11361 47256
rect -11297 47192 -6411 47256
rect -6347 47192 -6337 47256
rect -27097 43278 -26980 43318
rect -27097 43214 -27071 43278
rect -27007 43214 -26980 43278
rect -27097 43198 -26980 43214
rect -27097 43134 -27071 43198
rect -27007 43134 -26980 43198
rect -27097 43118 -26980 43134
rect -27097 43054 -27071 43118
rect -27007 43054 -26980 43118
rect -27097 43038 -26980 43054
rect -27097 42974 -27071 43038
rect -27007 42974 -26980 43038
rect -27097 42958 -26980 42974
rect -27097 42894 -27071 42958
rect -27007 42894 -26980 42958
rect -27097 42878 -26980 42894
rect -27097 42814 -27071 42878
rect -27007 42814 -26980 42878
rect -27097 42774 -26980 42814
rect -27092 42137 -26985 42174
rect -27092 42073 -27071 42137
rect -27007 42073 -26985 42137
rect -27092 42057 -26985 42073
rect -27092 41993 -27071 42057
rect -27007 41993 -26985 42057
rect -27092 41977 -26985 41993
rect -27092 41913 -27071 41977
rect -27007 41913 -26985 41977
rect -27092 41897 -26985 41913
rect -27092 41833 -27071 41897
rect -27007 41833 -26985 41897
rect -27092 41817 -26985 41833
rect -27092 41753 -27071 41817
rect -27007 41753 -26985 41817
rect -27092 41737 -26985 41753
rect -27092 41673 -27071 41737
rect -27007 41673 -26985 41737
rect -27092 41657 -26985 41673
rect -27092 41593 -27071 41657
rect -27007 41593 -26985 41657
rect -27092 41577 -26985 41593
rect -27092 41513 -27071 41577
rect -27007 41513 -26985 41577
rect -27092 41497 -26985 41513
rect -27092 41433 -27071 41497
rect -27007 41433 -26985 41497
rect -27092 41417 -26985 41433
rect -27092 41353 -27071 41417
rect -27007 41353 -26985 41417
rect -27092 41337 -26985 41353
rect -27092 41273 -27071 41337
rect -27007 41273 -26985 41337
rect -27092 41257 -26985 41273
rect -27092 41193 -27071 41257
rect -27007 41193 -26985 41257
rect -27092 41177 -26985 41193
rect -27092 41113 -27071 41177
rect -27007 41113 -26985 41177
rect -27092 41097 -26985 41113
rect -27092 41033 -27071 41097
rect -27007 41033 -26985 41097
rect -27092 40997 -26985 41033
rect -27087 40611 -26980 40648
rect -27087 40547 -27066 40611
rect -27002 40547 -26980 40611
rect -27087 40531 -26980 40547
rect -27087 40467 -27066 40531
rect -27002 40467 -26980 40531
rect -27087 40451 -26980 40467
rect -27087 40387 -27066 40451
rect -27002 40387 -26980 40451
rect -27087 40371 -26980 40387
rect -27087 40307 -27066 40371
rect -27002 40307 -26980 40371
rect -27087 40291 -26980 40307
rect -27087 40227 -27066 40291
rect -27002 40227 -26980 40291
rect -27087 40211 -26980 40227
rect -27087 40147 -27066 40211
rect -27002 40147 -26980 40211
rect -27087 40131 -26980 40147
rect -27087 40067 -27066 40131
rect -27002 40067 -26980 40131
rect -27087 40051 -26980 40067
rect -27087 39987 -27066 40051
rect -27002 39987 -26980 40051
rect -27087 39971 -26980 39987
rect -27087 39907 -27066 39971
rect -27002 39907 -26980 39971
rect -27087 39891 -26980 39907
rect -27087 39827 -27066 39891
rect -27002 39827 -26980 39891
rect -27087 39811 -26980 39827
rect -27087 39747 -27066 39811
rect -27002 39747 -26980 39811
rect -27087 39731 -26980 39747
rect -27087 39667 -27066 39731
rect -27002 39667 -26980 39731
rect -27087 39651 -26980 39667
rect -27087 39587 -27066 39651
rect -27002 39587 -26980 39651
rect -27087 39571 -26980 39587
rect -27087 39507 -27066 39571
rect -27002 39507 -26980 39571
rect -27087 39471 -26980 39507
rect -31822 39148 -31738 39171
rect -31822 39084 -31812 39148
rect -31748 39084 -31738 39148
rect -31822 39068 -31738 39084
rect -31822 39004 -31812 39068
rect -31748 39004 -31738 39068
rect -31822 38988 -31738 39004
rect -31822 38924 -31812 38988
rect -31748 38924 -31738 38988
rect -31822 38908 -31738 38924
rect -31822 38844 -31812 38908
rect -31748 38844 -31738 38908
rect -31822 38822 -31738 38844
rect -27092 39108 -26988 39125
rect -27092 39044 -27072 39108
rect -27008 39044 -26988 39108
rect -27092 39028 -26988 39044
rect -27092 38964 -27072 39028
rect -27008 38964 -26988 39028
rect -27092 38948 -26988 38964
rect -27092 38884 -27072 38948
rect -27008 38884 -26988 38948
rect -27092 38868 -26988 38884
rect -27092 38804 -27072 38868
rect -27008 38804 -26988 38868
rect -27092 38788 -26988 38804
rect -27092 38724 -27072 38788
rect -27008 38724 -26988 38788
rect -27092 38708 -26988 38724
rect -27092 38644 -27072 38708
rect -27008 38644 -26988 38708
rect -27092 38628 -26988 38644
rect -31821 38609 -31737 38618
rect -31821 38545 -31811 38609
rect -31747 38545 -31737 38609
rect -31821 38529 -31737 38545
rect -31821 38465 -31811 38529
rect -31747 38465 -31737 38529
rect -31821 38449 -31737 38465
rect -31821 38385 -31811 38449
rect -31747 38385 -31737 38449
rect -27092 38564 -27072 38628
rect -27008 38564 -26988 38628
rect -27092 38548 -26988 38564
rect -27092 38484 -27072 38548
rect -27008 38484 -26988 38548
rect -27092 38468 -26988 38484
rect -31821 38369 -31737 38385
rect -31821 38305 -31811 38369
rect -31747 38305 -31737 38369
rect -29624 38413 -29140 38418
rect -29624 38349 -29614 38413
rect -29550 38349 -29534 38413
rect -29470 38349 -29454 38413
rect -29390 38349 -29374 38413
rect -29310 38349 -29294 38413
rect -29230 38349 -29214 38413
rect -29150 38349 -29140 38413
rect -29624 38344 -29140 38349
rect -27092 38404 -27072 38468
rect -27008 38404 -26988 38468
rect -27092 38388 -26988 38404
rect -31821 38289 -31737 38305
rect -31821 38225 -31811 38289
rect -31747 38225 -31737 38289
rect -27092 38324 -27072 38388
rect -27008 38324 -26988 38388
rect -27092 38308 -26988 38324
rect -27092 38244 -27072 38308
rect -27008 38244 -26988 38308
rect -27092 38227 -26988 38244
rect -31821 38209 -31737 38225
rect -31821 38145 -31811 38209
rect -31747 38145 -31737 38209
rect -31821 38136 -31737 38145
rect -23498 37802 -23434 47192
rect 17965 46725 18051 46745
rect 17965 46661 17976 46725
rect 18040 46661 18051 46725
rect 17965 46645 18051 46661
rect -10497 46569 -10487 46633
rect -10423 46569 -6411 46633
rect -6347 46569 -6335 46633
rect 17965 46581 17976 46645
rect 18040 46581 18051 46645
rect 17965 46565 18051 46581
rect 17965 46501 17976 46565
rect 18040 46501 18051 46565
rect 17965 46485 18051 46501
rect 17965 46421 17976 46485
rect 18040 46421 18051 46485
rect 17965 46405 18051 46421
rect 17965 46341 17976 46405
rect 18040 46341 18051 46405
rect 17965 46325 18051 46341
rect -5934 46238 -5712 46279
rect -13479 43061 -13395 43066
rect -13479 42997 -13469 43061
rect -13405 42997 -9208 43061
rect -9144 42997 -9134 43061
rect -13479 42992 -13395 42997
rect -12703 42398 -12619 42403
rect -12703 42334 -12693 42398
rect -12629 42334 -10069 42398
rect -10005 42334 -9995 42398
rect -12703 42329 -12619 42334
rect -21501 42163 -21386 42190
rect -21501 42099 -21475 42163
rect -21411 42099 -21386 42163
rect -21501 42074 -21386 42099
rect -5934 39917 -5895 46238
rect -5967 39854 -5895 39917
rect -5751 39917 -5712 46238
rect 17965 46261 17976 46325
rect 18040 46261 18051 46325
rect 17965 46245 18051 46261
rect 17965 46181 17976 46245
rect 18040 46181 18051 46245
rect 17965 46161 18051 46181
rect 19053 46725 19139 46745
rect 19053 46661 19064 46725
rect 19128 46661 19139 46725
rect 19053 46645 19139 46661
rect 19053 46581 19064 46645
rect 19128 46581 19139 46645
rect 19053 46565 19139 46581
rect 19053 46501 19064 46565
rect 19128 46501 19139 46565
rect 19053 46485 19139 46501
rect 19053 46421 19064 46485
rect 19128 46421 19139 46485
rect 19053 46405 19139 46421
rect 19053 46341 19064 46405
rect 19128 46341 19139 46405
rect 19053 46325 19139 46341
rect 19053 46261 19064 46325
rect 19128 46261 19139 46325
rect 19053 46245 19139 46261
rect 19053 46181 19064 46245
rect 19128 46181 19139 46245
rect 19053 46161 19139 46181
rect 20141 46725 20227 46745
rect 20141 46661 20152 46725
rect 20216 46661 20227 46725
rect 20141 46645 20227 46661
rect 20141 46581 20152 46645
rect 20216 46581 20227 46645
rect 20141 46565 20227 46581
rect 20141 46501 20152 46565
rect 20216 46501 20227 46565
rect 20141 46485 20227 46501
rect 20141 46421 20152 46485
rect 20216 46421 20227 46485
rect 20141 46405 20227 46421
rect 20141 46341 20152 46405
rect 20216 46341 20227 46405
rect 20141 46325 20227 46341
rect 20141 46261 20152 46325
rect 20216 46261 20227 46325
rect 20141 46245 20227 46261
rect 20141 46181 20152 46245
rect 20216 46181 20227 46245
rect 20141 46161 20227 46181
rect 21229 46725 21315 46745
rect 21229 46661 21240 46725
rect 21304 46661 21315 46725
rect 21229 46645 21315 46661
rect 21229 46581 21240 46645
rect 21304 46581 21315 46645
rect 21229 46565 21315 46581
rect 21229 46501 21240 46565
rect 21304 46501 21315 46565
rect 21229 46485 21315 46501
rect 21229 46421 21240 46485
rect 21304 46421 21315 46485
rect 21229 46405 21315 46421
rect 21229 46341 21240 46405
rect 21304 46341 21315 46405
rect 21229 46325 21315 46341
rect 21229 46261 21240 46325
rect 21304 46261 21315 46325
rect 21229 46245 21315 46261
rect 21229 46181 21240 46245
rect 21304 46181 21315 46245
rect 21229 46161 21315 46181
rect 22317 46725 22403 46745
rect 22317 46661 22328 46725
rect 22392 46661 22403 46725
rect 22317 46645 22403 46661
rect 22317 46581 22328 46645
rect 22392 46581 22403 46645
rect 22317 46565 22403 46581
rect 22317 46501 22328 46565
rect 22392 46501 22403 46565
rect 22317 46485 22403 46501
rect 22317 46421 22328 46485
rect 22392 46421 22403 46485
rect 22317 46405 22403 46421
rect 22317 46341 22328 46405
rect 22392 46341 22403 46405
rect 22317 46325 22403 46341
rect 22317 46261 22328 46325
rect 22392 46261 22403 46325
rect 22317 46245 22403 46261
rect 22317 46181 22328 46245
rect 22392 46181 22403 46245
rect 22317 46161 22403 46181
rect 24493 46725 24579 46745
rect 24493 46661 24504 46725
rect 24568 46661 24579 46725
rect 24493 46645 24579 46661
rect 24493 46581 24504 46645
rect 24568 46581 24579 46645
rect 24493 46565 24579 46581
rect 24493 46501 24504 46565
rect 24568 46501 24579 46565
rect 24493 46485 24579 46501
rect 24493 46421 24504 46485
rect 24568 46421 24579 46485
rect 24493 46405 24579 46421
rect 24493 46341 24504 46405
rect 24568 46341 24579 46405
rect 24493 46325 24579 46341
rect 24493 46261 24504 46325
rect 24568 46261 24579 46325
rect 24493 46245 24579 46261
rect 24493 46181 24504 46245
rect 24568 46181 24579 46245
rect 24493 46161 24579 46181
rect 25581 46725 25667 46745
rect 25581 46661 25592 46725
rect 25656 46661 25667 46725
rect 25581 46645 25667 46661
rect 25581 46581 25592 46645
rect 25656 46581 25667 46645
rect 25581 46565 25667 46581
rect 25581 46501 25592 46565
rect 25656 46501 25667 46565
rect 25581 46485 25667 46501
rect 25581 46421 25592 46485
rect 25656 46421 25667 46485
rect 25581 46405 25667 46421
rect 25581 46341 25592 46405
rect 25656 46341 25667 46405
rect 25581 46325 25667 46341
rect 25581 46261 25592 46325
rect 25656 46261 25667 46325
rect 25581 46245 25667 46261
rect 25581 46181 25592 46245
rect 25656 46181 25667 46245
rect 25581 46161 25667 46181
rect 26669 46725 26755 46745
rect 26669 46661 26680 46725
rect 26744 46661 26755 46725
rect 26669 46645 26755 46661
rect 26669 46581 26680 46645
rect 26744 46581 26755 46645
rect 26669 46565 26755 46581
rect 26669 46501 26680 46565
rect 26744 46501 26755 46565
rect 26669 46485 26755 46501
rect 26669 46421 26680 46485
rect 26744 46421 26755 46485
rect 26669 46405 26755 46421
rect 26669 46341 26680 46405
rect 26744 46341 26755 46405
rect 26669 46325 26755 46341
rect 26669 46261 26680 46325
rect 26744 46261 26755 46325
rect 26669 46245 26755 46261
rect 26669 46181 26680 46245
rect 26744 46181 26755 46245
rect 26669 46161 26755 46181
rect 27757 46725 27843 46745
rect 27757 46661 27768 46725
rect 27832 46661 27843 46725
rect 27757 46645 27843 46661
rect 27757 46581 27768 46645
rect 27832 46581 27843 46645
rect 27757 46565 27843 46581
rect 27757 46501 27768 46565
rect 27832 46501 27843 46565
rect 27757 46485 27843 46501
rect 27757 46421 27768 46485
rect 27832 46421 27843 46485
rect 27757 46405 27843 46421
rect 27757 46341 27768 46405
rect 27832 46341 27843 46405
rect 27757 46325 27843 46341
rect 27757 46261 27768 46325
rect 27832 46261 27843 46325
rect 27757 46245 27843 46261
rect 27757 46181 27768 46245
rect 27832 46181 27843 46245
rect 27757 46161 27843 46181
rect 28845 46725 28931 46745
rect 28845 46661 28856 46725
rect 28920 46661 28931 46725
rect 28845 46645 28931 46661
rect 28845 46581 28856 46645
rect 28920 46581 28931 46645
rect 28845 46565 28931 46581
rect 28845 46501 28856 46565
rect 28920 46501 28931 46565
rect 28845 46485 28931 46501
rect 28845 46421 28856 46485
rect 28920 46421 28931 46485
rect 28845 46405 28931 46421
rect 28845 46341 28856 46405
rect 28920 46341 28931 46405
rect 28845 46325 28931 46341
rect 28845 46261 28856 46325
rect 28920 46261 28931 46325
rect 28845 46245 28931 46261
rect 28845 46181 28856 46245
rect 28920 46181 28931 46245
rect 28845 46161 28931 46181
rect 29933 46725 30019 46745
rect 29933 46661 29944 46725
rect 30008 46661 30019 46725
rect 29933 46645 30019 46661
rect 29933 46581 29944 46645
rect 30008 46581 30019 46645
rect 29933 46565 30019 46581
rect 29933 46501 29944 46565
rect 30008 46501 30019 46565
rect 29933 46485 30019 46501
rect 29933 46421 29944 46485
rect 30008 46421 30019 46485
rect 29933 46405 30019 46421
rect 29933 46341 29944 46405
rect 30008 46341 30019 46405
rect 29933 46325 30019 46341
rect 29933 46261 29944 46325
rect 30008 46261 30019 46325
rect 29933 46245 30019 46261
rect 29933 46181 29944 46245
rect 30008 46181 30019 46245
rect 29933 46161 30019 46181
rect 31021 46725 31107 46745
rect 31021 46661 31032 46725
rect 31096 46661 31107 46725
rect 31021 46645 31107 46661
rect 31021 46581 31032 46645
rect 31096 46581 31107 46645
rect 31021 46565 31107 46581
rect 31021 46501 31032 46565
rect 31096 46501 31107 46565
rect 31021 46485 31107 46501
rect 31021 46421 31032 46485
rect 31096 46421 31107 46485
rect 52756 46464 52992 55101
rect 31021 46405 31107 46421
rect 31021 46341 31032 46405
rect 31096 46341 31107 46405
rect 31021 46325 31107 46341
rect 31021 46261 31032 46325
rect 31096 46261 31107 46325
rect 40579 46375 40663 46380
rect 47769 46375 52992 46464
rect 40579 46371 52992 46375
rect 40579 46315 40593 46371
rect 40649 46315 52992 46371
rect 40579 46311 52992 46315
rect 40579 46306 40663 46311
rect 31021 46245 31107 46261
rect 31021 46181 31032 46245
rect 31096 46181 31107 46245
rect 47769 46228 52992 46311
rect 55186 50886 62907 51122
rect 31021 46161 31107 46181
rect 10170 46109 10561 46133
rect 334 45833 568 45849
rect 334 44329 379 45833
rect 523 44329 568 45833
rect 334 44313 568 44329
rect 342 41371 522 41388
rect -5751 39854 -5651 39917
rect -5967 39851 -5651 39854
rect 342 39867 360 41371
rect 504 39867 522 41371
rect -5967 39828 -138 39851
rect 342 39850 522 39867
rect 10170 39885 10213 46109
rect 10517 39885 10561 46109
rect 55186 45902 55422 50886
rect 41136 45819 41220 45824
rect 47769 45819 55422 45902
rect 41136 45815 55422 45819
rect 18221 45748 18339 45774
rect 18221 45684 18245 45748
rect 18309 45684 18339 45748
rect 18221 45659 18339 45684
rect 18766 45748 18884 45773
rect 18766 45684 18791 45748
rect 18855 45684 18884 45748
rect 18766 45658 18884 45684
rect 19308 45739 19426 45769
rect 19308 45675 19337 45739
rect 19401 45675 19426 45739
rect 19308 45654 19426 45675
rect 19856 45738 19974 45767
rect 19856 45674 19882 45738
rect 19946 45674 19974 45738
rect 19856 45652 19974 45674
rect 21486 45726 21598 45751
rect 21486 45662 21513 45726
rect 21577 45662 21598 45726
rect 21486 45637 21598 45662
rect 22033 45723 22142 45742
rect 22033 45659 22056 45723
rect 22120 45659 22142 45723
rect 22033 45637 22142 45659
rect 22575 45722 22696 45745
rect 22575 45658 22598 45722
rect 22662 45658 22696 45722
rect 22575 45633 22696 45658
rect 23114 45727 23237 45750
rect 23114 45663 23145 45727
rect 23209 45663 23237 45727
rect 23114 45634 23237 45663
rect 25837 45738 25955 45766
rect 25837 45674 25863 45738
rect 25927 45674 25955 45738
rect 25837 45651 25955 45674
rect 26381 45742 26499 45766
rect 26381 45678 26406 45742
rect 26470 45678 26499 45742
rect 26381 45651 26499 45678
rect 26920 45736 27038 45764
rect 26920 45672 26948 45736
rect 27012 45672 27038 45736
rect 26920 45649 27038 45672
rect 27479 45727 27597 45753
rect 27479 45663 27505 45727
rect 27569 45663 27597 45727
rect 27479 45638 27597 45663
rect 29103 45738 29221 45765
rect 29103 45674 29129 45738
rect 29193 45674 29221 45738
rect 29103 45650 29221 45674
rect 29645 45731 29763 45756
rect 29645 45667 29673 45731
rect 29737 45667 29763 45731
rect 29645 45641 29763 45667
rect 30198 45735 30316 45760
rect 30198 45671 30223 45735
rect 30287 45671 30316 45735
rect 30198 45645 30316 45671
rect 30728 45735 30846 45762
rect 41136 45759 41150 45815
rect 41206 45759 55422 45815
rect 41136 45755 55422 45759
rect 41136 45750 41220 45755
rect 30728 45671 30756 45735
rect 30820 45671 30846 45735
rect 30728 45647 30846 45671
rect 47769 45666 55422 45755
rect 57721 47147 62907 47383
rect 44744 45072 45316 45079
rect 18762 45008 18791 45072
rect 18855 45008 39775 45072
rect 39711 44991 39775 45008
rect 44744 45008 44758 45072
rect 44822 45008 44838 45072
rect 44902 45008 44918 45072
rect 44982 45008 44998 45072
rect 45062 45008 45078 45072
rect 45142 45008 45158 45072
rect 45222 45008 45238 45072
rect 45302 45008 45316 45072
rect 44744 45002 45316 45008
rect 40978 44991 41062 44996
rect 39711 44987 41062 44991
rect 39711 44931 40992 44987
rect 41048 44931 41062 44987
rect 39711 44927 41062 44931
rect 40978 44922 41062 44927
rect 46284 44939 46540 44944
rect 57721 44939 57957 47147
rect 46284 44929 57957 44939
rect 39547 44891 39631 44896
rect 25844 44827 25863 44891
rect 25927 44887 39631 44891
rect 25927 44831 39561 44887
rect 39617 44831 39631 44887
rect 25927 44827 39631 44831
rect 39547 44822 39631 44827
rect 46284 44713 46304 44929
rect 46520 44713 57957 44929
rect 39547 44701 39631 44706
rect 18231 44637 18245 44701
rect 18309 44697 39631 44701
rect 46284 44703 57957 44713
rect 46284 44698 46540 44703
rect 18309 44641 39561 44697
rect 39617 44641 39631 44697
rect 18309 44637 39631 44641
rect 39547 44632 39631 44637
rect 40878 44607 40962 44612
rect 39711 44603 40962 44607
rect 39711 44547 40892 44603
rect 40948 44547 40962 44603
rect 39711 44543 40962 44547
rect 39711 44526 39775 44543
rect 40878 44538 40962 44543
rect 26392 44462 26406 44526
rect 26470 44462 39775 44526
rect 41506 44526 41884 44532
rect 41506 44462 41543 44526
rect 41607 44462 41623 44526
rect 41687 44462 41703 44526
rect 41767 44462 41783 44526
rect 41847 44462 41884 44526
rect 41506 44457 41884 44462
rect 22587 43858 22597 43922
rect 22661 43858 39775 43922
rect 39711 43841 39775 43858
rect 44756 43921 45303 43930
rect 44756 43857 44797 43921
rect 44861 43857 44877 43921
rect 44941 43857 44957 43921
rect 45021 43857 45037 43921
rect 45101 43857 45117 43921
rect 45181 43857 45197 43921
rect 45261 43857 45303 43921
rect 44756 43849 45303 43857
rect 40978 43841 41062 43846
rect 39711 43837 41062 43841
rect 39711 43781 40992 43837
rect 41048 43781 41062 43837
rect 39711 43777 41062 43781
rect 40978 43772 41062 43777
rect 46272 43788 46528 43793
rect 46272 43778 62907 43788
rect 39547 43741 39631 43746
rect 30746 43677 30756 43741
rect 30820 43737 39631 43741
rect 30820 43681 39561 43737
rect 39617 43681 39631 43737
rect 30820 43677 39631 43681
rect 39547 43672 39631 43677
rect 46272 43562 46292 43778
rect 46508 43562 62907 43778
rect 39547 43551 39631 43556
rect 23135 43487 23145 43551
rect 23209 43547 39631 43551
rect 46272 43552 62907 43562
rect 46272 43547 46528 43552
rect 23209 43491 39561 43547
rect 39617 43491 39631 43547
rect 23209 43487 39631 43491
rect 39547 43482 39631 43487
rect 40878 43457 40962 43462
rect 39711 43453 40962 43457
rect 39711 43397 40892 43453
rect 40948 43397 40962 43453
rect 39711 43393 40962 43397
rect 39711 43376 39775 43393
rect 40878 43388 40962 43393
rect 30214 43375 39775 43376
rect 30212 43311 30222 43375
rect 30286 43312 39775 43375
rect 41504 43376 41882 43382
rect 41504 43312 41541 43376
rect 41605 43312 41621 43376
rect 41685 43312 41701 43376
rect 41765 43312 41781 43376
rect 41845 43312 41882 43376
rect 30286 43311 30296 43312
rect 41504 43307 41882 43312
rect 40579 42685 40663 42690
rect 47760 42685 57965 42777
rect 40579 42681 57965 42685
rect 40579 42625 40593 42681
rect 40649 42625 57965 42681
rect 40579 42621 57965 42625
rect 40579 42616 40663 42621
rect 47760 42541 57965 42621
rect 41136 42129 41220 42134
rect 47751 42129 55382 42223
rect 41136 42125 55382 42129
rect 41136 42069 41150 42125
rect 41206 42069 55382 42125
rect 41136 42065 55382 42069
rect 41136 42060 41220 42065
rect 47751 41987 55382 42065
rect 19872 41318 19882 41382
rect 19946 41318 39775 41382
rect 39711 41301 39775 41318
rect 44746 41379 45293 41388
rect 44746 41315 44787 41379
rect 44851 41315 44867 41379
rect 44931 41315 44947 41379
rect 45011 41315 45027 41379
rect 45091 41315 45107 41379
rect 45171 41315 45187 41379
rect 45251 41315 45293 41379
rect 44746 41307 45293 41315
rect 40978 41301 41062 41306
rect 39711 41297 41062 41301
rect 39711 41241 40992 41297
rect 41048 41241 41062 41297
rect 39711 41237 41062 41241
rect 40978 41232 41062 41237
rect 46130 41256 46386 41261
rect 46130 41246 53037 41256
rect 39547 41201 39631 41206
rect 26938 41137 26948 41201
rect 27012 41197 39631 41201
rect 27012 41141 39561 41197
rect 39617 41141 39631 41197
rect 27012 41137 39631 41141
rect 39547 41132 39631 41137
rect 46130 41030 46150 41246
rect 46366 41030 53037 41246
rect 46130 41020 53037 41030
rect 39547 41011 39631 41016
rect 46130 41015 46386 41020
rect 19305 40947 19337 41011
rect 19401 41007 39631 41011
rect 19401 40951 39561 41007
rect 39617 40951 39631 41007
rect 19401 40947 39631 40951
rect 39547 40942 39631 40947
rect 40878 40917 40962 40922
rect 39711 40913 40962 40917
rect 39711 40857 40892 40913
rect 40948 40857 40962 40913
rect 39711 40853 40962 40857
rect 39711 40836 39775 40853
rect 40878 40848 40962 40853
rect 27490 40772 27505 40836
rect 27569 40772 39775 40836
rect 41422 40835 41800 40841
rect 41422 40771 41459 40835
rect 41523 40771 41539 40835
rect 41603 40771 41619 40835
rect 41683 40771 41699 40835
rect 41763 40771 41800 40835
rect 41422 40766 41800 40771
rect 21503 40048 21513 40112
rect 21577 40048 39775 40112
rect 39711 40031 39775 40048
rect 44746 40109 45293 40118
rect 44746 40045 44787 40109
rect 44851 40045 44867 40109
rect 44931 40045 44947 40109
rect 45011 40045 45027 40109
rect 45091 40045 45107 40109
rect 45171 40045 45187 40109
rect 45251 40045 45293 40109
rect 44746 40037 45293 40045
rect 40978 40031 41062 40036
rect 39711 40027 41062 40031
rect 39711 39971 40992 40027
rect 41048 39971 41062 40027
rect 39711 39967 41062 39971
rect 40978 39962 41062 39967
rect 46101 39966 46357 39971
rect 46101 39956 50842 39966
rect 39547 39931 39631 39936
rect 10170 39862 10561 39885
rect 29663 39867 29673 39931
rect 29737 39927 39631 39931
rect 29737 39871 39561 39927
rect 39617 39871 39631 39927
rect 29737 39867 39631 39871
rect 39547 39862 39631 39867
rect -5967 39684 -5668 39828
rect -164 39684 -138 39828
rect 39547 39741 39631 39746
rect -5967 39661 -138 39684
rect 22047 39677 22057 39741
rect 22121 39737 39631 39741
rect 22121 39681 39561 39737
rect 39617 39681 39631 39737
rect 46101 39740 46121 39956
rect 46337 39740 50842 39956
rect 46101 39730 50842 39740
rect 46101 39725 46357 39730
rect 22121 39677 39631 39681
rect 39547 39672 39631 39677
rect -5967 39650 -5651 39661
rect 40878 39647 40962 39652
rect 39711 39643 40962 39647
rect 39711 39587 40892 39643
rect 40948 39587 40962 39643
rect 39711 39583 40962 39587
rect 39711 39566 39775 39583
rect 40878 39578 40962 39583
rect -18893 39502 -18797 39542
rect 29119 39502 29129 39566
rect 29193 39502 39775 39566
rect 41420 39566 41798 39572
rect 41420 39502 41457 39566
rect 41521 39502 41537 39566
rect 41601 39502 41617 39566
rect 41681 39502 41697 39566
rect 41761 39502 41798 39566
rect -18893 39438 -18877 39502
rect -18813 39438 -18797 39502
rect 41420 39497 41798 39502
rect -18893 39422 -18797 39438
rect -18893 39358 -18877 39422
rect -18813 39358 -18797 39422
rect -18893 39342 -18797 39358
rect -18893 39278 -18877 39342
rect -18813 39278 -18797 39342
rect -18893 39262 -18797 39278
rect -18893 39198 -18877 39262
rect -18813 39198 -18797 39262
rect -18893 39182 -18797 39198
rect -18893 39118 -18877 39182
rect -18813 39118 -18797 39182
rect -18893 39102 -18797 39118
rect -18893 39038 -18877 39102
rect -18813 39038 -18797 39102
rect -18893 39022 -18797 39038
rect -18893 38958 -18877 39022
rect -18813 38958 -18797 39022
rect -18893 38942 -18797 38958
rect -18893 38878 -18877 38942
rect -18813 38878 -18797 38942
rect 1473 38883 1537 38887
rect -18893 38862 -18797 38878
rect -18893 38798 -18877 38862
rect -18813 38798 -18797 38862
rect 1463 38874 1547 38883
rect 1463 38818 1477 38874
rect 1533 38818 1547 38874
rect 1463 38809 1547 38818
rect 2503 38873 2605 38886
rect 2503 38809 2522 38873
rect 2586 38809 2605 38873
rect -18893 38782 -18797 38798
rect -18893 38718 -18877 38782
rect -18813 38718 -18797 38782
rect -11723 38726 -11713 38790
rect -11649 38726 -4713 38790
rect -4649 38726 -4639 38790
rect -18893 38702 -18797 38718
rect -18893 38638 -18877 38702
rect -18813 38638 -18797 38702
rect -18893 38622 -18797 38638
rect -18893 38558 -18877 38622
rect -18813 38558 -18797 38622
rect -18893 38542 -18797 38558
rect -18893 38478 -18877 38542
rect -18813 38478 -18797 38542
rect -18893 38462 -18797 38478
rect -18893 38398 -18877 38462
rect -18813 38398 -18797 38462
rect -18893 38382 -18797 38398
rect -18893 38318 -18877 38382
rect -18813 38318 -18797 38382
rect -18893 38302 -18797 38318
rect -18893 38238 -18877 38302
rect -18813 38238 -18797 38302
rect -18893 38222 -18797 38238
rect -18893 38158 -18877 38222
rect -18813 38158 -18797 38222
rect -18893 38142 -18797 38158
rect -18893 38078 -18877 38142
rect -18813 38078 -18797 38142
rect -18893 38062 -18797 38078
rect -18893 37998 -18877 38062
rect -18813 37998 -18797 38062
rect -18893 37982 -18797 37998
rect -18893 37918 -18877 37982
rect -18813 37918 -18797 37982
rect -18893 37902 -18797 37918
rect -18893 37838 -18877 37902
rect -18813 37838 -18797 37902
rect -18893 37822 -18797 37838
rect -18893 37758 -18877 37822
rect -18813 37758 -18797 37822
rect -18893 37742 -18797 37758
rect -18893 37678 -18877 37742
rect -18813 37678 -18797 37742
rect -18893 37662 -18797 37678
rect -18893 37598 -18877 37662
rect -18813 37598 -18797 37662
rect -18893 37582 -18797 37598
rect -16012 38181 -15860 38546
rect -10912 38383 -10905 38447
rect -10841 38383 -4123 38447
rect -4059 38383 -4049 38447
rect -15226 38281 -14722 38299
rect -15226 38181 -15206 38281
rect -16012 37899 -15206 38181
rect -16012 37597 -15860 37899
rect -15226 37817 -15206 37899
rect -14742 37817 -14722 38281
rect 1473 37899 1537 38809
rect 2503 38793 2605 38809
rect 2503 38729 2522 38793
rect 2586 38729 2605 38793
rect 2503 38713 2605 38729
rect 2503 38649 2522 38713
rect 2586 38649 2605 38713
rect 2503 38637 2605 38649
rect 2505 38400 2624 38425
rect 2505 38336 2532 38400
rect 2596 38336 2624 38400
rect 13821 38372 13831 38436
rect 13895 38372 18245 38436
rect 18309 38372 18319 38436
rect 25853 38354 25863 38418
rect 25927 38354 32414 38418
rect 32478 38354 32488 38418
rect 2505 38320 2624 38336
rect 2505 38256 2532 38320
rect 2596 38256 2624 38320
rect 2505 38240 2624 38256
rect 2505 38176 2532 38240
rect 2596 38176 2624 38240
rect 2505 38160 2624 38176
rect 2505 38096 2532 38160
rect 2596 38096 2624 38160
rect 1996 38074 2060 38083
rect 2505 38080 2624 38096
rect 1986 38065 2070 38074
rect 1986 38009 2000 38065
rect 2056 38009 2070 38065
rect 1986 38000 2070 38009
rect 2505 38016 2532 38080
rect 2596 38016 2624 38080
rect -7732 37835 -7722 37899
rect -7658 37835 -2398 37899
rect -2334 37835 -760 37899
rect -696 37835 -686 37899
rect 1463 37835 1473 37899
rect 1537 37835 1547 37899
rect -15226 37799 -14722 37817
rect -35528 37569 -35272 37573
rect -57094 37558 -35272 37569
rect -57094 37342 -35508 37558
rect -35292 37342 -35272 37558
rect -18893 37518 -18877 37582
rect -18813 37518 -18797 37582
rect -18893 37502 -18797 37518
rect -18893 37438 -18877 37502
rect -18813 37438 -18797 37502
rect -18893 37422 -18797 37438
rect -18893 37358 -18877 37422
rect -18813 37358 -18797 37422
rect -57094 37333 -35272 37342
rect -35528 37327 -35272 37333
rect -27089 37341 -26985 37358
rect -29662 37323 -29133 37328
rect -29662 37259 -29630 37323
rect -29566 37259 -29550 37323
rect -29486 37259 -29470 37323
rect -29406 37259 -29390 37323
rect -29326 37259 -29310 37323
rect -29246 37259 -29230 37323
rect -29166 37259 -29133 37323
rect -29662 37254 -29133 37259
rect -27089 37277 -27069 37341
rect -27005 37277 -26985 37341
rect -27089 37261 -26985 37277
rect -27089 37197 -27069 37261
rect -27005 37197 -26985 37261
rect -27089 37181 -26985 37197
rect -27089 37117 -27069 37181
rect -27005 37117 -26985 37181
rect -27089 37101 -26985 37117
rect -27089 37037 -27069 37101
rect -27005 37037 -26985 37101
rect -27089 37021 -26985 37037
rect -27089 36957 -27069 37021
rect -27005 36957 -26985 37021
rect -27089 36941 -26985 36957
rect -27089 36877 -27069 36941
rect -27005 36877 -26985 36941
rect -27089 36861 -26985 36877
rect -27089 36797 -27069 36861
rect -27005 36797 -26985 36861
rect -27089 36781 -26985 36797
rect -27089 36717 -27069 36781
rect -27005 36717 -26985 36781
rect -27089 36701 -26985 36717
rect -27089 36637 -27069 36701
rect -27005 36637 -26985 36701
rect -27089 36621 -26985 36637
rect -27089 36557 -27069 36621
rect -27005 36557 -26985 36621
rect -27089 36541 -26985 36557
rect -27089 36477 -27069 36541
rect -27005 36477 -26985 36541
rect -27089 36460 -26985 36477
rect -18893 37342 -18797 37358
rect -18893 37278 -18877 37342
rect -18813 37278 -18797 37342
rect -8490 37307 -8480 37371
rect -8416 37307 -2815 37371
rect -2751 37370 -729 37371
rect -2751 37307 -760 37370
rect -770 37306 -760 37307
rect -696 37306 -686 37370
rect -18893 37262 -18797 37278
rect -18893 37198 -18877 37262
rect -18813 37198 -18797 37262
rect -18893 37182 -18797 37198
rect -18893 37118 -18877 37182
rect -18813 37118 -18797 37182
rect 1473 37134 1537 37835
rect 1996 37370 2060 38000
rect 2505 37991 2624 38016
rect 14576 37797 14586 37861
rect 14650 37797 18791 37861
rect 18855 37797 18865 37861
rect 26396 37774 26406 37838
rect 26470 37774 31824 37838
rect 31888 37774 31898 37838
rect 1986 37306 1996 37370
rect 2060 37306 2070 37370
rect -18893 37102 -18797 37118
rect -18893 37038 -18877 37102
rect -18813 37038 -18797 37102
rect 1463 37125 1547 37134
rect 1463 37069 1477 37125
rect 1533 37069 1547 37125
rect 1463 37060 1547 37069
rect -18893 37022 -18797 37038
rect -18893 36958 -18877 37022
rect -18813 36958 -18797 37022
rect -18893 36942 -18797 36958
rect -18893 36878 -18877 36942
rect -18813 36878 -18797 36942
rect -18893 36862 -18797 36878
rect -18893 36798 -18877 36862
rect -18813 36798 -18797 36862
rect -18893 36782 -18797 36798
rect -18893 36718 -18877 36782
rect -18813 36718 -18797 36782
rect -18893 36702 -18797 36718
rect -18893 36638 -18877 36702
rect -18813 36638 -18797 36702
rect -18893 36622 -18797 36638
rect -18893 36558 -18877 36622
rect -18813 36558 -18797 36622
rect -18893 36542 -18797 36558
rect -18893 36478 -18877 36542
rect -18813 36478 -18797 36542
rect -18893 36462 -18797 36478
rect -18893 36398 -18877 36462
rect -18813 36398 -18797 36462
rect -18893 36382 -18797 36398
rect -18893 36318 -18877 36382
rect -18813 36318 -18797 36382
rect 1996 36324 2060 37306
rect 15220 37246 15230 37310
rect 15294 37246 19337 37310
rect 19401 37246 19411 37310
rect 30746 37165 30756 37229
rect 30820 37165 31231 37229
rect 31295 37165 31305 37229
rect 2158 37135 2242 37154
rect 2158 37071 2168 37135
rect 2232 37071 2242 37135
rect 2158 37055 2242 37071
rect 2158 36991 2168 37055
rect 2232 36991 2242 37055
rect 2158 36975 2242 36991
rect 2158 36911 2168 36975
rect 2232 36911 2242 36975
rect 2158 36893 2242 36911
rect 2159 36651 2243 36673
rect 15980 36664 15990 36728
rect 16054 36664 19882 36728
rect 19946 36664 19956 36728
rect 2159 36587 2169 36651
rect 2233 36587 2243 36651
rect 6335 36597 6419 36602
rect 2159 36571 2243 36587
rect 2159 36507 2169 36571
rect 2233 36507 2243 36571
rect 2159 36491 2243 36507
rect 2159 36427 2169 36491
rect 2233 36427 2243 36491
rect 2159 36411 2243 36427
rect 2159 36347 2169 36411
rect 2233 36347 2243 36411
rect 2159 36331 2243 36347
rect -18893 36302 -18797 36318
rect -18893 36238 -18877 36302
rect -18813 36238 -18797 36302
rect 1986 36315 2070 36324
rect 1986 36259 2000 36315
rect 2056 36259 2070 36315
rect 1986 36250 2070 36259
rect 2159 36267 2169 36331
rect 2233 36267 2243 36331
rect 2159 36245 2243 36267
rect 2461 36593 6419 36597
rect 2461 36537 6349 36593
rect 6405 36537 6419 36593
rect 2461 36533 6419 36537
rect -18893 36222 -18797 36238
rect -27087 36124 -26986 36165
rect -27087 36060 -27069 36124
rect -27005 36060 -26986 36124
rect -18893 36158 -18877 36222
rect -18813 36158 -18797 36222
rect -18893 36119 -18797 36158
rect -27087 36044 -26986 36060
rect -27087 35980 -27069 36044
rect -27005 35980 -26986 36044
rect -27087 35964 -26986 35980
rect -27087 35900 -27069 35964
rect -27005 35900 -26986 35964
rect 2461 35941 2525 36533
rect 6335 36528 6419 36533
rect 30212 36529 30222 36593
rect 30286 36529 30584 36593
rect 30648 36529 30658 36593
rect 6345 36523 6409 36528
rect 6345 36258 6409 36264
rect 6335 36249 6419 36258
rect 6335 36193 6349 36249
rect 6405 36193 6419 36249
rect 6335 36184 6419 36193
rect 3122 36093 3241 36135
rect 3572 36094 3821 36099
rect 2928 36087 3353 36093
rect 2928 36031 2952 36087
rect 3008 36031 3032 36087
rect 3088 36031 3112 36087
rect 3168 36031 3192 36087
rect 3248 36031 3272 36087
rect 3328 36031 3353 36087
rect 2928 36025 3353 36031
rect 3572 36030 3584 36094
rect 3648 36030 3664 36094
rect 3728 36030 3744 36094
rect 3808 36030 3821 36094
rect 3572 36025 3821 36030
rect 5045 36093 5361 36109
rect 5045 36089 5091 36093
rect 5155 36089 5171 36093
rect 5235 36089 5251 36093
rect 5315 36089 5361 36093
rect 5045 36033 5055 36089
rect 5351 36033 5361 36089
rect 5045 36029 5091 36033
rect 5155 36029 5171 36033
rect 5235 36029 5251 36033
rect 5315 36029 5361 36033
rect -27087 35884 -26986 35900
rect -27087 35820 -27069 35884
rect -27005 35820 -26986 35884
rect -9218 35877 -9208 35941
rect -9144 35877 2525 35941
rect -27087 35804 -26986 35820
rect -27087 35740 -27069 35804
rect -27005 35740 -26986 35804
rect -27087 35724 -26986 35740
rect -27087 35660 -27069 35724
rect -27005 35660 -26986 35724
rect 3122 35672 3241 36025
rect 5045 36013 5361 36029
rect 5564 36094 5811 36102
rect 5564 36030 5575 36094
rect 5639 36030 5655 36094
rect 5719 36030 5735 36094
rect 5799 36030 5811 36094
rect 5564 36022 5811 36030
rect -27087 35644 -26986 35660
rect -27087 35580 -27069 35644
rect -27005 35580 -26986 35644
rect -27087 35564 -26986 35580
rect -27087 35500 -27069 35564
rect -27005 35500 -26986 35564
rect 3111 35644 3250 35672
rect 3111 35580 3148 35644
rect 3212 35580 3250 35644
rect 3111 35553 3250 35580
rect -27087 35484 -26986 35500
rect -27087 35420 -27069 35484
rect -27005 35420 -26986 35484
rect -27087 35404 -26986 35420
rect -27087 35340 -27069 35404
rect -27005 35340 -26986 35404
rect 6345 35351 6409 36184
rect 7503 36099 7622 36121
rect 6926 36086 7167 36094
rect 6926 36082 6974 36086
rect 7038 36082 7054 36086
rect 7118 36082 7167 36086
rect 6926 36026 6938 36082
rect 7154 36026 7167 36082
rect 6926 36022 6974 36026
rect 7038 36022 7054 36026
rect 7118 36022 7167 36026
rect 7373 36089 7691 36099
rect 7373 36033 7384 36089
rect 7440 36033 7464 36089
rect 7520 36033 7544 36089
rect 7600 36033 7624 36089
rect 7680 36033 7691 36089
rect 7373 36023 7691 36033
rect 8911 36088 9358 36098
rect 8911 36032 8946 36088
rect 9002 36032 9026 36088
rect 9082 36032 9106 36088
rect 9162 36032 9186 36088
rect 9242 36032 9266 36088
rect 9322 36032 9358 36088
rect 8911 36023 9358 36032
rect 9565 36089 9812 36096
rect 9565 36025 9576 36089
rect 9640 36025 9656 36089
rect 9720 36025 9736 36089
rect 9800 36025 9812 36089
rect 6926 36015 7167 36022
rect 7503 35641 7622 36023
rect 9070 35650 9189 36023
rect 9565 36018 9812 36025
rect 16711 35986 16721 36050
rect 16785 35986 23145 36050
rect 23209 35986 23219 36050
rect 29663 35906 29673 35970
rect 29737 35906 29990 35970
rect 30054 35906 30064 35970
rect 7493 35613 7632 35641
rect 7493 35549 7530 35613
rect 7594 35549 7632 35613
rect 7493 35522 7632 35549
rect 9060 35622 9199 35650
rect 9060 35558 9097 35622
rect 9161 35558 9199 35622
rect 9060 35531 9199 35558
rect -27087 35324 -26986 35340
rect -27087 35260 -27069 35324
rect -27005 35260 -26986 35324
rect -10079 35287 -10069 35351
rect -10005 35287 6409 35351
rect 17402 35279 17412 35343
rect 17476 35279 22598 35343
rect 22662 35279 22672 35343
rect -27087 35244 -26986 35260
rect -27087 35180 -27069 35244
rect -27005 35180 -26986 35244
rect 29119 35194 29129 35258
rect 29193 35194 29407 35258
rect 29471 35194 29481 35258
rect -27087 35164 -26986 35180
rect -27087 35100 -27069 35164
rect -27005 35100 -26986 35164
rect -27087 35084 -26986 35100
rect -27087 35020 -27069 35084
rect -27005 35020 -26986 35084
rect -27087 34980 -26986 35020
rect -27089 34686 -26990 34696
rect -27089 34622 -27072 34686
rect -27008 34622 -26990 34686
rect -9379 34676 -9295 34681
rect -27089 34606 -26990 34622
rect -13405 34612 -13395 34676
rect -13331 34672 -9295 34676
rect -13331 34616 -9365 34672
rect -9309 34616 -9295 34672
rect -13331 34612 -9295 34616
rect -9379 34607 -9295 34612
rect -27089 34542 -27072 34606
rect -27008 34542 -26990 34606
rect -27089 34526 -26990 34542
rect -27089 34462 -27072 34526
rect -27008 34462 -26990 34526
rect 18242 34519 18252 34583
rect 18316 34519 22056 34583
rect 22120 34519 22130 34583
rect -27089 34446 -26990 34462
rect 26938 34458 26948 34522
rect 27012 34458 28828 34522
rect 28892 34458 28902 34522
rect -27089 34382 -27072 34446
rect -27008 34382 -26990 34446
rect -27089 34366 -26990 34382
rect -27089 34302 -27072 34366
rect -27008 34302 -26990 34366
rect -27089 34286 -26990 34302
rect -27089 34222 -27072 34286
rect -27008 34222 -26990 34286
rect -27089 34206 -26990 34222
rect -27089 34142 -27072 34206
rect -27008 34142 -26990 34206
rect 5922 34195 6006 34200
rect -27089 34126 -26990 34142
rect -4723 34131 -4713 34195
rect -4649 34191 6006 34195
rect -4649 34135 5936 34191
rect 5992 34135 6006 34191
rect -4649 34131 6006 34135
rect 5922 34126 6006 34131
rect -27089 34062 -27072 34126
rect -27008 34062 -26990 34126
rect -27089 34046 -26990 34062
rect -27089 33982 -27072 34046
rect -27008 33982 -26990 34046
rect -27089 33966 -26990 33982
rect -27089 33902 -27072 33966
rect -27008 33902 -26990 33966
rect -27089 33886 -26990 33902
rect -27089 33822 -27072 33886
rect -27008 33822 -26990 33886
rect 6728 33850 6812 33855
rect -27089 33806 -26990 33822
rect -27089 33742 -27072 33806
rect -27008 33742 -26990 33806
rect -4133 33786 -4123 33850
rect -4059 33846 6812 33850
rect -4059 33790 6742 33846
rect 6798 33790 6812 33846
rect -4059 33786 6812 33790
rect 6728 33781 6812 33786
rect 27495 33749 27505 33813
rect 27569 33749 28315 33813
rect 28379 33749 28389 33813
rect -27089 33726 -26990 33742
rect -27089 33662 -27072 33726
rect -27008 33662 -26990 33726
rect 19245 33682 19255 33746
rect 19319 33682 21513 33746
rect 21577 33682 21588 33746
rect -27089 33646 -26990 33662
rect -27089 33582 -27072 33646
rect -27008 33582 -26990 33646
rect -27089 33566 -26990 33582
rect -27089 33502 -27072 33566
rect -27008 33502 -26990 33566
rect -27089 33493 -26990 33502
rect -21540 33551 -21434 33575
rect -21540 33487 -21518 33551
rect -21454 33487 -21434 33551
rect -21540 33466 -21434 33487
rect -6958 33179 -6874 33184
rect -15149 33115 -15139 33179
rect -15075 33175 -6874 33179
rect -15075 33119 -6944 33175
rect -6888 33119 -6874 33175
rect -15075 33115 -6874 33119
rect -6958 33110 -6874 33115
rect -27094 32864 -26995 32904
rect -27094 32800 -27077 32864
rect -27013 32800 -26995 32864
rect -27094 32784 -26995 32800
rect -27094 32720 -27077 32784
rect -27013 32720 -26995 32784
rect -27094 32704 -26995 32720
rect -27094 32640 -27077 32704
rect -27013 32640 -26995 32704
rect -27094 32624 -26995 32640
rect -27094 32560 -27077 32624
rect -27013 32560 -26995 32624
rect -27094 32544 -26995 32560
rect -27094 32480 -27077 32544
rect -27013 32480 -26995 32544
rect -27094 32464 -26995 32480
rect -27094 32400 -27077 32464
rect -27013 32400 -26995 32464
rect -27094 32360 -26995 32400
rect 7354 32352 7438 32357
rect 5307 32345 5391 32350
rect 5121 32341 5391 32345
rect 5121 32285 5321 32341
rect 5377 32285 5391 32341
rect 5121 32281 5391 32285
rect 7354 32348 7607 32352
rect 7354 32292 7368 32348
rect 7424 32292 7607 32348
rect 7354 32288 7607 32292
rect 7354 32283 7438 32288
rect 5307 32276 5391 32281
rect 4964 31452 5028 32173
rect 7702 31452 7766 32173
rect 7942 31811 8053 31841
rect 7942 31747 7965 31811
rect 8029 31747 8053 31811
rect 7942 31723 8053 31747
rect 4964 31375 5028 31388
rect 7702 31375 7766 31388
rect 11337 31327 11347 31391
rect 11411 31327 13831 31391
rect 13895 31327 13905 31391
rect 5702 31191 5766 31192
rect 3944 31123 4742 31187
rect 4941 31127 5766 31191
rect 3961 30389 4025 31123
rect 4325 30432 4440 30460
rect 4325 30368 4354 30432
rect 4418 30368 4440 30432
rect 5702 30394 5766 31127
rect 6964 31191 7028 31192
rect 6964 31127 7789 31191
rect 6964 30394 7028 31127
rect 7988 31123 8786 31187
rect 8300 30437 8415 30464
rect 4325 30342 4440 30368
rect 8300 30373 8328 30437
rect 8392 30373 8415 30437
rect 8705 30389 8769 31123
rect 11956 30708 11966 30772
rect 12030 30708 14586 30772
rect 14650 30708 14660 30772
rect 50606 30469 50842 39730
rect 52801 33632 53037 41020
rect 55146 37094 55382 41987
rect 57729 40402 57965 42541
rect 57729 40166 62907 40402
rect 55146 36858 62907 37094
rect 52801 33396 62907 33632
rect 8300 30348 8415 30373
rect 3298 30305 3418 30335
rect 3298 30241 3326 30305
rect 3390 30241 3418 30305
rect 3298 30212 3418 30241
rect 50606 30233 62907 30469
rect -12703 29752 -12619 29757
rect 1903 29752 1987 29757
rect -12703 29748 -3918 29752
rect -12703 29692 -12689 29748
rect -12633 29692 -3918 29748
rect -12703 29688 -3918 29692
rect -3854 29748 1987 29752
rect -3854 29692 1917 29748
rect 1973 29692 1987 29748
rect -3854 29688 1987 29692
rect -12703 29683 -12619 29688
rect 1903 29683 1987 29688
rect 3961 29389 4025 30187
rect 4328 29982 4609 30046
rect -13479 29329 -13395 29334
rect 1903 29329 1987 29334
rect -13479 29325 -5279 29329
rect -13479 29269 -13465 29325
rect -13409 29269 -5279 29325
rect -13479 29265 -5279 29269
rect -5215 29325 1987 29329
rect -5215 29269 1917 29325
rect 1973 29269 1987 29325
rect -5215 29265 1987 29269
rect -13479 29260 -13395 29265
rect 1903 29260 1987 29265
rect 3961 28389 4025 29187
rect 4328 28600 4392 29982
rect 5702 29394 5766 30192
rect 6964 29394 7028 30192
rect 8121 29982 8402 30046
rect 4701 28813 4765 29012
rect 4691 28804 4775 28813
rect 4691 28748 4705 28804
rect 4761 28748 4775 28804
rect 4691 28739 4775 28748
rect 4318 28593 4402 28600
rect 4318 28591 4579 28593
rect 4318 28535 4332 28591
rect 4388 28535 4579 28591
rect 4318 28529 4579 28535
rect 4318 28526 4402 28529
rect 5702 28394 5766 29192
rect 6964 28394 7028 29192
rect 7960 28851 8024 29021
rect 7950 28842 8034 28851
rect 7950 28786 7964 28842
rect 8020 28786 8034 28842
rect 7950 28777 8034 28786
rect 8338 28597 8402 29982
rect 8705 29389 8769 30187
rect 16692 29752 16811 29781
rect 16692 29688 16721 29752
rect 16785 29688 16811 29752
rect 16692 29659 16811 29688
rect 17378 29329 17506 29366
rect 17378 29265 17412 29329
rect 17476 29265 17506 29329
rect 17378 29232 17506 29265
rect 8328 28593 8412 28597
rect 8151 28588 8412 28593
rect 8151 28532 8342 28588
rect 8398 28532 8412 28588
rect 8151 28529 8412 28532
rect 8328 28523 8412 28529
rect 8705 28389 8769 29187
rect 10623 28740 10633 28804
rect 10697 28740 11966 28804
rect 12030 28740 12040 28804
rect -15722 28063 -15603 28103
rect -15722 27999 -15695 28063
rect -15631 27999 -15603 28063
rect -15722 27983 -15603 27999
rect -15722 27919 -15695 27983
rect -15631 27919 -15603 27983
rect -15722 27903 -15603 27919
rect -15722 27839 -15695 27903
rect -15631 27839 -15603 27903
rect -15722 27823 -15603 27839
rect -15722 27759 -15695 27823
rect -15631 27759 -15603 27823
rect -15722 27743 -15603 27759
rect -15722 27679 -15695 27743
rect -15631 27679 -15603 27743
rect -17645 27612 -17497 27649
rect -15722 27640 -15603 27679
rect -12399 28065 -12306 28081
rect -12399 28001 -12385 28065
rect -12321 28001 -12306 28065
rect -12399 27985 -12306 28001
rect -12399 27921 -12385 27985
rect -12321 27921 -12306 27985
rect -12399 27905 -12306 27921
rect -12399 27841 -12385 27905
rect -12321 27841 -12306 27905
rect -12399 27825 -12306 27841
rect -12399 27761 -12385 27825
rect -12321 27761 -12306 27825
rect -12399 27745 -12306 27761
rect -12399 27681 -12385 27745
rect -12321 27681 -12306 27745
rect -12399 27665 -12306 27681
rect -17645 27548 -17603 27612
rect -17539 27548 -17497 27612
rect -17645 27511 -17497 27548
rect -5309 27532 -5186 27565
rect -5309 27468 -5279 27532
rect -5215 27468 -5186 27532
rect -5309 27440 -5186 27468
rect 3961 27451 4025 28187
rect 5702 27451 5766 28192
rect -12404 27424 -12287 27432
rect -12404 27360 -12378 27424
rect -12314 27360 -12287 27424
rect 3961 27389 4764 27451
rect 3966 27387 4764 27389
rect 4966 27394 5766 27451
rect 6964 27451 7028 28192
rect 8705 27451 8769 28187
rect 6964 27394 7764 27451
rect 4966 27387 5764 27394
rect 6966 27387 7764 27394
rect 7966 27389 8769 27451
rect 7966 27387 8764 27389
rect -12404 27344 -12287 27360
rect -12404 27280 -12378 27344
rect -12314 27280 -12287 27344
rect -12404 27264 -12287 27280
rect -12404 27200 -12378 27264
rect -12314 27200 -12287 27264
rect -12404 27193 -12287 27200
rect -3948 26855 -3825 26889
rect -3948 26791 -3918 26855
rect -3854 26791 -3825 26855
rect -3948 26764 -3825 26791
rect -38200 26594 -34846 26616
rect -38200 26530 -38155 26594
rect -38091 26530 -38075 26594
rect -38011 26530 -37995 26594
rect -37931 26530 -37915 26594
rect -37851 26530 -37835 26594
rect -37771 26530 -37755 26594
rect -37691 26530 -37675 26594
rect -37611 26530 -37595 26594
rect -37531 26530 -37515 26594
rect -37451 26530 -37435 26594
rect -37371 26530 -37355 26594
rect -37291 26530 -37275 26594
rect -37211 26530 -37195 26594
rect -37131 26530 -37115 26594
rect -37051 26530 -37035 26594
rect -36971 26530 -36955 26594
rect -36891 26530 -36875 26594
rect -36811 26530 -36795 26594
rect -36731 26530 -36715 26594
rect -36651 26530 -36635 26594
rect -36571 26530 -36555 26594
rect -36491 26530 -36475 26594
rect -36411 26530 -36395 26594
rect -36331 26530 -36315 26594
rect -36251 26530 -36235 26594
rect -36171 26530 -36155 26594
rect -36091 26530 -36075 26594
rect -36011 26530 -35995 26594
rect -35931 26530 -35915 26594
rect -35851 26530 -35835 26594
rect -35771 26530 -35755 26594
rect -35691 26530 -35675 26594
rect -35611 26530 -35595 26594
rect -35531 26530 -35515 26594
rect -35451 26530 -35435 26594
rect -35371 26530 -35355 26594
rect -35291 26530 -35275 26594
rect -35211 26530 -35195 26594
rect -35131 26530 -35115 26594
rect -35051 26530 -35035 26594
rect -34971 26530 -34955 26594
rect -34891 26530 -34846 26594
rect -38200 26509 -34846 26530
rect -12406 26463 -12291 26491
rect -17645 26383 -17497 26420
rect -17645 26319 -17603 26383
rect -17539 26319 -17497 26383
rect -17645 26282 -17497 26319
rect -12406 26399 -12381 26463
rect -12317 26399 -12291 26463
rect 4966 26402 5030 27200
rect 7700 26402 7764 27200
rect -12406 26383 -12291 26399
rect -12406 26319 -12381 26383
rect -12317 26319 -12291 26383
rect -12406 26303 -12291 26319
rect -15735 26274 -15626 26286
rect -15735 26210 -15713 26274
rect -15649 26210 -15626 26274
rect -15735 26194 -15626 26210
rect -15735 26130 -15713 26194
rect -15649 26130 -15626 26194
rect -15735 26114 -15626 26130
rect -15735 26050 -15713 26114
rect -15649 26050 -15626 26114
rect -12406 26239 -12381 26303
rect -12317 26239 -12291 26303
rect 11337 26286 11347 26350
rect 11411 26286 11837 26350
rect 11901 26286 11911 26350
rect -12406 26223 -12291 26239
rect -12406 26159 -12381 26223
rect -12317 26159 -12291 26223
rect -12406 26143 -12291 26159
rect -12406 26079 -12381 26143
rect -12317 26079 -12291 26143
rect -12406 26052 -12291 26079
rect -15735 26039 -15626 26050
rect 19861 26009 19945 26014
rect 13840 25945 13850 26009
rect 13914 26005 25879 26009
rect 13914 25949 19875 26005
rect 19931 25949 25879 26005
rect 13914 25945 25879 25949
rect 25943 25945 25950 26009
rect 19861 25940 19945 25945
rect -12394 25821 -12311 25828
rect -19098 25799 -15505 25804
rect -19098 25575 -19084 25799
rect -18860 25575 -15505 25799
rect -12394 25765 -12381 25821
rect -12325 25765 -12311 25821
rect -12394 25741 -12311 25765
rect -12394 25685 -12381 25741
rect -12325 25685 -12311 25741
rect -13999 25664 -13915 25669
rect -13999 25660 -12544 25664
rect -13999 25604 -13985 25660
rect -13929 25604 -12544 25660
rect -13999 25600 -12544 25604
rect -13999 25595 -13915 25600
rect -19098 25571 -15505 25575
rect -18560 25570 -18327 25571
rect -25459 25480 -25359 25487
rect -25459 25416 -25441 25480
rect -25377 25416 -25359 25480
rect -25459 25400 -25359 25416
rect -25459 25336 -25441 25400
rect -25377 25336 -25359 25400
rect -25459 25320 -25359 25336
rect -25459 25256 -25441 25320
rect -25377 25256 -25359 25320
rect -25459 25240 -25359 25256
rect -25459 25176 -25441 25240
rect -25377 25176 -25359 25240
rect -40603 25171 -40347 25176
rect -57094 25161 -40347 25171
rect -25459 25170 -25359 25176
rect -15738 25420 -15505 25571
rect -15738 25364 -15708 25420
rect -15652 25364 -15505 25420
rect -15738 25340 -15505 25364
rect -12608 25419 -12544 25600
rect -12394 25661 -12311 25685
rect -12394 25605 -12381 25661
rect -12325 25605 -12311 25661
rect -12394 25599 -12311 25605
rect -12177 25600 -11324 25664
rect -11260 25600 -11250 25664
rect -12177 25419 -12113 25600
rect 19863 25598 19947 25603
rect 13256 25534 13266 25598
rect 13330 25594 26463 25598
rect 13330 25538 19877 25594
rect 19933 25538 26463 25594
rect 13330 25534 26463 25538
rect 26527 25534 26537 25598
rect 19863 25529 19947 25534
rect -12608 25355 -12113 25419
rect -15738 25284 -15708 25340
rect -15652 25284 -15505 25340
rect -15738 25260 -15505 25284
rect -15738 25204 -15708 25260
rect -15652 25204 -15505 25260
rect -15738 25180 -15505 25204
rect -57094 24945 -40583 25161
rect -40367 24945 -40347 25161
rect -15738 25124 -15708 25180
rect -15652 25124 -15505 25180
rect -15738 25100 -15505 25124
rect -15738 25044 -15708 25100
rect -15652 25044 -15505 25100
rect -15738 25011 -15505 25044
rect -17645 24970 -17497 25007
rect -57094 24935 -40347 24945
rect -40603 24930 -40347 24935
rect -25462 24941 -25355 24950
rect -25462 24877 -25441 24941
rect -25377 24877 -25355 24941
rect -25462 24861 -25355 24877
rect -17645 24906 -17603 24970
rect -17539 24906 -17497 24970
rect -17645 24869 -17497 24906
rect -14420 24872 -14336 24877
rect -25462 24797 -25441 24861
rect -25377 24797 -25355 24861
rect -14420 24868 -11977 24872
rect -14420 24812 -14406 24868
rect -14350 24812 -11977 24868
rect -14420 24808 -11977 24812
rect -11913 24808 -11903 24872
rect -14420 24803 -14336 24808
rect -25462 24781 -25355 24797
rect 7591 24784 7601 24848
rect 7665 24784 15230 24848
rect 15294 24784 15304 24848
rect -25462 24717 -25441 24781
rect -25377 24717 -25355 24781
rect -25462 24709 -25355 24717
rect -12403 24697 -12318 24717
rect -12403 24633 -12393 24697
rect -12329 24633 -12318 24697
rect -12403 24617 -12318 24633
rect -12403 24553 -12393 24617
rect -12329 24553 -12318 24617
rect -12403 24537 -12318 24553
rect -12403 24473 -12393 24537
rect -12329 24473 -12318 24537
rect -12403 24453 -12318 24473
rect 5705 24582 5793 24599
rect 5705 24518 5717 24582
rect 5781 24518 5793 24582
rect 7058 24592 7142 24597
rect 7256 24592 7266 24593
rect 7058 24588 7266 24592
rect 7058 24532 7072 24588
rect 7128 24532 7266 24588
rect 7058 24529 7266 24532
rect 7330 24529 7340 24593
rect 7058 24528 7290 24529
rect 7058 24523 7142 24528
rect 5705 24502 5793 24518
rect 5705 24438 5717 24502
rect 5781 24438 5793 24502
rect 8119 24466 8129 24530
rect 8193 24466 15990 24530
rect 16054 24466 16064 24530
rect 5705 24422 5793 24438
rect 5705 24358 5717 24422
rect 5781 24358 5793 24422
rect 5705 24342 5793 24358
rect 5705 24278 5717 24342
rect 5781 24278 5793 24342
rect 5705 24262 5793 24278
rect -12408 24233 -12306 24244
rect -12408 24169 -12389 24233
rect -12325 24169 -12306 24233
rect 5705 24198 5717 24262
rect 5781 24198 5793 24262
rect 5705 24181 5793 24198
rect -12408 24153 -12306 24169
rect -12408 24089 -12389 24153
rect -12325 24089 -12306 24153
rect 11073 24138 11080 24202
rect 11144 24138 19929 24202
rect -12408 24073 -12306 24089
rect -12408 24009 -12389 24073
rect -12325 24009 -12306 24073
rect -12408 23998 -12306 24009
rect -11334 23823 -11324 23887
rect -11260 23823 7266 23887
rect 7330 23823 19255 23887
rect 19319 23823 19329 23887
rect -17645 23741 -17497 23778
rect -17645 23677 -17603 23741
rect -17539 23677 -17497 23741
rect -17645 23640 -17497 23677
rect 7081 23648 7165 23657
rect -15735 23633 -15648 23642
rect -38192 23586 -34842 23610
rect -38192 23522 -38149 23586
rect -38085 23522 -38069 23586
rect -38005 23522 -37989 23586
rect -37925 23522 -37909 23586
rect -37845 23522 -37829 23586
rect -37765 23522 -37749 23586
rect -37685 23522 -37669 23586
rect -37605 23522 -37589 23586
rect -37525 23522 -37509 23586
rect -37445 23522 -37429 23586
rect -37365 23522 -37349 23586
rect -37285 23522 -37269 23586
rect -37205 23522 -37189 23586
rect -37125 23522 -37109 23586
rect -37045 23522 -37029 23586
rect -36965 23522 -36949 23586
rect -36885 23522 -36869 23586
rect -36805 23522 -36789 23586
rect -36725 23522 -36709 23586
rect -36645 23522 -36629 23586
rect -36565 23522 -36549 23586
rect -36485 23522 -36469 23586
rect -36405 23522 -36389 23586
rect -36325 23522 -36309 23586
rect -36245 23522 -36229 23586
rect -36165 23522 -36149 23586
rect -36085 23522 -36069 23586
rect -36005 23522 -35989 23586
rect -35925 23522 -35909 23586
rect -35845 23522 -35829 23586
rect -35765 23522 -35749 23586
rect -35685 23522 -35669 23586
rect -35605 23522 -35589 23586
rect -35525 23522 -35509 23586
rect -35445 23522 -35429 23586
rect -35365 23522 -35349 23586
rect -35285 23522 -35269 23586
rect -35205 23522 -35189 23586
rect -35125 23522 -35109 23586
rect -35045 23522 -35029 23586
rect -34965 23522 -34949 23586
rect -34885 23522 -34842 23586
rect -38192 23498 -34842 23522
rect -15735 23569 -15724 23633
rect -15660 23569 -15648 23633
rect 7081 23592 7095 23648
rect 7151 23592 7165 23648
rect 7081 23583 7165 23592
rect -15735 23553 -15648 23569
rect -15735 23489 -15724 23553
rect -15660 23489 -15648 23553
rect 7091 23518 7155 23583
rect -15735 23473 -15648 23489
rect -15735 23409 -15724 23473
rect -15660 23409 -15648 23473
rect -11987 23454 -11977 23518
rect -11913 23454 18252 23518
rect 18316 23454 18326 23518
rect -15735 23400 -15648 23409
rect 8777 23333 8953 23361
rect -12399 23259 -12309 23282
rect -12399 23195 -12386 23259
rect -12322 23195 -12309 23259
rect 8777 23269 8793 23333
rect 8857 23269 8873 23333
rect 8937 23269 8953 23333
rect 8777 23241 8953 23269
rect 19865 23210 19929 24138
rect 42846 24151 46200 24179
rect 42846 24087 42891 24151
rect 42955 24087 42971 24151
rect 43035 24087 43051 24151
rect 43115 24087 43131 24151
rect 43195 24087 43211 24151
rect 43275 24087 43291 24151
rect 43355 24087 43371 24151
rect 43435 24087 43451 24151
rect 43515 24087 43531 24151
rect 43595 24087 43611 24151
rect 43675 24087 43691 24151
rect 43755 24087 43771 24151
rect 43835 24087 43851 24151
rect 43915 24087 43931 24151
rect 43995 24087 44011 24151
rect 44075 24087 44091 24151
rect 44155 24087 44171 24151
rect 44235 24087 44251 24151
rect 44315 24087 44331 24151
rect 44395 24087 44411 24151
rect 44475 24087 44491 24151
rect 44555 24087 44571 24151
rect 44635 24087 44651 24151
rect 44715 24087 44731 24151
rect 44795 24087 44811 24151
rect 44875 24087 44891 24151
rect 44955 24087 44971 24151
rect 45035 24087 45051 24151
rect 45115 24087 45131 24151
rect 45195 24087 45211 24151
rect 45275 24087 45291 24151
rect 45355 24087 45371 24151
rect 45435 24087 45451 24151
rect 45515 24087 45531 24151
rect 45595 24087 45611 24151
rect 45675 24087 45691 24151
rect 45755 24087 45771 24151
rect 45835 24087 45851 24151
rect 45915 24087 45931 24151
rect 45995 24087 46011 24151
rect 46075 24087 46091 24151
rect 46155 24087 46200 24151
rect 42846 24060 46200 24087
rect 36045 24018 36148 24038
rect 36045 23954 36066 24018
rect 36130 23954 36148 24018
rect 36045 23934 36148 23954
rect 35126 23866 35241 23893
rect 35126 23802 35152 23866
rect 35216 23802 35241 23866
rect 35126 23772 35241 23802
rect 39336 23711 39430 23719
rect 39336 23675 39355 23711
rect 39411 23675 39430 23711
rect 37809 23583 37902 23616
rect 37809 23519 37823 23583
rect 37887 23519 37902 23583
rect 37809 23487 37902 23519
rect 39336 23611 39351 23675
rect 39415 23611 39430 23675
rect 39336 23595 39355 23611
rect 39411 23595 39430 23611
rect 39336 23531 39351 23595
rect 39415 23531 39430 23595
rect 39336 23495 39355 23531
rect 39411 23495 39430 23531
rect 39336 23488 39430 23495
rect -12399 23179 -12309 23195
rect -12399 23115 -12386 23179
rect -12322 23115 -12309 23179
rect -12399 23099 -12309 23115
rect -12399 23035 -12386 23099
rect -12322 23035 -12309 23099
rect 4770 23151 5253 23159
rect -12399 23019 -12309 23035
rect -12399 22955 -12386 23019
rect -12322 22955 -12309 23019
rect 2540 23063 2624 23068
rect 4770 23063 4819 23151
rect 2540 23059 4819 23063
rect 2540 23003 2554 23059
rect 2610 23003 4819 23059
rect 2540 22999 4819 23003
rect 2540 22994 2624 22999
rect -12399 22939 -12309 22955
rect -12399 22875 -12386 22939
rect -12322 22875 -12309 22939
rect 4770 22927 4819 22999
rect 5203 23063 5253 23151
rect 12578 23146 12588 23210
rect 12652 23146 27111 23210
rect 27175 23146 27186 23210
rect 37809 23182 37915 23199
rect 37809 23118 37830 23182
rect 37894 23118 37915 23182
rect 37809 23102 37915 23118
rect 10192 23063 10276 23068
rect 5203 22999 5718 23063
rect 5782 23059 10276 23063
rect 5782 23003 10206 23059
rect 10262 23003 10276 23059
rect 5782 22999 10276 23003
rect 5203 22927 5253 22999
rect 10192 22994 10276 22999
rect 37809 23038 37830 23102
rect 37894 23038 37915 23102
rect 37809 23022 37915 23038
rect 4770 22919 5253 22927
rect 11836 22916 11900 22979
rect 37809 22958 37830 23022
rect 37894 22958 37915 23022
rect 37809 22941 37915 22958
rect 39325 23188 39431 23205
rect 39325 23124 39346 23188
rect 39410 23124 39431 23188
rect 39325 23108 39431 23124
rect 39325 23044 39346 23108
rect 39410 23044 39431 23108
rect 39325 23028 39431 23044
rect 39325 22964 39346 23028
rect 39410 22964 39431 23028
rect 39325 22947 39431 22964
rect 11827 22915 11837 22916
rect -12399 22852 -12309 22875
rect 11466 22851 11476 22915
rect 11540 22852 11837 22915
rect 11901 22915 11911 22916
rect 11901 22852 14589 22915
rect 11540 22851 14589 22852
rect -12762 22724 -12087 22777
rect -16609 22660 -16599 22724
rect -16535 22713 8129 22724
rect -16535 22660 -12687 22713
rect -12151 22660 8129 22713
rect 8193 22660 8203 22724
rect -12401 22623 -12313 22629
rect -12401 22559 -12389 22623
rect -12325 22559 -12313 22623
rect -12401 22543 -12313 22559
rect -12401 22479 -12389 22543
rect -12325 22479 -12313 22543
rect -12401 22463 -12313 22479
rect -12401 22399 -12389 22463
rect -12325 22399 -12313 22463
rect -12401 22394 -12313 22399
rect -17046 22209 7601 22273
rect 7665 22209 7675 22273
rect -17046 21097 -16982 22209
rect 14525 22091 14589 22851
rect 15481 22851 16400 22915
rect 15481 22091 15545 22851
rect 14525 22027 15545 22091
rect 16336 22084 16400 22851
rect 17405 22851 18389 22915
rect 17405 22084 17469 22851
rect 18325 22493 18389 22851
rect 18900 22851 19930 22915
rect 18900 22493 18964 22851
rect 18325 22429 18964 22493
rect 16336 22020 17469 22084
rect 19866 21655 19930 22851
rect 36904 22809 37166 22815
rect 35090 22790 35290 22795
rect 36904 22790 36923 22809
rect 35090 22768 36923 22790
rect 35090 22632 35122 22768
rect 35258 22727 36923 22768
rect 35258 22671 35782 22727
rect 35838 22671 35862 22727
rect 35918 22671 35942 22727
rect 35998 22671 36923 22727
rect 35258 22632 36923 22671
rect 35090 22610 36923 22632
rect 35090 22605 35290 22610
rect 36904 22585 36923 22610
rect 37147 22585 37166 22809
rect 36904 22579 37166 22585
rect 47546 22734 47802 22739
rect 47546 22724 62907 22734
rect 47546 22508 47566 22724
rect 47782 22508 62907 22724
rect 47546 22498 62907 22508
rect 47546 22493 47802 22498
rect 39336 22385 39430 22393
rect 39336 22349 39355 22385
rect 39411 22349 39430 22385
rect 39336 22285 39351 22349
rect 39415 22285 39430 22349
rect 37816 22247 37906 22285
rect 37816 22183 37829 22247
rect 37893 22183 37906 22247
rect 37816 22146 37906 22183
rect 39336 22269 39355 22285
rect 39411 22269 39430 22285
rect 39336 22205 39351 22269
rect 39415 22205 39430 22269
rect 39336 22169 39355 22205
rect 39411 22169 39430 22205
rect 39336 22162 39430 22169
rect 37804 21794 37909 21828
rect 37804 21730 37824 21794
rect 37888 21730 37909 21794
rect 37804 21714 37909 21730
rect -981 21625 -897 21630
rect 6297 21625 6381 21630
rect -981 21621 6381 21625
rect -981 21565 -967 21621
rect -911 21565 6311 21621
rect 6367 21565 6381 21621
rect 12062 21591 12072 21655
rect 12136 21591 27657 21655
rect 27721 21591 27731 21655
rect 37804 21650 37824 21714
rect 37888 21650 37909 21714
rect 37804 21616 37909 21650
rect 39331 21822 39437 21839
rect 39331 21758 39352 21822
rect 39416 21758 39437 21822
rect 39331 21742 39437 21758
rect 39331 21678 39352 21742
rect 39416 21678 39437 21742
rect 39331 21662 39437 21678
rect -981 21561 6381 21565
rect -981 21556 -897 21561
rect 6297 21556 6381 21561
rect 35126 21585 35244 21615
rect 35126 21521 35152 21585
rect 35216 21521 35244 21585
rect 39331 21598 39352 21662
rect 39416 21598 39437 21662
rect 39331 21581 39437 21598
rect 35126 21488 35244 21521
rect 35457 21379 35564 21402
rect 35457 21315 35477 21379
rect 35541 21315 35564 21379
rect 35457 21293 35564 21315
rect 42844 21155 46198 21183
rect -27920 21033 6374 21097
rect 42844 21091 42889 21155
rect 42953 21091 42969 21155
rect 43033 21091 43049 21155
rect 43113 21091 43129 21155
rect 43193 21091 43209 21155
rect 43273 21091 43289 21155
rect 43353 21091 43369 21155
rect 43433 21091 43449 21155
rect 43513 21091 43529 21155
rect 43593 21091 43609 21155
rect 43673 21091 43689 21155
rect 43753 21091 43769 21155
rect 43833 21091 43849 21155
rect 43913 21091 43929 21155
rect 43993 21091 44009 21155
rect 44073 21091 44089 21155
rect 44153 21091 44169 21155
rect 44233 21091 44249 21155
rect 44313 21091 44329 21155
rect 44393 21091 44409 21155
rect 44473 21091 44489 21155
rect 44553 21091 44569 21155
rect 44633 21091 44649 21155
rect 44713 21091 44729 21155
rect 44793 21091 44809 21155
rect 44873 21091 44889 21155
rect 44953 21091 44969 21155
rect 45033 21091 45049 21155
rect 45113 21091 45129 21155
rect 45193 21091 45209 21155
rect 45273 21091 45289 21155
rect 45353 21091 45369 21155
rect 45433 21091 45449 21155
rect 45513 21091 45529 21155
rect 45593 21091 45609 21155
rect 45673 21091 45689 21155
rect 45753 21091 45769 21155
rect 45833 21091 45849 21155
rect 45913 21091 45929 21155
rect 45993 21091 46009 21155
rect 46073 21091 46089 21155
rect 46153 21091 46198 21155
rect 42844 21064 46198 21091
rect -38178 19058 -34851 19070
rect -38178 18994 -38147 19058
rect -38083 18994 -38067 19058
rect -38003 18994 -37987 19058
rect -37923 18994 -37907 19058
rect -37843 18994 -37827 19058
rect -37763 18994 -37747 19058
rect -37683 18994 -37667 19058
rect -37603 18994 -37587 19058
rect -37523 18994 -37507 19058
rect -37443 18994 -37427 19058
rect -37363 18994 -37347 19058
rect -37283 18994 -37267 19058
rect -37203 18994 -37187 19058
rect -37123 18994 -37107 19058
rect -37043 18994 -37027 19058
rect -36963 18994 -36947 19058
rect -36883 18994 -36867 19058
rect -36803 18994 -36787 19058
rect -36723 18994 -36707 19058
rect -36643 18994 -36627 19058
rect -36563 18994 -36547 19058
rect -36483 18994 -36467 19058
rect -36403 18994 -36387 19058
rect -36323 18994 -36307 19058
rect -36243 18994 -36227 19058
rect -36163 18994 -36147 19058
rect -36083 18994 -36067 19058
rect -36003 18994 -35987 19058
rect -35923 18994 -35907 19058
rect -35843 18994 -35827 19058
rect -35763 18994 -35747 19058
rect -35683 18994 -35667 19058
rect -35603 18994 -35587 19058
rect -35523 18994 -35507 19058
rect -35443 18994 -35427 19058
rect -35363 18994 -35347 19058
rect -35283 18994 -35267 19058
rect -35203 18994 -35187 19058
rect -35123 18994 -35107 19058
rect -35043 18994 -35027 19058
rect -34963 18994 -34947 19058
rect -34883 18994 -34851 19058
rect -38178 18982 -34851 18994
rect -40606 17630 -40350 17635
rect -57094 17620 -40350 17630
rect -57094 17404 -40586 17620
rect -40370 17404 -40350 17620
rect -57094 17394 -40350 17404
rect -40606 17389 -40350 17394
rect -38184 16063 -34842 16080
rect -38184 15999 -38145 16063
rect -38081 15999 -38065 16063
rect -38001 15999 -37985 16063
rect -37921 15999 -37905 16063
rect -37841 15999 -37825 16063
rect -37761 15999 -37745 16063
rect -37681 15999 -37665 16063
rect -37601 15999 -37585 16063
rect -37521 15999 -37505 16063
rect -37441 15999 -37425 16063
rect -37361 15999 -37345 16063
rect -37281 15999 -37265 16063
rect -37201 15999 -37185 16063
rect -37121 15999 -37105 16063
rect -37041 15999 -37025 16063
rect -36961 15999 -36945 16063
rect -36881 15999 -36865 16063
rect -36801 15999 -36785 16063
rect -36721 15999 -36705 16063
rect -36641 15999 -36625 16063
rect -36561 15999 -36545 16063
rect -36481 15999 -36465 16063
rect -36401 15999 -36385 16063
rect -36321 15999 -36305 16063
rect -36241 15999 -36225 16063
rect -36161 15999 -36145 16063
rect -36081 15999 -36065 16063
rect -36001 15999 -35985 16063
rect -35921 15999 -35905 16063
rect -35841 15999 -35825 16063
rect -35761 15999 -35745 16063
rect -35681 15999 -35665 16063
rect -35601 15999 -35585 16063
rect -35521 15999 -35505 16063
rect -35441 15999 -35425 16063
rect -35361 15999 -35345 16063
rect -35281 15999 -35265 16063
rect -35201 15999 -35185 16063
rect -35121 15999 -35105 16063
rect -35041 15999 -35025 16063
rect -34961 15999 -34945 16063
rect -34881 15999 -34842 16063
rect -38184 15982 -34842 15999
rect -27920 15446 -27856 21033
rect 6310 20962 6374 21033
rect 14678 21027 14762 21032
rect 12926 20963 12936 21027
rect 13000 21023 14762 21027
rect 13000 20967 14692 21023
rect 14748 20967 14762 21023
rect 13000 20963 14762 20967
rect 6300 20953 6384 20962
rect 14678 20958 14762 20963
rect 6300 20897 6314 20953
rect 6370 20897 6384 20953
rect 6300 20888 6384 20897
rect -981 20715 -897 20720
rect -24170 20711 -897 20715
rect -24170 20655 -967 20711
rect -911 20655 -897 20711
rect -24170 20651 -897 20655
rect -25462 17886 -25377 17927
rect -25462 17822 -25452 17886
rect -25388 17822 -25377 17886
rect -25462 17806 -25377 17822
rect -25462 17742 -25452 17806
rect -25388 17742 -25377 17806
rect -25462 17726 -25377 17742
rect -25462 17662 -25452 17726
rect -25388 17662 -25377 17726
rect -25462 17622 -25377 17662
rect -25460 17398 -25368 17409
rect -25460 17334 -25446 17398
rect -25382 17334 -25368 17398
rect -25460 17318 -25368 17334
rect -25460 17254 -25446 17318
rect -25382 17254 -25368 17318
rect -25460 17238 -25368 17254
rect -25460 17174 -25446 17238
rect -25382 17174 -25368 17238
rect -25460 17164 -25368 17174
rect -24170 16254 -24106 20651
rect -16609 20587 -16599 20651
rect -16535 20587 -16525 20651
rect -981 20646 -897 20651
rect -7442 20270 11080 20334
rect 11144 20270 11154 20334
rect -10445 17157 -10321 17194
rect -10445 17093 -10416 17157
rect -10352 17093 -10321 17157
rect -10445 17061 -10321 17093
rect -10425 16288 -10341 16293
rect -10785 16284 -10341 16288
rect -24180 16245 -24096 16254
rect -24180 16189 -24166 16245
rect -24110 16189 -24096 16245
rect -18719 16203 -17699 16267
rect -16119 16203 -15099 16267
rect -13519 16203 -12499 16267
rect -10785 16228 -10411 16284
rect -10355 16228 -10341 16284
rect -10785 16224 -10341 16228
rect -10425 16219 -10341 16224
rect -24180 16180 -24096 16189
rect -27930 15437 -27846 15446
rect -27930 15381 -27916 15437
rect -27860 15381 -27846 15437
rect -27930 15372 -27846 15381
rect -19071 14880 -19007 15900
rect -14194 15370 -14046 15407
rect -14194 15306 -14152 15370
rect -14088 15306 -14046 15370
rect -14194 15269 -14046 15306
rect -12197 14873 -12133 15893
rect -15965 14472 -15232 14536
rect -25527 14413 -25434 14451
rect -25527 14349 -25513 14413
rect -25449 14349 -25434 14413
rect -25527 14333 -25434 14349
rect -25527 14269 -25513 14333
rect -25449 14269 -25434 14333
rect -25527 14253 -25434 14269
rect -25527 14189 -25513 14253
rect -25449 14189 -25434 14253
rect -25527 14152 -25434 14189
rect -13074 14141 -12990 14146
rect -13331 14137 -12990 14141
rect -18240 14073 -18139 14097
rect -13331 14081 -13060 14137
rect -13004 14081 -12990 14137
rect -13331 14077 -12990 14081
rect -18240 14009 -18223 14073
rect -18159 14009 -18139 14073
rect -13074 14072 -12990 14077
rect -18240 13986 -18139 14009
rect -25528 13919 -25436 13930
rect -25528 13855 -25514 13919
rect -25450 13855 -25436 13919
rect -25528 13839 -25436 13855
rect -25528 13775 -25514 13839
rect -25450 13775 -25436 13839
rect -25528 13759 -25436 13775
rect -25528 13695 -25514 13759
rect -25450 13695 -25436 13759
rect -25528 13685 -25436 13695
rect -19071 12280 -19007 13300
rect -12197 12273 -12133 13293
rect -18722 11937 -17702 12001
rect -16122 11937 -15102 12001
rect -13522 11937 -12502 12001
rect -10999 10223 -10881 10250
rect -10999 10159 -10970 10223
rect -10906 10159 -10881 10223
rect -10999 10138 -10881 10159
rect -7442 9819 -7378 20270
rect -6759 19739 11476 19803
rect 11540 19739 11550 19803
rect -6759 10646 -6695 19739
rect 41 19513 125 19518
rect -2825 19449 -2815 19513
rect -2751 19509 125 19513
rect -2751 19453 55 19509
rect 111 19453 125 19509
rect -2751 19449 125 19453
rect -5289 18979 -5279 19043
rect -5215 18979 -5205 19043
rect -3928 18979 -3918 19043
rect -3854 18979 -3844 19043
rect -5279 18871 -5215 18979
rect -5279 18807 -4725 18871
rect -3918 18870 -3854 18979
rect -5815 15708 -5690 15744
rect -5815 15644 -5786 15708
rect -5722 15644 -5690 15708
rect -5815 15613 -5690 15644
rect -4789 14637 -4725 18807
rect -4448 18806 -3854 18870
rect -4789 14573 -4552 14637
rect -4912 14413 -4822 14451
rect -4912 14349 -4899 14413
rect -4835 14349 -4822 14413
rect -4912 14333 -4822 14349
rect -4912 14269 -4899 14333
rect -4835 14269 -4822 14333
rect -4912 14231 -4822 14269
rect -4914 14003 -4850 14011
rect -4927 13960 -4823 14003
rect -4927 13904 -4903 13960
rect -4847 13904 -4823 13960
rect -4927 13880 -4823 13904
rect -4927 13824 -4903 13880
rect -4847 13824 -4823 13880
rect -4927 13800 -4823 13824
rect -4927 13744 -4903 13800
rect -4847 13744 -4823 13800
rect -4927 13701 -4823 13744
rect -4914 13279 -4850 13701
rect -5014 13215 -4850 13279
rect -5717 10838 -5391 10843
rect -5014 10838 -4950 13215
rect -4616 12380 -4552 14573
rect -6172 10827 -5927 10838
rect -6172 10763 -6162 10827
rect -6098 10763 -6082 10827
rect -6018 10763 -6002 10827
rect -5938 10763 -5927 10827
rect -5735 10822 -4950 10838
rect -5735 10774 -5702 10822
rect -6172 10753 -5927 10763
rect -5717 10766 -5702 10774
rect -5646 10766 -5622 10822
rect -5566 10766 -5542 10822
rect -5486 10766 -5462 10822
rect -5406 10774 -4950 10822
rect -5406 10766 -5391 10774
rect -5717 10746 -5391 10766
rect -6759 10582 -6092 10646
rect -6156 10209 -6092 10582
rect -6166 10200 -6082 10209
rect -6166 10144 -6152 10200
rect -6096 10144 -6082 10200
rect -6166 10135 -6082 10144
rect -5371 10200 -5287 10209
rect -5371 10144 -5357 10200
rect -5301 10144 -5287 10200
rect -5371 10135 -5287 10144
rect -5361 9819 -5297 10135
rect -7442 9755 -5297 9819
rect -6177 9584 -5919 9597
rect -6177 9520 -6160 9584
rect -6096 9520 -6080 9584
rect -6016 9520 -6000 9584
rect -5936 9520 -5919 9584
rect -6177 9508 -5919 9520
rect -5718 9580 -5389 9600
rect -5718 9524 -5702 9580
rect -5646 9524 -5622 9580
rect -5566 9524 -5542 9580
rect -5486 9524 -5462 9580
rect -5406 9572 -5389 9580
rect -5014 9572 -4950 10774
rect -4789 12316 -4552 12380
rect -4789 10238 -4725 12316
rect -4448 10238 -4384 18806
rect -2815 18299 -2751 19449
rect 41 19444 125 19449
rect 23667 19382 23776 19404
rect 14661 19327 14777 19351
rect 14661 19263 14687 19327
rect 14751 19263 14777 19327
rect 23667 19318 23689 19382
rect 23753 19318 23776 19382
rect 23667 19292 23776 19318
rect 14661 19242 14777 19263
rect -766 19212 -682 19217
rect -2408 19148 -2398 19212
rect -2334 19208 -682 19212
rect -2334 19152 -752 19208
rect -696 19152 -682 19208
rect -2334 19148 -682 19152
rect -766 19143 -682 19148
rect 4847 19172 5204 19178
rect 3051 19106 3135 19111
rect 4847 19106 4873 19172
rect 3051 19102 4873 19106
rect 3051 19046 3065 19102
rect 3121 19046 4873 19102
rect 3051 19042 4873 19046
rect 3051 19037 3135 19042
rect 4847 19028 4873 19042
rect 5177 19106 5204 19172
rect 7075 19106 7159 19111
rect 8971 19106 9055 19111
rect 5177 19102 9089 19106
rect 5177 19046 7089 19102
rect 7145 19046 8985 19102
rect 9041 19046 9089 19102
rect 5177 19042 9089 19046
rect 10203 19058 10327 19083
rect 5177 19028 5204 19042
rect 7075 19037 7159 19042
rect 8971 19037 9055 19042
rect 4847 19022 5204 19028
rect 10203 18994 10232 19058
rect 10296 18994 10327 19058
rect 10203 18968 10327 18994
rect 20928 19062 21079 19106
rect 20928 18998 20971 19062
rect 21035 18998 21079 19062
rect 20928 18951 21079 18998
rect 5697 18910 5781 18915
rect 7696 18910 7780 18915
rect -1514 18846 -1504 18910
rect -1440 18906 7780 18910
rect -1440 18850 5711 18906
rect 5767 18850 7710 18906
rect 7766 18850 7780 18906
rect -1440 18846 7780 18850
rect 5697 18841 5781 18846
rect 7696 18841 7780 18846
rect 8239 18718 8373 18758
rect 4889 18651 4973 18656
rect 6887 18651 6971 18656
rect -1143 18587 -1133 18651
rect -1069 18647 6971 18651
rect -1069 18591 4903 18647
rect 4959 18591 6901 18647
rect 6957 18591 6971 18647
rect 8239 18654 8280 18718
rect 8344 18654 8373 18718
rect 13564 18688 13648 18693
rect 8239 18617 8373 18654
rect 12920 18624 12930 18688
rect 12994 18684 13648 18688
rect 12994 18628 13578 18684
rect 13634 18628 13648 18684
rect 12994 18624 13648 18628
rect 13564 18619 13648 18624
rect -1069 18587 6971 18591
rect 4889 18582 4973 18587
rect 6887 18582 6971 18587
rect 14105 18507 14115 18571
rect 14179 18507 14189 18571
rect 25604 18507 25614 18571
rect 25678 18507 25688 18571
rect 3697 18312 3781 18317
rect 9696 18312 9780 18317
rect -3509 18235 -2751 18299
rect -690 18248 -680 18312
rect -616 18308 9780 18312
rect -616 18252 3711 18308
rect 3767 18252 9710 18308
rect 9766 18252 9780 18308
rect -616 18248 9780 18252
rect 3697 18243 3781 18248
rect 9696 18243 9780 18248
rect -3509 16205 -3445 18235
rect 2888 18031 2972 18036
rect 8889 18031 8973 18036
rect -294 17967 -284 18031
rect -220 18027 8973 18031
rect -220 17971 2902 18027
rect 2958 17971 8903 18027
rect 8959 17971 8973 18027
rect -220 17967 8973 17971
rect 2888 17962 2972 17967
rect 8889 17962 8973 17967
rect -3221 17856 -2738 17864
rect -3221 17632 -3172 17856
rect -2788 17772 -2738 17856
rect 223 17772 307 17777
rect -2788 17768 307 17772
rect -2788 17712 237 17768
rect 293 17712 307 17768
rect -2788 17708 307 17712
rect -2788 17632 -2738 17708
rect 223 17703 307 17708
rect 14358 17699 14368 17763
rect 14432 17699 14442 17763
rect 25351 17700 25361 17764
rect 25425 17700 25435 17764
rect -3221 17624 -2738 17632
rect 14662 17542 14782 17566
rect -831 17525 -747 17530
rect -847 17521 981 17525
rect -847 17465 -817 17521
rect -761 17465 981 17521
rect -847 17461 981 17465
rect 1045 17461 1077 17525
rect 14662 17478 14689 17542
rect 14753 17478 14782 17542
rect -831 17456 -747 17461
rect 14662 17449 14782 17478
rect 23665 17552 23778 17575
rect 23665 17488 23689 17552
rect 23753 17488 23778 17552
rect 23665 17458 23778 17488
rect 4268 17289 4387 17313
rect 4268 17225 4295 17289
rect 4359 17225 4387 17289
rect 4268 17194 4387 17225
rect 6200 17289 6319 17314
rect 6200 17225 6227 17289
rect 6291 17225 6319 17289
rect 6200 17195 6319 17225
rect 13593 17083 13677 17088
rect 12946 17019 12956 17083
rect 13020 17079 13677 17083
rect 13020 17023 13607 17079
rect 13663 17023 13677 17079
rect 13020 17019 13677 17023
rect 13593 17014 13677 17019
rect 18 16414 11149 16451
rect 18 16413 263 16414
rect -2932 16270 263 16413
rect 11127 16270 11149 16414
rect -2932 16252 11149 16270
rect 18 16233 11149 16252
rect -3519 16141 -3509 16205
rect -3445 16141 -3435 16205
rect 18 16184 248 16233
rect 18 16162 197 16184
rect -3018 15454 -2934 15459
rect -3938 15390 -3928 15454
rect -3864 15450 -2934 15454
rect -3864 15394 -3004 15450
rect -2948 15394 -2934 15450
rect -3864 15390 -2934 15394
rect -3018 15385 -2934 15390
rect -3154 14970 -3051 15003
rect -3154 14906 -3135 14970
rect -3071 14906 -3051 14970
rect -3154 14890 -3051 14906
rect -3154 14826 -3135 14890
rect -3071 14826 -3051 14890
rect -3154 14810 -3051 14826
rect -3154 14746 -3135 14810
rect -3071 14746 -3051 14810
rect -3154 14714 -3051 14746
rect -3033 14644 -2949 14649
rect -3519 14580 -3509 14644
rect -3445 14640 -2949 14644
rect -3445 14584 -3019 14640
rect -2963 14584 -2949 14640
rect -3445 14580 -2949 14584
rect -3033 14575 -2949 14580
rect 18 13993 39 16162
rect -2956 13832 39 13993
rect -2608 13133 -2524 13142
rect -2608 13077 -2594 13133
rect -2538 13077 -2524 13133
rect -2608 13068 -2524 13077
rect -1818 13121 -1715 13138
rect -2895 12324 -2811 12333
rect -2895 12268 -2881 12324
rect -2825 12268 -2811 12324
rect -2895 12259 -2811 12268
rect -4799 10229 -4715 10238
rect -4799 10173 -4785 10229
rect -4729 10173 -4715 10229
rect -4799 10164 -4715 10173
rect -4458 10229 -4374 10238
rect -4458 10173 -4444 10229
rect -4388 10173 -4374 10229
rect -4458 10164 -4374 10173
rect -5406 9524 -4950 9572
rect -5718 9508 -4950 9524
rect -5718 9504 -5389 9508
rect -5014 8707 -4950 9508
rect -5014 8643 -3185 8707
rect -3121 8643 -3111 8707
rect -18719 8403 -17699 8467
rect -16119 8403 -15099 8467
rect -13519 8403 -12499 8467
rect -19071 7080 -19007 8100
rect -16791 7607 -16643 7644
rect -16791 7543 -16749 7607
rect -16685 7543 -16643 7607
rect -16791 7506 -16643 7543
rect -12197 7073 -12133 8093
rect -2885 7532 -2821 12259
rect -2598 8340 -2534 13068
rect -1818 13057 -1799 13121
rect -1735 13057 -1715 13121
rect -1818 13041 -1715 13057
rect -1818 12977 -1799 13041
rect -1735 12977 -1715 13041
rect -1818 12961 -1715 12977
rect -1818 12897 -1799 12961
rect -1735 12897 -1715 12961
rect -1818 12881 -1715 12897
rect -1818 12817 -1799 12881
rect -1735 12817 -1715 12881
rect -1818 12801 -1715 12817
rect -1818 12737 -1799 12801
rect -1735 12737 -1715 12801
rect -1818 12721 -1715 12737
rect -1508 12405 -1424 12414
rect -1508 12349 -1494 12405
rect -1438 12349 -1424 12405
rect -1508 12340 -1424 12349
rect -1936 11531 -1852 11540
rect -1936 11475 -1922 11531
rect -1866 11475 -1852 11531
rect -1936 11466 -1852 11475
rect -1769 11526 -1683 11534
rect -2222 10725 -2138 10734
rect -2222 10669 -2208 10725
rect -2152 10669 -2138 10725
rect -2222 10660 -2138 10669
rect -2212 9134 -2148 10660
rect -1926 9942 -1862 11466
rect -1769 11462 -1758 11526
rect -1694 11462 -1683 11526
rect -1769 11446 -1683 11462
rect -1769 11382 -1758 11446
rect -1694 11382 -1683 11446
rect -1769 11366 -1683 11382
rect -1769 11302 -1758 11366
rect -1694 11302 -1683 11366
rect -1769 11286 -1683 11302
rect -1769 11222 -1758 11286
rect -1694 11222 -1683 11286
rect -1769 11206 -1683 11222
rect -1769 11142 -1758 11206
rect -1694 11142 -1683 11206
rect -1769 11135 -1683 11142
rect -1498 10788 -1434 12340
rect -1508 10779 -1424 10788
rect -1508 10723 -1494 10779
rect -1438 10723 -1424 10779
rect -1508 10714 -1424 10723
rect -1936 9933 -1852 9942
rect -1936 9877 -1922 9933
rect -1866 9877 -1852 9933
rect -1936 9868 -1852 9877
rect -1769 9923 -1685 9935
rect -2222 9125 -2138 9134
rect -2222 9069 -2208 9125
rect -2152 9069 -2138 9125
rect -2222 9060 -2138 9069
rect -2608 8331 -2524 8340
rect -2608 8275 -2594 8331
rect -2538 8275 -2524 8331
rect -2608 8266 -2524 8275
rect -2895 7523 -2811 7532
rect -2895 7467 -2881 7523
rect -2825 7467 -2811 7523
rect -2895 7458 -2811 7467
rect -7224 7235 -6741 7248
rect -7224 7231 -7175 7235
rect -6791 7231 -6741 7235
rect -7224 7015 -7211 7231
rect -6755 7015 -6741 7231
rect -7224 7011 -7175 7015
rect -6791 7011 -6741 7015
rect -7224 6998 -6741 7011
rect -25531 6650 -25436 6674
rect -15965 6672 -15232 6736
rect -4927 6691 -4826 6700
rect -25531 6586 -25516 6650
rect -25452 6586 -25436 6650
rect -25531 6570 -25436 6586
rect -25531 6506 -25516 6570
rect -25452 6506 -25436 6570
rect -25531 6490 -25436 6506
rect -25531 6426 -25516 6490
rect -25452 6426 -25436 6490
rect -25531 6403 -25436 6426
rect -4927 6635 -4905 6691
rect -4849 6649 -4826 6691
rect -4849 6635 -3184 6649
rect -4927 6611 -3184 6635
rect -4927 6555 -4905 6611
rect -4849 6585 -3184 6611
rect -3120 6585 -3110 6649
rect -4849 6555 -4826 6585
rect -4927 6531 -4826 6555
rect -4927 6475 -4905 6531
rect -4849 6475 -4826 6531
rect -4927 6451 -4826 6475
rect -4927 6395 -4905 6451
rect -4849 6395 -4826 6451
rect -4927 6387 -4826 6395
rect -18271 6303 -18171 6328
rect -13085 6313 -13001 6318
rect -18271 6239 -18251 6303
rect -18187 6239 -18171 6303
rect -13326 6309 -13001 6313
rect -13326 6253 -13071 6309
rect -13015 6253 -13001 6309
rect -13326 6249 -13001 6253
rect -13085 6244 -13001 6249
rect -18271 6217 -18171 6239
rect -25532 6163 -25437 6179
rect -25532 6099 -25517 6163
rect -25453 6099 -25437 6163
rect -25532 6083 -25437 6099
rect -25532 6019 -25517 6083
rect -25453 6019 -25437 6083
rect -25532 6003 -25437 6019
rect -25532 5939 -25517 6003
rect -25453 5939 -25437 6003
rect -4917 6128 -4831 6168
rect -4917 6064 -4906 6128
rect -4842 6064 -4831 6128
rect -4917 6048 -4831 6064
rect -4917 5984 -4906 6048
rect -4842 5984 -4831 6048
rect -3060 6042 -2976 6047
rect -4917 5945 -4831 5984
rect -3938 5978 -3928 6042
rect -3864 6038 -2976 6042
rect -3864 5982 -3046 6038
rect -2990 5982 -2976 6038
rect -3864 5978 -2976 5982
rect -3060 5973 -2976 5978
rect -25532 5924 -25437 5939
rect -3203 5548 -3100 5582
rect -19071 4480 -19007 5500
rect -12197 4473 -12133 5493
rect -3203 5484 -3184 5548
rect -3120 5484 -3100 5548
rect -3203 5468 -3100 5484
rect -3203 5404 -3184 5468
rect -3120 5404 -3100 5468
rect -3203 5388 -3100 5404
rect -3203 5324 -3184 5388
rect -3120 5324 -3100 5388
rect -10766 5052 -10702 5314
rect -3203 5291 -3100 5324
rect -3519 5169 -3509 5233
rect -3445 5169 -3435 5233
rect -3038 5229 -2954 5238
rect -3038 5173 -3024 5229
rect -2968 5173 -2954 5229
rect -10776 5043 -10692 5052
rect -10776 4987 -10762 5043
rect -10706 4987 -10692 5043
rect -10776 4978 -10692 4987
rect -3509 4978 -3445 5169
rect -3038 5164 -2954 5173
rect -3031 4978 -2967 5164
rect -3509 4914 -2967 4978
rect -18722 4137 -17702 4201
rect -16122 4137 -15102 4201
rect -13522 4137 -12502 4201
rect -2885 -4979 -2821 7458
rect -2598 -4516 -2534 8266
rect -2212 -3981 -2148 9060
rect -1926 -3509 -1862 9868
rect -1769 9859 -1759 9923
rect -1695 9859 -1685 9923
rect -1769 9843 -1685 9859
rect -1769 9779 -1759 9843
rect -1695 9779 -1685 9843
rect -1769 9763 -1685 9779
rect -1769 9699 -1759 9763
rect -1695 9699 -1685 9763
rect -1769 9683 -1685 9699
rect -1769 9619 -1759 9683
rect -1695 9619 -1685 9683
rect -1769 9603 -1685 9619
rect -1769 9539 -1759 9603
rect -1695 9539 -1685 9603
rect -1769 9527 -1685 9539
rect -1498 9130 -1434 10714
rect 18 10666 39 13832
rect 175 10666 197 16162
rect 11229 16173 11409 16189
rect 11229 14437 11251 16173
rect 11387 15269 11409 16173
rect 23644 15788 23786 15820
rect 14655 15711 14781 15738
rect 14655 15647 14686 15711
rect 14750 15647 14781 15711
rect 23644 15724 23686 15788
rect 23750 15724 23786 15788
rect 23644 15685 23786 15724
rect 14655 15621 14781 15647
rect 20897 15496 21018 15526
rect 20897 15432 20928 15496
rect 20992 15432 21018 15496
rect 20897 15400 21018 15432
rect 11387 15228 13084 15269
rect 14680 15228 14764 15233
rect 11387 15164 12973 15228
rect 13037 15224 14764 15228
rect 13037 15168 14694 15224
rect 14750 15168 14764 15224
rect 13037 15164 14764 15168
rect 11387 15113 13084 15164
rect 14680 15159 14764 15164
rect 11387 14437 11409 15113
rect 11229 14421 11409 14437
rect 23664 13997 23769 14018
rect 14650 13965 14778 13997
rect 11247 13940 11394 13959
rect 11247 13884 11292 13940
rect 11348 13884 11394 13940
rect 11247 13860 11394 13884
rect 14650 13901 14685 13965
rect 14749 13901 14778 13965
rect 23664 13933 23686 13997
rect 23750 13933 23769 13997
rect 23664 13909 23769 13933
rect 14650 13860 14778 13901
rect 11247 13804 11292 13860
rect 11348 13804 11394 13860
rect 11247 13780 11394 13804
rect 11247 13724 11292 13780
rect 11348 13724 11394 13780
rect 11247 13700 11394 13724
rect 11247 13644 11292 13700
rect 11348 13644 11394 13700
rect 11247 13620 11394 13644
rect 11247 13572 11292 13620
rect 11246 13564 11292 13572
rect 11348 13572 11394 13620
rect 11348 13564 13075 13572
rect 11246 13540 13075 13564
rect 11246 13484 11292 13540
rect 11348 13528 13075 13540
rect 13626 13528 13710 13533
rect 11348 13484 13003 13528
rect 11246 13464 13003 13484
rect 13067 13524 13710 13528
rect 13067 13468 13640 13524
rect 13696 13468 13710 13524
rect 13067 13464 13710 13468
rect 11246 13460 13075 13464
rect 11246 13426 11292 13460
rect 11247 13404 11292 13426
rect 11348 13426 13075 13460
rect 13626 13459 13710 13464
rect 11348 13404 11394 13426
rect 11247 13380 11394 13404
rect 11247 13324 11292 13380
rect 11348 13324 11394 13380
rect 11247 13300 11394 13324
rect 11247 13244 11292 13300
rect 11348 13244 11394 13300
rect 11247 13220 11394 13244
rect 11247 13164 11292 13220
rect 11348 13164 11394 13220
rect 11247 13140 11394 13164
rect 11247 13084 11292 13140
rect 11348 13084 11394 13140
rect 14105 13107 14115 13171
rect 14179 13107 14189 13171
rect 11247 13060 11394 13084
rect 11247 13004 11292 13060
rect 11348 13004 11394 13060
rect 11247 12985 11394 13004
rect 14358 12299 14368 12363
rect 14432 12299 14442 12363
rect 14675 12180 14789 12202
rect 11233 12110 11408 12134
rect 11233 11334 11252 12110
rect 11388 11724 11408 12110
rect 14675 12116 14702 12180
rect 14766 12116 14789 12180
rect 14675 12087 14789 12116
rect 23667 12190 23779 12214
rect 23667 12126 23691 12190
rect 23755 12126 23779 12190
rect 23667 12098 23779 12126
rect 20945 11906 21080 11947
rect 20945 11842 20985 11906
rect 21049 11842 21080 11906
rect 20945 11804 21080 11842
rect 11388 11676 13124 11724
rect 13689 11676 13773 11681
rect 11388 11612 13001 11676
rect 13065 11672 13773 11676
rect 13065 11616 13703 11672
rect 13759 11616 13773 11672
rect 13065 11612 13773 11616
rect 11388 11560 13124 11612
rect 13689 11607 13773 11612
rect 11388 11334 11408 11560
rect 11233 11311 11408 11334
rect 18 10635 197 10666
rect 6473 10518 11228 10542
rect 6473 10374 6498 10518
rect 11202 10374 11228 10518
rect 6473 10351 11228 10374
rect 14666 10383 14780 10406
rect 14666 10319 14691 10383
rect 14755 10319 14780 10383
rect 14666 10290 14780 10319
rect 23664 10380 23783 10410
rect 23664 10316 23691 10380
rect 23755 10316 23783 10380
rect 23664 10286 23783 10316
rect 36043 9154 36151 9176
rect -1508 9121 -1424 9130
rect -1508 9065 -1494 9121
rect -1438 9065 -1424 9121
rect -1508 9056 -1424 9065
rect 36043 9090 36066 9154
rect 36130 9090 36151 9154
rect 36043 9064 36151 9090
rect -1768 8322 -1680 8335
rect -1768 8258 -1756 8322
rect -1692 8258 -1680 8322
rect -1768 8242 -1680 8258
rect -1768 8178 -1756 8242
rect -1692 8178 -1680 8242
rect -1768 8162 -1680 8178
rect -1768 8098 -1756 8162
rect -1692 8098 -1680 8162
rect -1768 8082 -1680 8098
rect -1768 8018 -1756 8082
rect -1692 8018 -1680 8082
rect -1768 8002 -1680 8018
rect -1768 7938 -1756 8002
rect -1692 7938 -1680 8002
rect -1768 7925 -1680 7938
rect -1498 7591 -1434 9056
rect 36888 8786 37150 8792
rect 36888 8705 36907 8786
rect 34644 8641 36907 8705
rect 34644 8336 34708 8641
rect 35459 8531 35583 8563
rect 36888 8562 36907 8641
rect 37131 8562 37150 8786
rect 36888 8556 37150 8562
rect 35459 8467 35489 8531
rect 35553 8467 35583 8531
rect 35459 8436 35583 8467
rect 36604 8469 36720 8498
rect 36604 8405 36631 8469
rect 36695 8405 36720 8469
rect 36604 8377 36720 8405
rect 34644 8288 35088 8336
rect 34644 8279 35098 8288
rect 34644 8272 35028 8279
rect -1508 7582 -1424 7591
rect -1508 7526 -1494 7582
rect -1438 7526 -1424 7582
rect -1508 7517 -1424 7526
rect -1498 7263 -1434 7517
rect -1508 7224 -1424 7263
rect -1508 7168 -1494 7224
rect -1438 7168 -1424 7224
rect -1508 7144 -1424 7168
rect -1508 7088 -1494 7144
rect -1438 7088 -1424 7144
rect -1508 7064 -1424 7088
rect -1508 7008 -1494 7064
rect -1438 7008 -1424 7064
rect -1508 6969 -1424 7008
rect 34644 7013 34708 8272
rect 35014 8223 35028 8272
rect 35084 8223 35098 8279
rect 35014 8214 35098 8223
rect 40011 8095 40269 8135
rect 38558 8033 39142 8083
rect 38558 7977 38582 8033
rect 38638 7977 39142 8033
rect 38558 7953 39142 7977
rect 38558 7897 38582 7953
rect 38638 7913 39142 7953
rect 40011 8039 40112 8095
rect 40168 8039 40269 8095
rect 40011 8015 40269 8039
rect 40011 7959 40112 8015
rect 40168 7959 40269 8015
rect 40011 7913 40269 7959
rect 38638 7897 40721 7913
rect 36007 7875 36581 7896
rect 36007 7819 36308 7875
rect 36364 7819 36388 7875
rect 36444 7819 36468 7875
rect 36524 7819 36581 7875
rect 38558 7843 40721 7897
rect 36007 7800 36581 7819
rect 35008 7223 35127 7253
rect 35008 7159 35028 7223
rect 35092 7188 35127 7223
rect 36007 7188 36103 7800
rect 38902 7673 40721 7843
rect 38558 7541 38659 7568
rect 38558 7477 38576 7541
rect 38640 7477 38659 7541
rect 38558 7461 38659 7477
rect 38558 7397 38576 7461
rect 38640 7397 38659 7461
rect 38558 7370 38659 7397
rect 36338 7334 37077 7349
rect 36338 7278 36378 7334
rect 36434 7278 36458 7334
rect 36514 7333 37077 7334
rect 36514 7278 36987 7333
rect 36338 7269 36987 7278
rect 37051 7269 37077 7333
rect 36338 7253 37077 7269
rect 35092 7159 36103 7188
rect 35008 7124 36103 7159
rect 35008 7123 35127 7124
rect -1498 6456 -1434 6969
rect 34644 6959 35091 7013
rect 34644 6950 35101 6959
rect 34644 6949 35031 6950
rect -1508 6447 -1424 6456
rect -1508 6391 -1494 6447
rect -1438 6391 -1424 6447
rect -1508 6382 -1424 6391
rect 34644 5623 34708 6949
rect 35017 6894 35031 6949
rect 35087 6894 35101 6950
rect 35017 6885 35101 6894
rect 36007 6816 36103 7124
rect 36007 6800 36442 6816
rect 36007 6786 36447 6800
rect 36007 6730 36366 6786
rect 36422 6730 36447 6786
rect 38902 6765 39142 7673
rect 40077 7554 40178 7581
rect 40077 7490 40095 7554
rect 40159 7490 40178 7554
rect 40077 7474 40178 7490
rect 40077 7410 40095 7474
rect 40159 7410 40178 7474
rect 40077 7383 40178 7410
rect 40481 7170 40721 7673
rect 42592 7219 45933 7237
rect 40481 7162 41274 7170
rect 40481 6938 40840 7162
rect 41224 6938 41274 7162
rect 42592 7155 42630 7219
rect 42694 7155 42710 7219
rect 42774 7155 42790 7219
rect 42854 7155 42870 7219
rect 42934 7155 42950 7219
rect 43014 7155 43030 7219
rect 43094 7155 43110 7219
rect 43174 7155 43190 7219
rect 43254 7155 43270 7219
rect 43334 7155 43350 7219
rect 43414 7155 43430 7219
rect 43494 7155 43510 7219
rect 43574 7155 43590 7219
rect 43654 7155 43670 7219
rect 43734 7155 43750 7219
rect 43814 7155 43830 7219
rect 43894 7155 43910 7219
rect 43974 7155 43990 7219
rect 44054 7155 44070 7219
rect 44134 7155 44150 7219
rect 44214 7155 44230 7219
rect 44294 7155 44310 7219
rect 44374 7155 44390 7219
rect 44454 7155 44470 7219
rect 44534 7155 44550 7219
rect 44614 7155 44630 7219
rect 44694 7155 44710 7219
rect 44774 7155 44790 7219
rect 44854 7155 44870 7219
rect 44934 7155 44950 7219
rect 45014 7155 45030 7219
rect 45094 7155 45110 7219
rect 45174 7155 45190 7219
rect 45254 7155 45270 7219
rect 45334 7155 45350 7219
rect 45414 7155 45430 7219
rect 45494 7155 45510 7219
rect 45574 7155 45590 7219
rect 45654 7155 45670 7219
rect 45734 7155 45750 7219
rect 45814 7155 45830 7219
rect 45894 7155 45933 7219
rect 42592 7138 45933 7155
rect 40481 6930 41274 6938
rect 40481 6797 40721 6930
rect 36007 6720 36447 6730
rect 36342 6716 36447 6720
rect 35000 5885 35108 5908
rect 35000 5821 35027 5885
rect 35091 5866 35108 5885
rect 35091 5821 35644 5866
rect 35000 5802 35644 5821
rect 35000 5796 35108 5802
rect 35580 5714 35644 5802
rect 36346 5727 36442 6716
rect 38541 6672 39142 6765
rect 38541 6616 38582 6672
rect 38638 6616 39142 6672
rect 38541 6525 39142 6616
rect 40076 6759 40721 6797
rect 40076 6703 40104 6759
rect 40160 6703 40721 6759
rect 40076 6679 40721 6703
rect 40076 6623 40104 6679
rect 40160 6623 40721 6679
rect 40076 6557 40721 6623
rect 36961 6249 37077 6270
rect 36961 6185 36987 6249
rect 37051 6185 37077 6249
rect 36961 6164 37077 6185
rect 38553 6210 38654 6237
rect 38553 6146 38571 6210
rect 38635 6146 38654 6210
rect 38553 6130 38654 6146
rect 38553 6066 38571 6130
rect 38635 6066 38654 6130
rect 38553 6039 38654 6066
rect 35934 5714 36442 5727
rect 35580 5703 36442 5714
rect 35580 5650 35991 5703
rect 35934 5647 35991 5650
rect 36047 5647 36071 5703
rect 36127 5647 36442 5703
rect 35934 5631 36442 5647
rect 34644 5567 35088 5623
rect 34644 5559 35098 5567
rect 34644 4288 34708 5559
rect 35014 5558 35098 5559
rect 35014 5502 35028 5558
rect 35084 5502 35098 5558
rect 35014 5493 35098 5502
rect 35934 4727 36030 5631
rect 38902 5395 39142 6525
rect 40082 6207 40183 6234
rect 40082 6143 40100 6207
rect 40164 6143 40183 6207
rect 40082 6127 40183 6143
rect 40082 6063 40100 6127
rect 40164 6063 40183 6127
rect 40082 6036 40183 6063
rect 40481 5416 40721 6557
rect 47463 5800 47719 5805
rect 47463 5790 62907 5800
rect 47463 5574 47483 5790
rect 47699 5574 62907 5790
rect 47463 5564 62907 5574
rect 47463 5559 47719 5564
rect 38561 5282 39142 5395
rect 38561 5226 38583 5282
rect 38639 5226 39142 5282
rect 36498 5161 37077 5177
rect 36498 5155 36987 5161
rect 36498 5099 36516 5155
rect 36572 5099 36596 5155
rect 36652 5099 36676 5155
rect 36732 5099 36987 5155
rect 36498 5097 36987 5099
rect 37051 5097 37077 5161
rect 38561 5155 39142 5226
rect 40088 5379 40721 5416
rect 40088 5323 40121 5379
rect 40177 5323 40721 5379
rect 40088 5299 40721 5323
rect 40088 5243 40121 5299
rect 40177 5243 40721 5299
rect 40088 5176 40721 5243
rect 36498 5081 37077 5097
rect 38552 4857 38653 4884
rect 38552 4793 38570 4857
rect 38634 4793 38653 4857
rect 38552 4777 38653 4793
rect 35934 4633 36445 4727
rect 38552 4713 38570 4777
rect 38634 4713 38653 4777
rect 38552 4686 38653 4713
rect 35934 4631 36537 4633
rect 36349 4612 36537 4631
rect 36349 4556 36368 4612
rect 36424 4556 36448 4612
rect 36504 4556 36537 4612
rect 36349 4537 36537 4556
rect 35014 4492 35119 4516
rect 35014 4428 35035 4492
rect 35099 4480 35119 4492
rect 36349 4480 36445 4537
rect 35099 4428 36445 4480
rect 35014 4416 36445 4428
rect 35014 4403 35119 4416
rect 34644 4224 35088 4288
rect 35014 4192 35088 4224
rect 35014 4183 35098 4192
rect 35014 4127 35028 4183
rect 35084 4127 35098 4183
rect 35014 4118 35098 4127
rect 36349 3627 36445 4416
rect 36962 4073 37078 4094
rect 36962 4009 36988 4073
rect 37052 4009 37078 4073
rect 36962 3988 37078 4009
rect 38902 3986 39142 5155
rect 40082 4835 40183 4862
rect 40082 4771 40100 4835
rect 40164 4771 40183 4835
rect 40082 4755 40183 4771
rect 40082 4691 40100 4755
rect 40164 4691 40183 4755
rect 40082 4664 40183 4691
rect 40481 4267 40721 5176
rect 40481 4259 41272 4267
rect 38548 3925 39142 3986
rect 38548 3869 38583 3925
rect 38639 3869 39142 3925
rect 38548 3845 39142 3869
rect 38548 3789 38583 3845
rect 38639 3818 39142 3845
rect 40015 4000 40255 4037
rect 40015 3944 40111 4000
rect 40167 3944 40255 4000
rect 40015 3920 40255 3944
rect 40015 3864 40111 3920
rect 40167 3864 40255 3920
rect 40015 3818 40255 3864
rect 40481 4035 40838 4259
rect 41222 4035 41272 4259
rect 42589 4220 45969 4238
rect 42589 4156 42607 4220
rect 42671 4156 42687 4220
rect 42751 4156 42767 4220
rect 42831 4156 42847 4220
rect 42911 4156 42927 4220
rect 42991 4156 43007 4220
rect 43071 4156 43087 4220
rect 43151 4156 43167 4220
rect 43231 4156 43247 4220
rect 43311 4156 43327 4220
rect 43391 4156 43407 4220
rect 43471 4156 43487 4220
rect 43551 4156 43567 4220
rect 43631 4156 43647 4220
rect 43711 4156 43727 4220
rect 43791 4156 43807 4220
rect 43871 4156 43887 4220
rect 43951 4156 43967 4220
rect 44031 4156 44047 4220
rect 44111 4156 44127 4220
rect 44191 4156 44207 4220
rect 44271 4156 44287 4220
rect 44351 4156 44367 4220
rect 44431 4156 44447 4220
rect 44511 4156 44527 4220
rect 44591 4156 44607 4220
rect 44671 4156 44687 4220
rect 44751 4156 44767 4220
rect 44831 4156 44847 4220
rect 44911 4156 44927 4220
rect 44991 4156 45007 4220
rect 45071 4156 45087 4220
rect 45151 4156 45167 4220
rect 45231 4156 45247 4220
rect 45311 4156 45327 4220
rect 45391 4156 45407 4220
rect 45471 4156 45487 4220
rect 45551 4156 45567 4220
rect 45631 4156 45647 4220
rect 45711 4156 45727 4220
rect 45791 4156 45807 4220
rect 45871 4156 45887 4220
rect 45951 4156 45969 4220
rect 42589 4139 45969 4156
rect 40481 4027 41272 4035
rect 40481 3818 40721 4027
rect 38639 3789 40721 3818
rect 38548 3746 40721 3789
rect 36349 3536 36448 3627
rect 38902 3578 40721 3746
rect 36349 3523 36496 3536
rect 36349 3467 36394 3523
rect 36450 3467 36496 3523
rect 36349 3454 36496 3467
rect 38555 3457 38656 3484
rect 35005 3122 35116 3144
rect 35005 3058 35031 3122
rect 35095 3113 35116 3122
rect 36359 3113 36423 3454
rect 38555 3393 38573 3457
rect 38637 3393 38656 3457
rect 38555 3377 38656 3393
rect 38555 3313 38573 3377
rect 38637 3313 38656 3377
rect 38555 3286 38656 3313
rect 40079 3451 40180 3478
rect 40079 3387 40097 3451
rect 40161 3387 40180 3451
rect 40079 3371 40180 3387
rect 40079 3307 40097 3371
rect 40161 3307 40180 3371
rect 40079 3280 40180 3307
rect 35095 3058 36423 3113
rect 35005 3049 36423 3058
rect 35005 3029 35116 3049
rect 40481 3045 40721 3578
rect 36043 2214 36151 2236
rect 36043 2150 36066 2214
rect 36130 2150 36151 2214
rect 36043 2124 36151 2150
rect 36888 1846 37150 1852
rect 36888 1765 36907 1846
rect 34644 1701 36907 1765
rect 34644 1396 34708 1701
rect 35459 1591 35583 1623
rect 36888 1622 36907 1701
rect 37131 1622 37150 1846
rect 36888 1616 37150 1622
rect 35459 1527 35489 1591
rect 35553 1527 35583 1591
rect 35459 1496 35583 1527
rect 36604 1529 36720 1558
rect 36604 1465 36631 1529
rect 36695 1465 36720 1529
rect 36604 1437 36720 1465
rect 34644 1348 35088 1396
rect 34644 1339 35098 1348
rect 34644 1332 35028 1339
rect 312 221 21117 237
rect 312 77 322 221
rect 21106 77 21117 221
rect 312 62 21117 77
rect 34644 73 34708 1332
rect 35014 1283 35028 1332
rect 35084 1283 35098 1339
rect 35014 1274 35098 1283
rect 40011 1155 40269 1195
rect 38558 1093 39142 1143
rect 38558 1037 38582 1093
rect 38638 1037 39142 1093
rect 38558 1013 39142 1037
rect 38558 957 38582 1013
rect 38638 973 39142 1013
rect 40011 1099 40112 1155
rect 40168 1099 40269 1155
rect 40011 1075 40269 1099
rect 40011 1019 40112 1075
rect 40168 1019 40269 1075
rect 40011 973 40269 1019
rect 38638 957 40721 973
rect 36007 935 36581 956
rect 36007 879 36308 935
rect 36364 879 36388 935
rect 36444 879 36468 935
rect 36524 879 36581 935
rect 38558 903 40721 957
rect 36007 860 36581 879
rect 35008 283 35127 313
rect 35008 219 35028 283
rect 35092 248 35127 283
rect 36007 248 36103 860
rect 38902 733 40721 903
rect 38558 601 38659 628
rect 38558 537 38576 601
rect 38640 537 38659 601
rect 38558 521 38659 537
rect 38558 457 38576 521
rect 38640 457 38659 521
rect 38558 430 38659 457
rect 36338 394 37077 409
rect 36338 338 36378 394
rect 36434 338 36458 394
rect 36514 393 37077 394
rect 36514 338 36987 393
rect 36338 329 36987 338
rect 37051 329 37077 393
rect 36338 313 37077 329
rect 35092 219 36103 248
rect 35008 184 36103 219
rect 35008 183 35127 184
rect 34644 19 35091 73
rect 34644 10 35101 19
rect 34644 9 35031 10
rect 34644 -1317 34708 9
rect 35017 -46 35031 9
rect 35087 -46 35101 10
rect 35017 -55 35101 -46
rect 36007 -124 36103 184
rect 36007 -140 36442 -124
rect 36007 -154 36447 -140
rect 36007 -210 36366 -154
rect 36422 -210 36447 -154
rect 38902 -175 39142 733
rect 40077 614 40178 641
rect 40077 550 40095 614
rect 40159 550 40178 614
rect 40077 534 40178 550
rect 40077 470 40095 534
rect 40159 470 40178 534
rect 40077 443 40178 470
rect 40481 230 40721 733
rect 42589 286 45940 314
rect 40481 222 41274 230
rect 40481 -2 40840 222
rect 41224 -2 41274 222
rect 42589 222 42632 286
rect 42696 222 42712 286
rect 42776 222 42792 286
rect 42856 222 42872 286
rect 42936 222 42952 286
rect 43016 222 43032 286
rect 43096 222 43112 286
rect 43176 222 43192 286
rect 43256 222 43272 286
rect 43336 222 43352 286
rect 43416 222 43432 286
rect 43496 222 43512 286
rect 43576 222 43592 286
rect 43656 222 43672 286
rect 43736 222 43752 286
rect 43816 222 43832 286
rect 43896 222 43912 286
rect 43976 222 43992 286
rect 44056 222 44072 286
rect 44136 222 44152 286
rect 44216 222 44232 286
rect 44296 222 44312 286
rect 44376 222 44392 286
rect 44456 222 44472 286
rect 44536 222 44552 286
rect 44616 222 44632 286
rect 44696 222 44712 286
rect 44776 222 44792 286
rect 44856 222 44872 286
rect 44936 222 44952 286
rect 45016 222 45032 286
rect 45096 222 45112 286
rect 45176 222 45192 286
rect 45256 222 45272 286
rect 45336 222 45352 286
rect 45416 222 45432 286
rect 45496 222 45512 286
rect 45576 222 45592 286
rect 45656 222 45672 286
rect 45736 222 45752 286
rect 45816 222 45832 286
rect 45896 222 45940 286
rect 42589 194 45940 222
rect 40481 -10 41274 -2
rect 40481 -143 40721 -10
rect 36007 -220 36447 -210
rect 36342 -224 36447 -220
rect 35000 -1055 35108 -1032
rect 35000 -1119 35027 -1055
rect 35091 -1074 35108 -1055
rect 35091 -1119 35644 -1074
rect 35000 -1138 35644 -1119
rect 35000 -1144 35108 -1138
rect 35580 -1226 35644 -1138
rect 36346 -1213 36442 -224
rect 38541 -268 39142 -175
rect 38541 -324 38582 -268
rect 38638 -324 39142 -268
rect 38541 -415 39142 -324
rect 40076 -181 40721 -143
rect 40076 -237 40104 -181
rect 40160 -237 40721 -181
rect 40076 -261 40721 -237
rect 40076 -317 40104 -261
rect 40160 -317 40721 -261
rect 40076 -383 40721 -317
rect 36961 -691 37077 -670
rect 36961 -755 36987 -691
rect 37051 -755 37077 -691
rect 36961 -776 37077 -755
rect 38553 -730 38654 -703
rect 38553 -794 38571 -730
rect 38635 -794 38654 -730
rect 38553 -810 38654 -794
rect 38553 -874 38571 -810
rect 38635 -874 38654 -810
rect 38553 -901 38654 -874
rect 35934 -1226 36442 -1213
rect 35580 -1237 36442 -1226
rect 35580 -1290 35991 -1237
rect 35934 -1293 35991 -1290
rect 36047 -1293 36071 -1237
rect 36127 -1293 36442 -1237
rect 35934 -1309 36442 -1293
rect 34644 -1373 35088 -1317
rect 34644 -1381 35098 -1373
rect 34644 -2652 34708 -1381
rect 35014 -1382 35098 -1381
rect 35014 -1438 35028 -1382
rect 35084 -1438 35098 -1382
rect 35014 -1447 35098 -1438
rect 35934 -2213 36030 -1309
rect 38902 -1545 39142 -415
rect 40082 -733 40183 -706
rect 40082 -797 40100 -733
rect 40164 -797 40183 -733
rect 40082 -813 40183 -797
rect 40082 -877 40100 -813
rect 40164 -877 40183 -813
rect 40082 -904 40183 -877
rect 40481 -1524 40721 -383
rect 47479 -1140 47735 -1135
rect 47479 -1150 62907 -1140
rect 47479 -1366 47499 -1150
rect 47715 -1366 62907 -1150
rect 47479 -1376 62907 -1366
rect 47479 -1381 47735 -1376
rect 38561 -1658 39142 -1545
rect 38561 -1714 38583 -1658
rect 38639 -1714 39142 -1658
rect 36498 -1779 37077 -1763
rect 36498 -1785 36987 -1779
rect 36498 -1841 36516 -1785
rect 36572 -1841 36596 -1785
rect 36652 -1841 36676 -1785
rect 36732 -1841 36987 -1785
rect 36498 -1843 36987 -1841
rect 37051 -1843 37077 -1779
rect 38561 -1785 39142 -1714
rect 40088 -1561 40721 -1524
rect 40088 -1617 40121 -1561
rect 40177 -1617 40721 -1561
rect 40088 -1641 40721 -1617
rect 40088 -1697 40121 -1641
rect 40177 -1697 40721 -1641
rect 40088 -1764 40721 -1697
rect 36498 -1859 37077 -1843
rect 38552 -2083 38653 -2056
rect 38552 -2147 38570 -2083
rect 38634 -2147 38653 -2083
rect 38552 -2163 38653 -2147
rect 35934 -2307 36445 -2213
rect 38552 -2227 38570 -2163
rect 38634 -2227 38653 -2163
rect 38552 -2254 38653 -2227
rect 35934 -2309 36537 -2307
rect 36349 -2328 36537 -2309
rect 36349 -2384 36368 -2328
rect 36424 -2384 36448 -2328
rect 36504 -2384 36537 -2328
rect 36349 -2403 36537 -2384
rect 35014 -2448 35119 -2424
rect 35014 -2512 35035 -2448
rect 35099 -2460 35119 -2448
rect 36349 -2460 36445 -2403
rect 35099 -2512 36445 -2460
rect 35014 -2524 36445 -2512
rect 35014 -2537 35119 -2524
rect 34644 -2716 35088 -2652
rect 35014 -2748 35088 -2716
rect 35014 -2757 35098 -2748
rect 35014 -2813 35028 -2757
rect 35084 -2813 35098 -2757
rect 35014 -2822 35098 -2813
rect 36349 -3313 36445 -2524
rect 36962 -2867 37078 -2846
rect 36962 -2931 36988 -2867
rect 37052 -2931 37078 -2867
rect 36962 -2952 37078 -2931
rect 38902 -2954 39142 -1785
rect 40082 -2105 40183 -2078
rect 40082 -2169 40100 -2105
rect 40164 -2169 40183 -2105
rect 40082 -2185 40183 -2169
rect 40082 -2249 40100 -2185
rect 40164 -2249 40183 -2185
rect 40082 -2276 40183 -2249
rect 40481 -2673 40721 -1764
rect 40481 -2681 41272 -2673
rect 38548 -3015 39142 -2954
rect 38548 -3071 38583 -3015
rect 38639 -3071 39142 -3015
rect 38548 -3095 39142 -3071
rect 38548 -3151 38583 -3095
rect 38639 -3122 39142 -3095
rect 40015 -2940 40255 -2903
rect 40015 -2996 40111 -2940
rect 40167 -2996 40255 -2940
rect 40015 -3020 40255 -2996
rect 40015 -3076 40111 -3020
rect 40167 -3076 40255 -3020
rect 40015 -3122 40255 -3076
rect 40481 -2905 40838 -2681
rect 41222 -2905 41272 -2681
rect 42577 -2720 45943 -2703
rect 42577 -2784 42588 -2720
rect 42652 -2784 42668 -2720
rect 42732 -2784 42748 -2720
rect 42812 -2784 42828 -2720
rect 42892 -2784 42908 -2720
rect 42972 -2784 42988 -2720
rect 43052 -2784 43068 -2720
rect 43132 -2784 43148 -2720
rect 43212 -2784 43228 -2720
rect 43292 -2784 43308 -2720
rect 43372 -2784 43388 -2720
rect 43452 -2784 43468 -2720
rect 43532 -2784 43548 -2720
rect 43612 -2784 43628 -2720
rect 43692 -2784 43708 -2720
rect 43772 -2784 43788 -2720
rect 43852 -2784 43868 -2720
rect 43932 -2784 43948 -2720
rect 44012 -2784 44028 -2720
rect 44092 -2784 44108 -2720
rect 44172 -2784 44188 -2720
rect 44252 -2784 44268 -2720
rect 44332 -2784 44348 -2720
rect 44412 -2784 44428 -2720
rect 44492 -2784 44508 -2720
rect 44572 -2784 44588 -2720
rect 44652 -2784 44668 -2720
rect 44732 -2784 44748 -2720
rect 44812 -2784 44828 -2720
rect 44892 -2784 44908 -2720
rect 44972 -2784 44988 -2720
rect 45052 -2784 45068 -2720
rect 45132 -2784 45148 -2720
rect 45212 -2784 45228 -2720
rect 45292 -2784 45308 -2720
rect 45372 -2784 45388 -2720
rect 45452 -2784 45468 -2720
rect 45532 -2784 45548 -2720
rect 45612 -2784 45628 -2720
rect 45692 -2784 45708 -2720
rect 45772 -2784 45788 -2720
rect 45852 -2784 45868 -2720
rect 45932 -2784 45943 -2720
rect 42577 -2801 45943 -2784
rect 40481 -2913 41272 -2905
rect 40481 -3122 40721 -2913
rect 38639 -3151 40721 -3122
rect 38548 -3194 40721 -3151
rect 36349 -3404 36448 -3313
rect 38902 -3362 40721 -3194
rect 36349 -3417 36496 -3404
rect 36349 -3473 36394 -3417
rect 36450 -3473 36496 -3417
rect 36349 -3486 36496 -3473
rect 38555 -3483 38656 -3456
rect -1926 -3573 21202 -3509
rect 21266 -3573 21276 -3509
rect 35005 -3818 35116 -3796
rect 35005 -3882 35031 -3818
rect 35095 -3827 35116 -3818
rect 36359 -3827 36423 -3486
rect 38555 -3547 38573 -3483
rect 38637 -3547 38656 -3483
rect 38555 -3563 38656 -3547
rect 38555 -3627 38573 -3563
rect 38637 -3627 38656 -3563
rect 38555 -3654 38656 -3627
rect 40079 -3489 40180 -3462
rect 40079 -3553 40097 -3489
rect 40161 -3553 40180 -3489
rect 40079 -3569 40180 -3553
rect 40079 -3633 40097 -3569
rect 40161 -3633 40180 -3569
rect 40079 -3660 40180 -3633
rect 35095 -3882 36423 -3827
rect 35005 -3891 36423 -3882
rect 35005 -3911 35116 -3891
rect 40481 -3895 40721 -3362
rect -2212 -4045 21202 -3981
rect 21266 -4045 21276 -3981
rect -2598 -4580 21202 -4516
rect 21266 -4580 21276 -4516
rect -2885 -5043 21202 -4979
rect 21266 -5043 21276 -4979
rect -3605 -6844 -3493 -6817
rect -3605 -6908 -3581 -6844
rect -3517 -6908 -3493 -6844
rect -3605 -6924 -3493 -6908
rect -3605 -6988 -3581 -6924
rect -3517 -6988 -3493 -6924
rect -3605 -7004 -3493 -6988
rect -3605 -7068 -3581 -7004
rect -3517 -7068 -3493 -7004
rect -3605 -7084 -3493 -7068
rect -3605 -7148 -3581 -7084
rect -3517 -7148 -3493 -7084
rect -3605 -7164 -3493 -7148
rect -3605 -7228 -3581 -7164
rect -3517 -7228 -3493 -7164
rect -3605 -7244 -3493 -7228
rect -3605 -7308 -3581 -7244
rect -3517 -7308 -3493 -7244
rect -3605 -7324 -3493 -7308
rect -3605 -7388 -3581 -7324
rect -3517 -7388 -3493 -7324
rect -3605 -7404 -3493 -7388
rect -3605 -7468 -3581 -7404
rect -3517 -7468 -3493 -7404
rect -3605 -7484 -3493 -7468
rect -3605 -7548 -3581 -7484
rect -3517 -7548 -3493 -7484
rect -3605 -7564 -3493 -7548
rect -3605 -7628 -3581 -7564
rect -3517 -7628 -3493 -7564
rect -3605 -7644 -3493 -7628
rect -3605 -7708 -3581 -7644
rect -3517 -7708 -3493 -7644
rect -3605 -7724 -3493 -7708
rect -3605 -7788 -3581 -7724
rect -3517 -7788 -3493 -7724
rect -3605 -7804 -3493 -7788
rect -3605 -7868 -3581 -7804
rect -3517 -7868 -3493 -7804
rect -3605 -7884 -3493 -7868
rect -3605 -7948 -3581 -7884
rect -3517 -7948 -3493 -7884
rect -3605 -7964 -3493 -7948
rect -3605 -8028 -3581 -7964
rect -3517 -8028 -3493 -7964
rect -3605 -8044 -3493 -8028
rect -3605 -8108 -3581 -8044
rect -3517 -8108 -3493 -8044
rect -3605 -8124 -3493 -8108
rect -3605 -8188 -3581 -8124
rect -3517 -8188 -3493 -8124
rect -3605 -8204 -3493 -8188
rect -3605 -8268 -3581 -8204
rect -3517 -8268 -3493 -8204
rect -3605 -8284 -3493 -8268
rect -3605 -8348 -3581 -8284
rect -3517 -8348 -3493 -8284
rect -3605 -8364 -3493 -8348
rect -3605 -8428 -3581 -8364
rect -3517 -8428 -3493 -8364
rect -3605 -8444 -3493 -8428
rect -3605 -8508 -3581 -8444
rect -3517 -8508 -3493 -8444
rect -3605 -8524 -3493 -8508
rect -3605 -8588 -3581 -8524
rect -3517 -8588 -3493 -8524
rect -3605 -8604 -3493 -8588
rect -3605 -8668 -3581 -8604
rect -3517 -8668 -3493 -8604
rect -3605 -8684 -3493 -8668
rect -3605 -8748 -3581 -8684
rect -3517 -8748 -3493 -8684
rect -3605 -8764 -3493 -8748
rect -3605 -8828 -3581 -8764
rect -3517 -8828 -3493 -8764
rect -3605 -8844 -3493 -8828
rect -3605 -8908 -3581 -8844
rect -3517 -8908 -3493 -8844
rect -3605 -8924 -3493 -8908
rect -3605 -8988 -3581 -8924
rect -3517 -8988 -3493 -8924
rect -3605 -9004 -3493 -8988
rect -3605 -9068 -3581 -9004
rect -3517 -9068 -3493 -9004
rect -3605 -9084 -3493 -9068
rect -3605 -9148 -3581 -9084
rect -3517 -9148 -3493 -9084
rect -3605 -9164 -3493 -9148
rect -3605 -9228 -3581 -9164
rect -3517 -9228 -3493 -9164
rect -3605 -9244 -3493 -9228
rect -3605 -9308 -3581 -9244
rect -3517 -9308 -3493 -9244
rect -3605 -9324 -3493 -9308
rect -3605 -9388 -3581 -9324
rect -3517 -9388 -3493 -9324
rect -3605 -9404 -3493 -9388
rect -3605 -9468 -3581 -9404
rect -3517 -9468 -3493 -9404
rect -3605 -9484 -3493 -9468
rect -3605 -9548 -3581 -9484
rect -3517 -9548 -3493 -9484
rect -3605 -9564 -3493 -9548
rect -3605 -9628 -3581 -9564
rect -3517 -9628 -3493 -9564
rect -3605 -9644 -3493 -9628
rect -3605 -9708 -3581 -9644
rect -3517 -9708 -3493 -9644
rect -3605 -9724 -3493 -9708
rect -3605 -9788 -3581 -9724
rect -3517 -9788 -3493 -9724
rect -3605 -9804 -3493 -9788
rect -3605 -9868 -3581 -9804
rect -3517 -9868 -3493 -9804
rect -3605 -9884 -3493 -9868
rect -3605 -9948 -3581 -9884
rect -3517 -9948 -3493 -9884
rect -3605 -9964 -3493 -9948
rect -3605 -10028 -3581 -9964
rect -3517 -10028 -3493 -9964
rect -3605 -10044 -3493 -10028
rect -3605 -10108 -3581 -10044
rect -3517 -10108 -3493 -10044
rect -3605 -10135 -3493 -10108
rect -610 -6851 -476 -6820
rect -610 -6915 -575 -6851
rect -511 -6915 -476 -6851
rect -610 -6931 -476 -6915
rect -610 -6995 -575 -6931
rect -511 -6995 -476 -6931
rect -610 -7011 -476 -6995
rect -610 -7075 -575 -7011
rect -511 -7075 -476 -7011
rect -610 -7091 -476 -7075
rect -610 -7155 -575 -7091
rect -511 -7155 -476 -7091
rect -610 -7171 -476 -7155
rect -610 -7235 -575 -7171
rect -511 -7235 -476 -7171
rect -610 -7251 -476 -7235
rect -610 -7315 -575 -7251
rect -511 -7315 -476 -7251
rect -610 -7331 -476 -7315
rect -610 -7395 -575 -7331
rect -511 -7395 -476 -7331
rect -610 -7411 -476 -7395
rect -610 -7475 -575 -7411
rect -511 -7475 -476 -7411
rect -610 -7491 -476 -7475
rect -610 -7555 -575 -7491
rect -511 -7555 -476 -7491
rect -610 -7571 -476 -7555
rect -610 -7635 -575 -7571
rect -511 -7635 -476 -7571
rect -610 -7651 -476 -7635
rect -610 -7715 -575 -7651
rect -511 -7715 -476 -7651
rect -610 -7731 -476 -7715
rect -610 -7795 -575 -7731
rect -511 -7795 -476 -7731
rect -610 -7811 -476 -7795
rect -610 -7875 -575 -7811
rect -511 -7875 -476 -7811
rect -610 -7891 -476 -7875
rect -610 -7955 -575 -7891
rect -511 -7955 -476 -7891
rect -610 -7971 -476 -7955
rect -610 -8035 -575 -7971
rect -511 -8035 -476 -7971
rect -610 -8051 -476 -8035
rect -610 -8115 -575 -8051
rect -511 -8115 -476 -8051
rect -610 -8131 -476 -8115
rect -610 -8195 -575 -8131
rect -511 -8195 -476 -8131
rect -610 -8211 -476 -8195
rect -610 -8275 -575 -8211
rect -511 -8275 -476 -8211
rect -610 -8291 -476 -8275
rect -610 -8355 -575 -8291
rect -511 -8355 -476 -8291
rect -610 -8371 -476 -8355
rect -610 -8435 -575 -8371
rect -511 -8435 -476 -8371
rect -610 -8451 -476 -8435
rect -610 -8515 -575 -8451
rect -511 -8515 -476 -8451
rect -610 -8531 -476 -8515
rect -610 -8595 -575 -8531
rect -511 -8595 -476 -8531
rect -610 -8611 -476 -8595
rect -610 -8675 -575 -8611
rect -511 -8675 -476 -8611
rect -610 -8691 -476 -8675
rect -610 -8755 -575 -8691
rect -511 -8755 -476 -8691
rect -610 -8771 -476 -8755
rect -610 -8835 -575 -8771
rect -511 -8835 -476 -8771
rect -610 -8851 -476 -8835
rect -610 -8915 -575 -8851
rect -511 -8915 -476 -8851
rect -610 -8931 -476 -8915
rect -610 -8995 -575 -8931
rect -511 -8995 -476 -8931
rect -610 -9011 -476 -8995
rect -610 -9075 -575 -9011
rect -511 -9075 -476 -9011
rect -610 -9091 -476 -9075
rect -610 -9155 -575 -9091
rect -511 -9155 -476 -9091
rect -610 -9171 -476 -9155
rect -610 -9235 -575 -9171
rect -511 -9235 -476 -9171
rect -610 -9251 -476 -9235
rect -610 -9315 -575 -9251
rect -511 -9315 -476 -9251
rect -610 -9331 -476 -9315
rect -610 -9395 -575 -9331
rect -511 -9395 -476 -9331
rect -610 -9411 -476 -9395
rect -610 -9475 -575 -9411
rect -511 -9475 -476 -9411
rect -610 -9491 -476 -9475
rect -610 -9555 -575 -9491
rect -511 -9555 -476 -9491
rect -610 -9571 -476 -9555
rect -610 -9635 -575 -9571
rect -511 -9635 -476 -9571
rect -610 -9651 -476 -9635
rect -610 -9715 -575 -9651
rect -511 -9715 -476 -9651
rect -610 -9731 -476 -9715
rect -610 -9795 -575 -9731
rect -511 -9795 -476 -9731
rect -610 -9811 -476 -9795
rect -610 -9875 -575 -9811
rect -511 -9875 -476 -9811
rect -610 -9891 -476 -9875
rect -610 -9955 -575 -9891
rect -511 -9955 -476 -9891
rect -610 -9971 -476 -9955
rect -610 -10035 -575 -9971
rect -511 -10035 -476 -9971
rect -610 -10051 -476 -10035
rect -610 -10115 -575 -10051
rect -511 -10115 -476 -10051
rect -610 -10145 -476 -10115
rect -2189 -12092 -1933 -12077
rect -2189 -12308 -2169 -12092
rect -1953 -12308 -1933 -12092
rect -2189 -12323 -1933 -12308
rect -2179 -18865 -1943 -12323
rect -2179 -19101 -885 -18865
rect -1121 -24022 -885 -19101
<< via3 >>
rect -16831 76688 -16767 76692
rect -16831 76632 -16827 76688
rect -16827 76632 -16771 76688
rect -16771 76632 -16767 76688
rect -16831 76628 -16767 76632
rect -16831 76608 -16767 76612
rect -16831 76552 -16827 76608
rect -16827 76552 -16771 76608
rect -16771 76552 -16767 76608
rect -16831 76548 -16767 76552
rect -16831 76528 -16767 76532
rect -16831 76472 -16827 76528
rect -16827 76472 -16771 76528
rect -16771 76472 -16767 76528
rect -16831 76468 -16767 76472
rect -16831 76448 -16767 76452
rect -16831 76392 -16827 76448
rect -16827 76392 -16771 76448
rect -16771 76392 -16767 76448
rect -16831 76388 -16767 76392
rect -16831 76368 -16767 76372
rect -16831 76312 -16827 76368
rect -16827 76312 -16771 76368
rect -16771 76312 -16767 76368
rect -16831 76308 -16767 76312
rect -16831 76288 -16767 76292
rect -16831 76232 -16827 76288
rect -16827 76232 -16771 76288
rect -16771 76232 -16767 76288
rect -16831 76228 -16767 76232
rect -16831 76208 -16767 76212
rect -16831 76152 -16827 76208
rect -16827 76152 -16771 76208
rect -16771 76152 -16767 76208
rect -16831 76148 -16767 76152
rect -16831 76128 -16767 76132
rect -16831 76072 -16827 76128
rect -16827 76072 -16771 76128
rect -16771 76072 -16767 76128
rect -16831 76068 -16767 76072
rect -16831 76048 -16767 76052
rect -16831 75992 -16827 76048
rect -16827 75992 -16771 76048
rect -16771 75992 -16767 76048
rect -16831 75988 -16767 75992
rect -16831 75968 -16767 75972
rect -16831 75912 -16827 75968
rect -16827 75912 -16771 75968
rect -16771 75912 -16767 75968
rect -16831 75908 -16767 75912
rect -16831 75888 -16767 75892
rect -16831 75832 -16827 75888
rect -16827 75832 -16771 75888
rect -16771 75832 -16767 75888
rect -16831 75828 -16767 75832
rect -16831 75808 -16767 75812
rect -16831 75752 -16827 75808
rect -16827 75752 -16771 75808
rect -16771 75752 -16767 75808
rect -16831 75748 -16767 75752
rect -16831 75728 -16767 75732
rect -16831 75672 -16827 75728
rect -16827 75672 -16771 75728
rect -16771 75672 -16767 75728
rect -16831 75668 -16767 75672
rect -16831 75648 -16767 75652
rect -16831 75592 -16827 75648
rect -16827 75592 -16771 75648
rect -16771 75592 -16767 75648
rect -16831 75588 -16767 75592
rect -16831 75568 -16767 75572
rect -16831 75512 -16827 75568
rect -16827 75512 -16771 75568
rect -16771 75512 -16767 75568
rect -16831 75508 -16767 75512
rect -16831 75488 -16767 75492
rect -16831 75432 -16827 75488
rect -16827 75432 -16771 75488
rect -16771 75432 -16767 75488
rect -16831 75428 -16767 75432
rect -16831 75408 -16767 75412
rect -16831 75352 -16827 75408
rect -16827 75352 -16771 75408
rect -16771 75352 -16767 75408
rect -16831 75348 -16767 75352
rect -16831 75328 -16767 75332
rect -16831 75272 -16827 75328
rect -16827 75272 -16771 75328
rect -16771 75272 -16767 75328
rect -16831 75268 -16767 75272
rect -16831 75248 -16767 75252
rect -16831 75192 -16827 75248
rect -16827 75192 -16771 75248
rect -16771 75192 -16767 75248
rect -16831 75188 -16767 75192
rect -16831 75168 -16767 75172
rect -16831 75112 -16827 75168
rect -16827 75112 -16771 75168
rect -16771 75112 -16767 75168
rect -16831 75108 -16767 75112
rect -16831 75088 -16767 75092
rect -16831 75032 -16827 75088
rect -16827 75032 -16771 75088
rect -16771 75032 -16767 75088
rect -16831 75028 -16767 75032
rect -16831 75008 -16767 75012
rect -16831 74952 -16827 75008
rect -16827 74952 -16771 75008
rect -16771 74952 -16767 75008
rect -16831 74948 -16767 74952
rect -16831 74928 -16767 74932
rect -16831 74872 -16827 74928
rect -16827 74872 -16771 74928
rect -16771 74872 -16767 74928
rect -16831 74868 -16767 74872
rect -16831 74848 -16767 74852
rect -16831 74792 -16827 74848
rect -16827 74792 -16771 74848
rect -16771 74792 -16767 74848
rect -16831 74788 -16767 74792
rect -16831 74768 -16767 74772
rect -16831 74712 -16827 74768
rect -16827 74712 -16771 74768
rect -16771 74712 -16767 74768
rect -16831 74708 -16767 74712
rect -16831 74688 -16767 74692
rect -16831 74632 -16827 74688
rect -16827 74632 -16771 74688
rect -16771 74632 -16767 74688
rect -16831 74628 -16767 74632
rect -16831 74608 -16767 74612
rect -16831 74552 -16827 74608
rect -16827 74552 -16771 74608
rect -16771 74552 -16767 74608
rect -16831 74548 -16767 74552
rect -16831 74528 -16767 74532
rect -16831 74472 -16827 74528
rect -16827 74472 -16771 74528
rect -16771 74472 -16767 74528
rect -16831 74468 -16767 74472
rect -16831 74448 -16767 74452
rect -16831 74392 -16827 74448
rect -16827 74392 -16771 74448
rect -16771 74392 -16767 74448
rect -16831 74388 -16767 74392
rect -16831 74368 -16767 74372
rect -16831 74312 -16827 74368
rect -16827 74312 -16771 74368
rect -16771 74312 -16767 74368
rect -16831 74308 -16767 74312
rect -16831 74288 -16767 74292
rect -16831 74232 -16827 74288
rect -16827 74232 -16771 74288
rect -16771 74232 -16767 74288
rect -16831 74228 -16767 74232
rect -16831 74208 -16767 74212
rect -16831 74152 -16827 74208
rect -16827 74152 -16771 74208
rect -16771 74152 -16767 74208
rect -16831 74148 -16767 74152
rect -16831 74128 -16767 74132
rect -16831 74072 -16827 74128
rect -16827 74072 -16771 74128
rect -16771 74072 -16767 74128
rect -16831 74068 -16767 74072
rect -16831 74048 -16767 74052
rect -16831 73992 -16827 74048
rect -16827 73992 -16771 74048
rect -16771 73992 -16767 74048
rect -16831 73988 -16767 73992
rect -16831 73968 -16767 73972
rect -16831 73912 -16827 73968
rect -16827 73912 -16771 73968
rect -16771 73912 -16767 73968
rect -16831 73908 -16767 73912
rect -16831 73888 -16767 73892
rect -16831 73832 -16827 73888
rect -16827 73832 -16771 73888
rect -16771 73832 -16767 73888
rect -16831 73828 -16767 73832
rect -16831 73808 -16767 73812
rect -16831 73752 -16827 73808
rect -16827 73752 -16771 73808
rect -16771 73752 -16767 73808
rect -16831 73748 -16767 73752
rect -16831 73728 -16767 73732
rect -16831 73672 -16827 73728
rect -16827 73672 -16771 73728
rect -16771 73672 -16767 73728
rect -16831 73668 -16767 73672
rect -16831 73648 -16767 73652
rect -16831 73592 -16827 73648
rect -16827 73592 -16771 73648
rect -16771 73592 -16767 73648
rect -16831 73588 -16767 73592
rect -16831 73568 -16767 73572
rect -16831 73512 -16827 73568
rect -16827 73512 -16771 73568
rect -16771 73512 -16767 73568
rect -16831 73508 -16767 73512
rect -16831 73488 -16767 73492
rect -16831 73432 -16827 73488
rect -16827 73432 -16771 73488
rect -16771 73432 -16767 73488
rect -16831 73428 -16767 73432
rect -13830 76694 -13766 76698
rect -13830 76638 -13826 76694
rect -13826 76638 -13770 76694
rect -13770 76638 -13766 76694
rect -13830 76634 -13766 76638
rect -13830 76614 -13766 76618
rect -13830 76558 -13826 76614
rect -13826 76558 -13770 76614
rect -13770 76558 -13766 76614
rect -13830 76554 -13766 76558
rect -13830 76534 -13766 76538
rect -13830 76478 -13826 76534
rect -13826 76478 -13770 76534
rect -13770 76478 -13766 76534
rect -13830 76474 -13766 76478
rect -13830 76454 -13766 76458
rect -13830 76398 -13826 76454
rect -13826 76398 -13770 76454
rect -13770 76398 -13766 76454
rect -13830 76394 -13766 76398
rect -13830 76374 -13766 76378
rect -13830 76318 -13826 76374
rect -13826 76318 -13770 76374
rect -13770 76318 -13766 76374
rect -13830 76314 -13766 76318
rect -13830 76294 -13766 76298
rect -13830 76238 -13826 76294
rect -13826 76238 -13770 76294
rect -13770 76238 -13766 76294
rect -13830 76234 -13766 76238
rect -13830 76214 -13766 76218
rect -13830 76158 -13826 76214
rect -13826 76158 -13770 76214
rect -13770 76158 -13766 76214
rect -13830 76154 -13766 76158
rect -13830 76134 -13766 76138
rect -13830 76078 -13826 76134
rect -13826 76078 -13770 76134
rect -13770 76078 -13766 76134
rect -13830 76074 -13766 76078
rect -13830 76054 -13766 76058
rect -13830 75998 -13826 76054
rect -13826 75998 -13770 76054
rect -13770 75998 -13766 76054
rect -13830 75994 -13766 75998
rect -13830 75974 -13766 75978
rect -13830 75918 -13826 75974
rect -13826 75918 -13770 75974
rect -13770 75918 -13766 75974
rect -13830 75914 -13766 75918
rect -13830 75894 -13766 75898
rect -13830 75838 -13826 75894
rect -13826 75838 -13770 75894
rect -13770 75838 -13766 75894
rect -13830 75834 -13766 75838
rect -13830 75814 -13766 75818
rect -13830 75758 -13826 75814
rect -13826 75758 -13770 75814
rect -13770 75758 -13766 75814
rect -13830 75754 -13766 75758
rect -13830 75734 -13766 75738
rect -13830 75678 -13826 75734
rect -13826 75678 -13770 75734
rect -13770 75678 -13766 75734
rect -13830 75674 -13766 75678
rect -13830 75654 -13766 75658
rect -13830 75598 -13826 75654
rect -13826 75598 -13770 75654
rect -13770 75598 -13766 75654
rect -13830 75594 -13766 75598
rect -13830 75574 -13766 75578
rect -13830 75518 -13826 75574
rect -13826 75518 -13770 75574
rect -13770 75518 -13766 75574
rect -13830 75514 -13766 75518
rect -13830 75494 -13766 75498
rect -13830 75438 -13826 75494
rect -13826 75438 -13770 75494
rect -13770 75438 -13766 75494
rect -13830 75434 -13766 75438
rect -13830 75414 -13766 75418
rect -13830 75358 -13826 75414
rect -13826 75358 -13770 75414
rect -13770 75358 -13766 75414
rect -13830 75354 -13766 75358
rect -13830 75334 -13766 75338
rect -13830 75278 -13826 75334
rect -13826 75278 -13770 75334
rect -13770 75278 -13766 75334
rect -13830 75274 -13766 75278
rect -13830 75254 -13766 75258
rect -13830 75198 -13826 75254
rect -13826 75198 -13770 75254
rect -13770 75198 -13766 75254
rect -13830 75194 -13766 75198
rect -13830 75174 -13766 75178
rect -13830 75118 -13826 75174
rect -13826 75118 -13770 75174
rect -13770 75118 -13766 75174
rect -13830 75114 -13766 75118
rect -13830 75094 -13766 75098
rect -13830 75038 -13826 75094
rect -13826 75038 -13770 75094
rect -13770 75038 -13766 75094
rect -13830 75034 -13766 75038
rect -13830 75014 -13766 75018
rect -13830 74958 -13826 75014
rect -13826 74958 -13770 75014
rect -13770 74958 -13766 75014
rect -13830 74954 -13766 74958
rect -13830 74934 -13766 74938
rect -13830 74878 -13826 74934
rect -13826 74878 -13770 74934
rect -13770 74878 -13766 74934
rect -13830 74874 -13766 74878
rect -13830 74854 -13766 74858
rect -13830 74798 -13826 74854
rect -13826 74798 -13770 74854
rect -13770 74798 -13766 74854
rect -13830 74794 -13766 74798
rect -13830 74774 -13766 74778
rect -13830 74718 -13826 74774
rect -13826 74718 -13770 74774
rect -13770 74718 -13766 74774
rect -13830 74714 -13766 74718
rect -13830 74694 -13766 74698
rect -13830 74638 -13826 74694
rect -13826 74638 -13770 74694
rect -13770 74638 -13766 74694
rect -13830 74634 -13766 74638
rect -13830 74614 -13766 74618
rect -13830 74558 -13826 74614
rect -13826 74558 -13770 74614
rect -13770 74558 -13766 74614
rect -13830 74554 -13766 74558
rect -13830 74534 -13766 74538
rect -13830 74478 -13826 74534
rect -13826 74478 -13770 74534
rect -13770 74478 -13766 74534
rect -13830 74474 -13766 74478
rect -13830 74454 -13766 74458
rect -13830 74398 -13826 74454
rect -13826 74398 -13770 74454
rect -13770 74398 -13766 74454
rect -13830 74394 -13766 74398
rect -13830 74374 -13766 74378
rect -13830 74318 -13826 74374
rect -13826 74318 -13770 74374
rect -13770 74318 -13766 74374
rect -13830 74314 -13766 74318
rect -13830 74294 -13766 74298
rect -13830 74238 -13826 74294
rect -13826 74238 -13770 74294
rect -13770 74238 -13766 74294
rect -13830 74234 -13766 74238
rect -13830 74214 -13766 74218
rect -13830 74158 -13826 74214
rect -13826 74158 -13770 74214
rect -13770 74158 -13766 74214
rect -13830 74154 -13766 74158
rect -13830 74134 -13766 74138
rect -13830 74078 -13826 74134
rect -13826 74078 -13770 74134
rect -13770 74078 -13766 74134
rect -13830 74074 -13766 74078
rect -13830 74054 -13766 74058
rect -13830 73998 -13826 74054
rect -13826 73998 -13770 74054
rect -13770 73998 -13766 74054
rect -13830 73994 -13766 73998
rect -13830 73974 -13766 73978
rect -13830 73918 -13826 73974
rect -13826 73918 -13770 73974
rect -13770 73918 -13766 73974
rect -13830 73914 -13766 73918
rect -13830 73894 -13766 73898
rect -13830 73838 -13826 73894
rect -13826 73838 -13770 73894
rect -13770 73838 -13766 73894
rect -13830 73834 -13766 73838
rect -13830 73814 -13766 73818
rect -13830 73758 -13826 73814
rect -13826 73758 -13770 73814
rect -13770 73758 -13766 73814
rect -13830 73754 -13766 73758
rect -13830 73734 -13766 73738
rect -13830 73678 -13826 73734
rect -13826 73678 -13770 73734
rect -13770 73678 -13766 73734
rect -13830 73674 -13766 73678
rect -13830 73654 -13766 73658
rect -13830 73598 -13826 73654
rect -13826 73598 -13770 73654
rect -13770 73598 -13766 73654
rect -13830 73594 -13766 73598
rect -13830 73574 -13766 73578
rect -13830 73518 -13826 73574
rect -13826 73518 -13770 73574
rect -13770 73518 -13766 73574
rect -13830 73514 -13766 73518
rect -13830 73494 -13766 73498
rect -13830 73438 -13826 73494
rect -13826 73438 -13770 73494
rect -13770 73438 -13766 73494
rect -13830 73434 -13766 73438
rect 11175 76674 11179 76694
rect 11179 76674 11235 76694
rect 11235 76674 11239 76694
rect 11175 76650 11239 76674
rect 11175 76630 11179 76650
rect 11179 76630 11235 76650
rect 11235 76630 11239 76650
rect 11175 76594 11179 76614
rect 11179 76594 11235 76614
rect 11235 76594 11239 76614
rect 11175 76570 11239 76594
rect 11175 76550 11179 76570
rect 11179 76550 11235 76570
rect 11235 76550 11239 76570
rect 11175 76514 11179 76534
rect 11179 76514 11235 76534
rect 11235 76514 11239 76534
rect 11175 76490 11239 76514
rect 11175 76470 11179 76490
rect 11179 76470 11235 76490
rect 11235 76470 11239 76490
rect 11175 76434 11179 76454
rect 11179 76434 11235 76454
rect 11235 76434 11239 76454
rect 11175 76410 11239 76434
rect 11175 76390 11179 76410
rect 11179 76390 11235 76410
rect 11235 76390 11239 76410
rect 11175 76354 11179 76374
rect 11179 76354 11235 76374
rect 11235 76354 11239 76374
rect 11175 76330 11239 76354
rect 11175 76310 11179 76330
rect 11179 76310 11235 76330
rect 11235 76310 11239 76330
rect 11175 76274 11179 76294
rect 11179 76274 11235 76294
rect 11235 76274 11239 76294
rect 11175 76250 11239 76274
rect 11175 76230 11179 76250
rect 11179 76230 11235 76250
rect 11235 76230 11239 76250
rect 11175 76194 11179 76214
rect 11179 76194 11235 76214
rect 11235 76194 11239 76214
rect 11175 76170 11239 76194
rect 11175 76150 11179 76170
rect 11179 76150 11235 76170
rect 11235 76150 11239 76170
rect 11175 76114 11179 76134
rect 11179 76114 11235 76134
rect 11235 76114 11239 76134
rect 11175 76090 11239 76114
rect 11175 76070 11179 76090
rect 11179 76070 11235 76090
rect 11235 76070 11239 76090
rect 11175 76034 11179 76054
rect 11179 76034 11235 76054
rect 11235 76034 11239 76054
rect 11175 76010 11239 76034
rect 11175 75990 11179 76010
rect 11179 75990 11235 76010
rect 11235 75990 11239 76010
rect 11175 75954 11179 75974
rect 11179 75954 11235 75974
rect 11235 75954 11239 75974
rect 11175 75930 11239 75954
rect 11175 75910 11179 75930
rect 11179 75910 11235 75930
rect 11235 75910 11239 75930
rect 11175 75874 11179 75894
rect 11179 75874 11235 75894
rect 11235 75874 11239 75894
rect 11175 75850 11239 75874
rect 11175 75830 11179 75850
rect 11179 75830 11235 75850
rect 11235 75830 11239 75850
rect 11175 75794 11179 75814
rect 11179 75794 11235 75814
rect 11235 75794 11239 75814
rect 11175 75770 11239 75794
rect 11175 75750 11179 75770
rect 11179 75750 11235 75770
rect 11235 75750 11239 75770
rect 11175 75714 11179 75734
rect 11179 75714 11235 75734
rect 11235 75714 11239 75734
rect 11175 75690 11239 75714
rect 11175 75670 11179 75690
rect 11179 75670 11235 75690
rect 11235 75670 11239 75690
rect 11175 75634 11179 75654
rect 11179 75634 11235 75654
rect 11235 75634 11239 75654
rect 11175 75610 11239 75634
rect 11175 75590 11179 75610
rect 11179 75590 11235 75610
rect 11235 75590 11239 75610
rect 11175 75554 11179 75574
rect 11179 75554 11235 75574
rect 11235 75554 11239 75574
rect 11175 75530 11239 75554
rect 11175 75510 11179 75530
rect 11179 75510 11235 75530
rect 11235 75510 11239 75530
rect 11175 75474 11179 75494
rect 11179 75474 11235 75494
rect 11235 75474 11239 75494
rect 11175 75450 11239 75474
rect 11175 75430 11179 75450
rect 11179 75430 11235 75450
rect 11235 75430 11239 75450
rect 11175 75394 11179 75414
rect 11179 75394 11235 75414
rect 11235 75394 11239 75414
rect 11175 75370 11239 75394
rect 11175 75350 11179 75370
rect 11179 75350 11235 75370
rect 11235 75350 11239 75370
rect 11175 75314 11179 75334
rect 11179 75314 11235 75334
rect 11235 75314 11239 75334
rect 11175 75290 11239 75314
rect 11175 75270 11179 75290
rect 11179 75270 11235 75290
rect 11235 75270 11239 75290
rect 11175 75234 11179 75254
rect 11179 75234 11235 75254
rect 11235 75234 11239 75254
rect 11175 75210 11239 75234
rect 11175 75190 11179 75210
rect 11179 75190 11235 75210
rect 11235 75190 11239 75210
rect 11175 75154 11179 75174
rect 11179 75154 11235 75174
rect 11235 75154 11239 75174
rect 11175 75130 11239 75154
rect 11175 75110 11179 75130
rect 11179 75110 11235 75130
rect 11235 75110 11239 75130
rect 11175 75074 11179 75094
rect 11179 75074 11235 75094
rect 11235 75074 11239 75094
rect 11175 75050 11239 75074
rect 11175 75030 11179 75050
rect 11179 75030 11235 75050
rect 11235 75030 11239 75050
rect 11175 74994 11179 75014
rect 11179 74994 11235 75014
rect 11235 74994 11239 75014
rect 11175 74970 11239 74994
rect 11175 74950 11179 74970
rect 11179 74950 11235 74970
rect 11235 74950 11239 74970
rect 11175 74914 11179 74934
rect 11179 74914 11235 74934
rect 11235 74914 11239 74934
rect 11175 74890 11239 74914
rect 11175 74870 11179 74890
rect 11179 74870 11235 74890
rect 11235 74870 11239 74890
rect 11175 74834 11179 74854
rect 11179 74834 11235 74854
rect 11235 74834 11239 74854
rect 11175 74810 11239 74834
rect 11175 74790 11179 74810
rect 11179 74790 11235 74810
rect 11235 74790 11239 74810
rect 11175 74754 11179 74774
rect 11179 74754 11235 74774
rect 11235 74754 11239 74774
rect 11175 74730 11239 74754
rect 11175 74710 11179 74730
rect 11179 74710 11235 74730
rect 11235 74710 11239 74730
rect 11175 74674 11179 74694
rect 11179 74674 11235 74694
rect 11235 74674 11239 74694
rect 11175 74650 11239 74674
rect 11175 74630 11179 74650
rect 11179 74630 11235 74650
rect 11235 74630 11239 74650
rect 11175 74594 11179 74614
rect 11179 74594 11235 74614
rect 11235 74594 11239 74614
rect 11175 74570 11239 74594
rect 11175 74550 11179 74570
rect 11179 74550 11235 74570
rect 11235 74550 11239 74570
rect 11175 74514 11179 74534
rect 11179 74514 11235 74534
rect 11235 74514 11239 74534
rect 11175 74490 11239 74514
rect 11175 74470 11179 74490
rect 11179 74470 11235 74490
rect 11235 74470 11239 74490
rect 11175 74434 11179 74454
rect 11179 74434 11235 74454
rect 11235 74434 11239 74454
rect 11175 74410 11239 74434
rect 11175 74390 11179 74410
rect 11179 74390 11235 74410
rect 11235 74390 11239 74410
rect 11175 74354 11179 74374
rect 11179 74354 11235 74374
rect 11235 74354 11239 74374
rect 11175 74330 11239 74354
rect 11175 74310 11179 74330
rect 11179 74310 11235 74330
rect 11235 74310 11239 74330
rect 11175 74274 11179 74294
rect 11179 74274 11235 74294
rect 11235 74274 11239 74294
rect 11175 74250 11239 74274
rect 11175 74230 11179 74250
rect 11179 74230 11235 74250
rect 11235 74230 11239 74250
rect 11175 74194 11179 74214
rect 11179 74194 11235 74214
rect 11235 74194 11239 74214
rect 11175 74170 11239 74194
rect 11175 74150 11179 74170
rect 11179 74150 11235 74170
rect 11235 74150 11239 74170
rect 11175 74114 11179 74134
rect 11179 74114 11235 74134
rect 11235 74114 11239 74134
rect 11175 74090 11239 74114
rect 11175 74070 11179 74090
rect 11179 74070 11235 74090
rect 11235 74070 11239 74090
rect 11175 74034 11179 74054
rect 11179 74034 11235 74054
rect 11235 74034 11239 74054
rect 11175 74010 11239 74034
rect 11175 73990 11179 74010
rect 11179 73990 11235 74010
rect 11235 73990 11239 74010
rect 11175 73954 11179 73974
rect 11179 73954 11235 73974
rect 11235 73954 11239 73974
rect 11175 73930 11239 73954
rect 11175 73910 11179 73930
rect 11179 73910 11235 73930
rect 11235 73910 11239 73930
rect 11175 73874 11179 73894
rect 11179 73874 11235 73894
rect 11235 73874 11239 73894
rect 11175 73850 11239 73874
rect 11175 73830 11179 73850
rect 11179 73830 11235 73850
rect 11235 73830 11239 73850
rect 11175 73794 11179 73814
rect 11179 73794 11235 73814
rect 11235 73794 11239 73814
rect 11175 73770 11239 73794
rect 11175 73750 11179 73770
rect 11179 73750 11235 73770
rect 11235 73750 11239 73770
rect 11175 73714 11179 73734
rect 11179 73714 11235 73734
rect 11235 73714 11239 73734
rect 11175 73690 11239 73714
rect 11175 73670 11179 73690
rect 11179 73670 11235 73690
rect 11235 73670 11239 73690
rect 11175 73634 11179 73654
rect 11179 73634 11235 73654
rect 11235 73634 11239 73654
rect 11175 73610 11239 73634
rect 11175 73590 11179 73610
rect 11179 73590 11235 73610
rect 11235 73590 11239 73610
rect 11175 73554 11179 73574
rect 11179 73554 11235 73574
rect 11235 73554 11239 73574
rect 11175 73530 11239 73554
rect 11175 73510 11179 73530
rect 11179 73510 11235 73530
rect 11235 73510 11239 73530
rect 11175 73474 11179 73494
rect 11179 73474 11235 73494
rect 11235 73474 11239 73494
rect 11175 73450 11239 73474
rect 11175 73430 11179 73450
rect 11179 73430 11235 73450
rect 11235 73430 11239 73450
rect 14176 76687 14180 76707
rect 14180 76687 14236 76707
rect 14236 76687 14240 76707
rect 14176 76663 14240 76687
rect 14176 76643 14180 76663
rect 14180 76643 14236 76663
rect 14236 76643 14240 76663
rect 14176 76607 14180 76627
rect 14180 76607 14236 76627
rect 14236 76607 14240 76627
rect 14176 76583 14240 76607
rect 14176 76563 14180 76583
rect 14180 76563 14236 76583
rect 14236 76563 14240 76583
rect 14176 76527 14180 76547
rect 14180 76527 14236 76547
rect 14236 76527 14240 76547
rect 14176 76503 14240 76527
rect 14176 76483 14180 76503
rect 14180 76483 14236 76503
rect 14236 76483 14240 76503
rect 14176 76447 14180 76467
rect 14180 76447 14236 76467
rect 14236 76447 14240 76467
rect 14176 76423 14240 76447
rect 14176 76403 14180 76423
rect 14180 76403 14236 76423
rect 14236 76403 14240 76423
rect 14176 76367 14180 76387
rect 14180 76367 14236 76387
rect 14236 76367 14240 76387
rect 14176 76343 14240 76367
rect 14176 76323 14180 76343
rect 14180 76323 14236 76343
rect 14236 76323 14240 76343
rect 14176 76287 14180 76307
rect 14180 76287 14236 76307
rect 14236 76287 14240 76307
rect 14176 76263 14240 76287
rect 14176 76243 14180 76263
rect 14180 76243 14236 76263
rect 14236 76243 14240 76263
rect 14176 76207 14180 76227
rect 14180 76207 14236 76227
rect 14236 76207 14240 76227
rect 14176 76183 14240 76207
rect 14176 76163 14180 76183
rect 14180 76163 14236 76183
rect 14236 76163 14240 76183
rect 14176 76127 14180 76147
rect 14180 76127 14236 76147
rect 14236 76127 14240 76147
rect 14176 76103 14240 76127
rect 14176 76083 14180 76103
rect 14180 76083 14236 76103
rect 14236 76083 14240 76103
rect 14176 76047 14180 76067
rect 14180 76047 14236 76067
rect 14236 76047 14240 76067
rect 14176 76023 14240 76047
rect 14176 76003 14180 76023
rect 14180 76003 14236 76023
rect 14236 76003 14240 76023
rect 14176 75967 14180 75987
rect 14180 75967 14236 75987
rect 14236 75967 14240 75987
rect 14176 75943 14240 75967
rect 14176 75923 14180 75943
rect 14180 75923 14236 75943
rect 14236 75923 14240 75943
rect 14176 75887 14180 75907
rect 14180 75887 14236 75907
rect 14236 75887 14240 75907
rect 14176 75863 14240 75887
rect 14176 75843 14180 75863
rect 14180 75843 14236 75863
rect 14236 75843 14240 75863
rect 14176 75807 14180 75827
rect 14180 75807 14236 75827
rect 14236 75807 14240 75827
rect 14176 75783 14240 75807
rect 14176 75763 14180 75783
rect 14180 75763 14236 75783
rect 14236 75763 14240 75783
rect 14176 75727 14180 75747
rect 14180 75727 14236 75747
rect 14236 75727 14240 75747
rect 14176 75703 14240 75727
rect 14176 75683 14180 75703
rect 14180 75683 14236 75703
rect 14236 75683 14240 75703
rect 14176 75647 14180 75667
rect 14180 75647 14236 75667
rect 14236 75647 14240 75667
rect 14176 75623 14240 75647
rect 14176 75603 14180 75623
rect 14180 75603 14236 75623
rect 14236 75603 14240 75623
rect 14176 75567 14180 75587
rect 14180 75567 14236 75587
rect 14236 75567 14240 75587
rect 14176 75543 14240 75567
rect 14176 75523 14180 75543
rect 14180 75523 14236 75543
rect 14236 75523 14240 75543
rect 14176 75487 14180 75507
rect 14180 75487 14236 75507
rect 14236 75487 14240 75507
rect 14176 75463 14240 75487
rect 14176 75443 14180 75463
rect 14180 75443 14236 75463
rect 14236 75443 14240 75463
rect 14176 75407 14180 75427
rect 14180 75407 14236 75427
rect 14236 75407 14240 75427
rect 14176 75383 14240 75407
rect 14176 75363 14180 75383
rect 14180 75363 14236 75383
rect 14236 75363 14240 75383
rect 14176 75327 14180 75347
rect 14180 75327 14236 75347
rect 14236 75327 14240 75347
rect 14176 75303 14240 75327
rect 14176 75283 14180 75303
rect 14180 75283 14236 75303
rect 14236 75283 14240 75303
rect 14176 75247 14180 75267
rect 14180 75247 14236 75267
rect 14236 75247 14240 75267
rect 14176 75223 14240 75247
rect 14176 75203 14180 75223
rect 14180 75203 14236 75223
rect 14236 75203 14240 75223
rect 14176 75167 14180 75187
rect 14180 75167 14236 75187
rect 14236 75167 14240 75187
rect 14176 75143 14240 75167
rect 14176 75123 14180 75143
rect 14180 75123 14236 75143
rect 14236 75123 14240 75143
rect 14176 75087 14180 75107
rect 14180 75087 14236 75107
rect 14236 75087 14240 75107
rect 14176 75063 14240 75087
rect 14176 75043 14180 75063
rect 14180 75043 14236 75063
rect 14236 75043 14240 75063
rect 14176 75007 14180 75027
rect 14180 75007 14236 75027
rect 14236 75007 14240 75027
rect 14176 74983 14240 75007
rect 14176 74963 14180 74983
rect 14180 74963 14236 74983
rect 14236 74963 14240 74983
rect 14176 74927 14180 74947
rect 14180 74927 14236 74947
rect 14236 74927 14240 74947
rect 14176 74903 14240 74927
rect 14176 74883 14180 74903
rect 14180 74883 14236 74903
rect 14236 74883 14240 74903
rect 14176 74847 14180 74867
rect 14180 74847 14236 74867
rect 14236 74847 14240 74867
rect 14176 74823 14240 74847
rect 14176 74803 14180 74823
rect 14180 74803 14236 74823
rect 14236 74803 14240 74823
rect 14176 74767 14180 74787
rect 14180 74767 14236 74787
rect 14236 74767 14240 74787
rect 14176 74743 14240 74767
rect 14176 74723 14180 74743
rect 14180 74723 14236 74743
rect 14236 74723 14240 74743
rect 14176 74687 14180 74707
rect 14180 74687 14236 74707
rect 14236 74687 14240 74707
rect 14176 74663 14240 74687
rect 14176 74643 14180 74663
rect 14180 74643 14236 74663
rect 14236 74643 14240 74663
rect 14176 74607 14180 74627
rect 14180 74607 14236 74627
rect 14236 74607 14240 74627
rect 14176 74583 14240 74607
rect 14176 74563 14180 74583
rect 14180 74563 14236 74583
rect 14236 74563 14240 74583
rect 14176 74527 14180 74547
rect 14180 74527 14236 74547
rect 14236 74527 14240 74547
rect 14176 74503 14240 74527
rect 14176 74483 14180 74503
rect 14180 74483 14236 74503
rect 14236 74483 14240 74503
rect 14176 74447 14180 74467
rect 14180 74447 14236 74467
rect 14236 74447 14240 74467
rect 14176 74423 14240 74447
rect 14176 74403 14180 74423
rect 14180 74403 14236 74423
rect 14236 74403 14240 74423
rect 14176 74367 14180 74387
rect 14180 74367 14236 74387
rect 14236 74367 14240 74387
rect 14176 74343 14240 74367
rect 14176 74323 14180 74343
rect 14180 74323 14236 74343
rect 14236 74323 14240 74343
rect 14176 74287 14180 74307
rect 14180 74287 14236 74307
rect 14236 74287 14240 74307
rect 14176 74263 14240 74287
rect 14176 74243 14180 74263
rect 14180 74243 14236 74263
rect 14236 74243 14240 74263
rect 14176 74207 14180 74227
rect 14180 74207 14236 74227
rect 14236 74207 14240 74227
rect 14176 74183 14240 74207
rect 14176 74163 14180 74183
rect 14180 74163 14236 74183
rect 14236 74163 14240 74183
rect 14176 74127 14180 74147
rect 14180 74127 14236 74147
rect 14236 74127 14240 74147
rect 14176 74103 14240 74127
rect 14176 74083 14180 74103
rect 14180 74083 14236 74103
rect 14236 74083 14240 74103
rect 14176 74047 14180 74067
rect 14180 74047 14236 74067
rect 14236 74047 14240 74067
rect 14176 74023 14240 74047
rect 14176 74003 14180 74023
rect 14180 74003 14236 74023
rect 14236 74003 14240 74023
rect 14176 73967 14180 73987
rect 14180 73967 14236 73987
rect 14236 73967 14240 73987
rect 14176 73943 14240 73967
rect 14176 73923 14180 73943
rect 14180 73923 14236 73943
rect 14236 73923 14240 73943
rect 14176 73887 14180 73907
rect 14180 73887 14236 73907
rect 14236 73887 14240 73907
rect 14176 73863 14240 73887
rect 14176 73843 14180 73863
rect 14180 73843 14236 73863
rect 14236 73843 14240 73863
rect 14176 73807 14180 73827
rect 14180 73807 14236 73827
rect 14236 73807 14240 73827
rect 14176 73783 14240 73807
rect 14176 73763 14180 73783
rect 14180 73763 14236 73783
rect 14236 73763 14240 73783
rect 14176 73727 14180 73747
rect 14180 73727 14236 73747
rect 14236 73727 14240 73747
rect 14176 73703 14240 73727
rect 14176 73683 14180 73703
rect 14180 73683 14236 73703
rect 14236 73683 14240 73703
rect 14176 73647 14180 73667
rect 14180 73647 14236 73667
rect 14236 73647 14240 73667
rect 14176 73623 14240 73647
rect 14176 73603 14180 73623
rect 14180 73603 14236 73623
rect 14236 73603 14240 73623
rect 14176 73567 14180 73587
rect 14180 73567 14236 73587
rect 14236 73567 14240 73587
rect 14176 73543 14240 73567
rect 14176 73523 14180 73543
rect 14180 73523 14236 73543
rect 14236 73523 14240 73543
rect 14176 73487 14180 73507
rect 14180 73487 14236 73507
rect 14236 73487 14240 73507
rect 14176 73463 14240 73487
rect 14176 73443 14180 73463
rect 14180 73443 14236 73463
rect 14236 73443 14240 73463
rect -16664 71798 -16600 71802
rect -16664 71742 -16660 71798
rect -16660 71742 -16604 71798
rect -16604 71742 -16600 71798
rect -16664 71738 -16600 71742
rect -15486 71794 -15422 71798
rect -15486 71738 -15482 71794
rect -15482 71738 -15426 71794
rect -15426 71738 -15422 71794
rect -15486 71734 -15422 71738
rect -15269 71801 -15205 71805
rect -15269 71745 -15265 71801
rect -15265 71745 -15209 71801
rect -15209 71745 -15205 71801
rect -15269 71741 -15205 71745
rect -14135 71798 -14071 71802
rect -14135 71742 -14131 71798
rect -14131 71742 -14075 71798
rect -14075 71742 -14071 71798
rect -14135 71738 -14071 71742
rect -16554 70294 -16490 70298
rect -16554 70238 -16550 70294
rect -16550 70238 -16494 70294
rect -16494 70238 -16490 70294
rect -16554 70234 -16490 70238
rect -15440 70280 -15376 70284
rect -15440 70224 -15436 70280
rect -15436 70224 -15380 70280
rect -15380 70224 -15376 70280
rect -15440 70220 -15376 70224
rect -15227 70281 -15163 70285
rect -15227 70225 -15223 70281
rect -15223 70225 -15167 70281
rect -15167 70225 -15163 70281
rect -15227 70221 -15163 70225
rect -14063 70281 -13999 70285
rect -14063 70225 -14059 70281
rect -14059 70225 -14003 70281
rect -14003 70225 -13999 70281
rect -14063 70221 -13999 70225
rect 36631 69270 36695 69334
rect 36066 68677 36130 68741
rect -15422 68488 -15358 68492
rect -15422 68432 -15418 68488
rect -15418 68432 -15362 68488
rect -15362 68432 -15358 68488
rect -15422 68428 -15358 68432
rect -15422 68408 -15358 68412
rect -15422 68352 -15418 68408
rect -15418 68352 -15362 68408
rect -15362 68352 -15358 68408
rect -15422 68348 -15358 68352
rect -15422 68328 -15358 68332
rect -15422 68272 -15418 68328
rect -15418 68272 -15362 68328
rect -15362 68272 -15358 68328
rect -15422 68268 -15358 68272
rect -15959 68251 -15895 68255
rect -15959 68195 -15955 68251
rect -15955 68195 -15899 68251
rect -15899 68195 -15895 68251
rect -15959 68191 -15895 68195
rect -15959 68171 -15895 68175
rect -15959 68115 -15955 68171
rect -15955 68115 -15899 68171
rect -15899 68115 -15895 68171
rect -15959 68111 -15895 68115
rect -15422 68248 -15358 68252
rect -15422 68192 -15418 68248
rect -15418 68192 -15362 68248
rect -15362 68192 -15358 68248
rect -15422 68188 -15358 68192
rect -14875 68254 -14811 68258
rect -14875 68198 -14871 68254
rect -14871 68198 -14815 68254
rect -14815 68198 -14811 68254
rect -14875 68194 -14811 68198
rect -14875 68174 -14811 68178
rect -14875 68118 -14871 68174
rect -14871 68118 -14815 68174
rect -14815 68118 -14811 68174
rect -14875 68114 -14811 68118
rect 35477 68017 35541 68081
rect -16577 67609 -16513 67613
rect -16577 67553 -16573 67609
rect -16573 67553 -16517 67609
rect -16517 67553 -16513 67609
rect -16577 67549 -16513 67553
rect -15422 67603 -15358 67607
rect -15422 67547 -15418 67603
rect -15418 67547 -15362 67603
rect -15362 67547 -15358 67603
rect -15422 67543 -15358 67547
rect -14304 67614 -14240 67618
rect -14304 67558 -14300 67614
rect -14300 67558 -14244 67614
rect -14244 67558 -14240 67614
rect -14304 67554 -14240 67558
rect -13096 66705 -13032 66769
rect -8073 66705 -8009 66769
rect -12315 66382 -12251 66446
rect -7266 66382 -7202 66446
rect -11305 65949 -11241 66013
rect -2673 65949 -2609 66013
rect -10536 65696 -10472 65760
rect -1866 65696 -1802 65760
rect -8073 65265 -8009 65329
rect -2673 65265 -2609 65329
rect -7266 65012 -7202 65076
rect -1866 65012 -1802 65076
rect 17431 64724 17495 64728
rect 17431 64668 17435 64724
rect 17435 64668 17491 64724
rect 17491 64668 17495 64724
rect 17431 64664 17495 64668
rect 17431 64644 17495 64648
rect 17431 64588 17435 64644
rect 17435 64588 17491 64644
rect 17491 64588 17495 64644
rect 17431 64584 17495 64588
rect 17431 64564 17495 64568
rect 17431 64508 17435 64564
rect 17435 64508 17491 64564
rect 17491 64508 17495 64564
rect 17431 64504 17495 64508
rect 17431 64484 17495 64488
rect 17431 64428 17435 64484
rect 17435 64428 17491 64484
rect 17491 64428 17495 64484
rect 17431 64424 17495 64428
rect 17431 64404 17495 64408
rect 17431 64348 17435 64404
rect 17435 64348 17491 64404
rect 17491 64348 17495 64404
rect 17431 64344 17495 64348
rect 17431 64324 17495 64328
rect 17431 64268 17435 64324
rect 17435 64268 17491 64324
rect 17491 64268 17495 64324
rect 17431 64264 17495 64268
rect 17431 64244 17495 64248
rect 17431 64188 17435 64244
rect 17435 64188 17491 64244
rect 17491 64188 17495 64244
rect 17431 64184 17495 64188
rect 23959 64724 24023 64728
rect 23959 64668 23963 64724
rect 23963 64668 24019 64724
rect 24019 64668 24023 64724
rect 23959 64664 24023 64668
rect 23959 64644 24023 64648
rect 23959 64588 23963 64644
rect 23963 64588 24019 64644
rect 24019 64588 24023 64644
rect 23959 64584 24023 64588
rect 23959 64564 24023 64568
rect 23959 64508 23963 64564
rect 23963 64508 24019 64564
rect 24019 64508 24023 64564
rect 23959 64504 24023 64508
rect 23959 64484 24023 64488
rect 23959 64428 23963 64484
rect 23963 64428 24019 64484
rect 24019 64428 24023 64484
rect 23959 64424 24023 64428
rect 23959 64404 24023 64408
rect 23959 64348 23963 64404
rect 23963 64348 24019 64404
rect 24019 64348 24023 64404
rect 23959 64344 24023 64348
rect 23959 64324 24023 64328
rect 23959 64268 23963 64324
rect 23963 64268 24019 64324
rect 24019 64268 24023 64324
rect 23959 64264 24023 64268
rect 23959 64244 24023 64248
rect 23959 64188 23963 64244
rect 23963 64188 24019 64244
rect 24019 64188 24023 64244
rect 23959 64184 24023 64188
rect 31575 64724 31639 64728
rect 31575 64668 31579 64724
rect 31579 64668 31635 64724
rect 31635 64668 31639 64724
rect 31575 64664 31639 64668
rect 31575 64644 31639 64648
rect 31575 64588 31579 64644
rect 31579 64588 31635 64644
rect 31635 64588 31639 64644
rect 31575 64584 31639 64588
rect 31575 64564 31639 64568
rect 31575 64508 31579 64564
rect 31579 64508 31635 64564
rect 31635 64508 31639 64564
rect 31575 64504 31639 64508
rect 31575 64484 31639 64488
rect 31575 64428 31579 64484
rect 31579 64428 31635 64484
rect 31635 64428 31639 64484
rect 31575 64424 31639 64428
rect 31575 64404 31639 64408
rect 31575 64348 31579 64404
rect 31579 64348 31635 64404
rect 31635 64348 31639 64404
rect 31575 64344 31639 64348
rect 31575 64324 31639 64328
rect 31575 64268 31579 64324
rect 31579 64268 31635 64324
rect 31635 64268 31639 64324
rect 31575 64264 31639 64268
rect 31575 64244 31639 64248
rect 31575 64188 31579 64244
rect 31579 64188 31635 64244
rect 31635 64188 31639 64244
rect 31575 64184 31639 64188
rect -11056 63229 -10752 63533
rect -10187 63338 -10123 63402
rect -9855 63398 -9791 63402
rect -9855 63342 -9851 63398
rect -9851 63342 -9795 63398
rect -9795 63342 -9791 63398
rect -9855 63338 -9791 63342
rect -9775 63398 -9711 63402
rect -9775 63342 -9771 63398
rect -9771 63342 -9715 63398
rect -9715 63342 -9711 63398
rect -9775 63338 -9711 63342
rect -9695 63398 -9631 63402
rect -9695 63342 -9691 63398
rect -9691 63342 -9635 63398
rect -9635 63342 -9631 63398
rect -9695 63338 -9631 63342
rect -9615 63398 -9551 63402
rect -9615 63342 -9611 63398
rect -9611 63342 -9555 63398
rect -9555 63342 -9551 63398
rect -9615 63338 -9551 63342
rect -9535 63398 -9471 63402
rect -9535 63342 -9531 63398
rect -9531 63342 -9475 63398
rect -9475 63342 -9471 63398
rect -9535 63338 -9471 63342
rect -8044 63400 -7980 63404
rect -8044 63344 -8040 63400
rect -8040 63344 -7984 63400
rect -7984 63344 -7980 63400
rect -8044 63340 -7980 63344
rect -7964 63400 -7900 63404
rect -7964 63344 -7960 63400
rect -7960 63344 -7904 63400
rect -7904 63344 -7900 63400
rect -7964 63340 -7900 63344
rect -7884 63400 -7820 63404
rect -7884 63344 -7880 63400
rect -7880 63344 -7824 63400
rect -7824 63344 -7820 63400
rect -7884 63340 -7820 63344
rect -7804 63400 -7740 63404
rect -7804 63344 -7800 63400
rect -7800 63344 -7744 63400
rect -7744 63344 -7740 63400
rect -7804 63340 -7740 63344
rect -7724 63400 -7660 63404
rect -7724 63344 -7720 63400
rect -7720 63344 -7664 63400
rect -7664 63344 -7660 63400
rect -7724 63340 -7660 63344
rect -6249 63396 -6185 63400
rect -6249 63340 -6245 63396
rect -6245 63340 -6189 63396
rect -6189 63340 -6185 63396
rect -6249 63336 -6185 63340
rect -6169 63396 -6105 63400
rect -6169 63340 -6165 63396
rect -6165 63340 -6109 63396
rect -6109 63340 -6105 63396
rect -6169 63336 -6105 63340
rect -6089 63396 -6025 63400
rect -6089 63340 -6085 63396
rect -6085 63340 -6029 63396
rect -6029 63340 -6025 63396
rect -6089 63336 -6025 63340
rect -6009 63396 -5945 63400
rect -6009 63340 -6005 63396
rect -6005 63340 -5949 63396
rect -5949 63340 -5945 63396
rect -6009 63336 -5945 63340
rect -5929 63396 -5865 63400
rect -5929 63340 -5925 63396
rect -5925 63340 -5869 63396
rect -5869 63340 -5865 63396
rect -5929 63336 -5865 63340
rect -4450 63394 -4386 63398
rect -4450 63338 -4446 63394
rect -4446 63338 -4390 63394
rect -4390 63338 -4386 63394
rect -4450 63334 -4386 63338
rect -4370 63394 -4306 63398
rect -4370 63338 -4366 63394
rect -4366 63338 -4310 63394
rect -4310 63338 -4306 63394
rect -4370 63334 -4306 63338
rect -4290 63394 -4226 63398
rect -4290 63338 -4286 63394
rect -4286 63338 -4230 63394
rect -4230 63338 -4226 63394
rect -4290 63334 -4226 63338
rect -4210 63394 -4146 63398
rect -4210 63338 -4206 63394
rect -4206 63338 -4150 63394
rect -4150 63338 -4146 63394
rect -4210 63334 -4146 63338
rect -4130 63394 -4066 63398
rect -4130 63338 -4126 63394
rect -4126 63338 -4070 63394
rect -4070 63338 -4066 63394
rect -4130 63334 -4066 63338
rect -2659 63398 -2595 63402
rect -2659 63342 -2655 63398
rect -2655 63342 -2599 63398
rect -2599 63342 -2595 63398
rect -2659 63338 -2595 63342
rect -2579 63398 -2515 63402
rect -2579 63342 -2575 63398
rect -2575 63342 -2519 63398
rect -2519 63342 -2515 63398
rect -2579 63338 -2515 63342
rect -2499 63398 -2435 63402
rect -2499 63342 -2495 63398
rect -2495 63342 -2439 63398
rect -2439 63342 -2435 63398
rect -2499 63338 -2435 63342
rect -2419 63398 -2355 63402
rect -2419 63342 -2415 63398
rect -2415 63342 -2359 63398
rect -2359 63342 -2355 63398
rect -2419 63338 -2355 63342
rect -2339 63398 -2275 63402
rect -2339 63342 -2335 63398
rect -2335 63342 -2279 63398
rect -2279 63342 -2275 63398
rect -2339 63338 -2275 63342
rect -857 63394 -793 63398
rect -857 63338 -853 63394
rect -853 63338 -797 63394
rect -797 63338 -793 63394
rect -857 63334 -793 63338
rect -777 63394 -713 63398
rect -777 63338 -773 63394
rect -773 63338 -717 63394
rect -717 63338 -713 63394
rect -777 63334 -713 63338
rect -697 63394 -633 63398
rect -697 63338 -693 63394
rect -693 63338 -637 63394
rect -637 63338 -633 63394
rect -697 63334 -633 63338
rect -617 63394 -553 63398
rect -617 63338 -613 63394
rect -613 63338 -557 63394
rect -557 63338 -553 63394
rect -617 63334 -553 63338
rect -537 63394 -473 63398
rect -537 63338 -533 63394
rect -533 63338 -477 63394
rect -477 63338 -473 63394
rect -537 63334 -473 63338
rect -6931 63194 -6707 63198
rect -6931 62978 -6927 63194
rect -6927 62978 -6711 63194
rect -6711 62978 -6707 63194
rect -6931 62974 -6707 62978
rect 790 63220 1254 63224
rect 790 63004 794 63220
rect 794 63004 1250 63220
rect 1250 63004 1254 63220
rect 790 63000 1254 63004
rect 17976 62721 18040 62725
rect 17976 62665 17980 62721
rect 17980 62665 18036 62721
rect 18036 62665 18040 62721
rect 17976 62661 18040 62665
rect 17976 62641 18040 62645
rect 17976 62585 17980 62641
rect 17980 62585 18036 62641
rect 18036 62585 18040 62641
rect 17976 62581 18040 62585
rect 17976 62561 18040 62565
rect 17976 62505 17980 62561
rect 17980 62505 18036 62561
rect 18036 62505 18040 62561
rect 17976 62501 18040 62505
rect 17976 62481 18040 62485
rect 17976 62425 17980 62481
rect 17980 62425 18036 62481
rect 18036 62425 18040 62481
rect 17976 62421 18040 62425
rect 17976 62401 18040 62405
rect 17976 62345 17980 62401
rect 17980 62345 18036 62401
rect 18036 62345 18040 62401
rect 17976 62341 18040 62345
rect 17976 62321 18040 62325
rect 17976 62265 17980 62321
rect 17980 62265 18036 62321
rect 18036 62265 18040 62321
rect 17976 62261 18040 62265
rect 17976 62241 18040 62245
rect 17976 62185 17980 62241
rect 17980 62185 18036 62241
rect 18036 62185 18040 62241
rect 17976 62181 18040 62185
rect 19064 62721 19128 62725
rect 19064 62665 19068 62721
rect 19068 62665 19124 62721
rect 19124 62665 19128 62721
rect 19064 62661 19128 62665
rect 19064 62641 19128 62645
rect 19064 62585 19068 62641
rect 19068 62585 19124 62641
rect 19124 62585 19128 62641
rect 19064 62581 19128 62585
rect 19064 62561 19128 62565
rect 19064 62505 19068 62561
rect 19068 62505 19124 62561
rect 19124 62505 19128 62561
rect 19064 62501 19128 62505
rect 19064 62481 19128 62485
rect 19064 62425 19068 62481
rect 19068 62425 19124 62481
rect 19124 62425 19128 62481
rect 19064 62421 19128 62425
rect 19064 62401 19128 62405
rect 19064 62345 19068 62401
rect 19068 62345 19124 62401
rect 19124 62345 19128 62401
rect 19064 62341 19128 62345
rect 19064 62321 19128 62325
rect 19064 62265 19068 62321
rect 19068 62265 19124 62321
rect 19124 62265 19128 62321
rect 19064 62261 19128 62265
rect 19064 62241 19128 62245
rect 19064 62185 19068 62241
rect 19068 62185 19124 62241
rect 19124 62185 19128 62241
rect 19064 62181 19128 62185
rect 21240 62721 21304 62725
rect 21240 62665 21244 62721
rect 21244 62665 21300 62721
rect 21300 62665 21304 62721
rect 21240 62661 21304 62665
rect 21240 62641 21304 62645
rect 21240 62585 21244 62641
rect 21244 62585 21300 62641
rect 21300 62585 21304 62641
rect 21240 62581 21304 62585
rect 21240 62561 21304 62565
rect 21240 62505 21244 62561
rect 21244 62505 21300 62561
rect 21300 62505 21304 62561
rect 21240 62501 21304 62505
rect 21240 62481 21304 62485
rect 21240 62425 21244 62481
rect 21244 62425 21300 62481
rect 21300 62425 21304 62481
rect 21240 62421 21304 62425
rect 21240 62401 21304 62405
rect 21240 62345 21244 62401
rect 21244 62345 21300 62401
rect 21300 62345 21304 62401
rect 21240 62341 21304 62345
rect 21240 62321 21304 62325
rect 21240 62265 21244 62321
rect 21244 62265 21300 62321
rect 21300 62265 21304 62321
rect 21240 62261 21304 62265
rect 21240 62241 21304 62245
rect 21240 62185 21244 62241
rect 21244 62185 21300 62241
rect 21300 62185 21304 62241
rect 21240 62181 21304 62185
rect 22328 62721 22392 62725
rect 22328 62665 22332 62721
rect 22332 62665 22388 62721
rect 22388 62665 22392 62721
rect 22328 62661 22392 62665
rect 22328 62641 22392 62645
rect 22328 62585 22332 62641
rect 22332 62585 22388 62641
rect 22388 62585 22392 62641
rect 22328 62581 22392 62585
rect 22328 62561 22392 62565
rect 22328 62505 22332 62561
rect 22332 62505 22388 62561
rect 22388 62505 22392 62561
rect 22328 62501 22392 62505
rect 22328 62481 22392 62485
rect 22328 62425 22332 62481
rect 22332 62425 22388 62481
rect 22388 62425 22392 62481
rect 22328 62421 22392 62425
rect 22328 62401 22392 62405
rect 22328 62345 22332 62401
rect 22332 62345 22388 62401
rect 22388 62345 22392 62401
rect 22328 62341 22392 62345
rect 22328 62321 22392 62325
rect 22328 62265 22332 62321
rect 22332 62265 22388 62321
rect 22388 62265 22392 62321
rect 22328 62261 22392 62265
rect 22328 62241 22392 62245
rect 22328 62185 22332 62241
rect 22332 62185 22388 62241
rect 22388 62185 22392 62241
rect 22328 62181 22392 62185
rect 23416 62721 23480 62725
rect 23416 62665 23420 62721
rect 23420 62665 23476 62721
rect 23476 62665 23480 62721
rect 23416 62661 23480 62665
rect 23416 62641 23480 62645
rect 23416 62585 23420 62641
rect 23420 62585 23476 62641
rect 23476 62585 23480 62641
rect 23416 62581 23480 62585
rect 23416 62561 23480 62565
rect 23416 62505 23420 62561
rect 23420 62505 23476 62561
rect 23476 62505 23480 62561
rect 23416 62501 23480 62505
rect 23416 62481 23480 62485
rect 23416 62425 23420 62481
rect 23420 62425 23476 62481
rect 23476 62425 23480 62481
rect 23416 62421 23480 62425
rect 23416 62401 23480 62405
rect 23416 62345 23420 62401
rect 23420 62345 23476 62401
rect 23476 62345 23480 62401
rect 23416 62341 23480 62345
rect 23416 62321 23480 62325
rect 23416 62265 23420 62321
rect 23420 62265 23476 62321
rect 23476 62265 23480 62321
rect 23416 62261 23480 62265
rect 23416 62241 23480 62245
rect 23416 62185 23420 62241
rect 23420 62185 23476 62241
rect 23476 62185 23480 62241
rect 23416 62181 23480 62185
rect 24504 62721 24568 62725
rect 24504 62665 24508 62721
rect 24508 62665 24564 62721
rect 24564 62665 24568 62721
rect 24504 62661 24568 62665
rect 24504 62641 24568 62645
rect 24504 62585 24508 62641
rect 24508 62585 24564 62641
rect 24564 62585 24568 62641
rect 24504 62581 24568 62585
rect 24504 62561 24568 62565
rect 24504 62505 24508 62561
rect 24508 62505 24564 62561
rect 24564 62505 24568 62561
rect 24504 62501 24568 62505
rect 24504 62481 24568 62485
rect 24504 62425 24508 62481
rect 24508 62425 24564 62481
rect 24564 62425 24568 62481
rect 24504 62421 24568 62425
rect 24504 62401 24568 62405
rect 24504 62345 24508 62401
rect 24508 62345 24564 62401
rect 24564 62345 24568 62401
rect 24504 62341 24568 62345
rect 24504 62321 24568 62325
rect 24504 62265 24508 62321
rect 24508 62265 24564 62321
rect 24564 62265 24568 62321
rect 24504 62261 24568 62265
rect 24504 62241 24568 62245
rect 24504 62185 24508 62241
rect 24508 62185 24564 62241
rect 24564 62185 24568 62241
rect 24504 62181 24568 62185
rect 25592 62721 25656 62725
rect 25592 62665 25596 62721
rect 25596 62665 25652 62721
rect 25652 62665 25656 62721
rect 25592 62661 25656 62665
rect 25592 62641 25656 62645
rect 25592 62585 25596 62641
rect 25596 62585 25652 62641
rect 25652 62585 25656 62641
rect 25592 62581 25656 62585
rect 25592 62561 25656 62565
rect 25592 62505 25596 62561
rect 25596 62505 25652 62561
rect 25652 62505 25656 62561
rect 25592 62501 25656 62505
rect 25592 62481 25656 62485
rect 25592 62425 25596 62481
rect 25596 62425 25652 62481
rect 25652 62425 25656 62481
rect 25592 62421 25656 62425
rect 25592 62401 25656 62405
rect 25592 62345 25596 62401
rect 25596 62345 25652 62401
rect 25652 62345 25656 62401
rect 25592 62341 25656 62345
rect 25592 62321 25656 62325
rect 25592 62265 25596 62321
rect 25596 62265 25652 62321
rect 25652 62265 25656 62321
rect 25592 62261 25656 62265
rect 25592 62241 25656 62245
rect 25592 62185 25596 62241
rect 25596 62185 25652 62241
rect 25652 62185 25656 62241
rect 25592 62181 25656 62185
rect 26680 62721 26744 62725
rect 26680 62665 26684 62721
rect 26684 62665 26740 62721
rect 26740 62665 26744 62721
rect 26680 62661 26744 62665
rect 26680 62641 26744 62645
rect 26680 62585 26684 62641
rect 26684 62585 26740 62641
rect 26740 62585 26744 62641
rect 26680 62581 26744 62585
rect 26680 62561 26744 62565
rect 26680 62505 26684 62561
rect 26684 62505 26740 62561
rect 26740 62505 26744 62561
rect 26680 62501 26744 62505
rect 26680 62481 26744 62485
rect 26680 62425 26684 62481
rect 26684 62425 26740 62481
rect 26740 62425 26744 62481
rect 26680 62421 26744 62425
rect 26680 62401 26744 62405
rect 26680 62345 26684 62401
rect 26684 62345 26740 62401
rect 26740 62345 26744 62401
rect 26680 62341 26744 62345
rect 26680 62321 26744 62325
rect 26680 62265 26684 62321
rect 26684 62265 26740 62321
rect 26740 62265 26744 62321
rect 26680 62261 26744 62265
rect 26680 62241 26744 62245
rect 26680 62185 26684 62241
rect 26684 62185 26740 62241
rect 26740 62185 26744 62241
rect 26680 62181 26744 62185
rect 28856 62721 28920 62725
rect 28856 62665 28860 62721
rect 28860 62665 28916 62721
rect 28916 62665 28920 62721
rect 28856 62661 28920 62665
rect 28856 62641 28920 62645
rect 28856 62585 28860 62641
rect 28860 62585 28916 62641
rect 28916 62585 28920 62641
rect 28856 62581 28920 62585
rect 28856 62561 28920 62565
rect 28856 62505 28860 62561
rect 28860 62505 28916 62561
rect 28916 62505 28920 62561
rect 28856 62501 28920 62505
rect 28856 62481 28920 62485
rect 28856 62425 28860 62481
rect 28860 62425 28916 62481
rect 28916 62425 28920 62481
rect 28856 62421 28920 62425
rect 28856 62401 28920 62405
rect 28856 62345 28860 62401
rect 28860 62345 28916 62401
rect 28916 62345 28920 62401
rect 28856 62341 28920 62345
rect 28856 62321 28920 62325
rect 28856 62265 28860 62321
rect 28860 62265 28916 62321
rect 28916 62265 28920 62321
rect 28856 62261 28920 62265
rect 28856 62241 28920 62245
rect 28856 62185 28860 62241
rect 28860 62185 28916 62241
rect 28916 62185 28920 62241
rect 28856 62181 28920 62185
rect 29944 62721 30008 62725
rect 29944 62665 29948 62721
rect 29948 62665 30004 62721
rect 30004 62665 30008 62721
rect 29944 62661 30008 62665
rect 29944 62641 30008 62645
rect 29944 62585 29948 62641
rect 29948 62585 30004 62641
rect 30004 62585 30008 62641
rect 29944 62581 30008 62585
rect 29944 62561 30008 62565
rect 29944 62505 29948 62561
rect 29948 62505 30004 62561
rect 30004 62505 30008 62561
rect 29944 62501 30008 62505
rect 29944 62481 30008 62485
rect 29944 62425 29948 62481
rect 29948 62425 30004 62481
rect 30004 62425 30008 62481
rect 29944 62421 30008 62425
rect 29944 62401 30008 62405
rect 29944 62345 29948 62401
rect 29948 62345 30004 62401
rect 30004 62345 30008 62401
rect 29944 62341 30008 62345
rect 29944 62321 30008 62325
rect 29944 62265 29948 62321
rect 29948 62265 30004 62321
rect 30004 62265 30008 62321
rect 29944 62261 30008 62265
rect 29944 62241 30008 62245
rect 29944 62185 29948 62241
rect 29948 62185 30004 62241
rect 30004 62185 30008 62241
rect 29944 62181 30008 62185
rect 31032 62721 31096 62725
rect 31032 62665 31036 62721
rect 31036 62665 31092 62721
rect 31092 62665 31096 62721
rect 31032 62661 31096 62665
rect 31032 62641 31096 62645
rect 31032 62585 31036 62641
rect 31036 62585 31092 62641
rect 31092 62585 31096 62641
rect 31032 62581 31096 62585
rect 31032 62561 31096 62565
rect 31032 62505 31036 62561
rect 31036 62505 31092 62561
rect 31092 62505 31096 62561
rect 31032 62501 31096 62505
rect 31032 62481 31096 62485
rect 31032 62425 31036 62481
rect 31036 62425 31092 62481
rect 31092 62425 31096 62481
rect 31032 62421 31096 62425
rect 31032 62401 31096 62405
rect 31032 62345 31036 62401
rect 31036 62345 31092 62401
rect 31092 62345 31096 62401
rect 31032 62341 31096 62345
rect 31032 62321 31096 62325
rect 31032 62265 31036 62321
rect 31036 62265 31092 62321
rect 31092 62265 31096 62321
rect 31032 62261 31096 62265
rect 31032 62241 31096 62245
rect 31032 62185 31036 62241
rect 31036 62185 31092 62241
rect 31092 62185 31096 62241
rect 31032 62181 31096 62185
rect -8557 54591 -8493 54595
rect -8557 54535 -8553 54591
rect -8553 54535 -8497 54591
rect -8497 54535 -8493 54591
rect -8557 54531 -8493 54535
rect -6866 54592 -6802 54596
rect -6866 54536 -6862 54592
rect -6862 54536 -6806 54592
rect -6806 54536 -6802 54592
rect -6866 54532 -6802 54536
rect -5161 54591 -5097 54595
rect -5161 54535 -5157 54591
rect -5157 54535 -5101 54591
rect -5101 54535 -5097 54591
rect -5161 54531 -5097 54535
rect -3365 54591 -3301 54595
rect -3365 54535 -3361 54591
rect -3361 54535 -3305 54591
rect -3305 54535 -3301 54591
rect -3365 54531 -3301 54535
rect -1536 54591 -1472 54595
rect -1536 54535 -1532 54591
rect -1532 54535 -1476 54591
rect -1476 54535 -1472 54591
rect -1536 54531 -1472 54535
rect -9695 54399 -9631 54403
rect -9695 54343 -9691 54399
rect -9691 54343 -9635 54399
rect -9635 54343 -9631 54399
rect -9695 54339 -9631 54343
rect -9615 54399 -9551 54403
rect -9615 54343 -9611 54399
rect -9611 54343 -9555 54399
rect -9555 54343 -9551 54399
rect -9615 54339 -9551 54343
rect -9535 54399 -9471 54403
rect -9535 54343 -9531 54399
rect -9531 54343 -9475 54399
rect -9475 54343 -9471 54399
rect -9535 54339 -9471 54343
rect -7900 54398 -7836 54402
rect -7900 54342 -7896 54398
rect -7896 54342 -7840 54398
rect -7840 54342 -7836 54398
rect -7900 54338 -7836 54342
rect -7820 54398 -7756 54402
rect -7820 54342 -7816 54398
rect -7816 54342 -7760 54398
rect -7760 54342 -7756 54398
rect -7820 54338 -7756 54342
rect -7740 54398 -7676 54402
rect -7740 54342 -7736 54398
rect -7736 54342 -7680 54398
rect -7680 54342 -7676 54398
rect -7740 54338 -7676 54342
rect -6100 54400 -6036 54404
rect -6100 54344 -6096 54400
rect -6096 54344 -6040 54400
rect -6040 54344 -6036 54400
rect -6100 54340 -6036 54344
rect -6020 54400 -5956 54404
rect -6020 54344 -6016 54400
rect -6016 54344 -5960 54400
rect -5960 54344 -5956 54400
rect -6020 54340 -5956 54344
rect -5940 54400 -5876 54404
rect -5940 54344 -5936 54400
rect -5936 54344 -5880 54400
rect -5880 54344 -5876 54400
rect -5940 54340 -5876 54344
rect -4302 54399 -4238 54403
rect -4302 54343 -4298 54399
rect -4298 54343 -4242 54399
rect -4242 54343 -4238 54399
rect -4302 54339 -4238 54343
rect -4222 54399 -4158 54403
rect -4222 54343 -4218 54399
rect -4218 54343 -4162 54399
rect -4162 54343 -4158 54399
rect -4222 54339 -4158 54343
rect -4142 54399 -4078 54403
rect -4142 54343 -4138 54399
rect -4138 54343 -4082 54399
rect -4082 54343 -4078 54399
rect -4142 54339 -4078 54343
rect -2504 54400 -2440 54404
rect -2504 54344 -2500 54400
rect -2500 54344 -2444 54400
rect -2444 54344 -2440 54400
rect -2504 54340 -2440 54344
rect -2424 54400 -2360 54404
rect -2424 54344 -2420 54400
rect -2420 54344 -2364 54400
rect -2364 54344 -2360 54400
rect -2424 54340 -2360 54344
rect -2344 54400 -2280 54404
rect -2344 54344 -2340 54400
rect -2340 54344 -2284 54400
rect -2284 54344 -2280 54400
rect -2344 54340 -2280 54344
rect -701 54399 -637 54403
rect -701 54343 -697 54399
rect -697 54343 -641 54399
rect -641 54343 -637 54399
rect -701 54339 -637 54343
rect -621 54399 -557 54403
rect -621 54343 -617 54399
rect -617 54343 -561 54399
rect -561 54343 -557 54399
rect -621 54339 -557 54343
rect -541 54399 -477 54403
rect -541 54343 -537 54399
rect -537 54343 -481 54399
rect -481 54343 -477 54399
rect -541 54339 -477 54343
rect 176 54400 240 54404
rect 176 54344 180 54400
rect 180 54344 236 54400
rect 236 54344 240 54400
rect 176 54340 240 54344
rect -7265 54019 -7201 54083
rect -1865 54019 -1801 54083
rect -8073 53766 -8009 53830
rect -2673 53766 -2609 53830
rect -10536 53338 -10472 53402
rect -1865 53338 -1801 53402
rect -11305 53082 -11241 53146
rect -2673 53082 -2609 53146
rect 361 60802 505 60806
rect 361 53146 365 60802
rect 365 53146 501 60802
rect 501 53146 505 60802
rect 361 53142 505 53146
rect -12315 52649 -12251 52713
rect -7265 52649 -7201 52713
rect -13096 52326 -13032 52390
rect -8073 52326 -8009 52390
rect -8844 51239 -8780 51243
rect -8844 51183 -8840 51239
rect -8840 51183 -8784 51239
rect -8784 51183 -8780 51239
rect -8844 51179 -8780 51183
rect -8844 51159 -8780 51163
rect -8844 51103 -8840 51159
rect -8840 51103 -8784 51159
rect -8784 51103 -8780 51159
rect -8844 51099 -8780 51103
rect -7722 51243 -7658 51247
rect -7722 51187 -7718 51243
rect -7718 51187 -7662 51243
rect -7662 51187 -7658 51243
rect -7722 51183 -7658 51187
rect -8844 51079 -8780 51083
rect -8844 51023 -8840 51079
rect -8840 51023 -8784 51079
rect -8784 51023 -8780 51079
rect -8844 51019 -8780 51023
rect -5660 51042 -3916 51046
rect -5660 50906 -5656 51042
rect -5656 50906 -3920 51042
rect -3920 50906 -3916 51042
rect -5660 50902 -3916 50906
rect -3341 51053 -2557 51057
rect -3341 50917 -3337 51053
rect -3337 50917 -2561 51053
rect -2561 50917 -2557 51053
rect -3341 50913 -2557 50917
rect -1642 51043 -778 51047
rect -1642 50907 -1638 51043
rect -1638 50907 -782 51043
rect -782 50907 -778 51043
rect -1642 50903 -778 50907
rect -8859 50772 -8795 50776
rect -8859 50716 -8855 50772
rect -8855 50716 -8799 50772
rect -8799 50716 -8795 50772
rect -8859 50712 -8795 50716
rect -8859 50692 -8795 50696
rect -8859 50636 -8855 50692
rect -8855 50636 -8799 50692
rect -8799 50636 -8795 50692
rect -8859 50632 -8795 50636
rect -8859 50612 -8795 50616
rect -19005 50532 -18941 50596
rect -8859 50556 -8855 50612
rect -8855 50556 -8799 50612
rect -8799 50556 -8795 50612
rect -8859 50552 -8795 50556
rect -8859 50532 -8795 50536
rect -8859 50476 -8855 50532
rect -8855 50476 -8799 50532
rect -8799 50476 -8795 50532
rect -8859 50472 -8795 50476
rect -8859 50452 -8795 50456
rect -8859 50396 -8855 50452
rect -8855 50396 -8799 50452
rect -8799 50396 -8795 50452
rect -8859 50392 -8795 50396
rect -8480 50437 -8416 50441
rect -8480 50381 -8476 50437
rect -8476 50381 -8420 50437
rect -8420 50381 -8416 50437
rect -8480 50377 -8416 50381
rect -8480 50008 -8416 50072
rect -27050 49716 -26986 49720
rect -27050 49660 -27046 49716
rect -27046 49660 -26990 49716
rect -26990 49660 -26986 49716
rect -27050 49656 -26986 49660
rect -26970 49716 -26906 49720
rect -26970 49660 -26966 49716
rect -26966 49660 -26910 49716
rect -26910 49660 -26906 49716
rect -26970 49656 -26906 49660
rect -26890 49716 -26826 49720
rect -26890 49660 -26886 49716
rect -26886 49660 -26830 49716
rect -26830 49660 -26826 49716
rect -26890 49656 -26826 49660
rect -26810 49716 -26746 49720
rect -26810 49660 -26806 49716
rect -26806 49660 -26750 49716
rect -26750 49660 -26746 49716
rect -26810 49656 -26746 49660
rect -7722 49360 -7658 49424
rect -25964 49174 -25900 49178
rect -25964 49118 -25960 49174
rect -25960 49118 -25904 49174
rect -25904 49118 -25900 49174
rect -25964 49114 -25900 49118
rect -25884 49174 -25820 49178
rect -25884 49118 -25880 49174
rect -25880 49118 -25824 49174
rect -25824 49118 -25820 49174
rect -25884 49114 -25820 49118
rect -25804 49174 -25740 49178
rect -25804 49118 -25800 49174
rect -25800 49118 -25744 49174
rect -25744 49118 -25740 49174
rect -25804 49114 -25740 49118
rect -25724 49174 -25660 49178
rect -25724 49118 -25720 49174
rect -25720 49118 -25664 49174
rect -25664 49118 -25660 49174
rect -25724 49114 -25660 49118
rect -5912 50716 -5768 50720
rect -5912 47780 -5908 50716
rect -5908 47780 -5772 50716
rect -5772 47780 -5768 50716
rect -5912 47776 -5768 47780
rect -51 47791 -47 50735
rect -47 47791 89 50735
rect 89 47791 93 50735
rect 10212 60814 10516 60818
rect 10212 47638 10216 60814
rect 10216 47638 10512 60814
rect 10512 47638 10516 60814
rect 10212 47634 10516 47638
rect 17431 60724 17495 60728
rect 17431 60668 17435 60724
rect 17435 60668 17491 60724
rect 17491 60668 17495 60724
rect 17431 60664 17495 60668
rect 17431 60644 17495 60648
rect 17431 60588 17435 60644
rect 17435 60588 17491 60644
rect 17491 60588 17495 60644
rect 17431 60584 17495 60588
rect 17431 60564 17495 60568
rect 17431 60508 17435 60564
rect 17435 60508 17491 60564
rect 17491 60508 17495 60564
rect 17431 60504 17495 60508
rect 17431 60484 17495 60488
rect 17431 60428 17435 60484
rect 17435 60428 17491 60484
rect 17491 60428 17495 60484
rect 17431 60424 17495 60428
rect 17431 60404 17495 60408
rect 17431 60348 17435 60404
rect 17435 60348 17491 60404
rect 17491 60348 17495 60404
rect 17431 60344 17495 60348
rect 17431 60324 17495 60328
rect 17431 60268 17435 60324
rect 17435 60268 17491 60324
rect 17491 60268 17495 60324
rect 17431 60264 17495 60268
rect 17431 60244 17495 60248
rect 17431 60188 17435 60244
rect 17435 60188 17491 60244
rect 17491 60188 17495 60244
rect 17431 60184 17495 60188
rect 18519 60724 18583 60728
rect 18519 60668 18523 60724
rect 18523 60668 18579 60724
rect 18579 60668 18583 60724
rect 18519 60664 18583 60668
rect 18519 60644 18583 60648
rect 18519 60588 18523 60644
rect 18523 60588 18579 60644
rect 18579 60588 18583 60644
rect 18519 60584 18583 60588
rect 18519 60564 18583 60568
rect 18519 60508 18523 60564
rect 18523 60508 18579 60564
rect 18579 60508 18583 60564
rect 18519 60504 18583 60508
rect 18519 60484 18583 60488
rect 18519 60428 18523 60484
rect 18523 60428 18579 60484
rect 18579 60428 18583 60484
rect 18519 60424 18583 60428
rect 18519 60404 18583 60408
rect 18519 60348 18523 60404
rect 18523 60348 18579 60404
rect 18579 60348 18583 60404
rect 18519 60344 18583 60348
rect 18519 60324 18583 60328
rect 18519 60268 18523 60324
rect 18523 60268 18579 60324
rect 18579 60268 18583 60324
rect 18519 60264 18583 60268
rect 18519 60244 18583 60248
rect 18519 60188 18523 60244
rect 18523 60188 18579 60244
rect 18579 60188 18583 60244
rect 18519 60184 18583 60188
rect 19607 60724 19671 60728
rect 19607 60668 19611 60724
rect 19611 60668 19667 60724
rect 19667 60668 19671 60724
rect 19607 60664 19671 60668
rect 19607 60644 19671 60648
rect 19607 60588 19611 60644
rect 19611 60588 19667 60644
rect 19667 60588 19671 60644
rect 19607 60584 19671 60588
rect 19607 60564 19671 60568
rect 19607 60508 19611 60564
rect 19611 60508 19667 60564
rect 19667 60508 19671 60564
rect 19607 60504 19671 60508
rect 19607 60484 19671 60488
rect 19607 60428 19611 60484
rect 19611 60428 19667 60484
rect 19667 60428 19671 60484
rect 19607 60424 19671 60428
rect 19607 60404 19671 60408
rect 19607 60348 19611 60404
rect 19611 60348 19667 60404
rect 19667 60348 19671 60404
rect 19607 60344 19671 60348
rect 19607 60324 19671 60328
rect 19607 60268 19611 60324
rect 19611 60268 19667 60324
rect 19667 60268 19671 60324
rect 19607 60264 19671 60268
rect 19607 60244 19671 60248
rect 19607 60188 19611 60244
rect 19611 60188 19667 60244
rect 19667 60188 19671 60244
rect 19607 60184 19671 60188
rect 20695 60724 20759 60728
rect 20695 60668 20699 60724
rect 20699 60668 20755 60724
rect 20755 60668 20759 60724
rect 20695 60664 20759 60668
rect 20695 60644 20759 60648
rect 20695 60588 20699 60644
rect 20699 60588 20755 60644
rect 20755 60588 20759 60644
rect 20695 60584 20759 60588
rect 20695 60564 20759 60568
rect 20695 60508 20699 60564
rect 20699 60508 20755 60564
rect 20755 60508 20759 60564
rect 20695 60504 20759 60508
rect 20695 60484 20759 60488
rect 20695 60428 20699 60484
rect 20699 60428 20755 60484
rect 20755 60428 20759 60484
rect 20695 60424 20759 60428
rect 20695 60404 20759 60408
rect 20695 60348 20699 60404
rect 20699 60348 20755 60404
rect 20755 60348 20759 60404
rect 20695 60344 20759 60348
rect 20695 60324 20759 60328
rect 20695 60268 20699 60324
rect 20699 60268 20755 60324
rect 20755 60268 20759 60324
rect 20695 60264 20759 60268
rect 20695 60244 20759 60248
rect 20695 60188 20699 60244
rect 20699 60188 20755 60244
rect 20755 60188 20759 60244
rect 20695 60184 20759 60188
rect 21783 60724 21847 60728
rect 21783 60668 21787 60724
rect 21787 60668 21843 60724
rect 21843 60668 21847 60724
rect 21783 60664 21847 60668
rect 21783 60644 21847 60648
rect 21783 60588 21787 60644
rect 21787 60588 21843 60644
rect 21843 60588 21847 60644
rect 21783 60584 21847 60588
rect 21783 60564 21847 60568
rect 21783 60508 21787 60564
rect 21787 60508 21843 60564
rect 21843 60508 21847 60564
rect 21783 60504 21847 60508
rect 21783 60484 21847 60488
rect 21783 60428 21787 60484
rect 21787 60428 21843 60484
rect 21843 60428 21847 60484
rect 21783 60424 21847 60428
rect 21783 60404 21847 60408
rect 21783 60348 21787 60404
rect 21787 60348 21843 60404
rect 21843 60348 21847 60404
rect 21783 60344 21847 60348
rect 21783 60324 21847 60328
rect 21783 60268 21787 60324
rect 21787 60268 21843 60324
rect 21843 60268 21847 60324
rect 21783 60264 21847 60268
rect 21783 60244 21847 60248
rect 21783 60188 21787 60244
rect 21787 60188 21843 60244
rect 21843 60188 21847 60244
rect 21783 60184 21847 60188
rect 22871 60724 22935 60728
rect 22871 60668 22875 60724
rect 22875 60668 22931 60724
rect 22931 60668 22935 60724
rect 22871 60664 22935 60668
rect 22871 60644 22935 60648
rect 22871 60588 22875 60644
rect 22875 60588 22931 60644
rect 22931 60588 22935 60644
rect 22871 60584 22935 60588
rect 22871 60564 22935 60568
rect 22871 60508 22875 60564
rect 22875 60508 22931 60564
rect 22931 60508 22935 60564
rect 22871 60504 22935 60508
rect 22871 60484 22935 60488
rect 22871 60428 22875 60484
rect 22875 60428 22931 60484
rect 22931 60428 22935 60484
rect 22871 60424 22935 60428
rect 22871 60404 22935 60408
rect 22871 60348 22875 60404
rect 22875 60348 22931 60404
rect 22931 60348 22935 60404
rect 22871 60344 22935 60348
rect 22871 60324 22935 60328
rect 22871 60268 22875 60324
rect 22875 60268 22931 60324
rect 22931 60268 22935 60324
rect 22871 60264 22935 60268
rect 22871 60244 22935 60248
rect 22871 60188 22875 60244
rect 22875 60188 22931 60244
rect 22931 60188 22935 60244
rect 22871 60184 22935 60188
rect 23959 60724 24023 60728
rect 23959 60668 23963 60724
rect 23963 60668 24019 60724
rect 24019 60668 24023 60724
rect 23959 60664 24023 60668
rect 23959 60644 24023 60648
rect 23959 60588 23963 60644
rect 23963 60588 24019 60644
rect 24019 60588 24023 60644
rect 23959 60584 24023 60588
rect 23959 60564 24023 60568
rect 23959 60508 23963 60564
rect 23963 60508 24019 60564
rect 24019 60508 24023 60564
rect 23959 60504 24023 60508
rect 23959 60484 24023 60488
rect 23959 60428 23963 60484
rect 23963 60428 24019 60484
rect 24019 60428 24023 60484
rect 23959 60424 24023 60428
rect 23959 60404 24023 60408
rect 23959 60348 23963 60404
rect 23963 60348 24019 60404
rect 24019 60348 24023 60404
rect 23959 60344 24023 60348
rect 23959 60324 24023 60328
rect 23959 60268 23963 60324
rect 23963 60268 24019 60324
rect 24019 60268 24023 60324
rect 23959 60264 24023 60268
rect 23959 60244 24023 60248
rect 23959 60188 23963 60244
rect 23963 60188 24019 60244
rect 24019 60188 24023 60244
rect 23959 60184 24023 60188
rect 25047 60724 25111 60728
rect 25047 60668 25051 60724
rect 25051 60668 25107 60724
rect 25107 60668 25111 60724
rect 25047 60664 25111 60668
rect 25047 60644 25111 60648
rect 25047 60588 25051 60644
rect 25051 60588 25107 60644
rect 25107 60588 25111 60644
rect 25047 60584 25111 60588
rect 25047 60564 25111 60568
rect 25047 60508 25051 60564
rect 25051 60508 25107 60564
rect 25107 60508 25111 60564
rect 25047 60504 25111 60508
rect 25047 60484 25111 60488
rect 25047 60428 25051 60484
rect 25051 60428 25107 60484
rect 25107 60428 25111 60484
rect 25047 60424 25111 60428
rect 25047 60404 25111 60408
rect 25047 60348 25051 60404
rect 25051 60348 25107 60404
rect 25107 60348 25111 60404
rect 25047 60344 25111 60348
rect 25047 60324 25111 60328
rect 25047 60268 25051 60324
rect 25051 60268 25107 60324
rect 25107 60268 25111 60324
rect 25047 60264 25111 60268
rect 25047 60244 25111 60248
rect 25047 60188 25051 60244
rect 25051 60188 25107 60244
rect 25107 60188 25111 60244
rect 25047 60184 25111 60188
rect 26135 60724 26199 60728
rect 26135 60668 26139 60724
rect 26139 60668 26195 60724
rect 26195 60668 26199 60724
rect 26135 60664 26199 60668
rect 26135 60644 26199 60648
rect 26135 60588 26139 60644
rect 26139 60588 26195 60644
rect 26195 60588 26199 60644
rect 26135 60584 26199 60588
rect 26135 60564 26199 60568
rect 26135 60508 26139 60564
rect 26139 60508 26195 60564
rect 26195 60508 26199 60564
rect 26135 60504 26199 60508
rect 26135 60484 26199 60488
rect 26135 60428 26139 60484
rect 26139 60428 26195 60484
rect 26195 60428 26199 60484
rect 26135 60424 26199 60428
rect 26135 60404 26199 60408
rect 26135 60348 26139 60404
rect 26139 60348 26195 60404
rect 26195 60348 26199 60404
rect 26135 60344 26199 60348
rect 26135 60324 26199 60328
rect 26135 60268 26139 60324
rect 26139 60268 26195 60324
rect 26195 60268 26199 60324
rect 26135 60264 26199 60268
rect 26135 60244 26199 60248
rect 26135 60188 26139 60244
rect 26139 60188 26195 60244
rect 26195 60188 26199 60244
rect 26135 60184 26199 60188
rect 27223 60724 27287 60728
rect 27223 60668 27227 60724
rect 27227 60668 27283 60724
rect 27283 60668 27287 60724
rect 27223 60664 27287 60668
rect 27223 60644 27287 60648
rect 27223 60588 27227 60644
rect 27227 60588 27283 60644
rect 27283 60588 27287 60644
rect 27223 60584 27287 60588
rect 27223 60564 27287 60568
rect 27223 60508 27227 60564
rect 27227 60508 27283 60564
rect 27283 60508 27287 60564
rect 27223 60504 27287 60508
rect 27223 60484 27287 60488
rect 27223 60428 27227 60484
rect 27227 60428 27283 60484
rect 27283 60428 27287 60484
rect 27223 60424 27287 60428
rect 27223 60404 27287 60408
rect 27223 60348 27227 60404
rect 27227 60348 27283 60404
rect 27283 60348 27287 60404
rect 27223 60344 27287 60348
rect 27223 60324 27287 60328
rect 27223 60268 27227 60324
rect 27227 60268 27283 60324
rect 27283 60268 27287 60324
rect 27223 60264 27287 60268
rect 27223 60244 27287 60248
rect 27223 60188 27227 60244
rect 27227 60188 27283 60244
rect 27283 60188 27287 60244
rect 27223 60184 27287 60188
rect 28311 60724 28375 60728
rect 28311 60668 28315 60724
rect 28315 60668 28371 60724
rect 28371 60668 28375 60724
rect 28311 60664 28375 60668
rect 28311 60644 28375 60648
rect 28311 60588 28315 60644
rect 28315 60588 28371 60644
rect 28371 60588 28375 60644
rect 28311 60584 28375 60588
rect 28311 60564 28375 60568
rect 28311 60508 28315 60564
rect 28315 60508 28371 60564
rect 28371 60508 28375 60564
rect 28311 60504 28375 60508
rect 28311 60484 28375 60488
rect 28311 60428 28315 60484
rect 28315 60428 28371 60484
rect 28371 60428 28375 60484
rect 28311 60424 28375 60428
rect 28311 60404 28375 60408
rect 28311 60348 28315 60404
rect 28315 60348 28371 60404
rect 28371 60348 28375 60404
rect 28311 60344 28375 60348
rect 28311 60324 28375 60328
rect 28311 60268 28315 60324
rect 28315 60268 28371 60324
rect 28371 60268 28375 60324
rect 28311 60264 28375 60268
rect 28311 60244 28375 60248
rect 28311 60188 28315 60244
rect 28315 60188 28371 60244
rect 28371 60188 28375 60244
rect 28311 60184 28375 60188
rect 29399 60724 29463 60728
rect 29399 60668 29403 60724
rect 29403 60668 29459 60724
rect 29459 60668 29463 60724
rect 29399 60664 29463 60668
rect 29399 60644 29463 60648
rect 29399 60588 29403 60644
rect 29403 60588 29459 60644
rect 29459 60588 29463 60644
rect 29399 60584 29463 60588
rect 29399 60564 29463 60568
rect 29399 60508 29403 60564
rect 29403 60508 29459 60564
rect 29459 60508 29463 60564
rect 29399 60504 29463 60508
rect 29399 60484 29463 60488
rect 29399 60428 29403 60484
rect 29403 60428 29459 60484
rect 29459 60428 29463 60484
rect 29399 60424 29463 60428
rect 29399 60404 29463 60408
rect 29399 60348 29403 60404
rect 29403 60348 29459 60404
rect 29459 60348 29463 60404
rect 29399 60344 29463 60348
rect 29399 60324 29463 60328
rect 29399 60268 29403 60324
rect 29403 60268 29459 60324
rect 29459 60268 29463 60324
rect 29399 60264 29463 60268
rect 29399 60244 29463 60248
rect 29399 60188 29403 60244
rect 29403 60188 29459 60244
rect 29459 60188 29463 60244
rect 29399 60184 29463 60188
rect 30487 60724 30551 60728
rect 30487 60668 30491 60724
rect 30491 60668 30547 60724
rect 30547 60668 30551 60724
rect 30487 60664 30551 60668
rect 30487 60644 30551 60648
rect 30487 60588 30491 60644
rect 30491 60588 30547 60644
rect 30547 60588 30551 60644
rect 30487 60584 30551 60588
rect 30487 60564 30551 60568
rect 30487 60508 30491 60564
rect 30491 60508 30547 60564
rect 30547 60508 30551 60564
rect 30487 60504 30551 60508
rect 30487 60484 30551 60488
rect 30487 60428 30491 60484
rect 30491 60428 30547 60484
rect 30547 60428 30551 60484
rect 30487 60424 30551 60428
rect 30487 60404 30551 60408
rect 30487 60348 30491 60404
rect 30491 60348 30547 60404
rect 30547 60348 30551 60404
rect 30487 60344 30551 60348
rect 30487 60324 30551 60328
rect 30487 60268 30491 60324
rect 30491 60268 30547 60324
rect 30547 60268 30551 60324
rect 30487 60264 30551 60268
rect 30487 60244 30551 60248
rect 30487 60188 30491 60244
rect 30491 60188 30547 60244
rect 30547 60188 30551 60244
rect 30487 60184 30551 60188
rect 31575 60724 31639 60728
rect 31575 60668 31579 60724
rect 31579 60668 31635 60724
rect 31635 60668 31639 60724
rect 31575 60664 31639 60668
rect 31575 60644 31639 60648
rect 31575 60588 31579 60644
rect 31579 60588 31635 60644
rect 31635 60588 31639 60644
rect 31575 60584 31639 60588
rect 31575 60564 31639 60568
rect 31575 60508 31579 60564
rect 31579 60508 31635 60564
rect 31635 60508 31639 60564
rect 31575 60504 31639 60508
rect 31575 60484 31639 60488
rect 31575 60428 31579 60484
rect 31579 60428 31635 60484
rect 31635 60428 31639 60484
rect 31575 60424 31639 60428
rect 31575 60404 31639 60408
rect 31575 60348 31579 60404
rect 31579 60348 31635 60404
rect 31635 60348 31639 60404
rect 31575 60344 31639 60348
rect 31575 60324 31639 60328
rect 31575 60268 31579 60324
rect 31579 60268 31635 60324
rect 31635 60268 31639 60324
rect 31575 60264 31639 60268
rect 31575 60244 31639 60248
rect 31575 60188 31579 60244
rect 31579 60188 31635 60244
rect 31635 60188 31639 60244
rect 31575 60184 31639 60188
rect 17976 58721 18040 58725
rect 17976 58665 17980 58721
rect 17980 58665 18036 58721
rect 18036 58665 18040 58721
rect 17976 58661 18040 58665
rect 17976 58641 18040 58645
rect 17976 58585 17980 58641
rect 17980 58585 18036 58641
rect 18036 58585 18040 58641
rect 17976 58581 18040 58585
rect 17976 58561 18040 58565
rect 17976 58505 17980 58561
rect 17980 58505 18036 58561
rect 18036 58505 18040 58561
rect 17976 58501 18040 58505
rect 17976 58481 18040 58485
rect 17976 58425 17980 58481
rect 17980 58425 18036 58481
rect 18036 58425 18040 58481
rect 17976 58421 18040 58425
rect 17976 58401 18040 58405
rect 17976 58345 17980 58401
rect 17980 58345 18036 58401
rect 18036 58345 18040 58401
rect 17976 58341 18040 58345
rect 17976 58321 18040 58325
rect 17976 58265 17980 58321
rect 17980 58265 18036 58321
rect 18036 58265 18040 58321
rect 17976 58261 18040 58265
rect 17976 58241 18040 58245
rect 17976 58185 17980 58241
rect 17980 58185 18036 58241
rect 18036 58185 18040 58241
rect 17976 58181 18040 58185
rect 19064 58721 19128 58725
rect 19064 58665 19068 58721
rect 19068 58665 19124 58721
rect 19124 58665 19128 58721
rect 19064 58661 19128 58665
rect 19064 58641 19128 58645
rect 19064 58585 19068 58641
rect 19068 58585 19124 58641
rect 19124 58585 19128 58641
rect 19064 58581 19128 58585
rect 19064 58561 19128 58565
rect 19064 58505 19068 58561
rect 19068 58505 19124 58561
rect 19124 58505 19128 58561
rect 19064 58501 19128 58505
rect 19064 58481 19128 58485
rect 19064 58425 19068 58481
rect 19068 58425 19124 58481
rect 19124 58425 19128 58481
rect 19064 58421 19128 58425
rect 19064 58401 19128 58405
rect 19064 58345 19068 58401
rect 19068 58345 19124 58401
rect 19124 58345 19128 58401
rect 19064 58341 19128 58345
rect 19064 58321 19128 58325
rect 19064 58265 19068 58321
rect 19068 58265 19124 58321
rect 19124 58265 19128 58321
rect 19064 58261 19128 58265
rect 19064 58241 19128 58245
rect 19064 58185 19068 58241
rect 19068 58185 19124 58241
rect 19124 58185 19128 58241
rect 19064 58181 19128 58185
rect 20152 58721 20216 58725
rect 20152 58665 20156 58721
rect 20156 58665 20212 58721
rect 20212 58665 20216 58721
rect 20152 58661 20216 58665
rect 20152 58641 20216 58645
rect 20152 58585 20156 58641
rect 20156 58585 20212 58641
rect 20212 58585 20216 58641
rect 20152 58581 20216 58585
rect 20152 58561 20216 58565
rect 20152 58505 20156 58561
rect 20156 58505 20212 58561
rect 20212 58505 20216 58561
rect 20152 58501 20216 58505
rect 20152 58481 20216 58485
rect 20152 58425 20156 58481
rect 20156 58425 20212 58481
rect 20212 58425 20216 58481
rect 20152 58421 20216 58425
rect 20152 58401 20216 58405
rect 20152 58345 20156 58401
rect 20156 58345 20212 58401
rect 20212 58345 20216 58401
rect 20152 58341 20216 58345
rect 20152 58321 20216 58325
rect 20152 58265 20156 58321
rect 20156 58265 20212 58321
rect 20212 58265 20216 58321
rect 20152 58261 20216 58265
rect 20152 58241 20216 58245
rect 20152 58185 20156 58241
rect 20156 58185 20212 58241
rect 20212 58185 20216 58241
rect 20152 58181 20216 58185
rect 21240 58721 21304 58725
rect 21240 58665 21244 58721
rect 21244 58665 21300 58721
rect 21300 58665 21304 58721
rect 21240 58661 21304 58665
rect 21240 58641 21304 58645
rect 21240 58585 21244 58641
rect 21244 58585 21300 58641
rect 21300 58585 21304 58641
rect 21240 58581 21304 58585
rect 21240 58561 21304 58565
rect 21240 58505 21244 58561
rect 21244 58505 21300 58561
rect 21300 58505 21304 58561
rect 21240 58501 21304 58505
rect 21240 58481 21304 58485
rect 21240 58425 21244 58481
rect 21244 58425 21300 58481
rect 21300 58425 21304 58481
rect 21240 58421 21304 58425
rect 21240 58401 21304 58405
rect 21240 58345 21244 58401
rect 21244 58345 21300 58401
rect 21300 58345 21304 58401
rect 21240 58341 21304 58345
rect 21240 58321 21304 58325
rect 21240 58265 21244 58321
rect 21244 58265 21300 58321
rect 21300 58265 21304 58321
rect 21240 58261 21304 58265
rect 21240 58241 21304 58245
rect 21240 58185 21244 58241
rect 21244 58185 21300 58241
rect 21300 58185 21304 58241
rect 21240 58181 21304 58185
rect 22328 58721 22392 58725
rect 22328 58665 22332 58721
rect 22332 58665 22388 58721
rect 22388 58665 22392 58721
rect 22328 58661 22392 58665
rect 22328 58641 22392 58645
rect 22328 58585 22332 58641
rect 22332 58585 22388 58641
rect 22388 58585 22392 58641
rect 22328 58581 22392 58585
rect 22328 58561 22392 58565
rect 22328 58505 22332 58561
rect 22332 58505 22388 58561
rect 22388 58505 22392 58561
rect 22328 58501 22392 58505
rect 22328 58481 22392 58485
rect 22328 58425 22332 58481
rect 22332 58425 22388 58481
rect 22388 58425 22392 58481
rect 22328 58421 22392 58425
rect 22328 58401 22392 58405
rect 22328 58345 22332 58401
rect 22332 58345 22388 58401
rect 22388 58345 22392 58401
rect 22328 58341 22392 58345
rect 22328 58321 22392 58325
rect 22328 58265 22332 58321
rect 22332 58265 22388 58321
rect 22388 58265 22392 58321
rect 22328 58261 22392 58265
rect 22328 58241 22392 58245
rect 22328 58185 22332 58241
rect 22332 58185 22388 58241
rect 22388 58185 22392 58241
rect 22328 58181 22392 58185
rect 23416 58721 23480 58725
rect 23416 58665 23420 58721
rect 23420 58665 23476 58721
rect 23476 58665 23480 58721
rect 23416 58661 23480 58665
rect 23416 58641 23480 58645
rect 23416 58585 23420 58641
rect 23420 58585 23476 58641
rect 23476 58585 23480 58641
rect 23416 58581 23480 58585
rect 23416 58561 23480 58565
rect 23416 58505 23420 58561
rect 23420 58505 23476 58561
rect 23476 58505 23480 58561
rect 23416 58501 23480 58505
rect 23416 58481 23480 58485
rect 23416 58425 23420 58481
rect 23420 58425 23476 58481
rect 23476 58425 23480 58481
rect 23416 58421 23480 58425
rect 23416 58401 23480 58405
rect 23416 58345 23420 58401
rect 23420 58345 23476 58401
rect 23476 58345 23480 58401
rect 23416 58341 23480 58345
rect 23416 58321 23480 58325
rect 23416 58265 23420 58321
rect 23420 58265 23476 58321
rect 23476 58265 23480 58321
rect 23416 58261 23480 58265
rect 23416 58241 23480 58245
rect 23416 58185 23420 58241
rect 23420 58185 23476 58241
rect 23476 58185 23480 58241
rect 23416 58181 23480 58185
rect 24504 58721 24568 58725
rect 24504 58665 24508 58721
rect 24508 58665 24564 58721
rect 24564 58665 24568 58721
rect 24504 58661 24568 58665
rect 24504 58641 24568 58645
rect 24504 58585 24508 58641
rect 24508 58585 24564 58641
rect 24564 58585 24568 58641
rect 24504 58581 24568 58585
rect 24504 58561 24568 58565
rect 24504 58505 24508 58561
rect 24508 58505 24564 58561
rect 24564 58505 24568 58561
rect 24504 58501 24568 58505
rect 24504 58481 24568 58485
rect 24504 58425 24508 58481
rect 24508 58425 24564 58481
rect 24564 58425 24568 58481
rect 24504 58421 24568 58425
rect 24504 58401 24568 58405
rect 24504 58345 24508 58401
rect 24508 58345 24564 58401
rect 24564 58345 24568 58401
rect 24504 58341 24568 58345
rect 24504 58321 24568 58325
rect 24504 58265 24508 58321
rect 24508 58265 24564 58321
rect 24564 58265 24568 58321
rect 24504 58261 24568 58265
rect 24504 58241 24568 58245
rect 24504 58185 24508 58241
rect 24508 58185 24564 58241
rect 24564 58185 24568 58241
rect 24504 58181 24568 58185
rect 25592 58721 25656 58725
rect 25592 58665 25596 58721
rect 25596 58665 25652 58721
rect 25652 58665 25656 58721
rect 25592 58661 25656 58665
rect 25592 58641 25656 58645
rect 25592 58585 25596 58641
rect 25596 58585 25652 58641
rect 25652 58585 25656 58641
rect 25592 58581 25656 58585
rect 25592 58561 25656 58565
rect 25592 58505 25596 58561
rect 25596 58505 25652 58561
rect 25652 58505 25656 58561
rect 25592 58501 25656 58505
rect 25592 58481 25656 58485
rect 25592 58425 25596 58481
rect 25596 58425 25652 58481
rect 25652 58425 25656 58481
rect 25592 58421 25656 58425
rect 25592 58401 25656 58405
rect 25592 58345 25596 58401
rect 25596 58345 25652 58401
rect 25652 58345 25656 58401
rect 25592 58341 25656 58345
rect 25592 58321 25656 58325
rect 25592 58265 25596 58321
rect 25596 58265 25652 58321
rect 25652 58265 25656 58321
rect 25592 58261 25656 58265
rect 25592 58241 25656 58245
rect 25592 58185 25596 58241
rect 25596 58185 25652 58241
rect 25652 58185 25656 58241
rect 25592 58181 25656 58185
rect 26680 58721 26744 58725
rect 26680 58665 26684 58721
rect 26684 58665 26740 58721
rect 26740 58665 26744 58721
rect 26680 58661 26744 58665
rect 26680 58641 26744 58645
rect 26680 58585 26684 58641
rect 26684 58585 26740 58641
rect 26740 58585 26744 58641
rect 26680 58581 26744 58585
rect 26680 58561 26744 58565
rect 26680 58505 26684 58561
rect 26684 58505 26740 58561
rect 26740 58505 26744 58561
rect 26680 58501 26744 58505
rect 26680 58481 26744 58485
rect 26680 58425 26684 58481
rect 26684 58425 26740 58481
rect 26740 58425 26744 58481
rect 26680 58421 26744 58425
rect 26680 58401 26744 58405
rect 26680 58345 26684 58401
rect 26684 58345 26740 58401
rect 26740 58345 26744 58401
rect 26680 58341 26744 58345
rect 26680 58321 26744 58325
rect 26680 58265 26684 58321
rect 26684 58265 26740 58321
rect 26740 58265 26744 58321
rect 26680 58261 26744 58265
rect 26680 58241 26744 58245
rect 26680 58185 26684 58241
rect 26684 58185 26740 58241
rect 26740 58185 26744 58241
rect 26680 58181 26744 58185
rect 27768 58721 27832 58725
rect 27768 58665 27772 58721
rect 27772 58665 27828 58721
rect 27828 58665 27832 58721
rect 27768 58661 27832 58665
rect 27768 58641 27832 58645
rect 27768 58585 27772 58641
rect 27772 58585 27828 58641
rect 27828 58585 27832 58641
rect 27768 58581 27832 58585
rect 27768 58561 27832 58565
rect 27768 58505 27772 58561
rect 27772 58505 27828 58561
rect 27828 58505 27832 58561
rect 27768 58501 27832 58505
rect 27768 58481 27832 58485
rect 27768 58425 27772 58481
rect 27772 58425 27828 58481
rect 27828 58425 27832 58481
rect 27768 58421 27832 58425
rect 27768 58401 27832 58405
rect 27768 58345 27772 58401
rect 27772 58345 27828 58401
rect 27828 58345 27832 58401
rect 27768 58341 27832 58345
rect 27768 58321 27832 58325
rect 27768 58265 27772 58321
rect 27772 58265 27828 58321
rect 27828 58265 27832 58321
rect 27768 58261 27832 58265
rect 27768 58241 27832 58245
rect 27768 58185 27772 58241
rect 27772 58185 27828 58241
rect 27828 58185 27832 58241
rect 27768 58181 27832 58185
rect 28856 58721 28920 58725
rect 28856 58665 28860 58721
rect 28860 58665 28916 58721
rect 28916 58665 28920 58721
rect 28856 58661 28920 58665
rect 28856 58641 28920 58645
rect 28856 58585 28860 58641
rect 28860 58585 28916 58641
rect 28916 58585 28920 58641
rect 28856 58581 28920 58585
rect 28856 58561 28920 58565
rect 28856 58505 28860 58561
rect 28860 58505 28916 58561
rect 28916 58505 28920 58561
rect 28856 58501 28920 58505
rect 28856 58481 28920 58485
rect 28856 58425 28860 58481
rect 28860 58425 28916 58481
rect 28916 58425 28920 58481
rect 28856 58421 28920 58425
rect 28856 58401 28920 58405
rect 28856 58345 28860 58401
rect 28860 58345 28916 58401
rect 28916 58345 28920 58401
rect 28856 58341 28920 58345
rect 28856 58321 28920 58325
rect 28856 58265 28860 58321
rect 28860 58265 28916 58321
rect 28916 58265 28920 58321
rect 28856 58261 28920 58265
rect 28856 58241 28920 58245
rect 28856 58185 28860 58241
rect 28860 58185 28916 58241
rect 28916 58185 28920 58241
rect 28856 58181 28920 58185
rect 29944 58721 30008 58725
rect 29944 58665 29948 58721
rect 29948 58665 30004 58721
rect 30004 58665 30008 58721
rect 29944 58661 30008 58665
rect 29944 58641 30008 58645
rect 29944 58585 29948 58641
rect 29948 58585 30004 58641
rect 30004 58585 30008 58641
rect 29944 58581 30008 58585
rect 29944 58561 30008 58565
rect 29944 58505 29948 58561
rect 29948 58505 30004 58561
rect 30004 58505 30008 58561
rect 29944 58501 30008 58505
rect 29944 58481 30008 58485
rect 29944 58425 29948 58481
rect 29948 58425 30004 58481
rect 30004 58425 30008 58481
rect 29944 58421 30008 58425
rect 29944 58401 30008 58405
rect 29944 58345 29948 58401
rect 29948 58345 30004 58401
rect 30004 58345 30008 58401
rect 29944 58341 30008 58345
rect 29944 58321 30008 58325
rect 29944 58265 29948 58321
rect 29948 58265 30004 58321
rect 30004 58265 30008 58321
rect 29944 58261 30008 58265
rect 29944 58241 30008 58245
rect 29944 58185 29948 58241
rect 29948 58185 30004 58241
rect 30004 58185 30008 58241
rect 29944 58181 30008 58185
rect 31032 58721 31096 58725
rect 31032 58665 31036 58721
rect 31036 58665 31092 58721
rect 31092 58665 31096 58721
rect 31032 58661 31096 58665
rect 31032 58641 31096 58645
rect 31032 58585 31036 58641
rect 31036 58585 31092 58641
rect 31092 58585 31096 58641
rect 31032 58581 31096 58585
rect 31032 58561 31096 58565
rect 31032 58505 31036 58561
rect 31036 58505 31092 58561
rect 31092 58505 31096 58561
rect 31032 58501 31096 58505
rect 31032 58481 31096 58485
rect 31032 58425 31036 58481
rect 31036 58425 31092 58481
rect 31092 58425 31096 58481
rect 31032 58421 31096 58425
rect 31032 58401 31096 58405
rect 31032 58345 31036 58401
rect 31036 58345 31092 58401
rect 31092 58345 31096 58401
rect 31032 58341 31096 58345
rect 31032 58321 31096 58325
rect 31032 58265 31036 58321
rect 31036 58265 31092 58321
rect 31092 58265 31096 58321
rect 31032 58261 31096 58265
rect 31032 58241 31096 58245
rect 31032 58185 31036 58241
rect 31036 58185 31092 58241
rect 31092 58185 31096 58241
rect 31032 58181 31096 58185
rect 17431 56724 17495 56728
rect 17431 56668 17435 56724
rect 17435 56668 17491 56724
rect 17491 56668 17495 56724
rect 17431 56664 17495 56668
rect 17431 56644 17495 56648
rect 17431 56588 17435 56644
rect 17435 56588 17491 56644
rect 17491 56588 17495 56644
rect 17431 56584 17495 56588
rect 17431 56564 17495 56568
rect 17431 56508 17435 56564
rect 17435 56508 17491 56564
rect 17491 56508 17495 56564
rect 17431 56504 17495 56508
rect 17431 56484 17495 56488
rect 17431 56428 17435 56484
rect 17435 56428 17491 56484
rect 17491 56428 17495 56484
rect 17431 56424 17495 56428
rect 17431 56404 17495 56408
rect 17431 56348 17435 56404
rect 17435 56348 17491 56404
rect 17491 56348 17495 56404
rect 17431 56344 17495 56348
rect 17431 56324 17495 56328
rect 17431 56268 17435 56324
rect 17435 56268 17491 56324
rect 17491 56268 17495 56324
rect 17431 56264 17495 56268
rect 17431 56244 17495 56248
rect 17431 56188 17435 56244
rect 17435 56188 17491 56244
rect 17491 56188 17495 56244
rect 17431 56184 17495 56188
rect 18519 56724 18583 56728
rect 18519 56668 18523 56724
rect 18523 56668 18579 56724
rect 18579 56668 18583 56724
rect 18519 56664 18583 56668
rect 18519 56644 18583 56648
rect 18519 56588 18523 56644
rect 18523 56588 18579 56644
rect 18579 56588 18583 56644
rect 18519 56584 18583 56588
rect 18519 56564 18583 56568
rect 18519 56508 18523 56564
rect 18523 56508 18579 56564
rect 18579 56508 18583 56564
rect 18519 56504 18583 56508
rect 18519 56484 18583 56488
rect 18519 56428 18523 56484
rect 18523 56428 18579 56484
rect 18579 56428 18583 56484
rect 18519 56424 18583 56428
rect 18519 56404 18583 56408
rect 18519 56348 18523 56404
rect 18523 56348 18579 56404
rect 18579 56348 18583 56404
rect 18519 56344 18583 56348
rect 18519 56324 18583 56328
rect 18519 56268 18523 56324
rect 18523 56268 18579 56324
rect 18579 56268 18583 56324
rect 18519 56264 18583 56268
rect 18519 56244 18583 56248
rect 18519 56188 18523 56244
rect 18523 56188 18579 56244
rect 18579 56188 18583 56244
rect 18519 56184 18583 56188
rect 19607 56724 19671 56728
rect 19607 56668 19611 56724
rect 19611 56668 19667 56724
rect 19667 56668 19671 56724
rect 19607 56664 19671 56668
rect 19607 56644 19671 56648
rect 19607 56588 19611 56644
rect 19611 56588 19667 56644
rect 19667 56588 19671 56644
rect 19607 56584 19671 56588
rect 19607 56564 19671 56568
rect 19607 56508 19611 56564
rect 19611 56508 19667 56564
rect 19667 56508 19671 56564
rect 19607 56504 19671 56508
rect 19607 56484 19671 56488
rect 19607 56428 19611 56484
rect 19611 56428 19667 56484
rect 19667 56428 19671 56484
rect 19607 56424 19671 56428
rect 19607 56404 19671 56408
rect 19607 56348 19611 56404
rect 19611 56348 19667 56404
rect 19667 56348 19671 56404
rect 19607 56344 19671 56348
rect 19607 56324 19671 56328
rect 19607 56268 19611 56324
rect 19611 56268 19667 56324
rect 19667 56268 19671 56324
rect 19607 56264 19671 56268
rect 19607 56244 19671 56248
rect 19607 56188 19611 56244
rect 19611 56188 19667 56244
rect 19667 56188 19671 56244
rect 19607 56184 19671 56188
rect 20695 56724 20759 56728
rect 20695 56668 20699 56724
rect 20699 56668 20755 56724
rect 20755 56668 20759 56724
rect 20695 56664 20759 56668
rect 20695 56644 20759 56648
rect 20695 56588 20699 56644
rect 20699 56588 20755 56644
rect 20755 56588 20759 56644
rect 20695 56584 20759 56588
rect 20695 56564 20759 56568
rect 20695 56508 20699 56564
rect 20699 56508 20755 56564
rect 20755 56508 20759 56564
rect 20695 56504 20759 56508
rect 20695 56484 20759 56488
rect 20695 56428 20699 56484
rect 20699 56428 20755 56484
rect 20755 56428 20759 56484
rect 20695 56424 20759 56428
rect 20695 56404 20759 56408
rect 20695 56348 20699 56404
rect 20699 56348 20755 56404
rect 20755 56348 20759 56404
rect 20695 56344 20759 56348
rect 20695 56324 20759 56328
rect 20695 56268 20699 56324
rect 20699 56268 20755 56324
rect 20755 56268 20759 56324
rect 20695 56264 20759 56268
rect 20695 56244 20759 56248
rect 20695 56188 20699 56244
rect 20699 56188 20755 56244
rect 20755 56188 20759 56244
rect 20695 56184 20759 56188
rect 21783 56724 21847 56728
rect 21783 56668 21787 56724
rect 21787 56668 21843 56724
rect 21843 56668 21847 56724
rect 21783 56664 21847 56668
rect 21783 56644 21847 56648
rect 21783 56588 21787 56644
rect 21787 56588 21843 56644
rect 21843 56588 21847 56644
rect 21783 56584 21847 56588
rect 21783 56564 21847 56568
rect 21783 56508 21787 56564
rect 21787 56508 21843 56564
rect 21843 56508 21847 56564
rect 21783 56504 21847 56508
rect 21783 56484 21847 56488
rect 21783 56428 21787 56484
rect 21787 56428 21843 56484
rect 21843 56428 21847 56484
rect 21783 56424 21847 56428
rect 21783 56404 21847 56408
rect 21783 56348 21787 56404
rect 21787 56348 21843 56404
rect 21843 56348 21847 56404
rect 21783 56344 21847 56348
rect 21783 56324 21847 56328
rect 21783 56268 21787 56324
rect 21787 56268 21843 56324
rect 21843 56268 21847 56324
rect 21783 56264 21847 56268
rect 21783 56244 21847 56248
rect 21783 56188 21787 56244
rect 21787 56188 21843 56244
rect 21843 56188 21847 56244
rect 21783 56184 21847 56188
rect 22871 56724 22935 56728
rect 22871 56668 22875 56724
rect 22875 56668 22931 56724
rect 22931 56668 22935 56724
rect 22871 56664 22935 56668
rect 22871 56644 22935 56648
rect 22871 56588 22875 56644
rect 22875 56588 22931 56644
rect 22931 56588 22935 56644
rect 22871 56584 22935 56588
rect 22871 56564 22935 56568
rect 22871 56508 22875 56564
rect 22875 56508 22931 56564
rect 22931 56508 22935 56564
rect 22871 56504 22935 56508
rect 22871 56484 22935 56488
rect 22871 56428 22875 56484
rect 22875 56428 22931 56484
rect 22931 56428 22935 56484
rect 22871 56424 22935 56428
rect 22871 56404 22935 56408
rect 22871 56348 22875 56404
rect 22875 56348 22931 56404
rect 22931 56348 22935 56404
rect 22871 56344 22935 56348
rect 22871 56324 22935 56328
rect 22871 56268 22875 56324
rect 22875 56268 22931 56324
rect 22931 56268 22935 56324
rect 22871 56264 22935 56268
rect 22871 56244 22935 56248
rect 22871 56188 22875 56244
rect 22875 56188 22931 56244
rect 22931 56188 22935 56244
rect 22871 56184 22935 56188
rect 23959 56724 24023 56728
rect 23959 56668 23963 56724
rect 23963 56668 24019 56724
rect 24019 56668 24023 56724
rect 23959 56664 24023 56668
rect 23959 56644 24023 56648
rect 23959 56588 23963 56644
rect 23963 56588 24019 56644
rect 24019 56588 24023 56644
rect 23959 56584 24023 56588
rect 23959 56564 24023 56568
rect 23959 56508 23963 56564
rect 23963 56508 24019 56564
rect 24019 56508 24023 56564
rect 23959 56504 24023 56508
rect 23959 56484 24023 56488
rect 23959 56428 23963 56484
rect 23963 56428 24019 56484
rect 24019 56428 24023 56484
rect 23959 56424 24023 56428
rect 23959 56404 24023 56408
rect 23959 56348 23963 56404
rect 23963 56348 24019 56404
rect 24019 56348 24023 56404
rect 23959 56344 24023 56348
rect 23959 56324 24023 56328
rect 23959 56268 23963 56324
rect 23963 56268 24019 56324
rect 24019 56268 24023 56324
rect 23959 56264 24023 56268
rect 23959 56244 24023 56248
rect 23959 56188 23963 56244
rect 23963 56188 24019 56244
rect 24019 56188 24023 56244
rect 23959 56184 24023 56188
rect 25047 56724 25111 56728
rect 25047 56668 25051 56724
rect 25051 56668 25107 56724
rect 25107 56668 25111 56724
rect 25047 56664 25111 56668
rect 25047 56644 25111 56648
rect 25047 56588 25051 56644
rect 25051 56588 25107 56644
rect 25107 56588 25111 56644
rect 25047 56584 25111 56588
rect 25047 56564 25111 56568
rect 25047 56508 25051 56564
rect 25051 56508 25107 56564
rect 25107 56508 25111 56564
rect 25047 56504 25111 56508
rect 25047 56484 25111 56488
rect 25047 56428 25051 56484
rect 25051 56428 25107 56484
rect 25107 56428 25111 56484
rect 25047 56424 25111 56428
rect 25047 56404 25111 56408
rect 25047 56348 25051 56404
rect 25051 56348 25107 56404
rect 25107 56348 25111 56404
rect 25047 56344 25111 56348
rect 25047 56324 25111 56328
rect 25047 56268 25051 56324
rect 25051 56268 25107 56324
rect 25107 56268 25111 56324
rect 25047 56264 25111 56268
rect 25047 56244 25111 56248
rect 25047 56188 25051 56244
rect 25051 56188 25107 56244
rect 25107 56188 25111 56244
rect 25047 56184 25111 56188
rect 26135 56724 26199 56728
rect 26135 56668 26139 56724
rect 26139 56668 26195 56724
rect 26195 56668 26199 56724
rect 26135 56664 26199 56668
rect 26135 56644 26199 56648
rect 26135 56588 26139 56644
rect 26139 56588 26195 56644
rect 26195 56588 26199 56644
rect 26135 56584 26199 56588
rect 26135 56564 26199 56568
rect 26135 56508 26139 56564
rect 26139 56508 26195 56564
rect 26195 56508 26199 56564
rect 26135 56504 26199 56508
rect 26135 56484 26199 56488
rect 26135 56428 26139 56484
rect 26139 56428 26195 56484
rect 26195 56428 26199 56484
rect 26135 56424 26199 56428
rect 26135 56404 26199 56408
rect 26135 56348 26139 56404
rect 26139 56348 26195 56404
rect 26195 56348 26199 56404
rect 26135 56344 26199 56348
rect 26135 56324 26199 56328
rect 26135 56268 26139 56324
rect 26139 56268 26195 56324
rect 26195 56268 26199 56324
rect 26135 56264 26199 56268
rect 26135 56244 26199 56248
rect 26135 56188 26139 56244
rect 26139 56188 26195 56244
rect 26195 56188 26199 56244
rect 26135 56184 26199 56188
rect 27223 56724 27287 56728
rect 27223 56668 27227 56724
rect 27227 56668 27283 56724
rect 27283 56668 27287 56724
rect 27223 56664 27287 56668
rect 27223 56644 27287 56648
rect 27223 56588 27227 56644
rect 27227 56588 27283 56644
rect 27283 56588 27287 56644
rect 27223 56584 27287 56588
rect 27223 56564 27287 56568
rect 27223 56508 27227 56564
rect 27227 56508 27283 56564
rect 27283 56508 27287 56564
rect 27223 56504 27287 56508
rect 27223 56484 27287 56488
rect 27223 56428 27227 56484
rect 27227 56428 27283 56484
rect 27283 56428 27287 56484
rect 27223 56424 27287 56428
rect 27223 56404 27287 56408
rect 27223 56348 27227 56404
rect 27227 56348 27283 56404
rect 27283 56348 27287 56404
rect 27223 56344 27287 56348
rect 27223 56324 27287 56328
rect 27223 56268 27227 56324
rect 27227 56268 27283 56324
rect 27283 56268 27287 56324
rect 27223 56264 27287 56268
rect 27223 56244 27287 56248
rect 27223 56188 27227 56244
rect 27227 56188 27283 56244
rect 27283 56188 27287 56244
rect 27223 56184 27287 56188
rect 28311 56724 28375 56728
rect 28311 56668 28315 56724
rect 28315 56668 28371 56724
rect 28371 56668 28375 56724
rect 28311 56664 28375 56668
rect 28311 56644 28375 56648
rect 28311 56588 28315 56644
rect 28315 56588 28371 56644
rect 28371 56588 28375 56644
rect 28311 56584 28375 56588
rect 28311 56564 28375 56568
rect 28311 56508 28315 56564
rect 28315 56508 28371 56564
rect 28371 56508 28375 56564
rect 28311 56504 28375 56508
rect 28311 56484 28375 56488
rect 28311 56428 28315 56484
rect 28315 56428 28371 56484
rect 28371 56428 28375 56484
rect 28311 56424 28375 56428
rect 28311 56404 28375 56408
rect 28311 56348 28315 56404
rect 28315 56348 28371 56404
rect 28371 56348 28375 56404
rect 28311 56344 28375 56348
rect 28311 56324 28375 56328
rect 28311 56268 28315 56324
rect 28315 56268 28371 56324
rect 28371 56268 28375 56324
rect 28311 56264 28375 56268
rect 28311 56244 28375 56248
rect 28311 56188 28315 56244
rect 28315 56188 28371 56244
rect 28371 56188 28375 56244
rect 28311 56184 28375 56188
rect 29399 56724 29463 56728
rect 29399 56668 29403 56724
rect 29403 56668 29459 56724
rect 29459 56668 29463 56724
rect 29399 56664 29463 56668
rect 29399 56644 29463 56648
rect 29399 56588 29403 56644
rect 29403 56588 29459 56644
rect 29459 56588 29463 56644
rect 29399 56584 29463 56588
rect 29399 56564 29463 56568
rect 29399 56508 29403 56564
rect 29403 56508 29459 56564
rect 29459 56508 29463 56564
rect 29399 56504 29463 56508
rect 29399 56484 29463 56488
rect 29399 56428 29403 56484
rect 29403 56428 29459 56484
rect 29459 56428 29463 56484
rect 29399 56424 29463 56428
rect 29399 56404 29463 56408
rect 29399 56348 29403 56404
rect 29403 56348 29459 56404
rect 29459 56348 29463 56404
rect 29399 56344 29463 56348
rect 29399 56324 29463 56328
rect 29399 56268 29403 56324
rect 29403 56268 29459 56324
rect 29459 56268 29463 56324
rect 29399 56264 29463 56268
rect 29399 56244 29463 56248
rect 29399 56188 29403 56244
rect 29403 56188 29459 56244
rect 29459 56188 29463 56244
rect 29399 56184 29463 56188
rect 30487 56724 30551 56728
rect 30487 56668 30491 56724
rect 30491 56668 30547 56724
rect 30547 56668 30551 56724
rect 30487 56664 30551 56668
rect 30487 56644 30551 56648
rect 30487 56588 30491 56644
rect 30491 56588 30547 56644
rect 30547 56588 30551 56644
rect 30487 56584 30551 56588
rect 30487 56564 30551 56568
rect 30487 56508 30491 56564
rect 30491 56508 30547 56564
rect 30547 56508 30551 56564
rect 30487 56504 30551 56508
rect 30487 56484 30551 56488
rect 30487 56428 30491 56484
rect 30491 56428 30547 56484
rect 30547 56428 30551 56484
rect 30487 56424 30551 56428
rect 30487 56404 30551 56408
rect 30487 56348 30491 56404
rect 30491 56348 30547 56404
rect 30547 56348 30551 56404
rect 30487 56344 30551 56348
rect 30487 56324 30551 56328
rect 30487 56268 30491 56324
rect 30491 56268 30547 56324
rect 30547 56268 30551 56324
rect 30487 56264 30551 56268
rect 30487 56244 30551 56248
rect 30487 56188 30491 56244
rect 30491 56188 30547 56244
rect 30547 56188 30551 56244
rect 30487 56184 30551 56188
rect 31575 56724 31639 56728
rect 31575 56668 31579 56724
rect 31579 56668 31635 56724
rect 31635 56668 31639 56724
rect 31575 56664 31639 56668
rect 31575 56644 31639 56648
rect 31575 56588 31579 56644
rect 31579 56588 31635 56644
rect 31635 56588 31639 56644
rect 31575 56584 31639 56588
rect 31575 56564 31639 56568
rect 31575 56508 31579 56564
rect 31579 56508 31635 56564
rect 31635 56508 31639 56564
rect 31575 56504 31639 56508
rect 31575 56484 31639 56488
rect 31575 56428 31579 56484
rect 31579 56428 31635 56484
rect 31635 56428 31639 56484
rect 31575 56424 31639 56428
rect 31575 56404 31639 56408
rect 31575 56348 31579 56404
rect 31579 56348 31635 56404
rect 31635 56348 31639 56404
rect 31575 56344 31639 56348
rect 31575 56324 31639 56328
rect 31575 56268 31579 56324
rect 31579 56268 31635 56324
rect 31635 56268 31639 56324
rect 31575 56264 31639 56268
rect 31575 56244 31639 56248
rect 31575 56188 31579 56244
rect 31579 56188 31635 56244
rect 31635 56188 31639 56244
rect 31575 56184 31639 56188
rect 17976 54721 18040 54725
rect 17976 54665 17980 54721
rect 17980 54665 18036 54721
rect 18036 54665 18040 54721
rect 17976 54661 18040 54665
rect 17976 54641 18040 54645
rect 17976 54585 17980 54641
rect 17980 54585 18036 54641
rect 18036 54585 18040 54641
rect 17976 54581 18040 54585
rect 17976 54561 18040 54565
rect 17976 54505 17980 54561
rect 17980 54505 18036 54561
rect 18036 54505 18040 54561
rect 17976 54501 18040 54505
rect 17976 54481 18040 54485
rect 17976 54425 17980 54481
rect 17980 54425 18036 54481
rect 18036 54425 18040 54481
rect 17976 54421 18040 54425
rect 17976 54401 18040 54405
rect 17976 54345 17980 54401
rect 17980 54345 18036 54401
rect 18036 54345 18040 54401
rect 17976 54341 18040 54345
rect 17976 54321 18040 54325
rect 17976 54265 17980 54321
rect 17980 54265 18036 54321
rect 18036 54265 18040 54321
rect 17976 54261 18040 54265
rect 17976 54241 18040 54245
rect 17976 54185 17980 54241
rect 17980 54185 18036 54241
rect 18036 54185 18040 54241
rect 17976 54181 18040 54185
rect 19064 54721 19128 54725
rect 19064 54665 19068 54721
rect 19068 54665 19124 54721
rect 19124 54665 19128 54721
rect 19064 54661 19128 54665
rect 19064 54641 19128 54645
rect 19064 54585 19068 54641
rect 19068 54585 19124 54641
rect 19124 54585 19128 54641
rect 19064 54581 19128 54585
rect 19064 54561 19128 54565
rect 19064 54505 19068 54561
rect 19068 54505 19124 54561
rect 19124 54505 19128 54561
rect 19064 54501 19128 54505
rect 19064 54481 19128 54485
rect 19064 54425 19068 54481
rect 19068 54425 19124 54481
rect 19124 54425 19128 54481
rect 19064 54421 19128 54425
rect 19064 54401 19128 54405
rect 19064 54345 19068 54401
rect 19068 54345 19124 54401
rect 19124 54345 19128 54401
rect 19064 54341 19128 54345
rect 19064 54321 19128 54325
rect 19064 54265 19068 54321
rect 19068 54265 19124 54321
rect 19124 54265 19128 54321
rect 19064 54261 19128 54265
rect 19064 54241 19128 54245
rect 19064 54185 19068 54241
rect 19068 54185 19124 54241
rect 19124 54185 19128 54241
rect 19064 54181 19128 54185
rect 20152 54721 20216 54725
rect 20152 54665 20156 54721
rect 20156 54665 20212 54721
rect 20212 54665 20216 54721
rect 20152 54661 20216 54665
rect 20152 54641 20216 54645
rect 20152 54585 20156 54641
rect 20156 54585 20212 54641
rect 20212 54585 20216 54641
rect 20152 54581 20216 54585
rect 20152 54561 20216 54565
rect 20152 54505 20156 54561
rect 20156 54505 20212 54561
rect 20212 54505 20216 54561
rect 20152 54501 20216 54505
rect 20152 54481 20216 54485
rect 20152 54425 20156 54481
rect 20156 54425 20212 54481
rect 20212 54425 20216 54481
rect 20152 54421 20216 54425
rect 20152 54401 20216 54405
rect 20152 54345 20156 54401
rect 20156 54345 20212 54401
rect 20212 54345 20216 54401
rect 20152 54341 20216 54345
rect 20152 54321 20216 54325
rect 20152 54265 20156 54321
rect 20156 54265 20212 54321
rect 20212 54265 20216 54321
rect 20152 54261 20216 54265
rect 20152 54241 20216 54245
rect 20152 54185 20156 54241
rect 20156 54185 20212 54241
rect 20212 54185 20216 54241
rect 20152 54181 20216 54185
rect 21240 54721 21304 54725
rect 21240 54665 21244 54721
rect 21244 54665 21300 54721
rect 21300 54665 21304 54721
rect 21240 54661 21304 54665
rect 21240 54641 21304 54645
rect 21240 54585 21244 54641
rect 21244 54585 21300 54641
rect 21300 54585 21304 54641
rect 21240 54581 21304 54585
rect 21240 54561 21304 54565
rect 21240 54505 21244 54561
rect 21244 54505 21300 54561
rect 21300 54505 21304 54561
rect 21240 54501 21304 54505
rect 21240 54481 21304 54485
rect 21240 54425 21244 54481
rect 21244 54425 21300 54481
rect 21300 54425 21304 54481
rect 21240 54421 21304 54425
rect 21240 54401 21304 54405
rect 21240 54345 21244 54401
rect 21244 54345 21300 54401
rect 21300 54345 21304 54401
rect 21240 54341 21304 54345
rect 21240 54321 21304 54325
rect 21240 54265 21244 54321
rect 21244 54265 21300 54321
rect 21300 54265 21304 54321
rect 21240 54261 21304 54265
rect 21240 54241 21304 54245
rect 21240 54185 21244 54241
rect 21244 54185 21300 54241
rect 21300 54185 21304 54241
rect 21240 54181 21304 54185
rect 22328 54721 22392 54725
rect 22328 54665 22332 54721
rect 22332 54665 22388 54721
rect 22388 54665 22392 54721
rect 22328 54661 22392 54665
rect 22328 54641 22392 54645
rect 22328 54585 22332 54641
rect 22332 54585 22388 54641
rect 22388 54585 22392 54641
rect 22328 54581 22392 54585
rect 22328 54561 22392 54565
rect 22328 54505 22332 54561
rect 22332 54505 22388 54561
rect 22388 54505 22392 54561
rect 22328 54501 22392 54505
rect 22328 54481 22392 54485
rect 22328 54425 22332 54481
rect 22332 54425 22388 54481
rect 22388 54425 22392 54481
rect 22328 54421 22392 54425
rect 22328 54401 22392 54405
rect 22328 54345 22332 54401
rect 22332 54345 22388 54401
rect 22388 54345 22392 54401
rect 22328 54341 22392 54345
rect 22328 54321 22392 54325
rect 22328 54265 22332 54321
rect 22332 54265 22388 54321
rect 22388 54265 22392 54321
rect 22328 54261 22392 54265
rect 22328 54241 22392 54245
rect 22328 54185 22332 54241
rect 22332 54185 22388 54241
rect 22388 54185 22392 54241
rect 22328 54181 22392 54185
rect 23416 54721 23480 54725
rect 23416 54665 23420 54721
rect 23420 54665 23476 54721
rect 23476 54665 23480 54721
rect 23416 54661 23480 54665
rect 23416 54641 23480 54645
rect 23416 54585 23420 54641
rect 23420 54585 23476 54641
rect 23476 54585 23480 54641
rect 23416 54581 23480 54585
rect 23416 54561 23480 54565
rect 23416 54505 23420 54561
rect 23420 54505 23476 54561
rect 23476 54505 23480 54561
rect 23416 54501 23480 54505
rect 23416 54481 23480 54485
rect 23416 54425 23420 54481
rect 23420 54425 23476 54481
rect 23476 54425 23480 54481
rect 23416 54421 23480 54425
rect 23416 54401 23480 54405
rect 23416 54345 23420 54401
rect 23420 54345 23476 54401
rect 23476 54345 23480 54401
rect 23416 54341 23480 54345
rect 23416 54321 23480 54325
rect 23416 54265 23420 54321
rect 23420 54265 23476 54321
rect 23476 54265 23480 54321
rect 23416 54261 23480 54265
rect 23416 54241 23480 54245
rect 23416 54185 23420 54241
rect 23420 54185 23476 54241
rect 23476 54185 23480 54241
rect 23416 54181 23480 54185
rect 24504 54721 24568 54725
rect 24504 54665 24508 54721
rect 24508 54665 24564 54721
rect 24564 54665 24568 54721
rect 24504 54661 24568 54665
rect 24504 54641 24568 54645
rect 24504 54585 24508 54641
rect 24508 54585 24564 54641
rect 24564 54585 24568 54641
rect 24504 54581 24568 54585
rect 24504 54561 24568 54565
rect 24504 54505 24508 54561
rect 24508 54505 24564 54561
rect 24564 54505 24568 54561
rect 24504 54501 24568 54505
rect 24504 54481 24568 54485
rect 24504 54425 24508 54481
rect 24508 54425 24564 54481
rect 24564 54425 24568 54481
rect 24504 54421 24568 54425
rect 24504 54401 24568 54405
rect 24504 54345 24508 54401
rect 24508 54345 24564 54401
rect 24564 54345 24568 54401
rect 24504 54341 24568 54345
rect 24504 54321 24568 54325
rect 24504 54265 24508 54321
rect 24508 54265 24564 54321
rect 24564 54265 24568 54321
rect 24504 54261 24568 54265
rect 24504 54241 24568 54245
rect 24504 54185 24508 54241
rect 24508 54185 24564 54241
rect 24564 54185 24568 54241
rect 24504 54181 24568 54185
rect 25592 54721 25656 54725
rect 25592 54665 25596 54721
rect 25596 54665 25652 54721
rect 25652 54665 25656 54721
rect 25592 54661 25656 54665
rect 25592 54641 25656 54645
rect 25592 54585 25596 54641
rect 25596 54585 25652 54641
rect 25652 54585 25656 54641
rect 25592 54581 25656 54585
rect 25592 54561 25656 54565
rect 25592 54505 25596 54561
rect 25596 54505 25652 54561
rect 25652 54505 25656 54561
rect 25592 54501 25656 54505
rect 25592 54481 25656 54485
rect 25592 54425 25596 54481
rect 25596 54425 25652 54481
rect 25652 54425 25656 54481
rect 25592 54421 25656 54425
rect 25592 54401 25656 54405
rect 25592 54345 25596 54401
rect 25596 54345 25652 54401
rect 25652 54345 25656 54401
rect 25592 54341 25656 54345
rect 25592 54321 25656 54325
rect 25592 54265 25596 54321
rect 25596 54265 25652 54321
rect 25652 54265 25656 54321
rect 25592 54261 25656 54265
rect 25592 54241 25656 54245
rect 25592 54185 25596 54241
rect 25596 54185 25652 54241
rect 25652 54185 25656 54241
rect 25592 54181 25656 54185
rect 26680 54721 26744 54725
rect 26680 54665 26684 54721
rect 26684 54665 26740 54721
rect 26740 54665 26744 54721
rect 26680 54661 26744 54665
rect 26680 54641 26744 54645
rect 26680 54585 26684 54641
rect 26684 54585 26740 54641
rect 26740 54585 26744 54641
rect 26680 54581 26744 54585
rect 26680 54561 26744 54565
rect 26680 54505 26684 54561
rect 26684 54505 26740 54561
rect 26740 54505 26744 54561
rect 26680 54501 26744 54505
rect 26680 54481 26744 54485
rect 26680 54425 26684 54481
rect 26684 54425 26740 54481
rect 26740 54425 26744 54481
rect 26680 54421 26744 54425
rect 26680 54401 26744 54405
rect 26680 54345 26684 54401
rect 26684 54345 26740 54401
rect 26740 54345 26744 54401
rect 26680 54341 26744 54345
rect 26680 54321 26744 54325
rect 26680 54265 26684 54321
rect 26684 54265 26740 54321
rect 26740 54265 26744 54321
rect 26680 54261 26744 54265
rect 26680 54241 26744 54245
rect 26680 54185 26684 54241
rect 26684 54185 26740 54241
rect 26740 54185 26744 54241
rect 26680 54181 26744 54185
rect 27768 54721 27832 54725
rect 27768 54665 27772 54721
rect 27772 54665 27828 54721
rect 27828 54665 27832 54721
rect 27768 54661 27832 54665
rect 27768 54641 27832 54645
rect 27768 54585 27772 54641
rect 27772 54585 27828 54641
rect 27828 54585 27832 54641
rect 27768 54581 27832 54585
rect 27768 54561 27832 54565
rect 27768 54505 27772 54561
rect 27772 54505 27828 54561
rect 27828 54505 27832 54561
rect 27768 54501 27832 54505
rect 27768 54481 27832 54485
rect 27768 54425 27772 54481
rect 27772 54425 27828 54481
rect 27828 54425 27832 54481
rect 27768 54421 27832 54425
rect 27768 54401 27832 54405
rect 27768 54345 27772 54401
rect 27772 54345 27828 54401
rect 27828 54345 27832 54401
rect 27768 54341 27832 54345
rect 27768 54321 27832 54325
rect 27768 54265 27772 54321
rect 27772 54265 27828 54321
rect 27828 54265 27832 54321
rect 27768 54261 27832 54265
rect 27768 54241 27832 54245
rect 27768 54185 27772 54241
rect 27772 54185 27828 54241
rect 27828 54185 27832 54241
rect 27768 54181 27832 54185
rect 28856 54721 28920 54725
rect 28856 54665 28860 54721
rect 28860 54665 28916 54721
rect 28916 54665 28920 54721
rect 28856 54661 28920 54665
rect 28856 54641 28920 54645
rect 28856 54585 28860 54641
rect 28860 54585 28916 54641
rect 28916 54585 28920 54641
rect 28856 54581 28920 54585
rect 28856 54561 28920 54565
rect 28856 54505 28860 54561
rect 28860 54505 28916 54561
rect 28916 54505 28920 54561
rect 28856 54501 28920 54505
rect 28856 54481 28920 54485
rect 28856 54425 28860 54481
rect 28860 54425 28916 54481
rect 28916 54425 28920 54481
rect 28856 54421 28920 54425
rect 28856 54401 28920 54405
rect 28856 54345 28860 54401
rect 28860 54345 28916 54401
rect 28916 54345 28920 54401
rect 28856 54341 28920 54345
rect 28856 54321 28920 54325
rect 28856 54265 28860 54321
rect 28860 54265 28916 54321
rect 28916 54265 28920 54321
rect 28856 54261 28920 54265
rect 28856 54241 28920 54245
rect 28856 54185 28860 54241
rect 28860 54185 28916 54241
rect 28916 54185 28920 54241
rect 28856 54181 28920 54185
rect 29944 54721 30008 54725
rect 29944 54665 29948 54721
rect 29948 54665 30004 54721
rect 30004 54665 30008 54721
rect 29944 54661 30008 54665
rect 29944 54641 30008 54645
rect 29944 54585 29948 54641
rect 29948 54585 30004 54641
rect 30004 54585 30008 54641
rect 29944 54581 30008 54585
rect 29944 54561 30008 54565
rect 29944 54505 29948 54561
rect 29948 54505 30004 54561
rect 30004 54505 30008 54561
rect 29944 54501 30008 54505
rect 29944 54481 30008 54485
rect 29944 54425 29948 54481
rect 29948 54425 30004 54481
rect 30004 54425 30008 54481
rect 29944 54421 30008 54425
rect 29944 54401 30008 54405
rect 29944 54345 29948 54401
rect 29948 54345 30004 54401
rect 30004 54345 30008 54401
rect 29944 54341 30008 54345
rect 29944 54321 30008 54325
rect 29944 54265 29948 54321
rect 29948 54265 30004 54321
rect 30004 54265 30008 54321
rect 29944 54261 30008 54265
rect 29944 54241 30008 54245
rect 29944 54185 29948 54241
rect 29948 54185 30004 54241
rect 30004 54185 30008 54241
rect 29944 54181 30008 54185
rect 31032 54721 31096 54725
rect 31032 54665 31036 54721
rect 31036 54665 31092 54721
rect 31092 54665 31096 54721
rect 31032 54661 31096 54665
rect 31032 54641 31096 54645
rect 31032 54585 31036 54641
rect 31036 54585 31092 54641
rect 31092 54585 31096 54641
rect 31032 54581 31096 54585
rect 31032 54561 31096 54565
rect 31032 54505 31036 54561
rect 31036 54505 31092 54561
rect 31092 54505 31096 54561
rect 31032 54501 31096 54505
rect 31032 54481 31096 54485
rect 31032 54425 31036 54481
rect 31036 54425 31092 54481
rect 31092 54425 31096 54481
rect 31032 54421 31096 54425
rect 31032 54401 31096 54405
rect 31032 54345 31036 54401
rect 31036 54345 31092 54401
rect 31092 54345 31096 54401
rect 31032 54341 31096 54345
rect 31032 54321 31096 54325
rect 31032 54265 31036 54321
rect 31036 54265 31092 54321
rect 31092 54265 31096 54321
rect 31032 54261 31096 54265
rect 31032 54241 31096 54245
rect 31032 54185 31036 54241
rect 31036 54185 31092 54241
rect 31092 54185 31096 54241
rect 31032 54181 31096 54185
rect 17431 52724 17495 52728
rect 17431 52668 17435 52724
rect 17435 52668 17491 52724
rect 17491 52668 17495 52724
rect 17431 52664 17495 52668
rect 17431 52644 17495 52648
rect 17431 52588 17435 52644
rect 17435 52588 17491 52644
rect 17491 52588 17495 52644
rect 17431 52584 17495 52588
rect 17431 52564 17495 52568
rect 17431 52508 17435 52564
rect 17435 52508 17491 52564
rect 17491 52508 17495 52564
rect 17431 52504 17495 52508
rect 17431 52484 17495 52488
rect 17431 52428 17435 52484
rect 17435 52428 17491 52484
rect 17491 52428 17495 52484
rect 17431 52424 17495 52428
rect 17431 52404 17495 52408
rect 17431 52348 17435 52404
rect 17435 52348 17491 52404
rect 17491 52348 17495 52404
rect 17431 52344 17495 52348
rect 17431 52324 17495 52328
rect 17431 52268 17435 52324
rect 17435 52268 17491 52324
rect 17491 52268 17495 52324
rect 17431 52264 17495 52268
rect 17431 52244 17495 52248
rect 17431 52188 17435 52244
rect 17435 52188 17491 52244
rect 17491 52188 17495 52244
rect 17431 52184 17495 52188
rect 18519 52724 18583 52728
rect 18519 52668 18523 52724
rect 18523 52668 18579 52724
rect 18579 52668 18583 52724
rect 18519 52664 18583 52668
rect 18519 52644 18583 52648
rect 18519 52588 18523 52644
rect 18523 52588 18579 52644
rect 18579 52588 18583 52644
rect 18519 52584 18583 52588
rect 18519 52564 18583 52568
rect 18519 52508 18523 52564
rect 18523 52508 18579 52564
rect 18579 52508 18583 52564
rect 18519 52504 18583 52508
rect 18519 52484 18583 52488
rect 18519 52428 18523 52484
rect 18523 52428 18579 52484
rect 18579 52428 18583 52484
rect 18519 52424 18583 52428
rect 18519 52404 18583 52408
rect 18519 52348 18523 52404
rect 18523 52348 18579 52404
rect 18579 52348 18583 52404
rect 18519 52344 18583 52348
rect 18519 52324 18583 52328
rect 18519 52268 18523 52324
rect 18523 52268 18579 52324
rect 18579 52268 18583 52324
rect 18519 52264 18583 52268
rect 18519 52244 18583 52248
rect 18519 52188 18523 52244
rect 18523 52188 18579 52244
rect 18579 52188 18583 52244
rect 18519 52184 18583 52188
rect 19607 52724 19671 52728
rect 19607 52668 19611 52724
rect 19611 52668 19667 52724
rect 19667 52668 19671 52724
rect 19607 52664 19671 52668
rect 19607 52644 19671 52648
rect 19607 52588 19611 52644
rect 19611 52588 19667 52644
rect 19667 52588 19671 52644
rect 19607 52584 19671 52588
rect 19607 52564 19671 52568
rect 19607 52508 19611 52564
rect 19611 52508 19667 52564
rect 19667 52508 19671 52564
rect 19607 52504 19671 52508
rect 19607 52484 19671 52488
rect 19607 52428 19611 52484
rect 19611 52428 19667 52484
rect 19667 52428 19671 52484
rect 19607 52424 19671 52428
rect 19607 52404 19671 52408
rect 19607 52348 19611 52404
rect 19611 52348 19667 52404
rect 19667 52348 19671 52404
rect 19607 52344 19671 52348
rect 19607 52324 19671 52328
rect 19607 52268 19611 52324
rect 19611 52268 19667 52324
rect 19667 52268 19671 52324
rect 19607 52264 19671 52268
rect 19607 52244 19671 52248
rect 19607 52188 19611 52244
rect 19611 52188 19667 52244
rect 19667 52188 19671 52244
rect 19607 52184 19671 52188
rect 20695 52724 20759 52728
rect 20695 52668 20699 52724
rect 20699 52668 20755 52724
rect 20755 52668 20759 52724
rect 20695 52664 20759 52668
rect 20695 52644 20759 52648
rect 20695 52588 20699 52644
rect 20699 52588 20755 52644
rect 20755 52588 20759 52644
rect 20695 52584 20759 52588
rect 20695 52564 20759 52568
rect 20695 52508 20699 52564
rect 20699 52508 20755 52564
rect 20755 52508 20759 52564
rect 20695 52504 20759 52508
rect 20695 52484 20759 52488
rect 20695 52428 20699 52484
rect 20699 52428 20755 52484
rect 20755 52428 20759 52484
rect 20695 52424 20759 52428
rect 20695 52404 20759 52408
rect 20695 52348 20699 52404
rect 20699 52348 20755 52404
rect 20755 52348 20759 52404
rect 20695 52344 20759 52348
rect 20695 52324 20759 52328
rect 20695 52268 20699 52324
rect 20699 52268 20755 52324
rect 20755 52268 20759 52324
rect 20695 52264 20759 52268
rect 20695 52244 20759 52248
rect 20695 52188 20699 52244
rect 20699 52188 20755 52244
rect 20755 52188 20759 52244
rect 20695 52184 20759 52188
rect 21783 52724 21847 52728
rect 21783 52668 21787 52724
rect 21787 52668 21843 52724
rect 21843 52668 21847 52724
rect 21783 52664 21847 52668
rect 21783 52644 21847 52648
rect 21783 52588 21787 52644
rect 21787 52588 21843 52644
rect 21843 52588 21847 52644
rect 21783 52584 21847 52588
rect 21783 52564 21847 52568
rect 21783 52508 21787 52564
rect 21787 52508 21843 52564
rect 21843 52508 21847 52564
rect 21783 52504 21847 52508
rect 21783 52484 21847 52488
rect 21783 52428 21787 52484
rect 21787 52428 21843 52484
rect 21843 52428 21847 52484
rect 21783 52424 21847 52428
rect 21783 52404 21847 52408
rect 21783 52348 21787 52404
rect 21787 52348 21843 52404
rect 21843 52348 21847 52404
rect 21783 52344 21847 52348
rect 21783 52324 21847 52328
rect 21783 52268 21787 52324
rect 21787 52268 21843 52324
rect 21843 52268 21847 52324
rect 21783 52264 21847 52268
rect 21783 52244 21847 52248
rect 21783 52188 21787 52244
rect 21787 52188 21843 52244
rect 21843 52188 21847 52244
rect 21783 52184 21847 52188
rect 22871 52724 22935 52728
rect 22871 52668 22875 52724
rect 22875 52668 22931 52724
rect 22931 52668 22935 52724
rect 22871 52664 22935 52668
rect 22871 52644 22935 52648
rect 22871 52588 22875 52644
rect 22875 52588 22931 52644
rect 22931 52588 22935 52644
rect 22871 52584 22935 52588
rect 22871 52564 22935 52568
rect 22871 52508 22875 52564
rect 22875 52508 22931 52564
rect 22931 52508 22935 52564
rect 22871 52504 22935 52508
rect 22871 52484 22935 52488
rect 22871 52428 22875 52484
rect 22875 52428 22931 52484
rect 22931 52428 22935 52484
rect 22871 52424 22935 52428
rect 22871 52404 22935 52408
rect 22871 52348 22875 52404
rect 22875 52348 22931 52404
rect 22931 52348 22935 52404
rect 22871 52344 22935 52348
rect 22871 52324 22935 52328
rect 22871 52268 22875 52324
rect 22875 52268 22931 52324
rect 22931 52268 22935 52324
rect 22871 52264 22935 52268
rect 22871 52244 22935 52248
rect 22871 52188 22875 52244
rect 22875 52188 22931 52244
rect 22931 52188 22935 52244
rect 22871 52184 22935 52188
rect 23959 52724 24023 52728
rect 23959 52668 23963 52724
rect 23963 52668 24019 52724
rect 24019 52668 24023 52724
rect 23959 52664 24023 52668
rect 23959 52644 24023 52648
rect 23959 52588 23963 52644
rect 23963 52588 24019 52644
rect 24019 52588 24023 52644
rect 23959 52584 24023 52588
rect 23959 52564 24023 52568
rect 23959 52508 23963 52564
rect 23963 52508 24019 52564
rect 24019 52508 24023 52564
rect 23959 52504 24023 52508
rect 23959 52484 24023 52488
rect 23959 52428 23963 52484
rect 23963 52428 24019 52484
rect 24019 52428 24023 52484
rect 23959 52424 24023 52428
rect 23959 52404 24023 52408
rect 23959 52348 23963 52404
rect 23963 52348 24019 52404
rect 24019 52348 24023 52404
rect 23959 52344 24023 52348
rect 23959 52324 24023 52328
rect 23959 52268 23963 52324
rect 23963 52268 24019 52324
rect 24019 52268 24023 52324
rect 23959 52264 24023 52268
rect 23959 52244 24023 52248
rect 23959 52188 23963 52244
rect 23963 52188 24019 52244
rect 24019 52188 24023 52244
rect 23959 52184 24023 52188
rect 25047 52724 25111 52728
rect 25047 52668 25051 52724
rect 25051 52668 25107 52724
rect 25107 52668 25111 52724
rect 25047 52664 25111 52668
rect 25047 52644 25111 52648
rect 25047 52588 25051 52644
rect 25051 52588 25107 52644
rect 25107 52588 25111 52644
rect 25047 52584 25111 52588
rect 25047 52564 25111 52568
rect 25047 52508 25051 52564
rect 25051 52508 25107 52564
rect 25107 52508 25111 52564
rect 25047 52504 25111 52508
rect 25047 52484 25111 52488
rect 25047 52428 25051 52484
rect 25051 52428 25107 52484
rect 25107 52428 25111 52484
rect 25047 52424 25111 52428
rect 25047 52404 25111 52408
rect 25047 52348 25051 52404
rect 25051 52348 25107 52404
rect 25107 52348 25111 52404
rect 25047 52344 25111 52348
rect 25047 52324 25111 52328
rect 25047 52268 25051 52324
rect 25051 52268 25107 52324
rect 25107 52268 25111 52324
rect 25047 52264 25111 52268
rect 25047 52244 25111 52248
rect 25047 52188 25051 52244
rect 25051 52188 25107 52244
rect 25107 52188 25111 52244
rect 25047 52184 25111 52188
rect 26135 52724 26199 52728
rect 26135 52668 26139 52724
rect 26139 52668 26195 52724
rect 26195 52668 26199 52724
rect 26135 52664 26199 52668
rect 26135 52644 26199 52648
rect 26135 52588 26139 52644
rect 26139 52588 26195 52644
rect 26195 52588 26199 52644
rect 26135 52584 26199 52588
rect 26135 52564 26199 52568
rect 26135 52508 26139 52564
rect 26139 52508 26195 52564
rect 26195 52508 26199 52564
rect 26135 52504 26199 52508
rect 26135 52484 26199 52488
rect 26135 52428 26139 52484
rect 26139 52428 26195 52484
rect 26195 52428 26199 52484
rect 26135 52424 26199 52428
rect 26135 52404 26199 52408
rect 26135 52348 26139 52404
rect 26139 52348 26195 52404
rect 26195 52348 26199 52404
rect 26135 52344 26199 52348
rect 26135 52324 26199 52328
rect 26135 52268 26139 52324
rect 26139 52268 26195 52324
rect 26195 52268 26199 52324
rect 26135 52264 26199 52268
rect 26135 52244 26199 52248
rect 26135 52188 26139 52244
rect 26139 52188 26195 52244
rect 26195 52188 26199 52244
rect 26135 52184 26199 52188
rect 27223 52724 27287 52728
rect 27223 52668 27227 52724
rect 27227 52668 27283 52724
rect 27283 52668 27287 52724
rect 27223 52664 27287 52668
rect 27223 52644 27287 52648
rect 27223 52588 27227 52644
rect 27227 52588 27283 52644
rect 27283 52588 27287 52644
rect 27223 52584 27287 52588
rect 27223 52564 27287 52568
rect 27223 52508 27227 52564
rect 27227 52508 27283 52564
rect 27283 52508 27287 52564
rect 27223 52504 27287 52508
rect 27223 52484 27287 52488
rect 27223 52428 27227 52484
rect 27227 52428 27283 52484
rect 27283 52428 27287 52484
rect 27223 52424 27287 52428
rect 27223 52404 27287 52408
rect 27223 52348 27227 52404
rect 27227 52348 27283 52404
rect 27283 52348 27287 52404
rect 27223 52344 27287 52348
rect 27223 52324 27287 52328
rect 27223 52268 27227 52324
rect 27227 52268 27283 52324
rect 27283 52268 27287 52324
rect 27223 52264 27287 52268
rect 27223 52244 27287 52248
rect 27223 52188 27227 52244
rect 27227 52188 27283 52244
rect 27283 52188 27287 52244
rect 27223 52184 27287 52188
rect 28311 52724 28375 52728
rect 28311 52668 28315 52724
rect 28315 52668 28371 52724
rect 28371 52668 28375 52724
rect 28311 52664 28375 52668
rect 28311 52644 28375 52648
rect 28311 52588 28315 52644
rect 28315 52588 28371 52644
rect 28371 52588 28375 52644
rect 28311 52584 28375 52588
rect 28311 52564 28375 52568
rect 28311 52508 28315 52564
rect 28315 52508 28371 52564
rect 28371 52508 28375 52564
rect 28311 52504 28375 52508
rect 28311 52484 28375 52488
rect 28311 52428 28315 52484
rect 28315 52428 28371 52484
rect 28371 52428 28375 52484
rect 28311 52424 28375 52428
rect 28311 52404 28375 52408
rect 28311 52348 28315 52404
rect 28315 52348 28371 52404
rect 28371 52348 28375 52404
rect 28311 52344 28375 52348
rect 28311 52324 28375 52328
rect 28311 52268 28315 52324
rect 28315 52268 28371 52324
rect 28371 52268 28375 52324
rect 28311 52264 28375 52268
rect 28311 52244 28375 52248
rect 28311 52188 28315 52244
rect 28315 52188 28371 52244
rect 28371 52188 28375 52244
rect 28311 52184 28375 52188
rect 29399 52724 29463 52728
rect 29399 52668 29403 52724
rect 29403 52668 29459 52724
rect 29459 52668 29463 52724
rect 29399 52664 29463 52668
rect 29399 52644 29463 52648
rect 29399 52588 29403 52644
rect 29403 52588 29459 52644
rect 29459 52588 29463 52644
rect 29399 52584 29463 52588
rect 29399 52564 29463 52568
rect 29399 52508 29403 52564
rect 29403 52508 29459 52564
rect 29459 52508 29463 52564
rect 29399 52504 29463 52508
rect 29399 52484 29463 52488
rect 29399 52428 29403 52484
rect 29403 52428 29459 52484
rect 29459 52428 29463 52484
rect 29399 52424 29463 52428
rect 29399 52404 29463 52408
rect 29399 52348 29403 52404
rect 29403 52348 29459 52404
rect 29459 52348 29463 52404
rect 29399 52344 29463 52348
rect 29399 52324 29463 52328
rect 29399 52268 29403 52324
rect 29403 52268 29459 52324
rect 29459 52268 29463 52324
rect 29399 52264 29463 52268
rect 29399 52244 29463 52248
rect 29399 52188 29403 52244
rect 29403 52188 29459 52244
rect 29459 52188 29463 52244
rect 29399 52184 29463 52188
rect 30487 52724 30551 52728
rect 30487 52668 30491 52724
rect 30491 52668 30547 52724
rect 30547 52668 30551 52724
rect 30487 52664 30551 52668
rect 30487 52644 30551 52648
rect 30487 52588 30491 52644
rect 30491 52588 30547 52644
rect 30547 52588 30551 52644
rect 30487 52584 30551 52588
rect 30487 52564 30551 52568
rect 30487 52508 30491 52564
rect 30491 52508 30547 52564
rect 30547 52508 30551 52564
rect 30487 52504 30551 52508
rect 30487 52484 30551 52488
rect 30487 52428 30491 52484
rect 30491 52428 30547 52484
rect 30547 52428 30551 52484
rect 30487 52424 30551 52428
rect 30487 52404 30551 52408
rect 30487 52348 30491 52404
rect 30491 52348 30547 52404
rect 30547 52348 30551 52404
rect 30487 52344 30551 52348
rect 30487 52324 30551 52328
rect 30487 52268 30491 52324
rect 30491 52268 30547 52324
rect 30547 52268 30551 52324
rect 30487 52264 30551 52268
rect 30487 52244 30551 52248
rect 30487 52188 30491 52244
rect 30491 52188 30547 52244
rect 30547 52188 30551 52244
rect 30487 52184 30551 52188
rect 31575 52724 31639 52728
rect 31575 52668 31579 52724
rect 31579 52668 31635 52724
rect 31635 52668 31639 52724
rect 31575 52664 31639 52668
rect 31575 52644 31639 52648
rect 31575 52588 31579 52644
rect 31579 52588 31635 52644
rect 31635 52588 31639 52644
rect 31575 52584 31639 52588
rect 31575 52564 31639 52568
rect 31575 52508 31579 52564
rect 31579 52508 31635 52564
rect 31635 52508 31639 52564
rect 31575 52504 31639 52508
rect 31575 52484 31639 52488
rect 31575 52428 31579 52484
rect 31579 52428 31635 52484
rect 31635 52428 31639 52484
rect 31575 52424 31639 52428
rect 31575 52404 31639 52408
rect 31575 52348 31579 52404
rect 31579 52348 31635 52404
rect 31635 52348 31639 52404
rect 31575 52344 31639 52348
rect 31575 52324 31639 52328
rect 31575 52268 31579 52324
rect 31579 52268 31635 52324
rect 31635 52268 31639 52324
rect 31575 52264 31639 52268
rect 31575 52244 31639 52248
rect 31575 52188 31579 52244
rect 31579 52188 31635 52244
rect 31635 52188 31639 52244
rect 31575 52184 31639 52188
rect 17976 50721 18040 50725
rect 17976 50665 17980 50721
rect 17980 50665 18036 50721
rect 18036 50665 18040 50721
rect 17976 50661 18040 50665
rect 17976 50641 18040 50645
rect 17976 50585 17980 50641
rect 17980 50585 18036 50641
rect 18036 50585 18040 50641
rect 17976 50581 18040 50585
rect 17976 50561 18040 50565
rect 17976 50505 17980 50561
rect 17980 50505 18036 50561
rect 18036 50505 18040 50561
rect 17976 50501 18040 50505
rect 17976 50481 18040 50485
rect 17976 50425 17980 50481
rect 17980 50425 18036 50481
rect 18036 50425 18040 50481
rect 17976 50421 18040 50425
rect 17976 50401 18040 50405
rect 17976 50345 17980 50401
rect 17980 50345 18036 50401
rect 18036 50345 18040 50401
rect 17976 50341 18040 50345
rect 17976 50321 18040 50325
rect 17976 50265 17980 50321
rect 17980 50265 18036 50321
rect 18036 50265 18040 50321
rect 17976 50261 18040 50265
rect 17976 50241 18040 50245
rect 17976 50185 17980 50241
rect 17980 50185 18036 50241
rect 18036 50185 18040 50241
rect 17976 50181 18040 50185
rect 20152 50721 20216 50725
rect 20152 50665 20156 50721
rect 20156 50665 20212 50721
rect 20212 50665 20216 50721
rect 20152 50661 20216 50665
rect 20152 50641 20216 50645
rect 20152 50585 20156 50641
rect 20156 50585 20212 50641
rect 20212 50585 20216 50641
rect 20152 50581 20216 50585
rect 20152 50561 20216 50565
rect 20152 50505 20156 50561
rect 20156 50505 20212 50561
rect 20212 50505 20216 50561
rect 20152 50501 20216 50505
rect 20152 50481 20216 50485
rect 20152 50425 20156 50481
rect 20156 50425 20212 50481
rect 20212 50425 20216 50481
rect 20152 50421 20216 50425
rect 20152 50401 20216 50405
rect 20152 50345 20156 50401
rect 20156 50345 20212 50401
rect 20212 50345 20216 50401
rect 20152 50341 20216 50345
rect 20152 50321 20216 50325
rect 20152 50265 20156 50321
rect 20156 50265 20212 50321
rect 20212 50265 20216 50321
rect 20152 50261 20216 50265
rect 20152 50241 20216 50245
rect 20152 50185 20156 50241
rect 20156 50185 20212 50241
rect 20212 50185 20216 50241
rect 20152 50181 20216 50185
rect 21240 50721 21304 50725
rect 21240 50665 21244 50721
rect 21244 50665 21300 50721
rect 21300 50665 21304 50721
rect 21240 50661 21304 50665
rect 21240 50641 21304 50645
rect 21240 50585 21244 50641
rect 21244 50585 21300 50641
rect 21300 50585 21304 50641
rect 21240 50581 21304 50585
rect 21240 50561 21304 50565
rect 21240 50505 21244 50561
rect 21244 50505 21300 50561
rect 21300 50505 21304 50561
rect 21240 50501 21304 50505
rect 21240 50481 21304 50485
rect 21240 50425 21244 50481
rect 21244 50425 21300 50481
rect 21300 50425 21304 50481
rect 21240 50421 21304 50425
rect 21240 50401 21304 50405
rect 21240 50345 21244 50401
rect 21244 50345 21300 50401
rect 21300 50345 21304 50401
rect 21240 50341 21304 50345
rect 21240 50321 21304 50325
rect 21240 50265 21244 50321
rect 21244 50265 21300 50321
rect 21300 50265 21304 50321
rect 21240 50261 21304 50265
rect 21240 50241 21304 50245
rect 21240 50185 21244 50241
rect 21244 50185 21300 50241
rect 21300 50185 21304 50241
rect 21240 50181 21304 50185
rect 23416 50721 23480 50725
rect 23416 50665 23420 50721
rect 23420 50665 23476 50721
rect 23476 50665 23480 50721
rect 23416 50661 23480 50665
rect 23416 50641 23480 50645
rect 23416 50585 23420 50641
rect 23420 50585 23476 50641
rect 23476 50585 23480 50641
rect 23416 50581 23480 50585
rect 23416 50561 23480 50565
rect 23416 50505 23420 50561
rect 23420 50505 23476 50561
rect 23476 50505 23480 50561
rect 23416 50501 23480 50505
rect 23416 50481 23480 50485
rect 23416 50425 23420 50481
rect 23420 50425 23476 50481
rect 23476 50425 23480 50481
rect 23416 50421 23480 50425
rect 23416 50401 23480 50405
rect 23416 50345 23420 50401
rect 23420 50345 23476 50401
rect 23476 50345 23480 50401
rect 23416 50341 23480 50345
rect 23416 50321 23480 50325
rect 23416 50265 23420 50321
rect 23420 50265 23476 50321
rect 23476 50265 23480 50321
rect 23416 50261 23480 50265
rect 23416 50241 23480 50245
rect 23416 50185 23420 50241
rect 23420 50185 23476 50241
rect 23476 50185 23480 50241
rect 23416 50181 23480 50185
rect 24504 50721 24568 50725
rect 24504 50665 24508 50721
rect 24508 50665 24564 50721
rect 24564 50665 24568 50721
rect 24504 50661 24568 50665
rect 24504 50641 24568 50645
rect 24504 50585 24508 50641
rect 24508 50585 24564 50641
rect 24564 50585 24568 50641
rect 24504 50581 24568 50585
rect 24504 50561 24568 50565
rect 24504 50505 24508 50561
rect 24508 50505 24564 50561
rect 24564 50505 24568 50561
rect 24504 50501 24568 50505
rect 24504 50481 24568 50485
rect 24504 50425 24508 50481
rect 24508 50425 24564 50481
rect 24564 50425 24568 50481
rect 24504 50421 24568 50425
rect 24504 50401 24568 50405
rect 24504 50345 24508 50401
rect 24508 50345 24564 50401
rect 24564 50345 24568 50401
rect 24504 50341 24568 50345
rect 24504 50321 24568 50325
rect 24504 50265 24508 50321
rect 24508 50265 24564 50321
rect 24564 50265 24568 50321
rect 24504 50261 24568 50265
rect 24504 50241 24568 50245
rect 24504 50185 24508 50241
rect 24508 50185 24564 50241
rect 24564 50185 24568 50241
rect 24504 50181 24568 50185
rect 25592 50721 25656 50725
rect 25592 50665 25596 50721
rect 25596 50665 25652 50721
rect 25652 50665 25656 50721
rect 25592 50661 25656 50665
rect 25592 50641 25656 50645
rect 25592 50585 25596 50641
rect 25596 50585 25652 50641
rect 25652 50585 25656 50641
rect 25592 50581 25656 50585
rect 25592 50561 25656 50565
rect 25592 50505 25596 50561
rect 25596 50505 25652 50561
rect 25652 50505 25656 50561
rect 25592 50501 25656 50505
rect 25592 50481 25656 50485
rect 25592 50425 25596 50481
rect 25596 50425 25652 50481
rect 25652 50425 25656 50481
rect 25592 50421 25656 50425
rect 25592 50401 25656 50405
rect 25592 50345 25596 50401
rect 25596 50345 25652 50401
rect 25652 50345 25656 50401
rect 25592 50341 25656 50345
rect 25592 50321 25656 50325
rect 25592 50265 25596 50321
rect 25596 50265 25652 50321
rect 25652 50265 25656 50321
rect 25592 50261 25656 50265
rect 25592 50241 25656 50245
rect 25592 50185 25596 50241
rect 25596 50185 25652 50241
rect 25652 50185 25656 50241
rect 25592 50181 25656 50185
rect 27768 50721 27832 50725
rect 27768 50665 27772 50721
rect 27772 50665 27828 50721
rect 27828 50665 27832 50721
rect 27768 50661 27832 50665
rect 27768 50641 27832 50645
rect 27768 50585 27772 50641
rect 27772 50585 27828 50641
rect 27828 50585 27832 50641
rect 27768 50581 27832 50585
rect 27768 50561 27832 50565
rect 27768 50505 27772 50561
rect 27772 50505 27828 50561
rect 27828 50505 27832 50561
rect 27768 50501 27832 50505
rect 27768 50481 27832 50485
rect 27768 50425 27772 50481
rect 27772 50425 27828 50481
rect 27828 50425 27832 50481
rect 27768 50421 27832 50425
rect 27768 50401 27832 50405
rect 27768 50345 27772 50401
rect 27772 50345 27828 50401
rect 27828 50345 27832 50401
rect 27768 50341 27832 50345
rect 27768 50321 27832 50325
rect 27768 50265 27772 50321
rect 27772 50265 27828 50321
rect 27828 50265 27832 50321
rect 27768 50261 27832 50265
rect 27768 50241 27832 50245
rect 27768 50185 27772 50241
rect 27772 50185 27828 50241
rect 27828 50185 27832 50241
rect 27768 50181 27832 50185
rect 28856 50721 28920 50725
rect 28856 50665 28860 50721
rect 28860 50665 28916 50721
rect 28916 50665 28920 50721
rect 28856 50661 28920 50665
rect 28856 50641 28920 50645
rect 28856 50585 28860 50641
rect 28860 50585 28916 50641
rect 28916 50585 28920 50641
rect 28856 50581 28920 50585
rect 28856 50561 28920 50565
rect 28856 50505 28860 50561
rect 28860 50505 28916 50561
rect 28916 50505 28920 50561
rect 28856 50501 28920 50505
rect 28856 50481 28920 50485
rect 28856 50425 28860 50481
rect 28860 50425 28916 50481
rect 28916 50425 28920 50481
rect 28856 50421 28920 50425
rect 28856 50401 28920 50405
rect 28856 50345 28860 50401
rect 28860 50345 28916 50401
rect 28916 50345 28920 50401
rect 28856 50341 28920 50345
rect 28856 50321 28920 50325
rect 28856 50265 28860 50321
rect 28860 50265 28916 50321
rect 28916 50265 28920 50321
rect 28856 50261 28920 50265
rect 28856 50241 28920 50245
rect 28856 50185 28860 50241
rect 28860 50185 28916 50241
rect 28916 50185 28920 50241
rect 28856 50181 28920 50185
rect 31032 50721 31096 50725
rect 31032 50665 31036 50721
rect 31036 50665 31092 50721
rect 31092 50665 31096 50721
rect 31032 50661 31096 50665
rect 31032 50641 31096 50645
rect 31032 50585 31036 50641
rect 31036 50585 31092 50641
rect 31092 50585 31096 50641
rect 31032 50581 31096 50585
rect 31032 50561 31096 50565
rect 31032 50505 31036 50561
rect 31036 50505 31092 50561
rect 31092 50505 31096 50561
rect 31032 50501 31096 50505
rect 31032 50481 31096 50485
rect 31032 50425 31036 50481
rect 31036 50425 31092 50481
rect 31092 50425 31096 50481
rect 31032 50421 31096 50425
rect 31032 50401 31096 50405
rect 31032 50345 31036 50401
rect 31036 50345 31092 50401
rect 31092 50345 31096 50401
rect 31032 50341 31096 50345
rect 31032 50321 31096 50325
rect 31032 50265 31036 50321
rect 31036 50265 31092 50321
rect 31092 50265 31096 50321
rect 31032 50261 31096 50265
rect 31032 50241 31096 50245
rect 31032 50185 31036 50241
rect 31036 50185 31092 50241
rect 31092 50185 31096 50241
rect 31032 50181 31096 50185
rect 17431 48724 17495 48728
rect 17431 48668 17435 48724
rect 17435 48668 17491 48724
rect 17491 48668 17495 48724
rect 17431 48664 17495 48668
rect 17431 48644 17495 48648
rect 17431 48588 17435 48644
rect 17435 48588 17491 48644
rect 17491 48588 17495 48644
rect 17431 48584 17495 48588
rect 17431 48564 17495 48568
rect 17431 48508 17435 48564
rect 17435 48508 17491 48564
rect 17491 48508 17495 48564
rect 17431 48504 17495 48508
rect 17431 48484 17495 48488
rect 17431 48428 17435 48484
rect 17435 48428 17491 48484
rect 17491 48428 17495 48484
rect 17431 48424 17495 48428
rect 17431 48404 17495 48408
rect 17431 48348 17435 48404
rect 17435 48348 17491 48404
rect 17491 48348 17495 48404
rect 17431 48344 17495 48348
rect 17431 48324 17495 48328
rect 17431 48268 17435 48324
rect 17435 48268 17491 48324
rect 17491 48268 17495 48324
rect 17431 48264 17495 48268
rect 17431 48244 17495 48248
rect 17431 48188 17435 48244
rect 17435 48188 17491 48244
rect 17491 48188 17495 48244
rect 17431 48184 17495 48188
rect 18519 48724 18583 48728
rect 18519 48668 18523 48724
rect 18523 48668 18579 48724
rect 18579 48668 18583 48724
rect 18519 48664 18583 48668
rect 18519 48644 18583 48648
rect 18519 48588 18523 48644
rect 18523 48588 18579 48644
rect 18579 48588 18583 48644
rect 18519 48584 18583 48588
rect 18519 48564 18583 48568
rect 18519 48508 18523 48564
rect 18523 48508 18579 48564
rect 18579 48508 18583 48564
rect 18519 48504 18583 48508
rect 18519 48484 18583 48488
rect 18519 48428 18523 48484
rect 18523 48428 18579 48484
rect 18579 48428 18583 48484
rect 18519 48424 18583 48428
rect 18519 48404 18583 48408
rect 18519 48348 18523 48404
rect 18523 48348 18579 48404
rect 18579 48348 18583 48404
rect 18519 48344 18583 48348
rect 18519 48324 18583 48328
rect 18519 48268 18523 48324
rect 18523 48268 18579 48324
rect 18579 48268 18583 48324
rect 18519 48264 18583 48268
rect 18519 48244 18583 48248
rect 18519 48188 18523 48244
rect 18523 48188 18579 48244
rect 18579 48188 18583 48244
rect 18519 48184 18583 48188
rect 19607 48724 19671 48728
rect 19607 48668 19611 48724
rect 19611 48668 19667 48724
rect 19667 48668 19671 48724
rect 19607 48664 19671 48668
rect 19607 48644 19671 48648
rect 19607 48588 19611 48644
rect 19611 48588 19667 48644
rect 19667 48588 19671 48644
rect 19607 48584 19671 48588
rect 19607 48564 19671 48568
rect 19607 48508 19611 48564
rect 19611 48508 19667 48564
rect 19667 48508 19671 48564
rect 19607 48504 19671 48508
rect 19607 48484 19671 48488
rect 19607 48428 19611 48484
rect 19611 48428 19667 48484
rect 19667 48428 19671 48484
rect 19607 48424 19671 48428
rect 19607 48404 19671 48408
rect 19607 48348 19611 48404
rect 19611 48348 19667 48404
rect 19667 48348 19671 48404
rect 19607 48344 19671 48348
rect 19607 48324 19671 48328
rect 19607 48268 19611 48324
rect 19611 48268 19667 48324
rect 19667 48268 19671 48324
rect 19607 48264 19671 48268
rect 19607 48244 19671 48248
rect 19607 48188 19611 48244
rect 19611 48188 19667 48244
rect 19667 48188 19671 48244
rect 19607 48184 19671 48188
rect 20695 48724 20759 48728
rect 20695 48668 20699 48724
rect 20699 48668 20755 48724
rect 20755 48668 20759 48724
rect 20695 48664 20759 48668
rect 20695 48644 20759 48648
rect 20695 48588 20699 48644
rect 20699 48588 20755 48644
rect 20755 48588 20759 48644
rect 20695 48584 20759 48588
rect 20695 48564 20759 48568
rect 20695 48508 20699 48564
rect 20699 48508 20755 48564
rect 20755 48508 20759 48564
rect 20695 48504 20759 48508
rect 20695 48484 20759 48488
rect 20695 48428 20699 48484
rect 20699 48428 20755 48484
rect 20755 48428 20759 48484
rect 20695 48424 20759 48428
rect 20695 48404 20759 48408
rect 20695 48348 20699 48404
rect 20699 48348 20755 48404
rect 20755 48348 20759 48404
rect 20695 48344 20759 48348
rect 20695 48324 20759 48328
rect 20695 48268 20699 48324
rect 20699 48268 20755 48324
rect 20755 48268 20759 48324
rect 20695 48264 20759 48268
rect 20695 48244 20759 48248
rect 20695 48188 20699 48244
rect 20699 48188 20755 48244
rect 20755 48188 20759 48244
rect 20695 48184 20759 48188
rect 21783 48724 21847 48728
rect 21783 48668 21787 48724
rect 21787 48668 21843 48724
rect 21843 48668 21847 48724
rect 21783 48664 21847 48668
rect 21783 48644 21847 48648
rect 21783 48588 21787 48644
rect 21787 48588 21843 48644
rect 21843 48588 21847 48644
rect 21783 48584 21847 48588
rect 21783 48564 21847 48568
rect 21783 48508 21787 48564
rect 21787 48508 21843 48564
rect 21843 48508 21847 48564
rect 21783 48504 21847 48508
rect 21783 48484 21847 48488
rect 21783 48428 21787 48484
rect 21787 48428 21843 48484
rect 21843 48428 21847 48484
rect 21783 48424 21847 48428
rect 21783 48404 21847 48408
rect 21783 48348 21787 48404
rect 21787 48348 21843 48404
rect 21843 48348 21847 48404
rect 21783 48344 21847 48348
rect 21783 48324 21847 48328
rect 21783 48268 21787 48324
rect 21787 48268 21843 48324
rect 21843 48268 21847 48324
rect 21783 48264 21847 48268
rect 21783 48244 21847 48248
rect 21783 48188 21787 48244
rect 21787 48188 21843 48244
rect 21843 48188 21847 48244
rect 21783 48184 21847 48188
rect 22871 48724 22935 48728
rect 22871 48668 22875 48724
rect 22875 48668 22931 48724
rect 22931 48668 22935 48724
rect 22871 48664 22935 48668
rect 22871 48644 22935 48648
rect 22871 48588 22875 48644
rect 22875 48588 22931 48644
rect 22931 48588 22935 48644
rect 22871 48584 22935 48588
rect 22871 48564 22935 48568
rect 22871 48508 22875 48564
rect 22875 48508 22931 48564
rect 22931 48508 22935 48564
rect 22871 48504 22935 48508
rect 22871 48484 22935 48488
rect 22871 48428 22875 48484
rect 22875 48428 22931 48484
rect 22931 48428 22935 48484
rect 22871 48424 22935 48428
rect 22871 48404 22935 48408
rect 22871 48348 22875 48404
rect 22875 48348 22931 48404
rect 22931 48348 22935 48404
rect 22871 48344 22935 48348
rect 22871 48324 22935 48328
rect 22871 48268 22875 48324
rect 22875 48268 22931 48324
rect 22931 48268 22935 48324
rect 22871 48264 22935 48268
rect 22871 48244 22935 48248
rect 22871 48188 22875 48244
rect 22875 48188 22931 48244
rect 22931 48188 22935 48244
rect 22871 48184 22935 48188
rect 23959 48724 24023 48728
rect 23959 48668 23963 48724
rect 23963 48668 24019 48724
rect 24019 48668 24023 48724
rect 23959 48664 24023 48668
rect 23959 48644 24023 48648
rect 23959 48588 23963 48644
rect 23963 48588 24019 48644
rect 24019 48588 24023 48644
rect 23959 48584 24023 48588
rect 23959 48564 24023 48568
rect 23959 48508 23963 48564
rect 23963 48508 24019 48564
rect 24019 48508 24023 48564
rect 23959 48504 24023 48508
rect 23959 48484 24023 48488
rect 23959 48428 23963 48484
rect 23963 48428 24019 48484
rect 24019 48428 24023 48484
rect 23959 48424 24023 48428
rect 23959 48404 24023 48408
rect 23959 48348 23963 48404
rect 23963 48348 24019 48404
rect 24019 48348 24023 48404
rect 23959 48344 24023 48348
rect 23959 48324 24023 48328
rect 23959 48268 23963 48324
rect 23963 48268 24019 48324
rect 24019 48268 24023 48324
rect 23959 48264 24023 48268
rect 23959 48244 24023 48248
rect 23959 48188 23963 48244
rect 23963 48188 24019 48244
rect 24019 48188 24023 48244
rect 23959 48184 24023 48188
rect 29399 48724 29463 48728
rect 29399 48668 29403 48724
rect 29403 48668 29459 48724
rect 29459 48668 29463 48724
rect 29399 48664 29463 48668
rect 29399 48644 29463 48648
rect 29399 48588 29403 48644
rect 29403 48588 29459 48644
rect 29459 48588 29463 48644
rect 29399 48584 29463 48588
rect 29399 48564 29463 48568
rect 29399 48508 29403 48564
rect 29403 48508 29459 48564
rect 29459 48508 29463 48564
rect 29399 48504 29463 48508
rect 29399 48484 29463 48488
rect 29399 48428 29403 48484
rect 29403 48428 29459 48484
rect 29459 48428 29463 48484
rect 29399 48424 29463 48428
rect 29399 48404 29463 48408
rect 29399 48348 29403 48404
rect 29403 48348 29459 48404
rect 29459 48348 29463 48404
rect 29399 48344 29463 48348
rect 29399 48324 29463 48328
rect 29399 48268 29403 48324
rect 29403 48268 29459 48324
rect 29459 48268 29463 48324
rect 29399 48264 29463 48268
rect 29399 48244 29463 48248
rect 29399 48188 29403 48244
rect 29403 48188 29459 48244
rect 29459 48188 29463 48244
rect 29399 48184 29463 48188
rect 30487 48724 30551 48728
rect 30487 48668 30491 48724
rect 30491 48668 30547 48724
rect 30547 48668 30551 48724
rect 30487 48664 30551 48668
rect 30487 48644 30551 48648
rect 30487 48588 30491 48644
rect 30491 48588 30547 48644
rect 30547 48588 30551 48644
rect 30487 48584 30551 48588
rect 30487 48564 30551 48568
rect 30487 48508 30491 48564
rect 30491 48508 30547 48564
rect 30547 48508 30551 48564
rect 30487 48504 30551 48508
rect 30487 48484 30551 48488
rect 30487 48428 30491 48484
rect 30491 48428 30547 48484
rect 30547 48428 30551 48484
rect 30487 48424 30551 48428
rect 30487 48404 30551 48408
rect 30487 48348 30491 48404
rect 30491 48348 30547 48404
rect 30547 48348 30551 48404
rect 30487 48344 30551 48348
rect 30487 48324 30551 48328
rect 30487 48268 30491 48324
rect 30491 48268 30547 48324
rect 30547 48268 30551 48324
rect 30487 48264 30551 48268
rect 30487 48244 30551 48248
rect 30487 48188 30491 48244
rect 30491 48188 30547 48244
rect 30547 48188 30551 48244
rect 30487 48184 30551 48188
rect 31575 48724 31639 48728
rect 31575 48668 31579 48724
rect 31579 48668 31635 48724
rect 31635 48668 31639 48724
rect 31575 48664 31639 48668
rect 31575 48644 31639 48648
rect 31575 48588 31579 48644
rect 31579 48588 31635 48644
rect 31635 48588 31639 48644
rect 31575 48584 31639 48588
rect 31575 48564 31639 48568
rect 31575 48508 31579 48564
rect 31579 48508 31635 48564
rect 31635 48508 31639 48564
rect 31575 48504 31639 48508
rect 31575 48484 31639 48488
rect 31575 48428 31579 48484
rect 31579 48428 31635 48484
rect 31635 48428 31639 48484
rect 31575 48424 31639 48428
rect 31575 48404 31639 48408
rect 31575 48348 31579 48404
rect 31579 48348 31635 48404
rect 31635 48348 31639 48404
rect 31575 48344 31639 48348
rect 31575 48324 31639 48328
rect 31575 48268 31579 48324
rect 31579 48268 31635 48324
rect 31635 48268 31639 48324
rect 31575 48264 31639 48268
rect 31575 48244 31639 48248
rect 31575 48188 31579 48244
rect 31579 48188 31635 48244
rect 31635 48188 31639 48244
rect 31575 48184 31639 48188
rect -11361 47192 -11297 47256
rect -6411 47192 -6347 47256
rect -27071 43274 -27007 43278
rect -27071 43218 -27067 43274
rect -27067 43218 -27011 43274
rect -27011 43218 -27007 43274
rect -27071 43214 -27007 43218
rect -27071 43194 -27007 43198
rect -27071 43138 -27067 43194
rect -27067 43138 -27011 43194
rect -27011 43138 -27007 43194
rect -27071 43134 -27007 43138
rect -27071 43114 -27007 43118
rect -27071 43058 -27067 43114
rect -27067 43058 -27011 43114
rect -27011 43058 -27007 43114
rect -27071 43054 -27007 43058
rect -27071 43034 -27007 43038
rect -27071 42978 -27067 43034
rect -27067 42978 -27011 43034
rect -27011 42978 -27007 43034
rect -27071 42974 -27007 42978
rect -27071 42954 -27007 42958
rect -27071 42898 -27067 42954
rect -27067 42898 -27011 42954
rect -27011 42898 -27007 42954
rect -27071 42894 -27007 42898
rect -27071 42874 -27007 42878
rect -27071 42818 -27067 42874
rect -27067 42818 -27011 42874
rect -27011 42818 -27007 42874
rect -27071 42814 -27007 42818
rect -27071 42133 -27007 42137
rect -27071 42077 -27067 42133
rect -27067 42077 -27011 42133
rect -27011 42077 -27007 42133
rect -27071 42073 -27007 42077
rect -27071 42053 -27007 42057
rect -27071 41997 -27067 42053
rect -27067 41997 -27011 42053
rect -27011 41997 -27007 42053
rect -27071 41993 -27007 41997
rect -27071 41973 -27007 41977
rect -27071 41917 -27067 41973
rect -27067 41917 -27011 41973
rect -27011 41917 -27007 41973
rect -27071 41913 -27007 41917
rect -27071 41893 -27007 41897
rect -27071 41837 -27067 41893
rect -27067 41837 -27011 41893
rect -27011 41837 -27007 41893
rect -27071 41833 -27007 41837
rect -27071 41813 -27007 41817
rect -27071 41757 -27067 41813
rect -27067 41757 -27011 41813
rect -27011 41757 -27007 41813
rect -27071 41753 -27007 41757
rect -27071 41733 -27007 41737
rect -27071 41677 -27067 41733
rect -27067 41677 -27011 41733
rect -27011 41677 -27007 41733
rect -27071 41673 -27007 41677
rect -27071 41653 -27007 41657
rect -27071 41597 -27067 41653
rect -27067 41597 -27011 41653
rect -27011 41597 -27007 41653
rect -27071 41593 -27007 41597
rect -27071 41573 -27007 41577
rect -27071 41517 -27067 41573
rect -27067 41517 -27011 41573
rect -27011 41517 -27007 41573
rect -27071 41513 -27007 41517
rect -27071 41493 -27007 41497
rect -27071 41437 -27067 41493
rect -27067 41437 -27011 41493
rect -27011 41437 -27007 41493
rect -27071 41433 -27007 41437
rect -27071 41413 -27007 41417
rect -27071 41357 -27067 41413
rect -27067 41357 -27011 41413
rect -27011 41357 -27007 41413
rect -27071 41353 -27007 41357
rect -27071 41333 -27007 41337
rect -27071 41277 -27067 41333
rect -27067 41277 -27011 41333
rect -27011 41277 -27007 41333
rect -27071 41273 -27007 41277
rect -27071 41253 -27007 41257
rect -27071 41197 -27067 41253
rect -27067 41197 -27011 41253
rect -27011 41197 -27007 41253
rect -27071 41193 -27007 41197
rect -27071 41173 -27007 41177
rect -27071 41117 -27067 41173
rect -27067 41117 -27011 41173
rect -27011 41117 -27007 41173
rect -27071 41113 -27007 41117
rect -27071 41093 -27007 41097
rect -27071 41037 -27067 41093
rect -27067 41037 -27011 41093
rect -27011 41037 -27007 41093
rect -27071 41033 -27007 41037
rect -27066 40607 -27002 40611
rect -27066 40551 -27062 40607
rect -27062 40551 -27006 40607
rect -27006 40551 -27002 40607
rect -27066 40547 -27002 40551
rect -27066 40527 -27002 40531
rect -27066 40471 -27062 40527
rect -27062 40471 -27006 40527
rect -27006 40471 -27002 40527
rect -27066 40467 -27002 40471
rect -27066 40447 -27002 40451
rect -27066 40391 -27062 40447
rect -27062 40391 -27006 40447
rect -27006 40391 -27002 40447
rect -27066 40387 -27002 40391
rect -27066 40367 -27002 40371
rect -27066 40311 -27062 40367
rect -27062 40311 -27006 40367
rect -27006 40311 -27002 40367
rect -27066 40307 -27002 40311
rect -27066 40287 -27002 40291
rect -27066 40231 -27062 40287
rect -27062 40231 -27006 40287
rect -27006 40231 -27002 40287
rect -27066 40227 -27002 40231
rect -27066 40207 -27002 40211
rect -27066 40151 -27062 40207
rect -27062 40151 -27006 40207
rect -27006 40151 -27002 40207
rect -27066 40147 -27002 40151
rect -27066 40127 -27002 40131
rect -27066 40071 -27062 40127
rect -27062 40071 -27006 40127
rect -27006 40071 -27002 40127
rect -27066 40067 -27002 40071
rect -27066 40047 -27002 40051
rect -27066 39991 -27062 40047
rect -27062 39991 -27006 40047
rect -27006 39991 -27002 40047
rect -27066 39987 -27002 39991
rect -27066 39967 -27002 39971
rect -27066 39911 -27062 39967
rect -27062 39911 -27006 39967
rect -27006 39911 -27002 39967
rect -27066 39907 -27002 39911
rect -27066 39887 -27002 39891
rect -27066 39831 -27062 39887
rect -27062 39831 -27006 39887
rect -27006 39831 -27002 39887
rect -27066 39827 -27002 39831
rect -27066 39807 -27002 39811
rect -27066 39751 -27062 39807
rect -27062 39751 -27006 39807
rect -27006 39751 -27002 39807
rect -27066 39747 -27002 39751
rect -27066 39727 -27002 39731
rect -27066 39671 -27062 39727
rect -27062 39671 -27006 39727
rect -27006 39671 -27002 39727
rect -27066 39667 -27002 39671
rect -27066 39647 -27002 39651
rect -27066 39591 -27062 39647
rect -27062 39591 -27006 39647
rect -27006 39591 -27002 39647
rect -27066 39587 -27002 39591
rect -27066 39567 -27002 39571
rect -27066 39511 -27062 39567
rect -27062 39511 -27006 39567
rect -27006 39511 -27002 39567
rect -27066 39507 -27002 39511
rect -31812 39144 -31748 39148
rect -31812 39088 -31808 39144
rect -31808 39088 -31752 39144
rect -31752 39088 -31748 39144
rect -31812 39084 -31748 39088
rect -31812 39064 -31748 39068
rect -31812 39008 -31808 39064
rect -31808 39008 -31752 39064
rect -31752 39008 -31748 39064
rect -31812 39004 -31748 39008
rect -31812 38984 -31748 38988
rect -31812 38928 -31808 38984
rect -31808 38928 -31752 38984
rect -31752 38928 -31748 38984
rect -31812 38924 -31748 38928
rect -31812 38904 -31748 38908
rect -31812 38848 -31808 38904
rect -31808 38848 -31752 38904
rect -31752 38848 -31748 38904
rect -31812 38844 -31748 38848
rect -27072 39104 -27008 39108
rect -27072 39048 -27068 39104
rect -27068 39048 -27012 39104
rect -27012 39048 -27008 39104
rect -27072 39044 -27008 39048
rect -27072 39024 -27008 39028
rect -27072 38968 -27068 39024
rect -27068 38968 -27012 39024
rect -27012 38968 -27008 39024
rect -27072 38964 -27008 38968
rect -27072 38944 -27008 38948
rect -27072 38888 -27068 38944
rect -27068 38888 -27012 38944
rect -27012 38888 -27008 38944
rect -27072 38884 -27008 38888
rect -27072 38864 -27008 38868
rect -27072 38808 -27068 38864
rect -27068 38808 -27012 38864
rect -27012 38808 -27008 38864
rect -27072 38804 -27008 38808
rect -27072 38784 -27008 38788
rect -27072 38728 -27068 38784
rect -27068 38728 -27012 38784
rect -27012 38728 -27008 38784
rect -27072 38724 -27008 38728
rect -27072 38704 -27008 38708
rect -27072 38648 -27068 38704
rect -27068 38648 -27012 38704
rect -27012 38648 -27008 38704
rect -27072 38644 -27008 38648
rect -31811 38605 -31747 38609
rect -31811 38549 -31807 38605
rect -31807 38549 -31751 38605
rect -31751 38549 -31747 38605
rect -31811 38545 -31747 38549
rect -31811 38525 -31747 38529
rect -31811 38469 -31807 38525
rect -31807 38469 -31751 38525
rect -31751 38469 -31747 38525
rect -31811 38465 -31747 38469
rect -31811 38445 -31747 38449
rect -31811 38389 -31807 38445
rect -31807 38389 -31751 38445
rect -31751 38389 -31747 38445
rect -31811 38385 -31747 38389
rect -27072 38624 -27008 38628
rect -27072 38568 -27068 38624
rect -27068 38568 -27012 38624
rect -27012 38568 -27008 38624
rect -27072 38564 -27008 38568
rect -27072 38544 -27008 38548
rect -27072 38488 -27068 38544
rect -27068 38488 -27012 38544
rect -27012 38488 -27008 38544
rect -27072 38484 -27008 38488
rect -31811 38365 -31747 38369
rect -31811 38309 -31807 38365
rect -31807 38309 -31751 38365
rect -31751 38309 -31747 38365
rect -31811 38305 -31747 38309
rect -29614 38409 -29550 38413
rect -29614 38353 -29610 38409
rect -29610 38353 -29554 38409
rect -29554 38353 -29550 38409
rect -29614 38349 -29550 38353
rect -29534 38409 -29470 38413
rect -29534 38353 -29530 38409
rect -29530 38353 -29474 38409
rect -29474 38353 -29470 38409
rect -29534 38349 -29470 38353
rect -29454 38409 -29390 38413
rect -29454 38353 -29450 38409
rect -29450 38353 -29394 38409
rect -29394 38353 -29390 38409
rect -29454 38349 -29390 38353
rect -29374 38409 -29310 38413
rect -29374 38353 -29370 38409
rect -29370 38353 -29314 38409
rect -29314 38353 -29310 38409
rect -29374 38349 -29310 38353
rect -29294 38409 -29230 38413
rect -29294 38353 -29290 38409
rect -29290 38353 -29234 38409
rect -29234 38353 -29230 38409
rect -29294 38349 -29230 38353
rect -29214 38409 -29150 38413
rect -29214 38353 -29210 38409
rect -29210 38353 -29154 38409
rect -29154 38353 -29150 38409
rect -29214 38349 -29150 38353
rect -27072 38464 -27008 38468
rect -27072 38408 -27068 38464
rect -27068 38408 -27012 38464
rect -27012 38408 -27008 38464
rect -27072 38404 -27008 38408
rect -31811 38285 -31747 38289
rect -31811 38229 -31807 38285
rect -31807 38229 -31751 38285
rect -31751 38229 -31747 38285
rect -31811 38225 -31747 38229
rect -27072 38384 -27008 38388
rect -27072 38328 -27068 38384
rect -27068 38328 -27012 38384
rect -27012 38328 -27008 38384
rect -27072 38324 -27008 38328
rect -27072 38304 -27008 38308
rect -27072 38248 -27068 38304
rect -27068 38248 -27012 38304
rect -27012 38248 -27008 38304
rect -27072 38244 -27008 38248
rect -31811 38205 -31747 38209
rect -31811 38149 -31807 38205
rect -31807 38149 -31751 38205
rect -31751 38149 -31747 38205
rect -31811 38145 -31747 38149
rect 17976 46721 18040 46725
rect 17976 46665 17980 46721
rect 17980 46665 18036 46721
rect 18036 46665 18040 46721
rect 17976 46661 18040 46665
rect -10487 46569 -10423 46633
rect -6411 46569 -6347 46633
rect 17976 46641 18040 46645
rect 17976 46585 17980 46641
rect 17980 46585 18036 46641
rect 18036 46585 18040 46641
rect 17976 46581 18040 46585
rect 17976 46561 18040 46565
rect 17976 46505 17980 46561
rect 17980 46505 18036 46561
rect 18036 46505 18040 46561
rect 17976 46501 18040 46505
rect 17976 46481 18040 46485
rect 17976 46425 17980 46481
rect 17980 46425 18036 46481
rect 18036 46425 18040 46481
rect 17976 46421 18040 46425
rect 17976 46401 18040 46405
rect 17976 46345 17980 46401
rect 17980 46345 18036 46401
rect 18036 46345 18040 46401
rect 17976 46341 18040 46345
rect -13469 43057 -13405 43061
rect -13469 43001 -13465 43057
rect -13465 43001 -13409 43057
rect -13409 43001 -13405 43057
rect -13469 42997 -13405 43001
rect -9208 42997 -9144 43061
rect -12693 42394 -12629 42398
rect -12693 42338 -12689 42394
rect -12689 42338 -12633 42394
rect -12633 42338 -12629 42394
rect -12693 42334 -12629 42338
rect -10069 42334 -10005 42398
rect -21475 42159 -21411 42163
rect -21475 42103 -21471 42159
rect -21471 42103 -21415 42159
rect -21415 42103 -21411 42159
rect -21475 42099 -21411 42103
rect -5895 46234 -5751 46238
rect -5895 39858 -5891 46234
rect -5891 39858 -5755 46234
rect -5755 39858 -5751 46234
rect 17976 46321 18040 46325
rect 17976 46265 17980 46321
rect 17980 46265 18036 46321
rect 18036 46265 18040 46321
rect 17976 46261 18040 46265
rect 17976 46241 18040 46245
rect 17976 46185 17980 46241
rect 17980 46185 18036 46241
rect 18036 46185 18040 46241
rect 17976 46181 18040 46185
rect 19064 46721 19128 46725
rect 19064 46665 19068 46721
rect 19068 46665 19124 46721
rect 19124 46665 19128 46721
rect 19064 46661 19128 46665
rect 19064 46641 19128 46645
rect 19064 46585 19068 46641
rect 19068 46585 19124 46641
rect 19124 46585 19128 46641
rect 19064 46581 19128 46585
rect 19064 46561 19128 46565
rect 19064 46505 19068 46561
rect 19068 46505 19124 46561
rect 19124 46505 19128 46561
rect 19064 46501 19128 46505
rect 19064 46481 19128 46485
rect 19064 46425 19068 46481
rect 19068 46425 19124 46481
rect 19124 46425 19128 46481
rect 19064 46421 19128 46425
rect 19064 46401 19128 46405
rect 19064 46345 19068 46401
rect 19068 46345 19124 46401
rect 19124 46345 19128 46401
rect 19064 46341 19128 46345
rect 19064 46321 19128 46325
rect 19064 46265 19068 46321
rect 19068 46265 19124 46321
rect 19124 46265 19128 46321
rect 19064 46261 19128 46265
rect 19064 46241 19128 46245
rect 19064 46185 19068 46241
rect 19068 46185 19124 46241
rect 19124 46185 19128 46241
rect 19064 46181 19128 46185
rect 20152 46721 20216 46725
rect 20152 46665 20156 46721
rect 20156 46665 20212 46721
rect 20212 46665 20216 46721
rect 20152 46661 20216 46665
rect 20152 46641 20216 46645
rect 20152 46585 20156 46641
rect 20156 46585 20212 46641
rect 20212 46585 20216 46641
rect 20152 46581 20216 46585
rect 20152 46561 20216 46565
rect 20152 46505 20156 46561
rect 20156 46505 20212 46561
rect 20212 46505 20216 46561
rect 20152 46501 20216 46505
rect 20152 46481 20216 46485
rect 20152 46425 20156 46481
rect 20156 46425 20212 46481
rect 20212 46425 20216 46481
rect 20152 46421 20216 46425
rect 20152 46401 20216 46405
rect 20152 46345 20156 46401
rect 20156 46345 20212 46401
rect 20212 46345 20216 46401
rect 20152 46341 20216 46345
rect 20152 46321 20216 46325
rect 20152 46265 20156 46321
rect 20156 46265 20212 46321
rect 20212 46265 20216 46321
rect 20152 46261 20216 46265
rect 20152 46241 20216 46245
rect 20152 46185 20156 46241
rect 20156 46185 20212 46241
rect 20212 46185 20216 46241
rect 20152 46181 20216 46185
rect 21240 46721 21304 46725
rect 21240 46665 21244 46721
rect 21244 46665 21300 46721
rect 21300 46665 21304 46721
rect 21240 46661 21304 46665
rect 21240 46641 21304 46645
rect 21240 46585 21244 46641
rect 21244 46585 21300 46641
rect 21300 46585 21304 46641
rect 21240 46581 21304 46585
rect 21240 46561 21304 46565
rect 21240 46505 21244 46561
rect 21244 46505 21300 46561
rect 21300 46505 21304 46561
rect 21240 46501 21304 46505
rect 21240 46481 21304 46485
rect 21240 46425 21244 46481
rect 21244 46425 21300 46481
rect 21300 46425 21304 46481
rect 21240 46421 21304 46425
rect 21240 46401 21304 46405
rect 21240 46345 21244 46401
rect 21244 46345 21300 46401
rect 21300 46345 21304 46401
rect 21240 46341 21304 46345
rect 21240 46321 21304 46325
rect 21240 46265 21244 46321
rect 21244 46265 21300 46321
rect 21300 46265 21304 46321
rect 21240 46261 21304 46265
rect 21240 46241 21304 46245
rect 21240 46185 21244 46241
rect 21244 46185 21300 46241
rect 21300 46185 21304 46241
rect 21240 46181 21304 46185
rect 22328 46721 22392 46725
rect 22328 46665 22332 46721
rect 22332 46665 22388 46721
rect 22388 46665 22392 46721
rect 22328 46661 22392 46665
rect 22328 46641 22392 46645
rect 22328 46585 22332 46641
rect 22332 46585 22388 46641
rect 22388 46585 22392 46641
rect 22328 46581 22392 46585
rect 22328 46561 22392 46565
rect 22328 46505 22332 46561
rect 22332 46505 22388 46561
rect 22388 46505 22392 46561
rect 22328 46501 22392 46505
rect 22328 46481 22392 46485
rect 22328 46425 22332 46481
rect 22332 46425 22388 46481
rect 22388 46425 22392 46481
rect 22328 46421 22392 46425
rect 22328 46401 22392 46405
rect 22328 46345 22332 46401
rect 22332 46345 22388 46401
rect 22388 46345 22392 46401
rect 22328 46341 22392 46345
rect 22328 46321 22392 46325
rect 22328 46265 22332 46321
rect 22332 46265 22388 46321
rect 22388 46265 22392 46321
rect 22328 46261 22392 46265
rect 22328 46241 22392 46245
rect 22328 46185 22332 46241
rect 22332 46185 22388 46241
rect 22388 46185 22392 46241
rect 22328 46181 22392 46185
rect 24504 46721 24568 46725
rect 24504 46665 24508 46721
rect 24508 46665 24564 46721
rect 24564 46665 24568 46721
rect 24504 46661 24568 46665
rect 24504 46641 24568 46645
rect 24504 46585 24508 46641
rect 24508 46585 24564 46641
rect 24564 46585 24568 46641
rect 24504 46581 24568 46585
rect 24504 46561 24568 46565
rect 24504 46505 24508 46561
rect 24508 46505 24564 46561
rect 24564 46505 24568 46561
rect 24504 46501 24568 46505
rect 24504 46481 24568 46485
rect 24504 46425 24508 46481
rect 24508 46425 24564 46481
rect 24564 46425 24568 46481
rect 24504 46421 24568 46425
rect 24504 46401 24568 46405
rect 24504 46345 24508 46401
rect 24508 46345 24564 46401
rect 24564 46345 24568 46401
rect 24504 46341 24568 46345
rect 24504 46321 24568 46325
rect 24504 46265 24508 46321
rect 24508 46265 24564 46321
rect 24564 46265 24568 46321
rect 24504 46261 24568 46265
rect 24504 46241 24568 46245
rect 24504 46185 24508 46241
rect 24508 46185 24564 46241
rect 24564 46185 24568 46241
rect 24504 46181 24568 46185
rect 25592 46721 25656 46725
rect 25592 46665 25596 46721
rect 25596 46665 25652 46721
rect 25652 46665 25656 46721
rect 25592 46661 25656 46665
rect 25592 46641 25656 46645
rect 25592 46585 25596 46641
rect 25596 46585 25652 46641
rect 25652 46585 25656 46641
rect 25592 46581 25656 46585
rect 25592 46561 25656 46565
rect 25592 46505 25596 46561
rect 25596 46505 25652 46561
rect 25652 46505 25656 46561
rect 25592 46501 25656 46505
rect 25592 46481 25656 46485
rect 25592 46425 25596 46481
rect 25596 46425 25652 46481
rect 25652 46425 25656 46481
rect 25592 46421 25656 46425
rect 25592 46401 25656 46405
rect 25592 46345 25596 46401
rect 25596 46345 25652 46401
rect 25652 46345 25656 46401
rect 25592 46341 25656 46345
rect 25592 46321 25656 46325
rect 25592 46265 25596 46321
rect 25596 46265 25652 46321
rect 25652 46265 25656 46321
rect 25592 46261 25656 46265
rect 25592 46241 25656 46245
rect 25592 46185 25596 46241
rect 25596 46185 25652 46241
rect 25652 46185 25656 46241
rect 25592 46181 25656 46185
rect 26680 46721 26744 46725
rect 26680 46665 26684 46721
rect 26684 46665 26740 46721
rect 26740 46665 26744 46721
rect 26680 46661 26744 46665
rect 26680 46641 26744 46645
rect 26680 46585 26684 46641
rect 26684 46585 26740 46641
rect 26740 46585 26744 46641
rect 26680 46581 26744 46585
rect 26680 46561 26744 46565
rect 26680 46505 26684 46561
rect 26684 46505 26740 46561
rect 26740 46505 26744 46561
rect 26680 46501 26744 46505
rect 26680 46481 26744 46485
rect 26680 46425 26684 46481
rect 26684 46425 26740 46481
rect 26740 46425 26744 46481
rect 26680 46421 26744 46425
rect 26680 46401 26744 46405
rect 26680 46345 26684 46401
rect 26684 46345 26740 46401
rect 26740 46345 26744 46401
rect 26680 46341 26744 46345
rect 26680 46321 26744 46325
rect 26680 46265 26684 46321
rect 26684 46265 26740 46321
rect 26740 46265 26744 46321
rect 26680 46261 26744 46265
rect 26680 46241 26744 46245
rect 26680 46185 26684 46241
rect 26684 46185 26740 46241
rect 26740 46185 26744 46241
rect 26680 46181 26744 46185
rect 27768 46721 27832 46725
rect 27768 46665 27772 46721
rect 27772 46665 27828 46721
rect 27828 46665 27832 46721
rect 27768 46661 27832 46665
rect 27768 46641 27832 46645
rect 27768 46585 27772 46641
rect 27772 46585 27828 46641
rect 27828 46585 27832 46641
rect 27768 46581 27832 46585
rect 27768 46561 27832 46565
rect 27768 46505 27772 46561
rect 27772 46505 27828 46561
rect 27828 46505 27832 46561
rect 27768 46501 27832 46505
rect 27768 46481 27832 46485
rect 27768 46425 27772 46481
rect 27772 46425 27828 46481
rect 27828 46425 27832 46481
rect 27768 46421 27832 46425
rect 27768 46401 27832 46405
rect 27768 46345 27772 46401
rect 27772 46345 27828 46401
rect 27828 46345 27832 46401
rect 27768 46341 27832 46345
rect 27768 46321 27832 46325
rect 27768 46265 27772 46321
rect 27772 46265 27828 46321
rect 27828 46265 27832 46321
rect 27768 46261 27832 46265
rect 27768 46241 27832 46245
rect 27768 46185 27772 46241
rect 27772 46185 27828 46241
rect 27828 46185 27832 46241
rect 27768 46181 27832 46185
rect 28856 46721 28920 46725
rect 28856 46665 28860 46721
rect 28860 46665 28916 46721
rect 28916 46665 28920 46721
rect 28856 46661 28920 46665
rect 28856 46641 28920 46645
rect 28856 46585 28860 46641
rect 28860 46585 28916 46641
rect 28916 46585 28920 46641
rect 28856 46581 28920 46585
rect 28856 46561 28920 46565
rect 28856 46505 28860 46561
rect 28860 46505 28916 46561
rect 28916 46505 28920 46561
rect 28856 46501 28920 46505
rect 28856 46481 28920 46485
rect 28856 46425 28860 46481
rect 28860 46425 28916 46481
rect 28916 46425 28920 46481
rect 28856 46421 28920 46425
rect 28856 46401 28920 46405
rect 28856 46345 28860 46401
rect 28860 46345 28916 46401
rect 28916 46345 28920 46401
rect 28856 46341 28920 46345
rect 28856 46321 28920 46325
rect 28856 46265 28860 46321
rect 28860 46265 28916 46321
rect 28916 46265 28920 46321
rect 28856 46261 28920 46265
rect 28856 46241 28920 46245
rect 28856 46185 28860 46241
rect 28860 46185 28916 46241
rect 28916 46185 28920 46241
rect 28856 46181 28920 46185
rect 29944 46721 30008 46725
rect 29944 46665 29948 46721
rect 29948 46665 30004 46721
rect 30004 46665 30008 46721
rect 29944 46661 30008 46665
rect 29944 46641 30008 46645
rect 29944 46585 29948 46641
rect 29948 46585 30004 46641
rect 30004 46585 30008 46641
rect 29944 46581 30008 46585
rect 29944 46561 30008 46565
rect 29944 46505 29948 46561
rect 29948 46505 30004 46561
rect 30004 46505 30008 46561
rect 29944 46501 30008 46505
rect 29944 46481 30008 46485
rect 29944 46425 29948 46481
rect 29948 46425 30004 46481
rect 30004 46425 30008 46481
rect 29944 46421 30008 46425
rect 29944 46401 30008 46405
rect 29944 46345 29948 46401
rect 29948 46345 30004 46401
rect 30004 46345 30008 46401
rect 29944 46341 30008 46345
rect 29944 46321 30008 46325
rect 29944 46265 29948 46321
rect 29948 46265 30004 46321
rect 30004 46265 30008 46321
rect 29944 46261 30008 46265
rect 29944 46241 30008 46245
rect 29944 46185 29948 46241
rect 29948 46185 30004 46241
rect 30004 46185 30008 46241
rect 29944 46181 30008 46185
rect 31032 46721 31096 46725
rect 31032 46665 31036 46721
rect 31036 46665 31092 46721
rect 31092 46665 31096 46721
rect 31032 46661 31096 46665
rect 31032 46641 31096 46645
rect 31032 46585 31036 46641
rect 31036 46585 31092 46641
rect 31092 46585 31096 46641
rect 31032 46581 31096 46585
rect 31032 46561 31096 46565
rect 31032 46505 31036 46561
rect 31036 46505 31092 46561
rect 31092 46505 31096 46561
rect 31032 46501 31096 46505
rect 31032 46481 31096 46485
rect 31032 46425 31036 46481
rect 31036 46425 31092 46481
rect 31092 46425 31096 46481
rect 31032 46421 31096 46425
rect 31032 46401 31096 46405
rect 31032 46345 31036 46401
rect 31036 46345 31092 46401
rect 31092 46345 31096 46401
rect 31032 46341 31096 46345
rect 31032 46321 31096 46325
rect 31032 46265 31036 46321
rect 31036 46265 31092 46321
rect 31092 46265 31096 46321
rect 31032 46261 31096 46265
rect 31032 46241 31096 46245
rect 31032 46185 31036 46241
rect 31036 46185 31092 46241
rect 31092 46185 31096 46241
rect 31032 46181 31096 46185
rect 379 45829 523 45833
rect 379 44333 383 45829
rect 383 44333 519 45829
rect 519 44333 523 45829
rect 379 44329 523 44333
rect -5895 39854 -5751 39858
rect 360 41367 504 41371
rect 360 39871 364 41367
rect 364 39871 500 41367
rect 500 39871 504 41367
rect 360 39867 504 39871
rect 10213 46105 10517 46109
rect 10213 39889 10217 46105
rect 10217 39889 10513 46105
rect 10513 39889 10517 46105
rect 10213 39885 10517 39889
rect 18245 45744 18309 45748
rect 18245 45688 18249 45744
rect 18249 45688 18305 45744
rect 18305 45688 18309 45744
rect 18245 45684 18309 45688
rect 18791 45744 18855 45748
rect 18791 45688 18795 45744
rect 18795 45688 18851 45744
rect 18851 45688 18855 45744
rect 18791 45684 18855 45688
rect 19337 45735 19401 45739
rect 19337 45679 19341 45735
rect 19341 45679 19397 45735
rect 19397 45679 19401 45735
rect 19337 45675 19401 45679
rect 19882 45734 19946 45738
rect 19882 45678 19886 45734
rect 19886 45678 19942 45734
rect 19942 45678 19946 45734
rect 19882 45674 19946 45678
rect 21513 45722 21577 45726
rect 21513 45666 21517 45722
rect 21517 45666 21573 45722
rect 21573 45666 21577 45722
rect 21513 45662 21577 45666
rect 22056 45719 22120 45723
rect 22056 45663 22060 45719
rect 22060 45663 22116 45719
rect 22116 45663 22120 45719
rect 22056 45659 22120 45663
rect 22598 45718 22662 45722
rect 22598 45662 22602 45718
rect 22602 45662 22658 45718
rect 22658 45662 22662 45718
rect 22598 45658 22662 45662
rect 23145 45723 23209 45727
rect 23145 45667 23149 45723
rect 23149 45667 23205 45723
rect 23205 45667 23209 45723
rect 23145 45663 23209 45667
rect 25863 45734 25927 45738
rect 25863 45678 25867 45734
rect 25867 45678 25923 45734
rect 25923 45678 25927 45734
rect 25863 45674 25927 45678
rect 26406 45738 26470 45742
rect 26406 45682 26410 45738
rect 26410 45682 26466 45738
rect 26466 45682 26470 45738
rect 26406 45678 26470 45682
rect 26948 45732 27012 45736
rect 26948 45676 26952 45732
rect 26952 45676 27008 45732
rect 27008 45676 27012 45732
rect 26948 45672 27012 45676
rect 27505 45723 27569 45727
rect 27505 45667 27509 45723
rect 27509 45667 27565 45723
rect 27565 45667 27569 45723
rect 27505 45663 27569 45667
rect 29129 45734 29193 45738
rect 29129 45678 29133 45734
rect 29133 45678 29189 45734
rect 29189 45678 29193 45734
rect 29129 45674 29193 45678
rect 29673 45727 29737 45731
rect 29673 45671 29677 45727
rect 29677 45671 29733 45727
rect 29733 45671 29737 45727
rect 29673 45667 29737 45671
rect 30223 45731 30287 45735
rect 30223 45675 30227 45731
rect 30227 45675 30283 45731
rect 30283 45675 30287 45731
rect 30223 45671 30287 45675
rect 30756 45731 30820 45735
rect 30756 45675 30760 45731
rect 30760 45675 30816 45731
rect 30816 45675 30820 45731
rect 30756 45671 30820 45675
rect 18791 45008 18855 45072
rect 44758 45068 44822 45072
rect 44758 45012 44762 45068
rect 44762 45012 44818 45068
rect 44818 45012 44822 45068
rect 44758 45008 44822 45012
rect 44838 45068 44902 45072
rect 44838 45012 44842 45068
rect 44842 45012 44898 45068
rect 44898 45012 44902 45068
rect 44838 45008 44902 45012
rect 44918 45068 44982 45072
rect 44918 45012 44922 45068
rect 44922 45012 44978 45068
rect 44978 45012 44982 45068
rect 44918 45008 44982 45012
rect 44998 45068 45062 45072
rect 44998 45012 45002 45068
rect 45002 45012 45058 45068
rect 45058 45012 45062 45068
rect 44998 45008 45062 45012
rect 45078 45068 45142 45072
rect 45078 45012 45082 45068
rect 45082 45012 45138 45068
rect 45138 45012 45142 45068
rect 45078 45008 45142 45012
rect 45158 45068 45222 45072
rect 45158 45012 45162 45068
rect 45162 45012 45218 45068
rect 45218 45012 45222 45068
rect 45158 45008 45222 45012
rect 45238 45068 45302 45072
rect 45238 45012 45242 45068
rect 45242 45012 45298 45068
rect 45298 45012 45302 45068
rect 45238 45008 45302 45012
rect 25863 44827 25927 44891
rect 18245 44637 18309 44701
rect 26406 44462 26470 44526
rect 41543 44522 41607 44526
rect 41543 44466 41547 44522
rect 41547 44466 41603 44522
rect 41603 44466 41607 44522
rect 41543 44462 41607 44466
rect 41623 44522 41687 44526
rect 41623 44466 41627 44522
rect 41627 44466 41683 44522
rect 41683 44466 41687 44522
rect 41623 44462 41687 44466
rect 41703 44522 41767 44526
rect 41703 44466 41707 44522
rect 41707 44466 41763 44522
rect 41763 44466 41767 44522
rect 41703 44462 41767 44466
rect 41783 44522 41847 44526
rect 41783 44466 41787 44522
rect 41787 44466 41843 44522
rect 41843 44466 41847 44522
rect 41783 44462 41847 44466
rect 22597 43858 22661 43922
rect 44797 43917 44861 43921
rect 44797 43861 44801 43917
rect 44801 43861 44857 43917
rect 44857 43861 44861 43917
rect 44797 43857 44861 43861
rect 44877 43917 44941 43921
rect 44877 43861 44881 43917
rect 44881 43861 44937 43917
rect 44937 43861 44941 43917
rect 44877 43857 44941 43861
rect 44957 43917 45021 43921
rect 44957 43861 44961 43917
rect 44961 43861 45017 43917
rect 45017 43861 45021 43917
rect 44957 43857 45021 43861
rect 45037 43917 45101 43921
rect 45037 43861 45041 43917
rect 45041 43861 45097 43917
rect 45097 43861 45101 43917
rect 45037 43857 45101 43861
rect 45117 43917 45181 43921
rect 45117 43861 45121 43917
rect 45121 43861 45177 43917
rect 45177 43861 45181 43917
rect 45117 43857 45181 43861
rect 45197 43917 45261 43921
rect 45197 43861 45201 43917
rect 45201 43861 45257 43917
rect 45257 43861 45261 43917
rect 45197 43857 45261 43861
rect 30756 43677 30820 43741
rect 23145 43487 23209 43551
rect 30222 43311 30286 43375
rect 41541 43372 41605 43376
rect 41541 43316 41545 43372
rect 41545 43316 41601 43372
rect 41601 43316 41605 43372
rect 41541 43312 41605 43316
rect 41621 43372 41685 43376
rect 41621 43316 41625 43372
rect 41625 43316 41681 43372
rect 41681 43316 41685 43372
rect 41621 43312 41685 43316
rect 41701 43372 41765 43376
rect 41701 43316 41705 43372
rect 41705 43316 41761 43372
rect 41761 43316 41765 43372
rect 41701 43312 41765 43316
rect 41781 43372 41845 43376
rect 41781 43316 41785 43372
rect 41785 43316 41841 43372
rect 41841 43316 41845 43372
rect 41781 43312 41845 43316
rect 19882 41318 19946 41382
rect 44787 41375 44851 41379
rect 44787 41319 44791 41375
rect 44791 41319 44847 41375
rect 44847 41319 44851 41375
rect 44787 41315 44851 41319
rect 44867 41375 44931 41379
rect 44867 41319 44871 41375
rect 44871 41319 44927 41375
rect 44927 41319 44931 41375
rect 44867 41315 44931 41319
rect 44947 41375 45011 41379
rect 44947 41319 44951 41375
rect 44951 41319 45007 41375
rect 45007 41319 45011 41375
rect 44947 41315 45011 41319
rect 45027 41375 45091 41379
rect 45027 41319 45031 41375
rect 45031 41319 45087 41375
rect 45087 41319 45091 41375
rect 45027 41315 45091 41319
rect 45107 41375 45171 41379
rect 45107 41319 45111 41375
rect 45111 41319 45167 41375
rect 45167 41319 45171 41375
rect 45107 41315 45171 41319
rect 45187 41375 45251 41379
rect 45187 41319 45191 41375
rect 45191 41319 45247 41375
rect 45247 41319 45251 41375
rect 45187 41315 45251 41319
rect 26948 41137 27012 41201
rect 19337 40947 19401 41011
rect 27505 40772 27569 40836
rect 41459 40831 41523 40835
rect 41459 40775 41463 40831
rect 41463 40775 41519 40831
rect 41519 40775 41523 40831
rect 41459 40771 41523 40775
rect 41539 40831 41603 40835
rect 41539 40775 41543 40831
rect 41543 40775 41599 40831
rect 41599 40775 41603 40831
rect 41539 40771 41603 40775
rect 41619 40831 41683 40835
rect 41619 40775 41623 40831
rect 41623 40775 41679 40831
rect 41679 40775 41683 40831
rect 41619 40771 41683 40775
rect 41699 40831 41763 40835
rect 41699 40775 41703 40831
rect 41703 40775 41759 40831
rect 41759 40775 41763 40831
rect 41699 40771 41763 40775
rect 21513 40048 21577 40112
rect 44787 40105 44851 40109
rect 44787 40049 44791 40105
rect 44791 40049 44847 40105
rect 44847 40049 44851 40105
rect 44787 40045 44851 40049
rect 44867 40105 44931 40109
rect 44867 40049 44871 40105
rect 44871 40049 44927 40105
rect 44927 40049 44931 40105
rect 44867 40045 44931 40049
rect 44947 40105 45011 40109
rect 44947 40049 44951 40105
rect 44951 40049 45007 40105
rect 45007 40049 45011 40105
rect 44947 40045 45011 40049
rect 45027 40105 45091 40109
rect 45027 40049 45031 40105
rect 45031 40049 45087 40105
rect 45087 40049 45091 40105
rect 45027 40045 45091 40049
rect 45107 40105 45171 40109
rect 45107 40049 45111 40105
rect 45111 40049 45167 40105
rect 45167 40049 45171 40105
rect 45107 40045 45171 40049
rect 45187 40105 45251 40109
rect 45187 40049 45191 40105
rect 45191 40049 45247 40105
rect 45247 40049 45251 40105
rect 45187 40045 45251 40049
rect 29673 39867 29737 39931
rect -5668 39824 -164 39828
rect -5668 39688 -5664 39824
rect -5664 39688 -168 39824
rect -168 39688 -164 39824
rect -5668 39684 -164 39688
rect 22057 39677 22121 39741
rect 29129 39502 29193 39566
rect 41457 39562 41521 39566
rect 41457 39506 41461 39562
rect 41461 39506 41517 39562
rect 41517 39506 41521 39562
rect 41457 39502 41521 39506
rect 41537 39562 41601 39566
rect 41537 39506 41541 39562
rect 41541 39506 41597 39562
rect 41597 39506 41601 39562
rect 41537 39502 41601 39506
rect 41617 39562 41681 39566
rect 41617 39506 41621 39562
rect 41621 39506 41677 39562
rect 41677 39506 41681 39562
rect 41617 39502 41681 39506
rect 41697 39562 41761 39566
rect 41697 39506 41701 39562
rect 41701 39506 41757 39562
rect 41757 39506 41761 39562
rect 41697 39502 41761 39506
rect -18877 39498 -18813 39502
rect -18877 39442 -18873 39498
rect -18873 39442 -18817 39498
rect -18817 39442 -18813 39498
rect -18877 39438 -18813 39442
rect -18877 39418 -18813 39422
rect -18877 39362 -18873 39418
rect -18873 39362 -18817 39418
rect -18817 39362 -18813 39418
rect -18877 39358 -18813 39362
rect -18877 39338 -18813 39342
rect -18877 39282 -18873 39338
rect -18873 39282 -18817 39338
rect -18817 39282 -18813 39338
rect -18877 39278 -18813 39282
rect -18877 39258 -18813 39262
rect -18877 39202 -18873 39258
rect -18873 39202 -18817 39258
rect -18817 39202 -18813 39258
rect -18877 39198 -18813 39202
rect -18877 39178 -18813 39182
rect -18877 39122 -18873 39178
rect -18873 39122 -18817 39178
rect -18817 39122 -18813 39178
rect -18877 39118 -18813 39122
rect -18877 39098 -18813 39102
rect -18877 39042 -18873 39098
rect -18873 39042 -18817 39098
rect -18817 39042 -18813 39098
rect -18877 39038 -18813 39042
rect -18877 39018 -18813 39022
rect -18877 38962 -18873 39018
rect -18873 38962 -18817 39018
rect -18817 38962 -18813 39018
rect -18877 38958 -18813 38962
rect -18877 38938 -18813 38942
rect -18877 38882 -18873 38938
rect -18873 38882 -18817 38938
rect -18817 38882 -18813 38938
rect -18877 38878 -18813 38882
rect -18877 38858 -18813 38862
rect -18877 38802 -18873 38858
rect -18873 38802 -18817 38858
rect -18817 38802 -18813 38858
rect -18877 38798 -18813 38802
rect 2522 38869 2586 38873
rect 2522 38813 2526 38869
rect 2526 38813 2582 38869
rect 2582 38813 2586 38869
rect 2522 38809 2586 38813
rect -18877 38778 -18813 38782
rect -18877 38722 -18873 38778
rect -18873 38722 -18817 38778
rect -18817 38722 -18813 38778
rect -18877 38718 -18813 38722
rect -11713 38726 -11649 38790
rect -4713 38726 -4649 38790
rect -18877 38698 -18813 38702
rect -18877 38642 -18873 38698
rect -18873 38642 -18817 38698
rect -18817 38642 -18813 38698
rect -18877 38638 -18813 38642
rect -18877 38618 -18813 38622
rect -18877 38562 -18873 38618
rect -18873 38562 -18817 38618
rect -18817 38562 -18813 38618
rect -18877 38558 -18813 38562
rect -18877 38538 -18813 38542
rect -18877 38482 -18873 38538
rect -18873 38482 -18817 38538
rect -18817 38482 -18813 38538
rect -18877 38478 -18813 38482
rect -18877 38458 -18813 38462
rect -18877 38402 -18873 38458
rect -18873 38402 -18817 38458
rect -18817 38402 -18813 38458
rect -18877 38398 -18813 38402
rect -18877 38378 -18813 38382
rect -18877 38322 -18873 38378
rect -18873 38322 -18817 38378
rect -18817 38322 -18813 38378
rect -18877 38318 -18813 38322
rect -18877 38298 -18813 38302
rect -18877 38242 -18873 38298
rect -18873 38242 -18817 38298
rect -18817 38242 -18813 38298
rect -18877 38238 -18813 38242
rect -18877 38218 -18813 38222
rect -18877 38162 -18873 38218
rect -18873 38162 -18817 38218
rect -18817 38162 -18813 38218
rect -18877 38158 -18813 38162
rect -18877 38138 -18813 38142
rect -18877 38082 -18873 38138
rect -18873 38082 -18817 38138
rect -18817 38082 -18813 38138
rect -18877 38078 -18813 38082
rect -18877 38058 -18813 38062
rect -18877 38002 -18873 38058
rect -18873 38002 -18817 38058
rect -18817 38002 -18813 38058
rect -18877 37998 -18813 38002
rect -18877 37978 -18813 37982
rect -18877 37922 -18873 37978
rect -18873 37922 -18817 37978
rect -18817 37922 -18813 37978
rect -18877 37918 -18813 37922
rect -18877 37898 -18813 37902
rect -18877 37842 -18873 37898
rect -18873 37842 -18817 37898
rect -18817 37842 -18813 37898
rect -18877 37838 -18813 37842
rect -18877 37818 -18813 37822
rect -18877 37762 -18873 37818
rect -18873 37762 -18817 37818
rect -18817 37762 -18813 37818
rect -18877 37758 -18813 37762
rect -18877 37738 -18813 37742
rect -18877 37682 -18873 37738
rect -18873 37682 -18817 37738
rect -18817 37682 -18813 37738
rect -18877 37678 -18813 37682
rect -18877 37658 -18813 37662
rect -18877 37602 -18873 37658
rect -18873 37602 -18817 37658
rect -18817 37602 -18813 37658
rect -18877 37598 -18813 37602
rect -10905 38383 -10841 38447
rect -4123 38383 -4059 38447
rect -15206 37817 -14742 38281
rect 2522 38789 2586 38793
rect 2522 38733 2526 38789
rect 2526 38733 2582 38789
rect 2582 38733 2586 38789
rect 2522 38729 2586 38733
rect 2522 38709 2586 38713
rect 2522 38653 2526 38709
rect 2526 38653 2582 38709
rect 2582 38653 2586 38709
rect 2522 38649 2586 38653
rect 2532 38396 2596 38400
rect 2532 38340 2536 38396
rect 2536 38340 2592 38396
rect 2592 38340 2596 38396
rect 2532 38336 2596 38340
rect 13831 38372 13895 38436
rect 18245 38372 18309 38436
rect 25863 38354 25927 38418
rect 32414 38354 32478 38418
rect 2532 38316 2596 38320
rect 2532 38260 2536 38316
rect 2536 38260 2592 38316
rect 2592 38260 2596 38316
rect 2532 38256 2596 38260
rect 2532 38236 2596 38240
rect 2532 38180 2536 38236
rect 2536 38180 2592 38236
rect 2592 38180 2596 38236
rect 2532 38176 2596 38180
rect 2532 38156 2596 38160
rect 2532 38100 2536 38156
rect 2536 38100 2592 38156
rect 2592 38100 2596 38156
rect 2532 38096 2596 38100
rect 2532 38076 2596 38080
rect 2532 38020 2536 38076
rect 2536 38020 2592 38076
rect 2592 38020 2596 38076
rect 2532 38016 2596 38020
rect -7722 37835 -7658 37899
rect -2398 37835 -2334 37899
rect -760 37835 -696 37899
rect 1473 37835 1537 37899
rect -18877 37578 -18813 37582
rect -18877 37522 -18873 37578
rect -18873 37522 -18817 37578
rect -18817 37522 -18813 37578
rect -18877 37518 -18813 37522
rect -18877 37498 -18813 37502
rect -18877 37442 -18873 37498
rect -18873 37442 -18817 37498
rect -18817 37442 -18813 37498
rect -18877 37438 -18813 37442
rect -18877 37418 -18813 37422
rect -18877 37362 -18873 37418
rect -18873 37362 -18817 37418
rect -18817 37362 -18813 37418
rect -18877 37358 -18813 37362
rect -29630 37319 -29566 37323
rect -29630 37263 -29626 37319
rect -29626 37263 -29570 37319
rect -29570 37263 -29566 37319
rect -29630 37259 -29566 37263
rect -29550 37319 -29486 37323
rect -29550 37263 -29546 37319
rect -29546 37263 -29490 37319
rect -29490 37263 -29486 37319
rect -29550 37259 -29486 37263
rect -29470 37319 -29406 37323
rect -29470 37263 -29466 37319
rect -29466 37263 -29410 37319
rect -29410 37263 -29406 37319
rect -29470 37259 -29406 37263
rect -29390 37319 -29326 37323
rect -29390 37263 -29386 37319
rect -29386 37263 -29330 37319
rect -29330 37263 -29326 37319
rect -29390 37259 -29326 37263
rect -29310 37319 -29246 37323
rect -29310 37263 -29306 37319
rect -29306 37263 -29250 37319
rect -29250 37263 -29246 37319
rect -29310 37259 -29246 37263
rect -29230 37319 -29166 37323
rect -29230 37263 -29226 37319
rect -29226 37263 -29170 37319
rect -29170 37263 -29166 37319
rect -29230 37259 -29166 37263
rect -27069 37337 -27005 37341
rect -27069 37281 -27065 37337
rect -27065 37281 -27009 37337
rect -27009 37281 -27005 37337
rect -27069 37277 -27005 37281
rect -27069 37257 -27005 37261
rect -27069 37201 -27065 37257
rect -27065 37201 -27009 37257
rect -27009 37201 -27005 37257
rect -27069 37197 -27005 37201
rect -27069 37177 -27005 37181
rect -27069 37121 -27065 37177
rect -27065 37121 -27009 37177
rect -27009 37121 -27005 37177
rect -27069 37117 -27005 37121
rect -27069 37097 -27005 37101
rect -27069 37041 -27065 37097
rect -27065 37041 -27009 37097
rect -27009 37041 -27005 37097
rect -27069 37037 -27005 37041
rect -27069 37017 -27005 37021
rect -27069 36961 -27065 37017
rect -27065 36961 -27009 37017
rect -27009 36961 -27005 37017
rect -27069 36957 -27005 36961
rect -27069 36937 -27005 36941
rect -27069 36881 -27065 36937
rect -27065 36881 -27009 36937
rect -27009 36881 -27005 36937
rect -27069 36877 -27005 36881
rect -27069 36857 -27005 36861
rect -27069 36801 -27065 36857
rect -27065 36801 -27009 36857
rect -27009 36801 -27005 36857
rect -27069 36797 -27005 36801
rect -27069 36777 -27005 36781
rect -27069 36721 -27065 36777
rect -27065 36721 -27009 36777
rect -27009 36721 -27005 36777
rect -27069 36717 -27005 36721
rect -27069 36697 -27005 36701
rect -27069 36641 -27065 36697
rect -27065 36641 -27009 36697
rect -27009 36641 -27005 36697
rect -27069 36637 -27005 36641
rect -27069 36617 -27005 36621
rect -27069 36561 -27065 36617
rect -27065 36561 -27009 36617
rect -27009 36561 -27005 36617
rect -27069 36557 -27005 36561
rect -27069 36537 -27005 36541
rect -27069 36481 -27065 36537
rect -27065 36481 -27009 36537
rect -27009 36481 -27005 36537
rect -27069 36477 -27005 36481
rect -18877 37338 -18813 37342
rect -18877 37282 -18873 37338
rect -18873 37282 -18817 37338
rect -18817 37282 -18813 37338
rect -18877 37278 -18813 37282
rect -8480 37307 -8416 37371
rect -2815 37307 -2751 37371
rect -760 37306 -696 37370
rect -18877 37258 -18813 37262
rect -18877 37202 -18873 37258
rect -18873 37202 -18817 37258
rect -18817 37202 -18813 37258
rect -18877 37198 -18813 37202
rect -18877 37178 -18813 37182
rect -18877 37122 -18873 37178
rect -18873 37122 -18817 37178
rect -18817 37122 -18813 37178
rect -18877 37118 -18813 37122
rect 14586 37797 14650 37861
rect 18791 37797 18855 37861
rect 26406 37774 26470 37838
rect 31824 37774 31888 37838
rect 1996 37306 2060 37370
rect -18877 37098 -18813 37102
rect -18877 37042 -18873 37098
rect -18873 37042 -18817 37098
rect -18817 37042 -18813 37098
rect -18877 37038 -18813 37042
rect -18877 37018 -18813 37022
rect -18877 36962 -18873 37018
rect -18873 36962 -18817 37018
rect -18817 36962 -18813 37018
rect -18877 36958 -18813 36962
rect -18877 36938 -18813 36942
rect -18877 36882 -18873 36938
rect -18873 36882 -18817 36938
rect -18817 36882 -18813 36938
rect -18877 36878 -18813 36882
rect -18877 36858 -18813 36862
rect -18877 36802 -18873 36858
rect -18873 36802 -18817 36858
rect -18817 36802 -18813 36858
rect -18877 36798 -18813 36802
rect -18877 36778 -18813 36782
rect -18877 36722 -18873 36778
rect -18873 36722 -18817 36778
rect -18817 36722 -18813 36778
rect -18877 36718 -18813 36722
rect -18877 36698 -18813 36702
rect -18877 36642 -18873 36698
rect -18873 36642 -18817 36698
rect -18817 36642 -18813 36698
rect -18877 36638 -18813 36642
rect -18877 36618 -18813 36622
rect -18877 36562 -18873 36618
rect -18873 36562 -18817 36618
rect -18817 36562 -18813 36618
rect -18877 36558 -18813 36562
rect -18877 36538 -18813 36542
rect -18877 36482 -18873 36538
rect -18873 36482 -18817 36538
rect -18817 36482 -18813 36538
rect -18877 36478 -18813 36482
rect -18877 36458 -18813 36462
rect -18877 36402 -18873 36458
rect -18873 36402 -18817 36458
rect -18817 36402 -18813 36458
rect -18877 36398 -18813 36402
rect -18877 36378 -18813 36382
rect -18877 36322 -18873 36378
rect -18873 36322 -18817 36378
rect -18817 36322 -18813 36378
rect -18877 36318 -18813 36322
rect 15230 37246 15294 37310
rect 19337 37246 19401 37310
rect 30756 37165 30820 37229
rect 31231 37165 31295 37229
rect 2168 37131 2232 37135
rect 2168 37075 2172 37131
rect 2172 37075 2228 37131
rect 2228 37075 2232 37131
rect 2168 37071 2232 37075
rect 2168 37051 2232 37055
rect 2168 36995 2172 37051
rect 2172 36995 2228 37051
rect 2228 36995 2232 37051
rect 2168 36991 2232 36995
rect 2168 36971 2232 36975
rect 2168 36915 2172 36971
rect 2172 36915 2228 36971
rect 2228 36915 2232 36971
rect 2168 36911 2232 36915
rect 15990 36664 16054 36728
rect 19882 36664 19946 36728
rect 2169 36647 2233 36651
rect 2169 36591 2173 36647
rect 2173 36591 2229 36647
rect 2229 36591 2233 36647
rect 2169 36587 2233 36591
rect 2169 36567 2233 36571
rect 2169 36511 2173 36567
rect 2173 36511 2229 36567
rect 2229 36511 2233 36567
rect 2169 36507 2233 36511
rect 2169 36487 2233 36491
rect 2169 36431 2173 36487
rect 2173 36431 2229 36487
rect 2229 36431 2233 36487
rect 2169 36427 2233 36431
rect 2169 36407 2233 36411
rect 2169 36351 2173 36407
rect 2173 36351 2229 36407
rect 2229 36351 2233 36407
rect 2169 36347 2233 36351
rect -18877 36298 -18813 36302
rect -18877 36242 -18873 36298
rect -18873 36242 -18817 36298
rect -18817 36242 -18813 36298
rect -18877 36238 -18813 36242
rect 2169 36327 2233 36331
rect 2169 36271 2173 36327
rect 2173 36271 2229 36327
rect 2229 36271 2233 36327
rect 2169 36267 2233 36271
rect -27069 36120 -27005 36124
rect -27069 36064 -27065 36120
rect -27065 36064 -27009 36120
rect -27009 36064 -27005 36120
rect -27069 36060 -27005 36064
rect -18877 36218 -18813 36222
rect -18877 36162 -18873 36218
rect -18873 36162 -18817 36218
rect -18817 36162 -18813 36218
rect -18877 36158 -18813 36162
rect -27069 36040 -27005 36044
rect -27069 35984 -27065 36040
rect -27065 35984 -27009 36040
rect -27009 35984 -27005 36040
rect -27069 35980 -27005 35984
rect -27069 35960 -27005 35964
rect -27069 35904 -27065 35960
rect -27065 35904 -27009 35960
rect -27009 35904 -27005 35960
rect -27069 35900 -27005 35904
rect 30222 36529 30286 36593
rect 30584 36529 30648 36593
rect 3584 36090 3648 36094
rect 3584 36034 3588 36090
rect 3588 36034 3644 36090
rect 3644 36034 3648 36090
rect 3584 36030 3648 36034
rect 3664 36090 3728 36094
rect 3664 36034 3668 36090
rect 3668 36034 3724 36090
rect 3724 36034 3728 36090
rect 3664 36030 3728 36034
rect 3744 36090 3808 36094
rect 3744 36034 3748 36090
rect 3748 36034 3804 36090
rect 3804 36034 3808 36090
rect 3744 36030 3808 36034
rect 5091 36089 5155 36093
rect 5171 36089 5235 36093
rect 5251 36089 5315 36093
rect 5091 36033 5111 36089
rect 5111 36033 5135 36089
rect 5135 36033 5155 36089
rect 5171 36033 5191 36089
rect 5191 36033 5215 36089
rect 5215 36033 5235 36089
rect 5251 36033 5271 36089
rect 5271 36033 5295 36089
rect 5295 36033 5315 36089
rect 5091 36029 5155 36033
rect 5171 36029 5235 36033
rect 5251 36029 5315 36033
rect -27069 35880 -27005 35884
rect -27069 35824 -27065 35880
rect -27065 35824 -27009 35880
rect -27009 35824 -27005 35880
rect -27069 35820 -27005 35824
rect -9208 35877 -9144 35941
rect -27069 35800 -27005 35804
rect -27069 35744 -27065 35800
rect -27065 35744 -27009 35800
rect -27009 35744 -27005 35800
rect -27069 35740 -27005 35744
rect -27069 35720 -27005 35724
rect -27069 35664 -27065 35720
rect -27065 35664 -27009 35720
rect -27009 35664 -27005 35720
rect -27069 35660 -27005 35664
rect 5575 36090 5639 36094
rect 5575 36034 5579 36090
rect 5579 36034 5635 36090
rect 5635 36034 5639 36090
rect 5575 36030 5639 36034
rect 5655 36090 5719 36094
rect 5655 36034 5659 36090
rect 5659 36034 5715 36090
rect 5715 36034 5719 36090
rect 5655 36030 5719 36034
rect 5735 36090 5799 36094
rect 5735 36034 5739 36090
rect 5739 36034 5795 36090
rect 5795 36034 5799 36090
rect 5735 36030 5799 36034
rect -27069 35640 -27005 35644
rect -27069 35584 -27065 35640
rect -27065 35584 -27009 35640
rect -27009 35584 -27005 35640
rect -27069 35580 -27005 35584
rect -27069 35560 -27005 35564
rect -27069 35504 -27065 35560
rect -27065 35504 -27009 35560
rect -27009 35504 -27005 35560
rect -27069 35500 -27005 35504
rect 3148 35580 3212 35644
rect -27069 35480 -27005 35484
rect -27069 35424 -27065 35480
rect -27065 35424 -27009 35480
rect -27009 35424 -27005 35480
rect -27069 35420 -27005 35424
rect -27069 35400 -27005 35404
rect -27069 35344 -27065 35400
rect -27065 35344 -27009 35400
rect -27009 35344 -27005 35400
rect -27069 35340 -27005 35344
rect 6974 36082 7038 36086
rect 7054 36082 7118 36086
rect 6974 36026 6994 36082
rect 6994 36026 7018 36082
rect 7018 36026 7038 36082
rect 7054 36026 7074 36082
rect 7074 36026 7098 36082
rect 7098 36026 7118 36082
rect 6974 36022 7038 36026
rect 7054 36022 7118 36026
rect 9576 36085 9640 36089
rect 9576 36029 9580 36085
rect 9580 36029 9636 36085
rect 9636 36029 9640 36085
rect 9576 36025 9640 36029
rect 9656 36085 9720 36089
rect 9656 36029 9660 36085
rect 9660 36029 9716 36085
rect 9716 36029 9720 36085
rect 9656 36025 9720 36029
rect 9736 36085 9800 36089
rect 9736 36029 9740 36085
rect 9740 36029 9796 36085
rect 9796 36029 9800 36085
rect 9736 36025 9800 36029
rect 16721 35986 16785 36050
rect 23145 35986 23209 36050
rect 29673 35906 29737 35970
rect 29990 35906 30054 35970
rect 7530 35549 7594 35613
rect 9097 35558 9161 35622
rect -27069 35320 -27005 35324
rect -27069 35264 -27065 35320
rect -27065 35264 -27009 35320
rect -27009 35264 -27005 35320
rect -27069 35260 -27005 35264
rect -10069 35287 -10005 35351
rect 17412 35279 17476 35343
rect 22598 35279 22662 35343
rect -27069 35240 -27005 35244
rect -27069 35184 -27065 35240
rect -27065 35184 -27009 35240
rect -27009 35184 -27005 35240
rect -27069 35180 -27005 35184
rect 29129 35194 29193 35258
rect 29407 35194 29471 35258
rect -27069 35160 -27005 35164
rect -27069 35104 -27065 35160
rect -27065 35104 -27009 35160
rect -27009 35104 -27005 35160
rect -27069 35100 -27005 35104
rect -27069 35080 -27005 35084
rect -27069 35024 -27065 35080
rect -27065 35024 -27009 35080
rect -27009 35024 -27005 35080
rect -27069 35020 -27005 35024
rect -27072 34682 -27008 34686
rect -27072 34626 -27068 34682
rect -27068 34626 -27012 34682
rect -27012 34626 -27008 34682
rect -27072 34622 -27008 34626
rect -13395 34612 -13331 34676
rect -27072 34602 -27008 34606
rect -27072 34546 -27068 34602
rect -27068 34546 -27012 34602
rect -27012 34546 -27008 34602
rect -27072 34542 -27008 34546
rect -27072 34522 -27008 34526
rect -27072 34466 -27068 34522
rect -27068 34466 -27012 34522
rect -27012 34466 -27008 34522
rect -27072 34462 -27008 34466
rect 18252 34519 18316 34583
rect 22056 34519 22120 34583
rect 26948 34458 27012 34522
rect 28828 34458 28892 34522
rect -27072 34442 -27008 34446
rect -27072 34386 -27068 34442
rect -27068 34386 -27012 34442
rect -27012 34386 -27008 34442
rect -27072 34382 -27008 34386
rect -27072 34362 -27008 34366
rect -27072 34306 -27068 34362
rect -27068 34306 -27012 34362
rect -27012 34306 -27008 34362
rect -27072 34302 -27008 34306
rect -27072 34282 -27008 34286
rect -27072 34226 -27068 34282
rect -27068 34226 -27012 34282
rect -27012 34226 -27008 34282
rect -27072 34222 -27008 34226
rect -27072 34202 -27008 34206
rect -27072 34146 -27068 34202
rect -27068 34146 -27012 34202
rect -27012 34146 -27008 34202
rect -27072 34142 -27008 34146
rect -4713 34131 -4649 34195
rect -27072 34122 -27008 34126
rect -27072 34066 -27068 34122
rect -27068 34066 -27012 34122
rect -27012 34066 -27008 34122
rect -27072 34062 -27008 34066
rect -27072 34042 -27008 34046
rect -27072 33986 -27068 34042
rect -27068 33986 -27012 34042
rect -27012 33986 -27008 34042
rect -27072 33982 -27008 33986
rect -27072 33962 -27008 33966
rect -27072 33906 -27068 33962
rect -27068 33906 -27012 33962
rect -27012 33906 -27008 33962
rect -27072 33902 -27008 33906
rect -27072 33882 -27008 33886
rect -27072 33826 -27068 33882
rect -27068 33826 -27012 33882
rect -27012 33826 -27008 33882
rect -27072 33822 -27008 33826
rect -27072 33802 -27008 33806
rect -27072 33746 -27068 33802
rect -27068 33746 -27012 33802
rect -27012 33746 -27008 33802
rect -27072 33742 -27008 33746
rect -4123 33786 -4059 33850
rect 27505 33749 27569 33813
rect 28315 33749 28379 33813
rect -27072 33722 -27008 33726
rect -27072 33666 -27068 33722
rect -27068 33666 -27012 33722
rect -27012 33666 -27008 33722
rect -27072 33662 -27008 33666
rect 19255 33682 19319 33746
rect 21513 33682 21577 33746
rect -27072 33642 -27008 33646
rect -27072 33586 -27068 33642
rect -27068 33586 -27012 33642
rect -27012 33586 -27008 33642
rect -27072 33582 -27008 33586
rect -27072 33562 -27008 33566
rect -27072 33506 -27068 33562
rect -27068 33506 -27012 33562
rect -27012 33506 -27008 33562
rect -27072 33502 -27008 33506
rect -21518 33547 -21454 33551
rect -21518 33491 -21514 33547
rect -21514 33491 -21458 33547
rect -21458 33491 -21454 33547
rect -21518 33487 -21454 33491
rect -15139 33115 -15075 33179
rect -27077 32860 -27013 32864
rect -27077 32804 -27073 32860
rect -27073 32804 -27017 32860
rect -27017 32804 -27013 32860
rect -27077 32800 -27013 32804
rect -27077 32780 -27013 32784
rect -27077 32724 -27073 32780
rect -27073 32724 -27017 32780
rect -27017 32724 -27013 32780
rect -27077 32720 -27013 32724
rect -27077 32700 -27013 32704
rect -27077 32644 -27073 32700
rect -27073 32644 -27017 32700
rect -27017 32644 -27013 32700
rect -27077 32640 -27013 32644
rect -27077 32620 -27013 32624
rect -27077 32564 -27073 32620
rect -27073 32564 -27017 32620
rect -27017 32564 -27013 32620
rect -27077 32560 -27013 32564
rect -27077 32540 -27013 32544
rect -27077 32484 -27073 32540
rect -27073 32484 -27017 32540
rect -27017 32484 -27013 32540
rect -27077 32480 -27013 32484
rect -27077 32460 -27013 32464
rect -27077 32404 -27073 32460
rect -27073 32404 -27017 32460
rect -27017 32404 -27013 32460
rect -27077 32400 -27013 32404
rect 7965 31807 8029 31811
rect 7965 31751 7969 31807
rect 7969 31751 8025 31807
rect 8025 31751 8029 31807
rect 7965 31747 8029 31751
rect 11347 31327 11411 31391
rect 13831 31327 13895 31391
rect 4354 30428 4418 30432
rect 4354 30372 4358 30428
rect 4358 30372 4414 30428
rect 4414 30372 4418 30428
rect 4354 30368 4418 30372
rect 8328 30433 8392 30437
rect 8328 30377 8332 30433
rect 8332 30377 8388 30433
rect 8388 30377 8392 30433
rect 8328 30373 8392 30377
rect 11966 30708 12030 30772
rect 14586 30708 14650 30772
rect 3326 30301 3390 30305
rect 3326 30245 3330 30301
rect 3330 30245 3386 30301
rect 3386 30245 3390 30301
rect 3326 30241 3390 30245
rect -3918 29688 -3854 29752
rect -5279 29265 -5215 29329
rect 16721 29748 16785 29752
rect 16721 29692 16725 29748
rect 16725 29692 16781 29748
rect 16781 29692 16785 29748
rect 16721 29688 16785 29692
rect 17412 29325 17476 29329
rect 17412 29269 17416 29325
rect 17416 29269 17472 29325
rect 17472 29269 17476 29325
rect 17412 29265 17476 29269
rect 10633 28740 10697 28804
rect 11966 28740 12030 28804
rect -15695 28059 -15631 28063
rect -15695 28003 -15691 28059
rect -15691 28003 -15635 28059
rect -15635 28003 -15631 28059
rect -15695 27999 -15631 28003
rect -15695 27979 -15631 27983
rect -15695 27923 -15691 27979
rect -15691 27923 -15635 27979
rect -15635 27923 -15631 27979
rect -15695 27919 -15631 27923
rect -15695 27899 -15631 27903
rect -15695 27843 -15691 27899
rect -15691 27843 -15635 27899
rect -15635 27843 -15631 27899
rect -15695 27839 -15631 27843
rect -15695 27819 -15631 27823
rect -15695 27763 -15691 27819
rect -15691 27763 -15635 27819
rect -15635 27763 -15631 27819
rect -15695 27759 -15631 27763
rect -15695 27739 -15631 27743
rect -15695 27683 -15691 27739
rect -15691 27683 -15635 27739
rect -15635 27683 -15631 27739
rect -15695 27679 -15631 27683
rect -12385 28061 -12321 28065
rect -12385 28005 -12381 28061
rect -12381 28005 -12325 28061
rect -12325 28005 -12321 28061
rect -12385 28001 -12321 28005
rect -12385 27981 -12321 27985
rect -12385 27925 -12381 27981
rect -12381 27925 -12325 27981
rect -12325 27925 -12321 27981
rect -12385 27921 -12321 27925
rect -12385 27901 -12321 27905
rect -12385 27845 -12381 27901
rect -12381 27845 -12325 27901
rect -12325 27845 -12321 27901
rect -12385 27841 -12321 27845
rect -12385 27821 -12321 27825
rect -12385 27765 -12381 27821
rect -12381 27765 -12325 27821
rect -12325 27765 -12321 27821
rect -12385 27761 -12321 27765
rect -12385 27741 -12321 27745
rect -12385 27685 -12381 27741
rect -12381 27685 -12325 27741
rect -12325 27685 -12321 27741
rect -12385 27681 -12321 27685
rect -17603 27608 -17539 27612
rect -17603 27552 -17599 27608
rect -17599 27552 -17543 27608
rect -17543 27552 -17539 27608
rect -17603 27548 -17539 27552
rect -5279 27528 -5215 27532
rect -5279 27472 -5275 27528
rect -5275 27472 -5219 27528
rect -5219 27472 -5215 27528
rect -5279 27468 -5215 27472
rect -12378 27420 -12314 27424
rect -12378 27364 -12374 27420
rect -12374 27364 -12318 27420
rect -12318 27364 -12314 27420
rect -12378 27360 -12314 27364
rect -12378 27340 -12314 27344
rect -12378 27284 -12374 27340
rect -12374 27284 -12318 27340
rect -12318 27284 -12314 27340
rect -12378 27280 -12314 27284
rect -12378 27260 -12314 27264
rect -12378 27204 -12374 27260
rect -12374 27204 -12318 27260
rect -12318 27204 -12314 27260
rect -12378 27200 -12314 27204
rect -3918 26851 -3854 26855
rect -3918 26795 -3914 26851
rect -3914 26795 -3858 26851
rect -3858 26795 -3854 26851
rect -3918 26791 -3854 26795
rect -38155 26590 -38091 26594
rect -38155 26534 -38151 26590
rect -38151 26534 -38095 26590
rect -38095 26534 -38091 26590
rect -38155 26530 -38091 26534
rect -38075 26590 -38011 26594
rect -38075 26534 -38071 26590
rect -38071 26534 -38015 26590
rect -38015 26534 -38011 26590
rect -38075 26530 -38011 26534
rect -37995 26590 -37931 26594
rect -37995 26534 -37991 26590
rect -37991 26534 -37935 26590
rect -37935 26534 -37931 26590
rect -37995 26530 -37931 26534
rect -37915 26590 -37851 26594
rect -37915 26534 -37911 26590
rect -37911 26534 -37855 26590
rect -37855 26534 -37851 26590
rect -37915 26530 -37851 26534
rect -37835 26590 -37771 26594
rect -37835 26534 -37831 26590
rect -37831 26534 -37775 26590
rect -37775 26534 -37771 26590
rect -37835 26530 -37771 26534
rect -37755 26590 -37691 26594
rect -37755 26534 -37751 26590
rect -37751 26534 -37695 26590
rect -37695 26534 -37691 26590
rect -37755 26530 -37691 26534
rect -37675 26590 -37611 26594
rect -37675 26534 -37671 26590
rect -37671 26534 -37615 26590
rect -37615 26534 -37611 26590
rect -37675 26530 -37611 26534
rect -37595 26590 -37531 26594
rect -37595 26534 -37591 26590
rect -37591 26534 -37535 26590
rect -37535 26534 -37531 26590
rect -37595 26530 -37531 26534
rect -37515 26590 -37451 26594
rect -37515 26534 -37511 26590
rect -37511 26534 -37455 26590
rect -37455 26534 -37451 26590
rect -37515 26530 -37451 26534
rect -37435 26590 -37371 26594
rect -37435 26534 -37431 26590
rect -37431 26534 -37375 26590
rect -37375 26534 -37371 26590
rect -37435 26530 -37371 26534
rect -37355 26590 -37291 26594
rect -37355 26534 -37351 26590
rect -37351 26534 -37295 26590
rect -37295 26534 -37291 26590
rect -37355 26530 -37291 26534
rect -37275 26590 -37211 26594
rect -37275 26534 -37271 26590
rect -37271 26534 -37215 26590
rect -37215 26534 -37211 26590
rect -37275 26530 -37211 26534
rect -37195 26590 -37131 26594
rect -37195 26534 -37191 26590
rect -37191 26534 -37135 26590
rect -37135 26534 -37131 26590
rect -37195 26530 -37131 26534
rect -37115 26590 -37051 26594
rect -37115 26534 -37111 26590
rect -37111 26534 -37055 26590
rect -37055 26534 -37051 26590
rect -37115 26530 -37051 26534
rect -37035 26590 -36971 26594
rect -37035 26534 -37031 26590
rect -37031 26534 -36975 26590
rect -36975 26534 -36971 26590
rect -37035 26530 -36971 26534
rect -36955 26590 -36891 26594
rect -36955 26534 -36951 26590
rect -36951 26534 -36895 26590
rect -36895 26534 -36891 26590
rect -36955 26530 -36891 26534
rect -36875 26590 -36811 26594
rect -36875 26534 -36871 26590
rect -36871 26534 -36815 26590
rect -36815 26534 -36811 26590
rect -36875 26530 -36811 26534
rect -36795 26590 -36731 26594
rect -36795 26534 -36791 26590
rect -36791 26534 -36735 26590
rect -36735 26534 -36731 26590
rect -36795 26530 -36731 26534
rect -36715 26590 -36651 26594
rect -36715 26534 -36711 26590
rect -36711 26534 -36655 26590
rect -36655 26534 -36651 26590
rect -36715 26530 -36651 26534
rect -36635 26590 -36571 26594
rect -36635 26534 -36631 26590
rect -36631 26534 -36575 26590
rect -36575 26534 -36571 26590
rect -36635 26530 -36571 26534
rect -36555 26590 -36491 26594
rect -36555 26534 -36551 26590
rect -36551 26534 -36495 26590
rect -36495 26534 -36491 26590
rect -36555 26530 -36491 26534
rect -36475 26590 -36411 26594
rect -36475 26534 -36471 26590
rect -36471 26534 -36415 26590
rect -36415 26534 -36411 26590
rect -36475 26530 -36411 26534
rect -36395 26590 -36331 26594
rect -36395 26534 -36391 26590
rect -36391 26534 -36335 26590
rect -36335 26534 -36331 26590
rect -36395 26530 -36331 26534
rect -36315 26590 -36251 26594
rect -36315 26534 -36311 26590
rect -36311 26534 -36255 26590
rect -36255 26534 -36251 26590
rect -36315 26530 -36251 26534
rect -36235 26590 -36171 26594
rect -36235 26534 -36231 26590
rect -36231 26534 -36175 26590
rect -36175 26534 -36171 26590
rect -36235 26530 -36171 26534
rect -36155 26590 -36091 26594
rect -36155 26534 -36151 26590
rect -36151 26534 -36095 26590
rect -36095 26534 -36091 26590
rect -36155 26530 -36091 26534
rect -36075 26590 -36011 26594
rect -36075 26534 -36071 26590
rect -36071 26534 -36015 26590
rect -36015 26534 -36011 26590
rect -36075 26530 -36011 26534
rect -35995 26590 -35931 26594
rect -35995 26534 -35991 26590
rect -35991 26534 -35935 26590
rect -35935 26534 -35931 26590
rect -35995 26530 -35931 26534
rect -35915 26590 -35851 26594
rect -35915 26534 -35911 26590
rect -35911 26534 -35855 26590
rect -35855 26534 -35851 26590
rect -35915 26530 -35851 26534
rect -35835 26590 -35771 26594
rect -35835 26534 -35831 26590
rect -35831 26534 -35775 26590
rect -35775 26534 -35771 26590
rect -35835 26530 -35771 26534
rect -35755 26590 -35691 26594
rect -35755 26534 -35751 26590
rect -35751 26534 -35695 26590
rect -35695 26534 -35691 26590
rect -35755 26530 -35691 26534
rect -35675 26590 -35611 26594
rect -35675 26534 -35671 26590
rect -35671 26534 -35615 26590
rect -35615 26534 -35611 26590
rect -35675 26530 -35611 26534
rect -35595 26590 -35531 26594
rect -35595 26534 -35591 26590
rect -35591 26534 -35535 26590
rect -35535 26534 -35531 26590
rect -35595 26530 -35531 26534
rect -35515 26590 -35451 26594
rect -35515 26534 -35511 26590
rect -35511 26534 -35455 26590
rect -35455 26534 -35451 26590
rect -35515 26530 -35451 26534
rect -35435 26590 -35371 26594
rect -35435 26534 -35431 26590
rect -35431 26534 -35375 26590
rect -35375 26534 -35371 26590
rect -35435 26530 -35371 26534
rect -35355 26590 -35291 26594
rect -35355 26534 -35351 26590
rect -35351 26534 -35295 26590
rect -35295 26534 -35291 26590
rect -35355 26530 -35291 26534
rect -35275 26590 -35211 26594
rect -35275 26534 -35271 26590
rect -35271 26534 -35215 26590
rect -35215 26534 -35211 26590
rect -35275 26530 -35211 26534
rect -35195 26590 -35131 26594
rect -35195 26534 -35191 26590
rect -35191 26534 -35135 26590
rect -35135 26534 -35131 26590
rect -35195 26530 -35131 26534
rect -35115 26590 -35051 26594
rect -35115 26534 -35111 26590
rect -35111 26534 -35055 26590
rect -35055 26534 -35051 26590
rect -35115 26530 -35051 26534
rect -35035 26590 -34971 26594
rect -35035 26534 -35031 26590
rect -35031 26534 -34975 26590
rect -34975 26534 -34971 26590
rect -35035 26530 -34971 26534
rect -34955 26590 -34891 26594
rect -34955 26534 -34951 26590
rect -34951 26534 -34895 26590
rect -34895 26534 -34891 26590
rect -34955 26530 -34891 26534
rect -17603 26379 -17539 26383
rect -17603 26323 -17599 26379
rect -17599 26323 -17543 26379
rect -17543 26323 -17539 26379
rect -17603 26319 -17539 26323
rect -12381 26459 -12317 26463
rect -12381 26403 -12377 26459
rect -12377 26403 -12321 26459
rect -12321 26403 -12317 26459
rect -12381 26399 -12317 26403
rect -12381 26379 -12317 26383
rect -12381 26323 -12377 26379
rect -12377 26323 -12321 26379
rect -12321 26323 -12317 26379
rect -12381 26319 -12317 26323
rect -15713 26270 -15649 26274
rect -15713 26214 -15709 26270
rect -15709 26214 -15653 26270
rect -15653 26214 -15649 26270
rect -15713 26210 -15649 26214
rect -15713 26190 -15649 26194
rect -15713 26134 -15709 26190
rect -15709 26134 -15653 26190
rect -15653 26134 -15649 26190
rect -15713 26130 -15649 26134
rect -15713 26110 -15649 26114
rect -15713 26054 -15709 26110
rect -15709 26054 -15653 26110
rect -15653 26054 -15649 26110
rect -15713 26050 -15649 26054
rect -12381 26299 -12317 26303
rect -12381 26243 -12377 26299
rect -12377 26243 -12321 26299
rect -12321 26243 -12317 26299
rect -12381 26239 -12317 26243
rect 11347 26286 11411 26350
rect 11837 26286 11901 26350
rect -12381 26219 -12317 26223
rect -12381 26163 -12377 26219
rect -12377 26163 -12321 26219
rect -12321 26163 -12317 26219
rect -12381 26159 -12317 26163
rect -12381 26139 -12317 26143
rect -12381 26083 -12377 26139
rect -12377 26083 -12321 26139
rect -12321 26083 -12317 26139
rect -12381 26079 -12317 26083
rect 13850 25945 13914 26009
rect 25879 25945 25943 26009
rect -19084 25575 -18860 25799
rect -25441 25476 -25377 25480
rect -25441 25420 -25437 25476
rect -25437 25420 -25381 25476
rect -25381 25420 -25377 25476
rect -25441 25416 -25377 25420
rect -25441 25396 -25377 25400
rect -25441 25340 -25437 25396
rect -25437 25340 -25381 25396
rect -25381 25340 -25377 25396
rect -25441 25336 -25377 25340
rect -25441 25316 -25377 25320
rect -25441 25260 -25437 25316
rect -25437 25260 -25381 25316
rect -25381 25260 -25377 25316
rect -25441 25256 -25377 25260
rect -25441 25236 -25377 25240
rect -25441 25180 -25437 25236
rect -25437 25180 -25381 25236
rect -25381 25180 -25377 25236
rect -25441 25176 -25377 25180
rect -11324 25600 -11260 25664
rect 13266 25534 13330 25598
rect 26463 25534 26527 25598
rect -25441 24937 -25377 24941
rect -25441 24881 -25437 24937
rect -25437 24881 -25381 24937
rect -25381 24881 -25377 24937
rect -25441 24877 -25377 24881
rect -17603 24966 -17539 24970
rect -17603 24910 -17599 24966
rect -17599 24910 -17543 24966
rect -17543 24910 -17539 24966
rect -17603 24906 -17539 24910
rect -25441 24857 -25377 24861
rect -25441 24801 -25437 24857
rect -25437 24801 -25381 24857
rect -25381 24801 -25377 24857
rect -25441 24797 -25377 24801
rect -11977 24808 -11913 24872
rect 7601 24784 7665 24848
rect 15230 24784 15294 24848
rect -25441 24777 -25377 24781
rect -25441 24721 -25437 24777
rect -25437 24721 -25381 24777
rect -25381 24721 -25377 24777
rect -25441 24717 -25377 24721
rect -12393 24693 -12329 24697
rect -12393 24637 -12389 24693
rect -12389 24637 -12333 24693
rect -12333 24637 -12329 24693
rect -12393 24633 -12329 24637
rect -12393 24613 -12329 24617
rect -12393 24557 -12389 24613
rect -12389 24557 -12333 24613
rect -12333 24557 -12329 24613
rect -12393 24553 -12329 24557
rect -12393 24533 -12329 24537
rect -12393 24477 -12389 24533
rect -12389 24477 -12333 24533
rect -12333 24477 -12329 24533
rect -12393 24473 -12329 24477
rect 5717 24578 5781 24582
rect 5717 24522 5721 24578
rect 5721 24522 5777 24578
rect 5777 24522 5781 24578
rect 5717 24518 5781 24522
rect 7266 24529 7330 24593
rect 5717 24498 5781 24502
rect 5717 24442 5721 24498
rect 5721 24442 5777 24498
rect 5777 24442 5781 24498
rect 5717 24438 5781 24442
rect 8129 24466 8193 24530
rect 15990 24466 16054 24530
rect 5717 24418 5781 24422
rect 5717 24362 5721 24418
rect 5721 24362 5777 24418
rect 5777 24362 5781 24418
rect 5717 24358 5781 24362
rect 5717 24338 5781 24342
rect 5717 24282 5721 24338
rect 5721 24282 5777 24338
rect 5777 24282 5781 24338
rect 5717 24278 5781 24282
rect -12389 24229 -12325 24233
rect -12389 24173 -12385 24229
rect -12385 24173 -12329 24229
rect -12329 24173 -12325 24229
rect -12389 24169 -12325 24173
rect 5717 24258 5781 24262
rect 5717 24202 5721 24258
rect 5721 24202 5777 24258
rect 5777 24202 5781 24258
rect 5717 24198 5781 24202
rect -12389 24149 -12325 24153
rect -12389 24093 -12385 24149
rect -12385 24093 -12329 24149
rect -12329 24093 -12325 24149
rect -12389 24089 -12325 24093
rect 11080 24138 11144 24202
rect -12389 24069 -12325 24073
rect -12389 24013 -12385 24069
rect -12385 24013 -12329 24069
rect -12329 24013 -12325 24069
rect -12389 24009 -12325 24013
rect -11324 23823 -11260 23887
rect 7266 23823 7330 23887
rect 19255 23823 19319 23887
rect -17603 23737 -17539 23741
rect -17603 23681 -17599 23737
rect -17599 23681 -17543 23737
rect -17543 23681 -17539 23737
rect -17603 23677 -17539 23681
rect -38149 23582 -38085 23586
rect -38149 23526 -38145 23582
rect -38145 23526 -38089 23582
rect -38089 23526 -38085 23582
rect -38149 23522 -38085 23526
rect -38069 23582 -38005 23586
rect -38069 23526 -38065 23582
rect -38065 23526 -38009 23582
rect -38009 23526 -38005 23582
rect -38069 23522 -38005 23526
rect -37989 23582 -37925 23586
rect -37989 23526 -37985 23582
rect -37985 23526 -37929 23582
rect -37929 23526 -37925 23582
rect -37989 23522 -37925 23526
rect -37909 23582 -37845 23586
rect -37909 23526 -37905 23582
rect -37905 23526 -37849 23582
rect -37849 23526 -37845 23582
rect -37909 23522 -37845 23526
rect -37829 23582 -37765 23586
rect -37829 23526 -37825 23582
rect -37825 23526 -37769 23582
rect -37769 23526 -37765 23582
rect -37829 23522 -37765 23526
rect -37749 23582 -37685 23586
rect -37749 23526 -37745 23582
rect -37745 23526 -37689 23582
rect -37689 23526 -37685 23582
rect -37749 23522 -37685 23526
rect -37669 23582 -37605 23586
rect -37669 23526 -37665 23582
rect -37665 23526 -37609 23582
rect -37609 23526 -37605 23582
rect -37669 23522 -37605 23526
rect -37589 23582 -37525 23586
rect -37589 23526 -37585 23582
rect -37585 23526 -37529 23582
rect -37529 23526 -37525 23582
rect -37589 23522 -37525 23526
rect -37509 23582 -37445 23586
rect -37509 23526 -37505 23582
rect -37505 23526 -37449 23582
rect -37449 23526 -37445 23582
rect -37509 23522 -37445 23526
rect -37429 23582 -37365 23586
rect -37429 23526 -37425 23582
rect -37425 23526 -37369 23582
rect -37369 23526 -37365 23582
rect -37429 23522 -37365 23526
rect -37349 23582 -37285 23586
rect -37349 23526 -37345 23582
rect -37345 23526 -37289 23582
rect -37289 23526 -37285 23582
rect -37349 23522 -37285 23526
rect -37269 23582 -37205 23586
rect -37269 23526 -37265 23582
rect -37265 23526 -37209 23582
rect -37209 23526 -37205 23582
rect -37269 23522 -37205 23526
rect -37189 23582 -37125 23586
rect -37189 23526 -37185 23582
rect -37185 23526 -37129 23582
rect -37129 23526 -37125 23582
rect -37189 23522 -37125 23526
rect -37109 23582 -37045 23586
rect -37109 23526 -37105 23582
rect -37105 23526 -37049 23582
rect -37049 23526 -37045 23582
rect -37109 23522 -37045 23526
rect -37029 23582 -36965 23586
rect -37029 23526 -37025 23582
rect -37025 23526 -36969 23582
rect -36969 23526 -36965 23582
rect -37029 23522 -36965 23526
rect -36949 23582 -36885 23586
rect -36949 23526 -36945 23582
rect -36945 23526 -36889 23582
rect -36889 23526 -36885 23582
rect -36949 23522 -36885 23526
rect -36869 23582 -36805 23586
rect -36869 23526 -36865 23582
rect -36865 23526 -36809 23582
rect -36809 23526 -36805 23582
rect -36869 23522 -36805 23526
rect -36789 23582 -36725 23586
rect -36789 23526 -36785 23582
rect -36785 23526 -36729 23582
rect -36729 23526 -36725 23582
rect -36789 23522 -36725 23526
rect -36709 23582 -36645 23586
rect -36709 23526 -36705 23582
rect -36705 23526 -36649 23582
rect -36649 23526 -36645 23582
rect -36709 23522 -36645 23526
rect -36629 23582 -36565 23586
rect -36629 23526 -36625 23582
rect -36625 23526 -36569 23582
rect -36569 23526 -36565 23582
rect -36629 23522 -36565 23526
rect -36549 23582 -36485 23586
rect -36549 23526 -36545 23582
rect -36545 23526 -36489 23582
rect -36489 23526 -36485 23582
rect -36549 23522 -36485 23526
rect -36469 23582 -36405 23586
rect -36469 23526 -36465 23582
rect -36465 23526 -36409 23582
rect -36409 23526 -36405 23582
rect -36469 23522 -36405 23526
rect -36389 23582 -36325 23586
rect -36389 23526 -36385 23582
rect -36385 23526 -36329 23582
rect -36329 23526 -36325 23582
rect -36389 23522 -36325 23526
rect -36309 23582 -36245 23586
rect -36309 23526 -36305 23582
rect -36305 23526 -36249 23582
rect -36249 23526 -36245 23582
rect -36309 23522 -36245 23526
rect -36229 23582 -36165 23586
rect -36229 23526 -36225 23582
rect -36225 23526 -36169 23582
rect -36169 23526 -36165 23582
rect -36229 23522 -36165 23526
rect -36149 23582 -36085 23586
rect -36149 23526 -36145 23582
rect -36145 23526 -36089 23582
rect -36089 23526 -36085 23582
rect -36149 23522 -36085 23526
rect -36069 23582 -36005 23586
rect -36069 23526 -36065 23582
rect -36065 23526 -36009 23582
rect -36009 23526 -36005 23582
rect -36069 23522 -36005 23526
rect -35989 23582 -35925 23586
rect -35989 23526 -35985 23582
rect -35985 23526 -35929 23582
rect -35929 23526 -35925 23582
rect -35989 23522 -35925 23526
rect -35909 23582 -35845 23586
rect -35909 23526 -35905 23582
rect -35905 23526 -35849 23582
rect -35849 23526 -35845 23582
rect -35909 23522 -35845 23526
rect -35829 23582 -35765 23586
rect -35829 23526 -35825 23582
rect -35825 23526 -35769 23582
rect -35769 23526 -35765 23582
rect -35829 23522 -35765 23526
rect -35749 23582 -35685 23586
rect -35749 23526 -35745 23582
rect -35745 23526 -35689 23582
rect -35689 23526 -35685 23582
rect -35749 23522 -35685 23526
rect -35669 23582 -35605 23586
rect -35669 23526 -35665 23582
rect -35665 23526 -35609 23582
rect -35609 23526 -35605 23582
rect -35669 23522 -35605 23526
rect -35589 23582 -35525 23586
rect -35589 23526 -35585 23582
rect -35585 23526 -35529 23582
rect -35529 23526 -35525 23582
rect -35589 23522 -35525 23526
rect -35509 23582 -35445 23586
rect -35509 23526 -35505 23582
rect -35505 23526 -35449 23582
rect -35449 23526 -35445 23582
rect -35509 23522 -35445 23526
rect -35429 23582 -35365 23586
rect -35429 23526 -35425 23582
rect -35425 23526 -35369 23582
rect -35369 23526 -35365 23582
rect -35429 23522 -35365 23526
rect -35349 23582 -35285 23586
rect -35349 23526 -35345 23582
rect -35345 23526 -35289 23582
rect -35289 23526 -35285 23582
rect -35349 23522 -35285 23526
rect -35269 23582 -35205 23586
rect -35269 23526 -35265 23582
rect -35265 23526 -35209 23582
rect -35209 23526 -35205 23582
rect -35269 23522 -35205 23526
rect -35189 23582 -35125 23586
rect -35189 23526 -35185 23582
rect -35185 23526 -35129 23582
rect -35129 23526 -35125 23582
rect -35189 23522 -35125 23526
rect -35109 23582 -35045 23586
rect -35109 23526 -35105 23582
rect -35105 23526 -35049 23582
rect -35049 23526 -35045 23582
rect -35109 23522 -35045 23526
rect -35029 23582 -34965 23586
rect -35029 23526 -35025 23582
rect -35025 23526 -34969 23582
rect -34969 23526 -34965 23582
rect -35029 23522 -34965 23526
rect -34949 23582 -34885 23586
rect -34949 23526 -34945 23582
rect -34945 23526 -34889 23582
rect -34889 23526 -34885 23582
rect -34949 23522 -34885 23526
rect -15724 23629 -15660 23633
rect -15724 23573 -15720 23629
rect -15720 23573 -15664 23629
rect -15664 23573 -15660 23629
rect -15724 23569 -15660 23573
rect -15724 23549 -15660 23553
rect -15724 23493 -15720 23549
rect -15720 23493 -15664 23549
rect -15664 23493 -15660 23549
rect -15724 23489 -15660 23493
rect -15724 23469 -15660 23473
rect -15724 23413 -15720 23469
rect -15720 23413 -15664 23469
rect -15664 23413 -15660 23469
rect -15724 23409 -15660 23413
rect -11977 23454 -11913 23518
rect 18252 23454 18316 23518
rect -12386 23255 -12322 23259
rect -12386 23199 -12382 23255
rect -12382 23199 -12326 23255
rect -12326 23199 -12322 23255
rect -12386 23195 -12322 23199
rect 8793 23329 8857 23333
rect 8793 23273 8797 23329
rect 8797 23273 8853 23329
rect 8853 23273 8857 23329
rect 8793 23269 8857 23273
rect 8873 23329 8937 23333
rect 8873 23273 8877 23329
rect 8877 23273 8933 23329
rect 8933 23273 8937 23329
rect 8873 23269 8937 23273
rect 42891 24147 42955 24151
rect 42891 24091 42895 24147
rect 42895 24091 42951 24147
rect 42951 24091 42955 24147
rect 42891 24087 42955 24091
rect 42971 24147 43035 24151
rect 42971 24091 42975 24147
rect 42975 24091 43031 24147
rect 43031 24091 43035 24147
rect 42971 24087 43035 24091
rect 43051 24147 43115 24151
rect 43051 24091 43055 24147
rect 43055 24091 43111 24147
rect 43111 24091 43115 24147
rect 43051 24087 43115 24091
rect 43131 24147 43195 24151
rect 43131 24091 43135 24147
rect 43135 24091 43191 24147
rect 43191 24091 43195 24147
rect 43131 24087 43195 24091
rect 43211 24147 43275 24151
rect 43211 24091 43215 24147
rect 43215 24091 43271 24147
rect 43271 24091 43275 24147
rect 43211 24087 43275 24091
rect 43291 24147 43355 24151
rect 43291 24091 43295 24147
rect 43295 24091 43351 24147
rect 43351 24091 43355 24147
rect 43291 24087 43355 24091
rect 43371 24147 43435 24151
rect 43371 24091 43375 24147
rect 43375 24091 43431 24147
rect 43431 24091 43435 24147
rect 43371 24087 43435 24091
rect 43451 24147 43515 24151
rect 43451 24091 43455 24147
rect 43455 24091 43511 24147
rect 43511 24091 43515 24147
rect 43451 24087 43515 24091
rect 43531 24147 43595 24151
rect 43531 24091 43535 24147
rect 43535 24091 43591 24147
rect 43591 24091 43595 24147
rect 43531 24087 43595 24091
rect 43611 24147 43675 24151
rect 43611 24091 43615 24147
rect 43615 24091 43671 24147
rect 43671 24091 43675 24147
rect 43611 24087 43675 24091
rect 43691 24147 43755 24151
rect 43691 24091 43695 24147
rect 43695 24091 43751 24147
rect 43751 24091 43755 24147
rect 43691 24087 43755 24091
rect 43771 24147 43835 24151
rect 43771 24091 43775 24147
rect 43775 24091 43831 24147
rect 43831 24091 43835 24147
rect 43771 24087 43835 24091
rect 43851 24147 43915 24151
rect 43851 24091 43855 24147
rect 43855 24091 43911 24147
rect 43911 24091 43915 24147
rect 43851 24087 43915 24091
rect 43931 24147 43995 24151
rect 43931 24091 43935 24147
rect 43935 24091 43991 24147
rect 43991 24091 43995 24147
rect 43931 24087 43995 24091
rect 44011 24147 44075 24151
rect 44011 24091 44015 24147
rect 44015 24091 44071 24147
rect 44071 24091 44075 24147
rect 44011 24087 44075 24091
rect 44091 24147 44155 24151
rect 44091 24091 44095 24147
rect 44095 24091 44151 24147
rect 44151 24091 44155 24147
rect 44091 24087 44155 24091
rect 44171 24147 44235 24151
rect 44171 24091 44175 24147
rect 44175 24091 44231 24147
rect 44231 24091 44235 24147
rect 44171 24087 44235 24091
rect 44251 24147 44315 24151
rect 44251 24091 44255 24147
rect 44255 24091 44311 24147
rect 44311 24091 44315 24147
rect 44251 24087 44315 24091
rect 44331 24147 44395 24151
rect 44331 24091 44335 24147
rect 44335 24091 44391 24147
rect 44391 24091 44395 24147
rect 44331 24087 44395 24091
rect 44411 24147 44475 24151
rect 44411 24091 44415 24147
rect 44415 24091 44471 24147
rect 44471 24091 44475 24147
rect 44411 24087 44475 24091
rect 44491 24147 44555 24151
rect 44491 24091 44495 24147
rect 44495 24091 44551 24147
rect 44551 24091 44555 24147
rect 44491 24087 44555 24091
rect 44571 24147 44635 24151
rect 44571 24091 44575 24147
rect 44575 24091 44631 24147
rect 44631 24091 44635 24147
rect 44571 24087 44635 24091
rect 44651 24147 44715 24151
rect 44651 24091 44655 24147
rect 44655 24091 44711 24147
rect 44711 24091 44715 24147
rect 44651 24087 44715 24091
rect 44731 24147 44795 24151
rect 44731 24091 44735 24147
rect 44735 24091 44791 24147
rect 44791 24091 44795 24147
rect 44731 24087 44795 24091
rect 44811 24147 44875 24151
rect 44811 24091 44815 24147
rect 44815 24091 44871 24147
rect 44871 24091 44875 24147
rect 44811 24087 44875 24091
rect 44891 24147 44955 24151
rect 44891 24091 44895 24147
rect 44895 24091 44951 24147
rect 44951 24091 44955 24147
rect 44891 24087 44955 24091
rect 44971 24147 45035 24151
rect 44971 24091 44975 24147
rect 44975 24091 45031 24147
rect 45031 24091 45035 24147
rect 44971 24087 45035 24091
rect 45051 24147 45115 24151
rect 45051 24091 45055 24147
rect 45055 24091 45111 24147
rect 45111 24091 45115 24147
rect 45051 24087 45115 24091
rect 45131 24147 45195 24151
rect 45131 24091 45135 24147
rect 45135 24091 45191 24147
rect 45191 24091 45195 24147
rect 45131 24087 45195 24091
rect 45211 24147 45275 24151
rect 45211 24091 45215 24147
rect 45215 24091 45271 24147
rect 45271 24091 45275 24147
rect 45211 24087 45275 24091
rect 45291 24147 45355 24151
rect 45291 24091 45295 24147
rect 45295 24091 45351 24147
rect 45351 24091 45355 24147
rect 45291 24087 45355 24091
rect 45371 24147 45435 24151
rect 45371 24091 45375 24147
rect 45375 24091 45431 24147
rect 45431 24091 45435 24147
rect 45371 24087 45435 24091
rect 45451 24147 45515 24151
rect 45451 24091 45455 24147
rect 45455 24091 45511 24147
rect 45511 24091 45515 24147
rect 45451 24087 45515 24091
rect 45531 24147 45595 24151
rect 45531 24091 45535 24147
rect 45535 24091 45591 24147
rect 45591 24091 45595 24147
rect 45531 24087 45595 24091
rect 45611 24147 45675 24151
rect 45611 24091 45615 24147
rect 45615 24091 45671 24147
rect 45671 24091 45675 24147
rect 45611 24087 45675 24091
rect 45691 24147 45755 24151
rect 45691 24091 45695 24147
rect 45695 24091 45751 24147
rect 45751 24091 45755 24147
rect 45691 24087 45755 24091
rect 45771 24147 45835 24151
rect 45771 24091 45775 24147
rect 45775 24091 45831 24147
rect 45831 24091 45835 24147
rect 45771 24087 45835 24091
rect 45851 24147 45915 24151
rect 45851 24091 45855 24147
rect 45855 24091 45911 24147
rect 45911 24091 45915 24147
rect 45851 24087 45915 24091
rect 45931 24147 45995 24151
rect 45931 24091 45935 24147
rect 45935 24091 45991 24147
rect 45991 24091 45995 24147
rect 45931 24087 45995 24091
rect 46011 24147 46075 24151
rect 46011 24091 46015 24147
rect 46015 24091 46071 24147
rect 46071 24091 46075 24147
rect 46011 24087 46075 24091
rect 46091 24147 46155 24151
rect 46091 24091 46095 24147
rect 46095 24091 46151 24147
rect 46151 24091 46155 24147
rect 46091 24087 46155 24091
rect 36066 24014 36130 24018
rect 36066 23958 36070 24014
rect 36070 23958 36126 24014
rect 36126 23958 36130 24014
rect 36066 23954 36130 23958
rect 35152 23862 35216 23866
rect 35152 23806 35156 23862
rect 35156 23806 35212 23862
rect 35212 23806 35216 23862
rect 35152 23802 35216 23806
rect 37823 23579 37887 23583
rect 37823 23523 37827 23579
rect 37827 23523 37883 23579
rect 37883 23523 37887 23579
rect 37823 23519 37887 23523
rect 39351 23655 39355 23675
rect 39355 23655 39411 23675
rect 39411 23655 39415 23675
rect 39351 23631 39415 23655
rect 39351 23611 39355 23631
rect 39355 23611 39411 23631
rect 39411 23611 39415 23631
rect 39351 23575 39355 23595
rect 39355 23575 39411 23595
rect 39411 23575 39415 23595
rect 39351 23551 39415 23575
rect 39351 23531 39355 23551
rect 39355 23531 39411 23551
rect 39411 23531 39415 23551
rect -12386 23175 -12322 23179
rect -12386 23119 -12382 23175
rect -12382 23119 -12326 23175
rect -12326 23119 -12322 23175
rect -12386 23115 -12322 23119
rect -12386 23095 -12322 23099
rect -12386 23039 -12382 23095
rect -12382 23039 -12326 23095
rect -12326 23039 -12322 23095
rect -12386 23035 -12322 23039
rect -12386 23015 -12322 23019
rect -12386 22959 -12382 23015
rect -12382 22959 -12326 23015
rect -12326 22959 -12322 23015
rect -12386 22955 -12322 22959
rect -12386 22935 -12322 22939
rect -12386 22879 -12382 22935
rect -12382 22879 -12326 22935
rect -12326 22879 -12322 22935
rect -12386 22875 -12322 22879
rect 4819 22927 5203 23151
rect 12588 23146 12652 23210
rect 27111 23146 27175 23210
rect 37830 23178 37894 23182
rect 37830 23122 37834 23178
rect 37834 23122 37890 23178
rect 37890 23122 37894 23178
rect 37830 23118 37894 23122
rect 5718 22999 5782 23063
rect 37830 23098 37894 23102
rect 37830 23042 37834 23098
rect 37834 23042 37890 23098
rect 37890 23042 37894 23098
rect 37830 23038 37894 23042
rect 37830 23018 37894 23022
rect 37830 22962 37834 23018
rect 37834 22962 37890 23018
rect 37890 22962 37894 23018
rect 37830 22958 37894 22962
rect 39346 23184 39410 23188
rect 39346 23128 39350 23184
rect 39350 23128 39406 23184
rect 39406 23128 39410 23184
rect 39346 23124 39410 23128
rect 39346 23104 39410 23108
rect 39346 23048 39350 23104
rect 39350 23048 39406 23104
rect 39406 23048 39410 23104
rect 39346 23044 39410 23048
rect 39346 23024 39410 23028
rect 39346 22968 39350 23024
rect 39350 22968 39406 23024
rect 39406 22968 39410 23024
rect 39346 22964 39410 22968
rect 11476 22851 11540 22915
rect 11837 22852 11901 22916
rect -16599 22660 -16535 22724
rect 8129 22660 8193 22724
rect -12389 22619 -12325 22623
rect -12389 22563 -12385 22619
rect -12385 22563 -12329 22619
rect -12329 22563 -12325 22619
rect -12389 22559 -12325 22563
rect -12389 22539 -12325 22543
rect -12389 22483 -12385 22539
rect -12385 22483 -12329 22539
rect -12329 22483 -12325 22539
rect -12389 22479 -12325 22483
rect -12389 22459 -12325 22463
rect -12389 22403 -12385 22459
rect -12385 22403 -12329 22459
rect -12329 22403 -12325 22459
rect -12389 22399 -12325 22403
rect 7601 22209 7665 22273
rect 36923 22585 37147 22809
rect 39351 22329 39355 22349
rect 39355 22329 39411 22349
rect 39411 22329 39415 22349
rect 39351 22305 39415 22329
rect 39351 22285 39355 22305
rect 39355 22285 39411 22305
rect 39411 22285 39415 22305
rect 37829 22243 37893 22247
rect 37829 22187 37833 22243
rect 37833 22187 37889 22243
rect 37889 22187 37893 22243
rect 37829 22183 37893 22187
rect 39351 22249 39355 22269
rect 39355 22249 39411 22269
rect 39411 22249 39415 22269
rect 39351 22225 39415 22249
rect 39351 22205 39355 22225
rect 39355 22205 39411 22225
rect 39411 22205 39415 22225
rect 37824 21790 37888 21794
rect 37824 21734 37828 21790
rect 37828 21734 37884 21790
rect 37884 21734 37888 21790
rect 37824 21730 37888 21734
rect 12072 21591 12136 21655
rect 27657 21591 27721 21655
rect 37824 21710 37888 21714
rect 37824 21654 37828 21710
rect 37828 21654 37884 21710
rect 37884 21654 37888 21710
rect 37824 21650 37888 21654
rect 39352 21818 39416 21822
rect 39352 21762 39356 21818
rect 39356 21762 39412 21818
rect 39412 21762 39416 21818
rect 39352 21758 39416 21762
rect 39352 21738 39416 21742
rect 39352 21682 39356 21738
rect 39356 21682 39412 21738
rect 39412 21682 39416 21738
rect 39352 21678 39416 21682
rect 35152 21581 35216 21585
rect 35152 21525 35156 21581
rect 35156 21525 35212 21581
rect 35212 21525 35216 21581
rect 35152 21521 35216 21525
rect 39352 21658 39416 21662
rect 39352 21602 39356 21658
rect 39356 21602 39412 21658
rect 39412 21602 39416 21658
rect 39352 21598 39416 21602
rect 35477 21375 35541 21379
rect 35477 21319 35481 21375
rect 35481 21319 35537 21375
rect 35537 21319 35541 21375
rect 35477 21315 35541 21319
rect 42889 21151 42953 21155
rect 42889 21095 42893 21151
rect 42893 21095 42949 21151
rect 42949 21095 42953 21151
rect 42889 21091 42953 21095
rect 42969 21151 43033 21155
rect 42969 21095 42973 21151
rect 42973 21095 43029 21151
rect 43029 21095 43033 21151
rect 42969 21091 43033 21095
rect 43049 21151 43113 21155
rect 43049 21095 43053 21151
rect 43053 21095 43109 21151
rect 43109 21095 43113 21151
rect 43049 21091 43113 21095
rect 43129 21151 43193 21155
rect 43129 21095 43133 21151
rect 43133 21095 43189 21151
rect 43189 21095 43193 21151
rect 43129 21091 43193 21095
rect 43209 21151 43273 21155
rect 43209 21095 43213 21151
rect 43213 21095 43269 21151
rect 43269 21095 43273 21151
rect 43209 21091 43273 21095
rect 43289 21151 43353 21155
rect 43289 21095 43293 21151
rect 43293 21095 43349 21151
rect 43349 21095 43353 21151
rect 43289 21091 43353 21095
rect 43369 21151 43433 21155
rect 43369 21095 43373 21151
rect 43373 21095 43429 21151
rect 43429 21095 43433 21151
rect 43369 21091 43433 21095
rect 43449 21151 43513 21155
rect 43449 21095 43453 21151
rect 43453 21095 43509 21151
rect 43509 21095 43513 21151
rect 43449 21091 43513 21095
rect 43529 21151 43593 21155
rect 43529 21095 43533 21151
rect 43533 21095 43589 21151
rect 43589 21095 43593 21151
rect 43529 21091 43593 21095
rect 43609 21151 43673 21155
rect 43609 21095 43613 21151
rect 43613 21095 43669 21151
rect 43669 21095 43673 21151
rect 43609 21091 43673 21095
rect 43689 21151 43753 21155
rect 43689 21095 43693 21151
rect 43693 21095 43749 21151
rect 43749 21095 43753 21151
rect 43689 21091 43753 21095
rect 43769 21151 43833 21155
rect 43769 21095 43773 21151
rect 43773 21095 43829 21151
rect 43829 21095 43833 21151
rect 43769 21091 43833 21095
rect 43849 21151 43913 21155
rect 43849 21095 43853 21151
rect 43853 21095 43909 21151
rect 43909 21095 43913 21151
rect 43849 21091 43913 21095
rect 43929 21151 43993 21155
rect 43929 21095 43933 21151
rect 43933 21095 43989 21151
rect 43989 21095 43993 21151
rect 43929 21091 43993 21095
rect 44009 21151 44073 21155
rect 44009 21095 44013 21151
rect 44013 21095 44069 21151
rect 44069 21095 44073 21151
rect 44009 21091 44073 21095
rect 44089 21151 44153 21155
rect 44089 21095 44093 21151
rect 44093 21095 44149 21151
rect 44149 21095 44153 21151
rect 44089 21091 44153 21095
rect 44169 21151 44233 21155
rect 44169 21095 44173 21151
rect 44173 21095 44229 21151
rect 44229 21095 44233 21151
rect 44169 21091 44233 21095
rect 44249 21151 44313 21155
rect 44249 21095 44253 21151
rect 44253 21095 44309 21151
rect 44309 21095 44313 21151
rect 44249 21091 44313 21095
rect 44329 21151 44393 21155
rect 44329 21095 44333 21151
rect 44333 21095 44389 21151
rect 44389 21095 44393 21151
rect 44329 21091 44393 21095
rect 44409 21151 44473 21155
rect 44409 21095 44413 21151
rect 44413 21095 44469 21151
rect 44469 21095 44473 21151
rect 44409 21091 44473 21095
rect 44489 21151 44553 21155
rect 44489 21095 44493 21151
rect 44493 21095 44549 21151
rect 44549 21095 44553 21151
rect 44489 21091 44553 21095
rect 44569 21151 44633 21155
rect 44569 21095 44573 21151
rect 44573 21095 44629 21151
rect 44629 21095 44633 21151
rect 44569 21091 44633 21095
rect 44649 21151 44713 21155
rect 44649 21095 44653 21151
rect 44653 21095 44709 21151
rect 44709 21095 44713 21151
rect 44649 21091 44713 21095
rect 44729 21151 44793 21155
rect 44729 21095 44733 21151
rect 44733 21095 44789 21151
rect 44789 21095 44793 21151
rect 44729 21091 44793 21095
rect 44809 21151 44873 21155
rect 44809 21095 44813 21151
rect 44813 21095 44869 21151
rect 44869 21095 44873 21151
rect 44809 21091 44873 21095
rect 44889 21151 44953 21155
rect 44889 21095 44893 21151
rect 44893 21095 44949 21151
rect 44949 21095 44953 21151
rect 44889 21091 44953 21095
rect 44969 21151 45033 21155
rect 44969 21095 44973 21151
rect 44973 21095 45029 21151
rect 45029 21095 45033 21151
rect 44969 21091 45033 21095
rect 45049 21151 45113 21155
rect 45049 21095 45053 21151
rect 45053 21095 45109 21151
rect 45109 21095 45113 21151
rect 45049 21091 45113 21095
rect 45129 21151 45193 21155
rect 45129 21095 45133 21151
rect 45133 21095 45189 21151
rect 45189 21095 45193 21151
rect 45129 21091 45193 21095
rect 45209 21151 45273 21155
rect 45209 21095 45213 21151
rect 45213 21095 45269 21151
rect 45269 21095 45273 21151
rect 45209 21091 45273 21095
rect 45289 21151 45353 21155
rect 45289 21095 45293 21151
rect 45293 21095 45349 21151
rect 45349 21095 45353 21151
rect 45289 21091 45353 21095
rect 45369 21151 45433 21155
rect 45369 21095 45373 21151
rect 45373 21095 45429 21151
rect 45429 21095 45433 21151
rect 45369 21091 45433 21095
rect 45449 21151 45513 21155
rect 45449 21095 45453 21151
rect 45453 21095 45509 21151
rect 45509 21095 45513 21151
rect 45449 21091 45513 21095
rect 45529 21151 45593 21155
rect 45529 21095 45533 21151
rect 45533 21095 45589 21151
rect 45589 21095 45593 21151
rect 45529 21091 45593 21095
rect 45609 21151 45673 21155
rect 45609 21095 45613 21151
rect 45613 21095 45669 21151
rect 45669 21095 45673 21151
rect 45609 21091 45673 21095
rect 45689 21151 45753 21155
rect 45689 21095 45693 21151
rect 45693 21095 45749 21151
rect 45749 21095 45753 21151
rect 45689 21091 45753 21095
rect 45769 21151 45833 21155
rect 45769 21095 45773 21151
rect 45773 21095 45829 21151
rect 45829 21095 45833 21151
rect 45769 21091 45833 21095
rect 45849 21151 45913 21155
rect 45849 21095 45853 21151
rect 45853 21095 45909 21151
rect 45909 21095 45913 21151
rect 45849 21091 45913 21095
rect 45929 21151 45993 21155
rect 45929 21095 45933 21151
rect 45933 21095 45989 21151
rect 45989 21095 45993 21151
rect 45929 21091 45993 21095
rect 46009 21151 46073 21155
rect 46009 21095 46013 21151
rect 46013 21095 46069 21151
rect 46069 21095 46073 21151
rect 46009 21091 46073 21095
rect 46089 21151 46153 21155
rect 46089 21095 46093 21151
rect 46093 21095 46149 21151
rect 46149 21095 46153 21151
rect 46089 21091 46153 21095
rect -38147 19054 -38083 19058
rect -38147 18998 -38143 19054
rect -38143 18998 -38087 19054
rect -38087 18998 -38083 19054
rect -38147 18994 -38083 18998
rect -38067 19054 -38003 19058
rect -38067 18998 -38063 19054
rect -38063 18998 -38007 19054
rect -38007 18998 -38003 19054
rect -38067 18994 -38003 18998
rect -37987 19054 -37923 19058
rect -37987 18998 -37983 19054
rect -37983 18998 -37927 19054
rect -37927 18998 -37923 19054
rect -37987 18994 -37923 18998
rect -37907 19054 -37843 19058
rect -37907 18998 -37903 19054
rect -37903 18998 -37847 19054
rect -37847 18998 -37843 19054
rect -37907 18994 -37843 18998
rect -37827 19054 -37763 19058
rect -37827 18998 -37823 19054
rect -37823 18998 -37767 19054
rect -37767 18998 -37763 19054
rect -37827 18994 -37763 18998
rect -37747 19054 -37683 19058
rect -37747 18998 -37743 19054
rect -37743 18998 -37687 19054
rect -37687 18998 -37683 19054
rect -37747 18994 -37683 18998
rect -37667 19054 -37603 19058
rect -37667 18998 -37663 19054
rect -37663 18998 -37607 19054
rect -37607 18998 -37603 19054
rect -37667 18994 -37603 18998
rect -37587 19054 -37523 19058
rect -37587 18998 -37583 19054
rect -37583 18998 -37527 19054
rect -37527 18998 -37523 19054
rect -37587 18994 -37523 18998
rect -37507 19054 -37443 19058
rect -37507 18998 -37503 19054
rect -37503 18998 -37447 19054
rect -37447 18998 -37443 19054
rect -37507 18994 -37443 18998
rect -37427 19054 -37363 19058
rect -37427 18998 -37423 19054
rect -37423 18998 -37367 19054
rect -37367 18998 -37363 19054
rect -37427 18994 -37363 18998
rect -37347 19054 -37283 19058
rect -37347 18998 -37343 19054
rect -37343 18998 -37287 19054
rect -37287 18998 -37283 19054
rect -37347 18994 -37283 18998
rect -37267 19054 -37203 19058
rect -37267 18998 -37263 19054
rect -37263 18998 -37207 19054
rect -37207 18998 -37203 19054
rect -37267 18994 -37203 18998
rect -37187 19054 -37123 19058
rect -37187 18998 -37183 19054
rect -37183 18998 -37127 19054
rect -37127 18998 -37123 19054
rect -37187 18994 -37123 18998
rect -37107 19054 -37043 19058
rect -37107 18998 -37103 19054
rect -37103 18998 -37047 19054
rect -37047 18998 -37043 19054
rect -37107 18994 -37043 18998
rect -37027 19054 -36963 19058
rect -37027 18998 -37023 19054
rect -37023 18998 -36967 19054
rect -36967 18998 -36963 19054
rect -37027 18994 -36963 18998
rect -36947 19054 -36883 19058
rect -36947 18998 -36943 19054
rect -36943 18998 -36887 19054
rect -36887 18998 -36883 19054
rect -36947 18994 -36883 18998
rect -36867 19054 -36803 19058
rect -36867 18998 -36863 19054
rect -36863 18998 -36807 19054
rect -36807 18998 -36803 19054
rect -36867 18994 -36803 18998
rect -36787 19054 -36723 19058
rect -36787 18998 -36783 19054
rect -36783 18998 -36727 19054
rect -36727 18998 -36723 19054
rect -36787 18994 -36723 18998
rect -36707 19054 -36643 19058
rect -36707 18998 -36703 19054
rect -36703 18998 -36647 19054
rect -36647 18998 -36643 19054
rect -36707 18994 -36643 18998
rect -36627 19054 -36563 19058
rect -36627 18998 -36623 19054
rect -36623 18998 -36567 19054
rect -36567 18998 -36563 19054
rect -36627 18994 -36563 18998
rect -36547 19054 -36483 19058
rect -36547 18998 -36543 19054
rect -36543 18998 -36487 19054
rect -36487 18998 -36483 19054
rect -36547 18994 -36483 18998
rect -36467 19054 -36403 19058
rect -36467 18998 -36463 19054
rect -36463 18998 -36407 19054
rect -36407 18998 -36403 19054
rect -36467 18994 -36403 18998
rect -36387 19054 -36323 19058
rect -36387 18998 -36383 19054
rect -36383 18998 -36327 19054
rect -36327 18998 -36323 19054
rect -36387 18994 -36323 18998
rect -36307 19054 -36243 19058
rect -36307 18998 -36303 19054
rect -36303 18998 -36247 19054
rect -36247 18998 -36243 19054
rect -36307 18994 -36243 18998
rect -36227 19054 -36163 19058
rect -36227 18998 -36223 19054
rect -36223 18998 -36167 19054
rect -36167 18998 -36163 19054
rect -36227 18994 -36163 18998
rect -36147 19054 -36083 19058
rect -36147 18998 -36143 19054
rect -36143 18998 -36087 19054
rect -36087 18998 -36083 19054
rect -36147 18994 -36083 18998
rect -36067 19054 -36003 19058
rect -36067 18998 -36063 19054
rect -36063 18998 -36007 19054
rect -36007 18998 -36003 19054
rect -36067 18994 -36003 18998
rect -35987 19054 -35923 19058
rect -35987 18998 -35983 19054
rect -35983 18998 -35927 19054
rect -35927 18998 -35923 19054
rect -35987 18994 -35923 18998
rect -35907 19054 -35843 19058
rect -35907 18998 -35903 19054
rect -35903 18998 -35847 19054
rect -35847 18998 -35843 19054
rect -35907 18994 -35843 18998
rect -35827 19054 -35763 19058
rect -35827 18998 -35823 19054
rect -35823 18998 -35767 19054
rect -35767 18998 -35763 19054
rect -35827 18994 -35763 18998
rect -35747 19054 -35683 19058
rect -35747 18998 -35743 19054
rect -35743 18998 -35687 19054
rect -35687 18998 -35683 19054
rect -35747 18994 -35683 18998
rect -35667 19054 -35603 19058
rect -35667 18998 -35663 19054
rect -35663 18998 -35607 19054
rect -35607 18998 -35603 19054
rect -35667 18994 -35603 18998
rect -35587 19054 -35523 19058
rect -35587 18998 -35583 19054
rect -35583 18998 -35527 19054
rect -35527 18998 -35523 19054
rect -35587 18994 -35523 18998
rect -35507 19054 -35443 19058
rect -35507 18998 -35503 19054
rect -35503 18998 -35447 19054
rect -35447 18998 -35443 19054
rect -35507 18994 -35443 18998
rect -35427 19054 -35363 19058
rect -35427 18998 -35423 19054
rect -35423 18998 -35367 19054
rect -35367 18998 -35363 19054
rect -35427 18994 -35363 18998
rect -35347 19054 -35283 19058
rect -35347 18998 -35343 19054
rect -35343 18998 -35287 19054
rect -35287 18998 -35283 19054
rect -35347 18994 -35283 18998
rect -35267 19054 -35203 19058
rect -35267 18998 -35263 19054
rect -35263 18998 -35207 19054
rect -35207 18998 -35203 19054
rect -35267 18994 -35203 18998
rect -35187 19054 -35123 19058
rect -35187 18998 -35183 19054
rect -35183 18998 -35127 19054
rect -35127 18998 -35123 19054
rect -35187 18994 -35123 18998
rect -35107 19054 -35043 19058
rect -35107 18998 -35103 19054
rect -35103 18998 -35047 19054
rect -35047 18998 -35043 19054
rect -35107 18994 -35043 18998
rect -35027 19054 -34963 19058
rect -35027 18998 -35023 19054
rect -35023 18998 -34967 19054
rect -34967 18998 -34963 19054
rect -35027 18994 -34963 18998
rect -34947 19054 -34883 19058
rect -34947 18998 -34943 19054
rect -34943 18998 -34887 19054
rect -34887 18998 -34883 19054
rect -34947 18994 -34883 18998
rect -38145 16059 -38081 16063
rect -38145 16003 -38141 16059
rect -38141 16003 -38085 16059
rect -38085 16003 -38081 16059
rect -38145 15999 -38081 16003
rect -38065 16059 -38001 16063
rect -38065 16003 -38061 16059
rect -38061 16003 -38005 16059
rect -38005 16003 -38001 16059
rect -38065 15999 -38001 16003
rect -37985 16059 -37921 16063
rect -37985 16003 -37981 16059
rect -37981 16003 -37925 16059
rect -37925 16003 -37921 16059
rect -37985 15999 -37921 16003
rect -37905 16059 -37841 16063
rect -37905 16003 -37901 16059
rect -37901 16003 -37845 16059
rect -37845 16003 -37841 16059
rect -37905 15999 -37841 16003
rect -37825 16059 -37761 16063
rect -37825 16003 -37821 16059
rect -37821 16003 -37765 16059
rect -37765 16003 -37761 16059
rect -37825 15999 -37761 16003
rect -37745 16059 -37681 16063
rect -37745 16003 -37741 16059
rect -37741 16003 -37685 16059
rect -37685 16003 -37681 16059
rect -37745 15999 -37681 16003
rect -37665 16059 -37601 16063
rect -37665 16003 -37661 16059
rect -37661 16003 -37605 16059
rect -37605 16003 -37601 16059
rect -37665 15999 -37601 16003
rect -37585 16059 -37521 16063
rect -37585 16003 -37581 16059
rect -37581 16003 -37525 16059
rect -37525 16003 -37521 16059
rect -37585 15999 -37521 16003
rect -37505 16059 -37441 16063
rect -37505 16003 -37501 16059
rect -37501 16003 -37445 16059
rect -37445 16003 -37441 16059
rect -37505 15999 -37441 16003
rect -37425 16059 -37361 16063
rect -37425 16003 -37421 16059
rect -37421 16003 -37365 16059
rect -37365 16003 -37361 16059
rect -37425 15999 -37361 16003
rect -37345 16059 -37281 16063
rect -37345 16003 -37341 16059
rect -37341 16003 -37285 16059
rect -37285 16003 -37281 16059
rect -37345 15999 -37281 16003
rect -37265 16059 -37201 16063
rect -37265 16003 -37261 16059
rect -37261 16003 -37205 16059
rect -37205 16003 -37201 16059
rect -37265 15999 -37201 16003
rect -37185 16059 -37121 16063
rect -37185 16003 -37181 16059
rect -37181 16003 -37125 16059
rect -37125 16003 -37121 16059
rect -37185 15999 -37121 16003
rect -37105 16059 -37041 16063
rect -37105 16003 -37101 16059
rect -37101 16003 -37045 16059
rect -37045 16003 -37041 16059
rect -37105 15999 -37041 16003
rect -37025 16059 -36961 16063
rect -37025 16003 -37021 16059
rect -37021 16003 -36965 16059
rect -36965 16003 -36961 16059
rect -37025 15999 -36961 16003
rect -36945 16059 -36881 16063
rect -36945 16003 -36941 16059
rect -36941 16003 -36885 16059
rect -36885 16003 -36881 16059
rect -36945 15999 -36881 16003
rect -36865 16059 -36801 16063
rect -36865 16003 -36861 16059
rect -36861 16003 -36805 16059
rect -36805 16003 -36801 16059
rect -36865 15999 -36801 16003
rect -36785 16059 -36721 16063
rect -36785 16003 -36781 16059
rect -36781 16003 -36725 16059
rect -36725 16003 -36721 16059
rect -36785 15999 -36721 16003
rect -36705 16059 -36641 16063
rect -36705 16003 -36701 16059
rect -36701 16003 -36645 16059
rect -36645 16003 -36641 16059
rect -36705 15999 -36641 16003
rect -36625 16059 -36561 16063
rect -36625 16003 -36621 16059
rect -36621 16003 -36565 16059
rect -36565 16003 -36561 16059
rect -36625 15999 -36561 16003
rect -36545 16059 -36481 16063
rect -36545 16003 -36541 16059
rect -36541 16003 -36485 16059
rect -36485 16003 -36481 16059
rect -36545 15999 -36481 16003
rect -36465 16059 -36401 16063
rect -36465 16003 -36461 16059
rect -36461 16003 -36405 16059
rect -36405 16003 -36401 16059
rect -36465 15999 -36401 16003
rect -36385 16059 -36321 16063
rect -36385 16003 -36381 16059
rect -36381 16003 -36325 16059
rect -36325 16003 -36321 16059
rect -36385 15999 -36321 16003
rect -36305 16059 -36241 16063
rect -36305 16003 -36301 16059
rect -36301 16003 -36245 16059
rect -36245 16003 -36241 16059
rect -36305 15999 -36241 16003
rect -36225 16059 -36161 16063
rect -36225 16003 -36221 16059
rect -36221 16003 -36165 16059
rect -36165 16003 -36161 16059
rect -36225 15999 -36161 16003
rect -36145 16059 -36081 16063
rect -36145 16003 -36141 16059
rect -36141 16003 -36085 16059
rect -36085 16003 -36081 16059
rect -36145 15999 -36081 16003
rect -36065 16059 -36001 16063
rect -36065 16003 -36061 16059
rect -36061 16003 -36005 16059
rect -36005 16003 -36001 16059
rect -36065 15999 -36001 16003
rect -35985 16059 -35921 16063
rect -35985 16003 -35981 16059
rect -35981 16003 -35925 16059
rect -35925 16003 -35921 16059
rect -35985 15999 -35921 16003
rect -35905 16059 -35841 16063
rect -35905 16003 -35901 16059
rect -35901 16003 -35845 16059
rect -35845 16003 -35841 16059
rect -35905 15999 -35841 16003
rect -35825 16059 -35761 16063
rect -35825 16003 -35821 16059
rect -35821 16003 -35765 16059
rect -35765 16003 -35761 16059
rect -35825 15999 -35761 16003
rect -35745 16059 -35681 16063
rect -35745 16003 -35741 16059
rect -35741 16003 -35685 16059
rect -35685 16003 -35681 16059
rect -35745 15999 -35681 16003
rect -35665 16059 -35601 16063
rect -35665 16003 -35661 16059
rect -35661 16003 -35605 16059
rect -35605 16003 -35601 16059
rect -35665 15999 -35601 16003
rect -35585 16059 -35521 16063
rect -35585 16003 -35581 16059
rect -35581 16003 -35525 16059
rect -35525 16003 -35521 16059
rect -35585 15999 -35521 16003
rect -35505 16059 -35441 16063
rect -35505 16003 -35501 16059
rect -35501 16003 -35445 16059
rect -35445 16003 -35441 16059
rect -35505 15999 -35441 16003
rect -35425 16059 -35361 16063
rect -35425 16003 -35421 16059
rect -35421 16003 -35365 16059
rect -35365 16003 -35361 16059
rect -35425 15999 -35361 16003
rect -35345 16059 -35281 16063
rect -35345 16003 -35341 16059
rect -35341 16003 -35285 16059
rect -35285 16003 -35281 16059
rect -35345 15999 -35281 16003
rect -35265 16059 -35201 16063
rect -35265 16003 -35261 16059
rect -35261 16003 -35205 16059
rect -35205 16003 -35201 16059
rect -35265 15999 -35201 16003
rect -35185 16059 -35121 16063
rect -35185 16003 -35181 16059
rect -35181 16003 -35125 16059
rect -35125 16003 -35121 16059
rect -35185 15999 -35121 16003
rect -35105 16059 -35041 16063
rect -35105 16003 -35101 16059
rect -35101 16003 -35045 16059
rect -35045 16003 -35041 16059
rect -35105 15999 -35041 16003
rect -35025 16059 -34961 16063
rect -35025 16003 -35021 16059
rect -35021 16003 -34965 16059
rect -34965 16003 -34961 16059
rect -35025 15999 -34961 16003
rect -34945 16059 -34881 16063
rect -34945 16003 -34941 16059
rect -34941 16003 -34885 16059
rect -34885 16003 -34881 16059
rect -34945 15999 -34881 16003
rect 12936 20963 13000 21027
rect -25452 17882 -25388 17886
rect -25452 17826 -25448 17882
rect -25448 17826 -25392 17882
rect -25392 17826 -25388 17882
rect -25452 17822 -25388 17826
rect -25452 17802 -25388 17806
rect -25452 17746 -25448 17802
rect -25448 17746 -25392 17802
rect -25392 17746 -25388 17802
rect -25452 17742 -25388 17746
rect -25452 17722 -25388 17726
rect -25452 17666 -25448 17722
rect -25448 17666 -25392 17722
rect -25392 17666 -25388 17722
rect -25452 17662 -25388 17666
rect -25446 17394 -25382 17398
rect -25446 17338 -25442 17394
rect -25442 17338 -25386 17394
rect -25386 17338 -25382 17394
rect -25446 17334 -25382 17338
rect -25446 17314 -25382 17318
rect -25446 17258 -25442 17314
rect -25442 17258 -25386 17314
rect -25386 17258 -25382 17314
rect -25446 17254 -25382 17258
rect -25446 17234 -25382 17238
rect -25446 17178 -25442 17234
rect -25442 17178 -25386 17234
rect -25386 17178 -25382 17234
rect -25446 17174 -25382 17178
rect -16599 20587 -16535 20651
rect 11080 20270 11144 20334
rect -10416 17153 -10352 17157
rect -10416 17097 -10412 17153
rect -10412 17097 -10356 17153
rect -10356 17097 -10352 17153
rect -10416 17093 -10352 17097
rect -14152 15366 -14088 15370
rect -14152 15310 -14148 15366
rect -14148 15310 -14092 15366
rect -14092 15310 -14088 15366
rect -14152 15306 -14088 15310
rect -25513 14409 -25449 14413
rect -25513 14353 -25509 14409
rect -25509 14353 -25453 14409
rect -25453 14353 -25449 14409
rect -25513 14349 -25449 14353
rect -25513 14329 -25449 14333
rect -25513 14273 -25509 14329
rect -25509 14273 -25453 14329
rect -25453 14273 -25449 14329
rect -25513 14269 -25449 14273
rect -25513 14249 -25449 14253
rect -25513 14193 -25509 14249
rect -25509 14193 -25453 14249
rect -25453 14193 -25449 14249
rect -25513 14189 -25449 14193
rect -18223 14069 -18159 14073
rect -18223 14013 -18219 14069
rect -18219 14013 -18163 14069
rect -18163 14013 -18159 14069
rect -18223 14009 -18159 14013
rect -25514 13915 -25450 13919
rect -25514 13859 -25510 13915
rect -25510 13859 -25454 13915
rect -25454 13859 -25450 13915
rect -25514 13855 -25450 13859
rect -25514 13835 -25450 13839
rect -25514 13779 -25510 13835
rect -25510 13779 -25454 13835
rect -25454 13779 -25450 13835
rect -25514 13775 -25450 13779
rect -25514 13755 -25450 13759
rect -25514 13699 -25510 13755
rect -25510 13699 -25454 13755
rect -25454 13699 -25450 13755
rect -25514 13695 -25450 13699
rect -10970 10219 -10906 10223
rect -10970 10163 -10966 10219
rect -10966 10163 -10910 10219
rect -10910 10163 -10906 10219
rect -10970 10159 -10906 10163
rect 11476 19739 11540 19803
rect -2815 19449 -2751 19513
rect -5279 18979 -5215 19043
rect -3918 18979 -3854 19043
rect -5786 15704 -5722 15708
rect -5786 15648 -5782 15704
rect -5782 15648 -5726 15704
rect -5726 15648 -5722 15704
rect -5786 15644 -5722 15648
rect -4899 14409 -4835 14413
rect -4899 14353 -4895 14409
rect -4895 14353 -4839 14409
rect -4839 14353 -4835 14409
rect -4899 14349 -4835 14353
rect -4899 14329 -4835 14333
rect -4899 14273 -4895 14329
rect -4895 14273 -4839 14329
rect -4839 14273 -4835 14329
rect -4899 14269 -4835 14273
rect -6162 10823 -6098 10827
rect -6162 10767 -6158 10823
rect -6158 10767 -6102 10823
rect -6102 10767 -6098 10823
rect -6162 10763 -6098 10767
rect -6082 10823 -6018 10827
rect -6082 10767 -6078 10823
rect -6078 10767 -6022 10823
rect -6022 10767 -6018 10823
rect -6082 10763 -6018 10767
rect -6002 10823 -5938 10827
rect -6002 10767 -5998 10823
rect -5998 10767 -5942 10823
rect -5942 10767 -5938 10823
rect -6002 10763 -5938 10767
rect -6160 9580 -6096 9584
rect -6160 9524 -6156 9580
rect -6156 9524 -6100 9580
rect -6100 9524 -6096 9580
rect -6160 9520 -6096 9524
rect -6080 9580 -6016 9584
rect -6080 9524 -6076 9580
rect -6076 9524 -6020 9580
rect -6020 9524 -6016 9580
rect -6080 9520 -6016 9524
rect -6000 9580 -5936 9584
rect -6000 9524 -5996 9580
rect -5996 9524 -5940 9580
rect -5940 9524 -5936 9580
rect -6000 9520 -5936 9524
rect 14687 19323 14751 19327
rect 14687 19267 14691 19323
rect 14691 19267 14747 19323
rect 14747 19267 14751 19323
rect 14687 19263 14751 19267
rect 23689 19378 23753 19382
rect 23689 19322 23693 19378
rect 23693 19322 23749 19378
rect 23749 19322 23753 19378
rect 23689 19318 23753 19322
rect -2398 19148 -2334 19212
rect 4873 19168 5177 19172
rect 4873 19032 4877 19168
rect 4877 19032 5173 19168
rect 5173 19032 5177 19168
rect 4873 19028 5177 19032
rect 10232 19054 10296 19058
rect 10232 18998 10236 19054
rect 10236 18998 10292 19054
rect 10292 18998 10296 19054
rect 10232 18994 10296 18998
rect 20971 19058 21035 19062
rect 20971 19002 20975 19058
rect 20975 19002 21031 19058
rect 21031 19002 21035 19058
rect 20971 18998 21035 19002
rect -1504 18846 -1440 18910
rect -1133 18587 -1069 18651
rect 8280 18714 8344 18718
rect 8280 18658 8284 18714
rect 8284 18658 8340 18714
rect 8340 18658 8344 18714
rect 8280 18654 8344 18658
rect 12930 18624 12994 18688
rect 14115 18507 14179 18571
rect 25614 18507 25678 18571
rect -680 18248 -616 18312
rect -284 17967 -220 18031
rect -3172 17632 -2788 17856
rect 14368 17699 14432 17763
rect 25361 17700 25425 17764
rect 981 17461 1045 17525
rect 14689 17538 14753 17542
rect 14689 17482 14693 17538
rect 14693 17482 14749 17538
rect 14749 17482 14753 17538
rect 14689 17478 14753 17482
rect 23689 17548 23753 17552
rect 23689 17492 23693 17548
rect 23693 17492 23749 17548
rect 23749 17492 23753 17548
rect 23689 17488 23753 17492
rect 4295 17285 4359 17289
rect 4295 17229 4299 17285
rect 4299 17229 4355 17285
rect 4355 17229 4359 17285
rect 4295 17225 4359 17229
rect 6227 17285 6291 17289
rect 6227 17229 6231 17285
rect 6231 17229 6287 17285
rect 6287 17229 6291 17285
rect 6227 17225 6291 17229
rect 12956 17019 13020 17083
rect 263 16410 11127 16414
rect 263 16274 267 16410
rect 267 16274 11123 16410
rect 11123 16274 11127 16410
rect 263 16270 11127 16274
rect -3509 16141 -3445 16205
rect -3928 15390 -3864 15454
rect -3135 14966 -3071 14970
rect -3135 14910 -3131 14966
rect -3131 14910 -3075 14966
rect -3075 14910 -3071 14966
rect -3135 14906 -3071 14910
rect -3135 14886 -3071 14890
rect -3135 14830 -3131 14886
rect -3131 14830 -3075 14886
rect -3075 14830 -3071 14886
rect -3135 14826 -3071 14830
rect -3135 14806 -3071 14810
rect -3135 14750 -3131 14806
rect -3131 14750 -3075 14806
rect -3075 14750 -3071 14806
rect -3135 14746 -3071 14750
rect -3509 14580 -3445 14644
rect -3185 8643 -3121 8707
rect -16749 7603 -16685 7607
rect -16749 7547 -16745 7603
rect -16745 7547 -16689 7603
rect -16689 7547 -16685 7603
rect -16749 7543 -16685 7547
rect -1799 13117 -1735 13121
rect -1799 13061 -1795 13117
rect -1795 13061 -1739 13117
rect -1739 13061 -1735 13117
rect -1799 13057 -1735 13061
rect -1799 13037 -1735 13041
rect -1799 12981 -1795 13037
rect -1795 12981 -1739 13037
rect -1739 12981 -1735 13037
rect -1799 12977 -1735 12981
rect -1799 12957 -1735 12961
rect -1799 12901 -1795 12957
rect -1795 12901 -1739 12957
rect -1739 12901 -1735 12957
rect -1799 12897 -1735 12901
rect -1799 12877 -1735 12881
rect -1799 12821 -1795 12877
rect -1795 12821 -1739 12877
rect -1739 12821 -1735 12877
rect -1799 12817 -1735 12821
rect -1799 12797 -1735 12801
rect -1799 12741 -1795 12797
rect -1795 12741 -1739 12797
rect -1739 12741 -1735 12797
rect -1799 12737 -1735 12741
rect -1758 11522 -1694 11526
rect -1758 11466 -1754 11522
rect -1754 11466 -1698 11522
rect -1698 11466 -1694 11522
rect -1758 11462 -1694 11466
rect -1758 11442 -1694 11446
rect -1758 11386 -1754 11442
rect -1754 11386 -1698 11442
rect -1698 11386 -1694 11442
rect -1758 11382 -1694 11386
rect -1758 11362 -1694 11366
rect -1758 11306 -1754 11362
rect -1754 11306 -1698 11362
rect -1698 11306 -1694 11362
rect -1758 11302 -1694 11306
rect -1758 11282 -1694 11286
rect -1758 11226 -1754 11282
rect -1754 11226 -1698 11282
rect -1698 11226 -1694 11282
rect -1758 11222 -1694 11226
rect -1758 11202 -1694 11206
rect -1758 11146 -1754 11202
rect -1754 11146 -1698 11202
rect -1698 11146 -1694 11202
rect -1758 11142 -1694 11146
rect -7175 7231 -6791 7235
rect -7175 7015 -6791 7231
rect -7175 7011 -6791 7015
rect -25516 6646 -25452 6650
rect -25516 6590 -25512 6646
rect -25512 6590 -25456 6646
rect -25456 6590 -25452 6646
rect -25516 6586 -25452 6590
rect -25516 6566 -25452 6570
rect -25516 6510 -25512 6566
rect -25512 6510 -25456 6566
rect -25456 6510 -25452 6566
rect -25516 6506 -25452 6510
rect -25516 6486 -25452 6490
rect -25516 6430 -25512 6486
rect -25512 6430 -25456 6486
rect -25456 6430 -25452 6486
rect -25516 6426 -25452 6430
rect -3184 6585 -3120 6649
rect -18251 6299 -18187 6303
rect -18251 6243 -18247 6299
rect -18247 6243 -18191 6299
rect -18191 6243 -18187 6299
rect -18251 6239 -18187 6243
rect -25517 6159 -25453 6163
rect -25517 6103 -25513 6159
rect -25513 6103 -25457 6159
rect -25457 6103 -25453 6159
rect -25517 6099 -25453 6103
rect -25517 6079 -25453 6083
rect -25517 6023 -25513 6079
rect -25513 6023 -25457 6079
rect -25457 6023 -25453 6079
rect -25517 6019 -25453 6023
rect -25517 5999 -25453 6003
rect -25517 5943 -25513 5999
rect -25513 5943 -25457 5999
rect -25457 5943 -25453 5999
rect -25517 5939 -25453 5943
rect -4906 6124 -4842 6128
rect -4906 6068 -4902 6124
rect -4902 6068 -4846 6124
rect -4846 6068 -4842 6124
rect -4906 6064 -4842 6068
rect -4906 6044 -4842 6048
rect -4906 5988 -4902 6044
rect -4902 5988 -4846 6044
rect -4846 5988 -4842 6044
rect -4906 5984 -4842 5988
rect -3928 5978 -3864 6042
rect -3184 5544 -3120 5548
rect -3184 5488 -3180 5544
rect -3180 5488 -3124 5544
rect -3124 5488 -3120 5544
rect -3184 5484 -3120 5488
rect -3184 5464 -3120 5468
rect -3184 5408 -3180 5464
rect -3180 5408 -3124 5464
rect -3124 5408 -3120 5464
rect -3184 5404 -3120 5408
rect -3184 5384 -3120 5388
rect -3184 5328 -3180 5384
rect -3180 5328 -3124 5384
rect -3124 5328 -3120 5384
rect -3184 5324 -3120 5328
rect -3509 5169 -3445 5233
rect -1759 9919 -1695 9923
rect -1759 9863 -1755 9919
rect -1755 9863 -1699 9919
rect -1699 9863 -1695 9919
rect -1759 9859 -1695 9863
rect -1759 9839 -1695 9843
rect -1759 9783 -1755 9839
rect -1755 9783 -1699 9839
rect -1699 9783 -1695 9839
rect -1759 9779 -1695 9783
rect -1759 9759 -1695 9763
rect -1759 9703 -1755 9759
rect -1755 9703 -1699 9759
rect -1699 9703 -1695 9759
rect -1759 9699 -1695 9703
rect -1759 9679 -1695 9683
rect -1759 9623 -1755 9679
rect -1755 9623 -1699 9679
rect -1699 9623 -1695 9679
rect -1759 9619 -1695 9623
rect -1759 9599 -1695 9603
rect -1759 9543 -1755 9599
rect -1755 9543 -1699 9599
rect -1699 9543 -1695 9599
rect -1759 9539 -1695 9543
rect 14686 15707 14750 15711
rect 14686 15651 14690 15707
rect 14690 15651 14746 15707
rect 14746 15651 14750 15707
rect 14686 15647 14750 15651
rect 23686 15784 23750 15788
rect 23686 15728 23690 15784
rect 23690 15728 23746 15784
rect 23746 15728 23750 15784
rect 23686 15724 23750 15728
rect 20928 15492 20992 15496
rect 20928 15436 20932 15492
rect 20932 15436 20988 15492
rect 20988 15436 20992 15492
rect 20928 15432 20992 15436
rect 12973 15164 13037 15228
rect 14685 13961 14749 13965
rect 14685 13905 14689 13961
rect 14689 13905 14745 13961
rect 14745 13905 14749 13961
rect 14685 13901 14749 13905
rect 23686 13993 23750 13997
rect 23686 13937 23690 13993
rect 23690 13937 23746 13993
rect 23746 13937 23750 13993
rect 23686 13933 23750 13937
rect 13003 13464 13067 13528
rect 14115 13107 14179 13171
rect 14368 12299 14432 12363
rect 14702 12176 14766 12180
rect 14702 12120 14706 12176
rect 14706 12120 14762 12176
rect 14762 12120 14766 12176
rect 14702 12116 14766 12120
rect 23691 12186 23755 12190
rect 23691 12130 23695 12186
rect 23695 12130 23751 12186
rect 23751 12130 23755 12186
rect 23691 12126 23755 12130
rect 20985 11902 21049 11906
rect 20985 11846 20989 11902
rect 20989 11846 21045 11902
rect 21045 11846 21049 11902
rect 20985 11842 21049 11846
rect 13001 11612 13065 11676
rect 6498 10514 11202 10518
rect 6498 10378 6502 10514
rect 6502 10378 11198 10514
rect 11198 10378 11202 10514
rect 6498 10374 11202 10378
rect 14691 10379 14755 10383
rect 14691 10323 14695 10379
rect 14695 10323 14751 10379
rect 14751 10323 14755 10379
rect 14691 10319 14755 10323
rect 23691 10376 23755 10380
rect 23691 10320 23695 10376
rect 23695 10320 23751 10376
rect 23751 10320 23755 10376
rect 23691 10316 23755 10320
rect 36066 9150 36130 9154
rect 36066 9094 36070 9150
rect 36070 9094 36126 9150
rect 36126 9094 36130 9150
rect 36066 9090 36130 9094
rect -1756 8318 -1692 8322
rect -1756 8262 -1752 8318
rect -1752 8262 -1696 8318
rect -1696 8262 -1692 8318
rect -1756 8258 -1692 8262
rect -1756 8238 -1692 8242
rect -1756 8182 -1752 8238
rect -1752 8182 -1696 8238
rect -1696 8182 -1692 8238
rect -1756 8178 -1692 8182
rect -1756 8158 -1692 8162
rect -1756 8102 -1752 8158
rect -1752 8102 -1696 8158
rect -1696 8102 -1692 8158
rect -1756 8098 -1692 8102
rect -1756 8078 -1692 8082
rect -1756 8022 -1752 8078
rect -1752 8022 -1696 8078
rect -1696 8022 -1692 8078
rect -1756 8018 -1692 8022
rect -1756 7998 -1692 8002
rect -1756 7942 -1752 7998
rect -1752 7942 -1696 7998
rect -1696 7942 -1692 7998
rect -1756 7938 -1692 7942
rect 36907 8562 37131 8786
rect 35489 8527 35553 8531
rect 35489 8471 35493 8527
rect 35493 8471 35549 8527
rect 35549 8471 35553 8527
rect 35489 8467 35553 8471
rect 36631 8465 36695 8469
rect 36631 8409 36635 8465
rect 36635 8409 36691 8465
rect 36691 8409 36695 8465
rect 36631 8405 36695 8409
rect 35028 7219 35092 7223
rect 35028 7163 35032 7219
rect 35032 7163 35088 7219
rect 35088 7163 35092 7219
rect 38576 7537 38640 7541
rect 38576 7481 38580 7537
rect 38580 7481 38636 7537
rect 38636 7481 38640 7537
rect 38576 7477 38640 7481
rect 38576 7457 38640 7461
rect 38576 7401 38580 7457
rect 38580 7401 38636 7457
rect 38636 7401 38640 7457
rect 38576 7397 38640 7401
rect 36987 7269 37051 7333
rect 35028 7159 35092 7163
rect 40095 7550 40159 7554
rect 40095 7494 40099 7550
rect 40099 7494 40155 7550
rect 40155 7494 40159 7550
rect 40095 7490 40159 7494
rect 40095 7470 40159 7474
rect 40095 7414 40099 7470
rect 40099 7414 40155 7470
rect 40155 7414 40159 7470
rect 40095 7410 40159 7414
rect 40840 6938 41224 7162
rect 42630 7215 42694 7219
rect 42630 7159 42634 7215
rect 42634 7159 42690 7215
rect 42690 7159 42694 7215
rect 42630 7155 42694 7159
rect 42710 7215 42774 7219
rect 42710 7159 42714 7215
rect 42714 7159 42770 7215
rect 42770 7159 42774 7215
rect 42710 7155 42774 7159
rect 42790 7215 42854 7219
rect 42790 7159 42794 7215
rect 42794 7159 42850 7215
rect 42850 7159 42854 7215
rect 42790 7155 42854 7159
rect 42870 7215 42934 7219
rect 42870 7159 42874 7215
rect 42874 7159 42930 7215
rect 42930 7159 42934 7215
rect 42870 7155 42934 7159
rect 42950 7215 43014 7219
rect 42950 7159 42954 7215
rect 42954 7159 43010 7215
rect 43010 7159 43014 7215
rect 42950 7155 43014 7159
rect 43030 7215 43094 7219
rect 43030 7159 43034 7215
rect 43034 7159 43090 7215
rect 43090 7159 43094 7215
rect 43030 7155 43094 7159
rect 43110 7215 43174 7219
rect 43110 7159 43114 7215
rect 43114 7159 43170 7215
rect 43170 7159 43174 7215
rect 43110 7155 43174 7159
rect 43190 7215 43254 7219
rect 43190 7159 43194 7215
rect 43194 7159 43250 7215
rect 43250 7159 43254 7215
rect 43190 7155 43254 7159
rect 43270 7215 43334 7219
rect 43270 7159 43274 7215
rect 43274 7159 43330 7215
rect 43330 7159 43334 7215
rect 43270 7155 43334 7159
rect 43350 7215 43414 7219
rect 43350 7159 43354 7215
rect 43354 7159 43410 7215
rect 43410 7159 43414 7215
rect 43350 7155 43414 7159
rect 43430 7215 43494 7219
rect 43430 7159 43434 7215
rect 43434 7159 43490 7215
rect 43490 7159 43494 7215
rect 43430 7155 43494 7159
rect 43510 7215 43574 7219
rect 43510 7159 43514 7215
rect 43514 7159 43570 7215
rect 43570 7159 43574 7215
rect 43510 7155 43574 7159
rect 43590 7215 43654 7219
rect 43590 7159 43594 7215
rect 43594 7159 43650 7215
rect 43650 7159 43654 7215
rect 43590 7155 43654 7159
rect 43670 7215 43734 7219
rect 43670 7159 43674 7215
rect 43674 7159 43730 7215
rect 43730 7159 43734 7215
rect 43670 7155 43734 7159
rect 43750 7215 43814 7219
rect 43750 7159 43754 7215
rect 43754 7159 43810 7215
rect 43810 7159 43814 7215
rect 43750 7155 43814 7159
rect 43830 7215 43894 7219
rect 43830 7159 43834 7215
rect 43834 7159 43890 7215
rect 43890 7159 43894 7215
rect 43830 7155 43894 7159
rect 43910 7215 43974 7219
rect 43910 7159 43914 7215
rect 43914 7159 43970 7215
rect 43970 7159 43974 7215
rect 43910 7155 43974 7159
rect 43990 7215 44054 7219
rect 43990 7159 43994 7215
rect 43994 7159 44050 7215
rect 44050 7159 44054 7215
rect 43990 7155 44054 7159
rect 44070 7215 44134 7219
rect 44070 7159 44074 7215
rect 44074 7159 44130 7215
rect 44130 7159 44134 7215
rect 44070 7155 44134 7159
rect 44150 7215 44214 7219
rect 44150 7159 44154 7215
rect 44154 7159 44210 7215
rect 44210 7159 44214 7215
rect 44150 7155 44214 7159
rect 44230 7215 44294 7219
rect 44230 7159 44234 7215
rect 44234 7159 44290 7215
rect 44290 7159 44294 7215
rect 44230 7155 44294 7159
rect 44310 7215 44374 7219
rect 44310 7159 44314 7215
rect 44314 7159 44370 7215
rect 44370 7159 44374 7215
rect 44310 7155 44374 7159
rect 44390 7215 44454 7219
rect 44390 7159 44394 7215
rect 44394 7159 44450 7215
rect 44450 7159 44454 7215
rect 44390 7155 44454 7159
rect 44470 7215 44534 7219
rect 44470 7159 44474 7215
rect 44474 7159 44530 7215
rect 44530 7159 44534 7215
rect 44470 7155 44534 7159
rect 44550 7215 44614 7219
rect 44550 7159 44554 7215
rect 44554 7159 44610 7215
rect 44610 7159 44614 7215
rect 44550 7155 44614 7159
rect 44630 7215 44694 7219
rect 44630 7159 44634 7215
rect 44634 7159 44690 7215
rect 44690 7159 44694 7215
rect 44630 7155 44694 7159
rect 44710 7215 44774 7219
rect 44710 7159 44714 7215
rect 44714 7159 44770 7215
rect 44770 7159 44774 7215
rect 44710 7155 44774 7159
rect 44790 7215 44854 7219
rect 44790 7159 44794 7215
rect 44794 7159 44850 7215
rect 44850 7159 44854 7215
rect 44790 7155 44854 7159
rect 44870 7215 44934 7219
rect 44870 7159 44874 7215
rect 44874 7159 44930 7215
rect 44930 7159 44934 7215
rect 44870 7155 44934 7159
rect 44950 7215 45014 7219
rect 44950 7159 44954 7215
rect 44954 7159 45010 7215
rect 45010 7159 45014 7215
rect 44950 7155 45014 7159
rect 45030 7215 45094 7219
rect 45030 7159 45034 7215
rect 45034 7159 45090 7215
rect 45090 7159 45094 7215
rect 45030 7155 45094 7159
rect 45110 7215 45174 7219
rect 45110 7159 45114 7215
rect 45114 7159 45170 7215
rect 45170 7159 45174 7215
rect 45110 7155 45174 7159
rect 45190 7215 45254 7219
rect 45190 7159 45194 7215
rect 45194 7159 45250 7215
rect 45250 7159 45254 7215
rect 45190 7155 45254 7159
rect 45270 7215 45334 7219
rect 45270 7159 45274 7215
rect 45274 7159 45330 7215
rect 45330 7159 45334 7215
rect 45270 7155 45334 7159
rect 45350 7215 45414 7219
rect 45350 7159 45354 7215
rect 45354 7159 45410 7215
rect 45410 7159 45414 7215
rect 45350 7155 45414 7159
rect 45430 7215 45494 7219
rect 45430 7159 45434 7215
rect 45434 7159 45490 7215
rect 45490 7159 45494 7215
rect 45430 7155 45494 7159
rect 45510 7215 45574 7219
rect 45510 7159 45514 7215
rect 45514 7159 45570 7215
rect 45570 7159 45574 7215
rect 45510 7155 45574 7159
rect 45590 7215 45654 7219
rect 45590 7159 45594 7215
rect 45594 7159 45650 7215
rect 45650 7159 45654 7215
rect 45590 7155 45654 7159
rect 45670 7215 45734 7219
rect 45670 7159 45674 7215
rect 45674 7159 45730 7215
rect 45730 7159 45734 7215
rect 45670 7155 45734 7159
rect 45750 7215 45814 7219
rect 45750 7159 45754 7215
rect 45754 7159 45810 7215
rect 45810 7159 45814 7215
rect 45750 7155 45814 7159
rect 45830 7215 45894 7219
rect 45830 7159 45834 7215
rect 45834 7159 45890 7215
rect 45890 7159 45894 7215
rect 45830 7155 45894 7159
rect 35027 5881 35091 5885
rect 35027 5825 35031 5881
rect 35031 5825 35087 5881
rect 35087 5825 35091 5881
rect 35027 5821 35091 5825
rect 36987 6245 37051 6249
rect 36987 6189 36991 6245
rect 36991 6189 37047 6245
rect 37047 6189 37051 6245
rect 36987 6185 37051 6189
rect 38571 6206 38635 6210
rect 38571 6150 38575 6206
rect 38575 6150 38631 6206
rect 38631 6150 38635 6206
rect 38571 6146 38635 6150
rect 38571 6126 38635 6130
rect 38571 6070 38575 6126
rect 38575 6070 38631 6126
rect 38631 6070 38635 6126
rect 38571 6066 38635 6070
rect 40100 6203 40164 6207
rect 40100 6147 40104 6203
rect 40104 6147 40160 6203
rect 40160 6147 40164 6203
rect 40100 6143 40164 6147
rect 40100 6123 40164 6127
rect 40100 6067 40104 6123
rect 40104 6067 40160 6123
rect 40160 6067 40164 6123
rect 40100 6063 40164 6067
rect 36987 5097 37051 5161
rect 38570 4853 38634 4857
rect 38570 4797 38574 4853
rect 38574 4797 38630 4853
rect 38630 4797 38634 4853
rect 38570 4793 38634 4797
rect 38570 4773 38634 4777
rect 38570 4717 38574 4773
rect 38574 4717 38630 4773
rect 38630 4717 38634 4773
rect 38570 4713 38634 4717
rect 35035 4488 35099 4492
rect 35035 4432 35039 4488
rect 35039 4432 35095 4488
rect 35095 4432 35099 4488
rect 35035 4428 35099 4432
rect 36988 4069 37052 4073
rect 36988 4013 36992 4069
rect 36992 4013 37048 4069
rect 37048 4013 37052 4069
rect 36988 4009 37052 4013
rect 40100 4831 40164 4835
rect 40100 4775 40104 4831
rect 40104 4775 40160 4831
rect 40160 4775 40164 4831
rect 40100 4771 40164 4775
rect 40100 4751 40164 4755
rect 40100 4695 40104 4751
rect 40104 4695 40160 4751
rect 40160 4695 40164 4751
rect 40100 4691 40164 4695
rect 40838 4035 41222 4259
rect 42607 4216 42671 4220
rect 42607 4160 42611 4216
rect 42611 4160 42667 4216
rect 42667 4160 42671 4216
rect 42607 4156 42671 4160
rect 42687 4216 42751 4220
rect 42687 4160 42691 4216
rect 42691 4160 42747 4216
rect 42747 4160 42751 4216
rect 42687 4156 42751 4160
rect 42767 4216 42831 4220
rect 42767 4160 42771 4216
rect 42771 4160 42827 4216
rect 42827 4160 42831 4216
rect 42767 4156 42831 4160
rect 42847 4216 42911 4220
rect 42847 4160 42851 4216
rect 42851 4160 42907 4216
rect 42907 4160 42911 4216
rect 42847 4156 42911 4160
rect 42927 4216 42991 4220
rect 42927 4160 42931 4216
rect 42931 4160 42987 4216
rect 42987 4160 42991 4216
rect 42927 4156 42991 4160
rect 43007 4216 43071 4220
rect 43007 4160 43011 4216
rect 43011 4160 43067 4216
rect 43067 4160 43071 4216
rect 43007 4156 43071 4160
rect 43087 4216 43151 4220
rect 43087 4160 43091 4216
rect 43091 4160 43147 4216
rect 43147 4160 43151 4216
rect 43087 4156 43151 4160
rect 43167 4216 43231 4220
rect 43167 4160 43171 4216
rect 43171 4160 43227 4216
rect 43227 4160 43231 4216
rect 43167 4156 43231 4160
rect 43247 4216 43311 4220
rect 43247 4160 43251 4216
rect 43251 4160 43307 4216
rect 43307 4160 43311 4216
rect 43247 4156 43311 4160
rect 43327 4216 43391 4220
rect 43327 4160 43331 4216
rect 43331 4160 43387 4216
rect 43387 4160 43391 4216
rect 43327 4156 43391 4160
rect 43407 4216 43471 4220
rect 43407 4160 43411 4216
rect 43411 4160 43467 4216
rect 43467 4160 43471 4216
rect 43407 4156 43471 4160
rect 43487 4216 43551 4220
rect 43487 4160 43491 4216
rect 43491 4160 43547 4216
rect 43547 4160 43551 4216
rect 43487 4156 43551 4160
rect 43567 4216 43631 4220
rect 43567 4160 43571 4216
rect 43571 4160 43627 4216
rect 43627 4160 43631 4216
rect 43567 4156 43631 4160
rect 43647 4216 43711 4220
rect 43647 4160 43651 4216
rect 43651 4160 43707 4216
rect 43707 4160 43711 4216
rect 43647 4156 43711 4160
rect 43727 4216 43791 4220
rect 43727 4160 43731 4216
rect 43731 4160 43787 4216
rect 43787 4160 43791 4216
rect 43727 4156 43791 4160
rect 43807 4216 43871 4220
rect 43807 4160 43811 4216
rect 43811 4160 43867 4216
rect 43867 4160 43871 4216
rect 43807 4156 43871 4160
rect 43887 4216 43951 4220
rect 43887 4160 43891 4216
rect 43891 4160 43947 4216
rect 43947 4160 43951 4216
rect 43887 4156 43951 4160
rect 43967 4216 44031 4220
rect 43967 4160 43971 4216
rect 43971 4160 44027 4216
rect 44027 4160 44031 4216
rect 43967 4156 44031 4160
rect 44047 4216 44111 4220
rect 44047 4160 44051 4216
rect 44051 4160 44107 4216
rect 44107 4160 44111 4216
rect 44047 4156 44111 4160
rect 44127 4216 44191 4220
rect 44127 4160 44131 4216
rect 44131 4160 44187 4216
rect 44187 4160 44191 4216
rect 44127 4156 44191 4160
rect 44207 4216 44271 4220
rect 44207 4160 44211 4216
rect 44211 4160 44267 4216
rect 44267 4160 44271 4216
rect 44207 4156 44271 4160
rect 44287 4216 44351 4220
rect 44287 4160 44291 4216
rect 44291 4160 44347 4216
rect 44347 4160 44351 4216
rect 44287 4156 44351 4160
rect 44367 4216 44431 4220
rect 44367 4160 44371 4216
rect 44371 4160 44427 4216
rect 44427 4160 44431 4216
rect 44367 4156 44431 4160
rect 44447 4216 44511 4220
rect 44447 4160 44451 4216
rect 44451 4160 44507 4216
rect 44507 4160 44511 4216
rect 44447 4156 44511 4160
rect 44527 4216 44591 4220
rect 44527 4160 44531 4216
rect 44531 4160 44587 4216
rect 44587 4160 44591 4216
rect 44527 4156 44591 4160
rect 44607 4216 44671 4220
rect 44607 4160 44611 4216
rect 44611 4160 44667 4216
rect 44667 4160 44671 4216
rect 44607 4156 44671 4160
rect 44687 4216 44751 4220
rect 44687 4160 44691 4216
rect 44691 4160 44747 4216
rect 44747 4160 44751 4216
rect 44687 4156 44751 4160
rect 44767 4216 44831 4220
rect 44767 4160 44771 4216
rect 44771 4160 44827 4216
rect 44827 4160 44831 4216
rect 44767 4156 44831 4160
rect 44847 4216 44911 4220
rect 44847 4160 44851 4216
rect 44851 4160 44907 4216
rect 44907 4160 44911 4216
rect 44847 4156 44911 4160
rect 44927 4216 44991 4220
rect 44927 4160 44931 4216
rect 44931 4160 44987 4216
rect 44987 4160 44991 4216
rect 44927 4156 44991 4160
rect 45007 4216 45071 4220
rect 45007 4160 45011 4216
rect 45011 4160 45067 4216
rect 45067 4160 45071 4216
rect 45007 4156 45071 4160
rect 45087 4216 45151 4220
rect 45087 4160 45091 4216
rect 45091 4160 45147 4216
rect 45147 4160 45151 4216
rect 45087 4156 45151 4160
rect 45167 4216 45231 4220
rect 45167 4160 45171 4216
rect 45171 4160 45227 4216
rect 45227 4160 45231 4216
rect 45167 4156 45231 4160
rect 45247 4216 45311 4220
rect 45247 4160 45251 4216
rect 45251 4160 45307 4216
rect 45307 4160 45311 4216
rect 45247 4156 45311 4160
rect 45327 4216 45391 4220
rect 45327 4160 45331 4216
rect 45331 4160 45387 4216
rect 45387 4160 45391 4216
rect 45327 4156 45391 4160
rect 45407 4216 45471 4220
rect 45407 4160 45411 4216
rect 45411 4160 45467 4216
rect 45467 4160 45471 4216
rect 45407 4156 45471 4160
rect 45487 4216 45551 4220
rect 45487 4160 45491 4216
rect 45491 4160 45547 4216
rect 45547 4160 45551 4216
rect 45487 4156 45551 4160
rect 45567 4216 45631 4220
rect 45567 4160 45571 4216
rect 45571 4160 45627 4216
rect 45627 4160 45631 4216
rect 45567 4156 45631 4160
rect 45647 4216 45711 4220
rect 45647 4160 45651 4216
rect 45651 4160 45707 4216
rect 45707 4160 45711 4216
rect 45647 4156 45711 4160
rect 45727 4216 45791 4220
rect 45727 4160 45731 4216
rect 45731 4160 45787 4216
rect 45787 4160 45791 4216
rect 45727 4156 45791 4160
rect 45807 4216 45871 4220
rect 45807 4160 45811 4216
rect 45811 4160 45867 4216
rect 45867 4160 45871 4216
rect 45807 4156 45871 4160
rect 45887 4216 45951 4220
rect 45887 4160 45891 4216
rect 45891 4160 45947 4216
rect 45947 4160 45951 4216
rect 45887 4156 45951 4160
rect 35031 3118 35095 3122
rect 35031 3062 35035 3118
rect 35035 3062 35091 3118
rect 35091 3062 35095 3118
rect 38573 3453 38637 3457
rect 38573 3397 38577 3453
rect 38577 3397 38633 3453
rect 38633 3397 38637 3453
rect 38573 3393 38637 3397
rect 38573 3373 38637 3377
rect 38573 3317 38577 3373
rect 38577 3317 38633 3373
rect 38633 3317 38637 3373
rect 38573 3313 38637 3317
rect 40097 3447 40161 3451
rect 40097 3391 40101 3447
rect 40101 3391 40157 3447
rect 40157 3391 40161 3447
rect 40097 3387 40161 3391
rect 40097 3367 40161 3371
rect 40097 3311 40101 3367
rect 40101 3311 40157 3367
rect 40157 3311 40161 3367
rect 40097 3307 40161 3311
rect 35031 3058 35095 3062
rect 36066 2210 36130 2214
rect 36066 2154 36070 2210
rect 36070 2154 36126 2210
rect 36126 2154 36130 2210
rect 36066 2150 36130 2154
rect 36907 1622 37131 1846
rect 35489 1587 35553 1591
rect 35489 1531 35493 1587
rect 35493 1531 35549 1587
rect 35549 1531 35553 1587
rect 35489 1527 35553 1531
rect 36631 1525 36695 1529
rect 36631 1469 36635 1525
rect 36635 1469 36691 1525
rect 36691 1469 36695 1525
rect 36631 1465 36695 1469
rect 322 217 21106 221
rect 322 81 326 217
rect 326 81 21102 217
rect 21102 81 21106 217
rect 322 77 21106 81
rect 35028 279 35092 283
rect 35028 223 35032 279
rect 35032 223 35088 279
rect 35088 223 35092 279
rect 38576 597 38640 601
rect 38576 541 38580 597
rect 38580 541 38636 597
rect 38636 541 38640 597
rect 38576 537 38640 541
rect 38576 517 38640 521
rect 38576 461 38580 517
rect 38580 461 38636 517
rect 38636 461 38640 517
rect 38576 457 38640 461
rect 36987 329 37051 393
rect 35028 219 35092 223
rect 40095 610 40159 614
rect 40095 554 40099 610
rect 40099 554 40155 610
rect 40155 554 40159 610
rect 40095 550 40159 554
rect 40095 530 40159 534
rect 40095 474 40099 530
rect 40099 474 40155 530
rect 40155 474 40159 530
rect 40095 470 40159 474
rect 40840 -2 41224 222
rect 42632 282 42696 286
rect 42632 226 42636 282
rect 42636 226 42692 282
rect 42692 226 42696 282
rect 42632 222 42696 226
rect 42712 282 42776 286
rect 42712 226 42716 282
rect 42716 226 42772 282
rect 42772 226 42776 282
rect 42712 222 42776 226
rect 42792 282 42856 286
rect 42792 226 42796 282
rect 42796 226 42852 282
rect 42852 226 42856 282
rect 42792 222 42856 226
rect 42872 282 42936 286
rect 42872 226 42876 282
rect 42876 226 42932 282
rect 42932 226 42936 282
rect 42872 222 42936 226
rect 42952 282 43016 286
rect 42952 226 42956 282
rect 42956 226 43012 282
rect 43012 226 43016 282
rect 42952 222 43016 226
rect 43032 282 43096 286
rect 43032 226 43036 282
rect 43036 226 43092 282
rect 43092 226 43096 282
rect 43032 222 43096 226
rect 43112 282 43176 286
rect 43112 226 43116 282
rect 43116 226 43172 282
rect 43172 226 43176 282
rect 43112 222 43176 226
rect 43192 282 43256 286
rect 43192 226 43196 282
rect 43196 226 43252 282
rect 43252 226 43256 282
rect 43192 222 43256 226
rect 43272 282 43336 286
rect 43272 226 43276 282
rect 43276 226 43332 282
rect 43332 226 43336 282
rect 43272 222 43336 226
rect 43352 282 43416 286
rect 43352 226 43356 282
rect 43356 226 43412 282
rect 43412 226 43416 282
rect 43352 222 43416 226
rect 43432 282 43496 286
rect 43432 226 43436 282
rect 43436 226 43492 282
rect 43492 226 43496 282
rect 43432 222 43496 226
rect 43512 282 43576 286
rect 43512 226 43516 282
rect 43516 226 43572 282
rect 43572 226 43576 282
rect 43512 222 43576 226
rect 43592 282 43656 286
rect 43592 226 43596 282
rect 43596 226 43652 282
rect 43652 226 43656 282
rect 43592 222 43656 226
rect 43672 282 43736 286
rect 43672 226 43676 282
rect 43676 226 43732 282
rect 43732 226 43736 282
rect 43672 222 43736 226
rect 43752 282 43816 286
rect 43752 226 43756 282
rect 43756 226 43812 282
rect 43812 226 43816 282
rect 43752 222 43816 226
rect 43832 282 43896 286
rect 43832 226 43836 282
rect 43836 226 43892 282
rect 43892 226 43896 282
rect 43832 222 43896 226
rect 43912 282 43976 286
rect 43912 226 43916 282
rect 43916 226 43972 282
rect 43972 226 43976 282
rect 43912 222 43976 226
rect 43992 282 44056 286
rect 43992 226 43996 282
rect 43996 226 44052 282
rect 44052 226 44056 282
rect 43992 222 44056 226
rect 44072 282 44136 286
rect 44072 226 44076 282
rect 44076 226 44132 282
rect 44132 226 44136 282
rect 44072 222 44136 226
rect 44152 282 44216 286
rect 44152 226 44156 282
rect 44156 226 44212 282
rect 44212 226 44216 282
rect 44152 222 44216 226
rect 44232 282 44296 286
rect 44232 226 44236 282
rect 44236 226 44292 282
rect 44292 226 44296 282
rect 44232 222 44296 226
rect 44312 282 44376 286
rect 44312 226 44316 282
rect 44316 226 44372 282
rect 44372 226 44376 282
rect 44312 222 44376 226
rect 44392 282 44456 286
rect 44392 226 44396 282
rect 44396 226 44452 282
rect 44452 226 44456 282
rect 44392 222 44456 226
rect 44472 282 44536 286
rect 44472 226 44476 282
rect 44476 226 44532 282
rect 44532 226 44536 282
rect 44472 222 44536 226
rect 44552 282 44616 286
rect 44552 226 44556 282
rect 44556 226 44612 282
rect 44612 226 44616 282
rect 44552 222 44616 226
rect 44632 282 44696 286
rect 44632 226 44636 282
rect 44636 226 44692 282
rect 44692 226 44696 282
rect 44632 222 44696 226
rect 44712 282 44776 286
rect 44712 226 44716 282
rect 44716 226 44772 282
rect 44772 226 44776 282
rect 44712 222 44776 226
rect 44792 282 44856 286
rect 44792 226 44796 282
rect 44796 226 44852 282
rect 44852 226 44856 282
rect 44792 222 44856 226
rect 44872 282 44936 286
rect 44872 226 44876 282
rect 44876 226 44932 282
rect 44932 226 44936 282
rect 44872 222 44936 226
rect 44952 282 45016 286
rect 44952 226 44956 282
rect 44956 226 45012 282
rect 45012 226 45016 282
rect 44952 222 45016 226
rect 45032 282 45096 286
rect 45032 226 45036 282
rect 45036 226 45092 282
rect 45092 226 45096 282
rect 45032 222 45096 226
rect 45112 282 45176 286
rect 45112 226 45116 282
rect 45116 226 45172 282
rect 45172 226 45176 282
rect 45112 222 45176 226
rect 45192 282 45256 286
rect 45192 226 45196 282
rect 45196 226 45252 282
rect 45252 226 45256 282
rect 45192 222 45256 226
rect 45272 282 45336 286
rect 45272 226 45276 282
rect 45276 226 45332 282
rect 45332 226 45336 282
rect 45272 222 45336 226
rect 45352 282 45416 286
rect 45352 226 45356 282
rect 45356 226 45412 282
rect 45412 226 45416 282
rect 45352 222 45416 226
rect 45432 282 45496 286
rect 45432 226 45436 282
rect 45436 226 45492 282
rect 45492 226 45496 282
rect 45432 222 45496 226
rect 45512 282 45576 286
rect 45512 226 45516 282
rect 45516 226 45572 282
rect 45572 226 45576 282
rect 45512 222 45576 226
rect 45592 282 45656 286
rect 45592 226 45596 282
rect 45596 226 45652 282
rect 45652 226 45656 282
rect 45592 222 45656 226
rect 45672 282 45736 286
rect 45672 226 45676 282
rect 45676 226 45732 282
rect 45732 226 45736 282
rect 45672 222 45736 226
rect 45752 282 45816 286
rect 45752 226 45756 282
rect 45756 226 45812 282
rect 45812 226 45816 282
rect 45752 222 45816 226
rect 45832 282 45896 286
rect 45832 226 45836 282
rect 45836 226 45892 282
rect 45892 226 45896 282
rect 45832 222 45896 226
rect 35027 -1059 35091 -1055
rect 35027 -1115 35031 -1059
rect 35031 -1115 35087 -1059
rect 35087 -1115 35091 -1059
rect 35027 -1119 35091 -1115
rect 36987 -695 37051 -691
rect 36987 -751 36991 -695
rect 36991 -751 37047 -695
rect 37047 -751 37051 -695
rect 36987 -755 37051 -751
rect 38571 -734 38635 -730
rect 38571 -790 38575 -734
rect 38575 -790 38631 -734
rect 38631 -790 38635 -734
rect 38571 -794 38635 -790
rect 38571 -814 38635 -810
rect 38571 -870 38575 -814
rect 38575 -870 38631 -814
rect 38631 -870 38635 -814
rect 38571 -874 38635 -870
rect 40100 -737 40164 -733
rect 40100 -793 40104 -737
rect 40104 -793 40160 -737
rect 40160 -793 40164 -737
rect 40100 -797 40164 -793
rect 40100 -817 40164 -813
rect 40100 -873 40104 -817
rect 40104 -873 40160 -817
rect 40160 -873 40164 -817
rect 40100 -877 40164 -873
rect 36987 -1843 37051 -1779
rect 38570 -2087 38634 -2083
rect 38570 -2143 38574 -2087
rect 38574 -2143 38630 -2087
rect 38630 -2143 38634 -2087
rect 38570 -2147 38634 -2143
rect 38570 -2167 38634 -2163
rect 38570 -2223 38574 -2167
rect 38574 -2223 38630 -2167
rect 38630 -2223 38634 -2167
rect 38570 -2227 38634 -2223
rect 35035 -2452 35099 -2448
rect 35035 -2508 35039 -2452
rect 35039 -2508 35095 -2452
rect 35095 -2508 35099 -2452
rect 35035 -2512 35099 -2508
rect 36988 -2871 37052 -2867
rect 36988 -2927 36992 -2871
rect 36992 -2927 37048 -2871
rect 37048 -2927 37052 -2871
rect 36988 -2931 37052 -2927
rect 40100 -2109 40164 -2105
rect 40100 -2165 40104 -2109
rect 40104 -2165 40160 -2109
rect 40160 -2165 40164 -2109
rect 40100 -2169 40164 -2165
rect 40100 -2189 40164 -2185
rect 40100 -2245 40104 -2189
rect 40104 -2245 40160 -2189
rect 40160 -2245 40164 -2189
rect 40100 -2249 40164 -2245
rect 40838 -2905 41222 -2681
rect 42588 -2724 42652 -2720
rect 42588 -2780 42592 -2724
rect 42592 -2780 42648 -2724
rect 42648 -2780 42652 -2724
rect 42588 -2784 42652 -2780
rect 42668 -2724 42732 -2720
rect 42668 -2780 42672 -2724
rect 42672 -2780 42728 -2724
rect 42728 -2780 42732 -2724
rect 42668 -2784 42732 -2780
rect 42748 -2724 42812 -2720
rect 42748 -2780 42752 -2724
rect 42752 -2780 42808 -2724
rect 42808 -2780 42812 -2724
rect 42748 -2784 42812 -2780
rect 42828 -2724 42892 -2720
rect 42828 -2780 42832 -2724
rect 42832 -2780 42888 -2724
rect 42888 -2780 42892 -2724
rect 42828 -2784 42892 -2780
rect 42908 -2724 42972 -2720
rect 42908 -2780 42912 -2724
rect 42912 -2780 42968 -2724
rect 42968 -2780 42972 -2724
rect 42908 -2784 42972 -2780
rect 42988 -2724 43052 -2720
rect 42988 -2780 42992 -2724
rect 42992 -2780 43048 -2724
rect 43048 -2780 43052 -2724
rect 42988 -2784 43052 -2780
rect 43068 -2724 43132 -2720
rect 43068 -2780 43072 -2724
rect 43072 -2780 43128 -2724
rect 43128 -2780 43132 -2724
rect 43068 -2784 43132 -2780
rect 43148 -2724 43212 -2720
rect 43148 -2780 43152 -2724
rect 43152 -2780 43208 -2724
rect 43208 -2780 43212 -2724
rect 43148 -2784 43212 -2780
rect 43228 -2724 43292 -2720
rect 43228 -2780 43232 -2724
rect 43232 -2780 43288 -2724
rect 43288 -2780 43292 -2724
rect 43228 -2784 43292 -2780
rect 43308 -2724 43372 -2720
rect 43308 -2780 43312 -2724
rect 43312 -2780 43368 -2724
rect 43368 -2780 43372 -2724
rect 43308 -2784 43372 -2780
rect 43388 -2724 43452 -2720
rect 43388 -2780 43392 -2724
rect 43392 -2780 43448 -2724
rect 43448 -2780 43452 -2724
rect 43388 -2784 43452 -2780
rect 43468 -2724 43532 -2720
rect 43468 -2780 43472 -2724
rect 43472 -2780 43528 -2724
rect 43528 -2780 43532 -2724
rect 43468 -2784 43532 -2780
rect 43548 -2724 43612 -2720
rect 43548 -2780 43552 -2724
rect 43552 -2780 43608 -2724
rect 43608 -2780 43612 -2724
rect 43548 -2784 43612 -2780
rect 43628 -2724 43692 -2720
rect 43628 -2780 43632 -2724
rect 43632 -2780 43688 -2724
rect 43688 -2780 43692 -2724
rect 43628 -2784 43692 -2780
rect 43708 -2724 43772 -2720
rect 43708 -2780 43712 -2724
rect 43712 -2780 43768 -2724
rect 43768 -2780 43772 -2724
rect 43708 -2784 43772 -2780
rect 43788 -2724 43852 -2720
rect 43788 -2780 43792 -2724
rect 43792 -2780 43848 -2724
rect 43848 -2780 43852 -2724
rect 43788 -2784 43852 -2780
rect 43868 -2724 43932 -2720
rect 43868 -2780 43872 -2724
rect 43872 -2780 43928 -2724
rect 43928 -2780 43932 -2724
rect 43868 -2784 43932 -2780
rect 43948 -2724 44012 -2720
rect 43948 -2780 43952 -2724
rect 43952 -2780 44008 -2724
rect 44008 -2780 44012 -2724
rect 43948 -2784 44012 -2780
rect 44028 -2724 44092 -2720
rect 44028 -2780 44032 -2724
rect 44032 -2780 44088 -2724
rect 44088 -2780 44092 -2724
rect 44028 -2784 44092 -2780
rect 44108 -2724 44172 -2720
rect 44108 -2780 44112 -2724
rect 44112 -2780 44168 -2724
rect 44168 -2780 44172 -2724
rect 44108 -2784 44172 -2780
rect 44188 -2724 44252 -2720
rect 44188 -2780 44192 -2724
rect 44192 -2780 44248 -2724
rect 44248 -2780 44252 -2724
rect 44188 -2784 44252 -2780
rect 44268 -2724 44332 -2720
rect 44268 -2780 44272 -2724
rect 44272 -2780 44328 -2724
rect 44328 -2780 44332 -2724
rect 44268 -2784 44332 -2780
rect 44348 -2724 44412 -2720
rect 44348 -2780 44352 -2724
rect 44352 -2780 44408 -2724
rect 44408 -2780 44412 -2724
rect 44348 -2784 44412 -2780
rect 44428 -2724 44492 -2720
rect 44428 -2780 44432 -2724
rect 44432 -2780 44488 -2724
rect 44488 -2780 44492 -2724
rect 44428 -2784 44492 -2780
rect 44508 -2724 44572 -2720
rect 44508 -2780 44512 -2724
rect 44512 -2780 44568 -2724
rect 44568 -2780 44572 -2724
rect 44508 -2784 44572 -2780
rect 44588 -2724 44652 -2720
rect 44588 -2780 44592 -2724
rect 44592 -2780 44648 -2724
rect 44648 -2780 44652 -2724
rect 44588 -2784 44652 -2780
rect 44668 -2724 44732 -2720
rect 44668 -2780 44672 -2724
rect 44672 -2780 44728 -2724
rect 44728 -2780 44732 -2724
rect 44668 -2784 44732 -2780
rect 44748 -2724 44812 -2720
rect 44748 -2780 44752 -2724
rect 44752 -2780 44808 -2724
rect 44808 -2780 44812 -2724
rect 44748 -2784 44812 -2780
rect 44828 -2724 44892 -2720
rect 44828 -2780 44832 -2724
rect 44832 -2780 44888 -2724
rect 44888 -2780 44892 -2724
rect 44828 -2784 44892 -2780
rect 44908 -2724 44972 -2720
rect 44908 -2780 44912 -2724
rect 44912 -2780 44968 -2724
rect 44968 -2780 44972 -2724
rect 44908 -2784 44972 -2780
rect 44988 -2724 45052 -2720
rect 44988 -2780 44992 -2724
rect 44992 -2780 45048 -2724
rect 45048 -2780 45052 -2724
rect 44988 -2784 45052 -2780
rect 45068 -2724 45132 -2720
rect 45068 -2780 45072 -2724
rect 45072 -2780 45128 -2724
rect 45128 -2780 45132 -2724
rect 45068 -2784 45132 -2780
rect 45148 -2724 45212 -2720
rect 45148 -2780 45152 -2724
rect 45152 -2780 45208 -2724
rect 45208 -2780 45212 -2724
rect 45148 -2784 45212 -2780
rect 45228 -2724 45292 -2720
rect 45228 -2780 45232 -2724
rect 45232 -2780 45288 -2724
rect 45288 -2780 45292 -2724
rect 45228 -2784 45292 -2780
rect 45308 -2724 45372 -2720
rect 45308 -2780 45312 -2724
rect 45312 -2780 45368 -2724
rect 45368 -2780 45372 -2724
rect 45308 -2784 45372 -2780
rect 45388 -2724 45452 -2720
rect 45388 -2780 45392 -2724
rect 45392 -2780 45448 -2724
rect 45448 -2780 45452 -2724
rect 45388 -2784 45452 -2780
rect 45468 -2724 45532 -2720
rect 45468 -2780 45472 -2724
rect 45472 -2780 45528 -2724
rect 45528 -2780 45532 -2724
rect 45468 -2784 45532 -2780
rect 45548 -2724 45612 -2720
rect 45548 -2780 45552 -2724
rect 45552 -2780 45608 -2724
rect 45608 -2780 45612 -2724
rect 45548 -2784 45612 -2780
rect 45628 -2724 45692 -2720
rect 45628 -2780 45632 -2724
rect 45632 -2780 45688 -2724
rect 45688 -2780 45692 -2724
rect 45628 -2784 45692 -2780
rect 45708 -2724 45772 -2720
rect 45708 -2780 45712 -2724
rect 45712 -2780 45768 -2724
rect 45768 -2780 45772 -2724
rect 45708 -2784 45772 -2780
rect 45788 -2724 45852 -2720
rect 45788 -2780 45792 -2724
rect 45792 -2780 45848 -2724
rect 45848 -2780 45852 -2724
rect 45788 -2784 45852 -2780
rect 45868 -2724 45932 -2720
rect 45868 -2780 45872 -2724
rect 45872 -2780 45928 -2724
rect 45928 -2780 45932 -2724
rect 45868 -2784 45932 -2780
rect 21202 -3573 21266 -3509
rect 35031 -3822 35095 -3818
rect 35031 -3878 35035 -3822
rect 35035 -3878 35091 -3822
rect 35091 -3878 35095 -3822
rect 38573 -3487 38637 -3483
rect 38573 -3543 38577 -3487
rect 38577 -3543 38633 -3487
rect 38633 -3543 38637 -3487
rect 38573 -3547 38637 -3543
rect 38573 -3567 38637 -3563
rect 38573 -3623 38577 -3567
rect 38577 -3623 38633 -3567
rect 38633 -3623 38637 -3567
rect 38573 -3627 38637 -3623
rect 40097 -3493 40161 -3489
rect 40097 -3549 40101 -3493
rect 40101 -3549 40157 -3493
rect 40157 -3549 40161 -3493
rect 40097 -3553 40161 -3549
rect 40097 -3573 40161 -3569
rect 40097 -3629 40101 -3573
rect 40101 -3629 40157 -3573
rect 40157 -3629 40161 -3573
rect 40097 -3633 40161 -3629
rect 35031 -3882 35095 -3878
rect 21202 -4045 21266 -3981
rect 21202 -4580 21266 -4516
rect 21202 -5043 21266 -4979
rect -3581 -6848 -3517 -6844
rect -3581 -6904 -3577 -6848
rect -3577 -6904 -3521 -6848
rect -3521 -6904 -3517 -6848
rect -3581 -6908 -3517 -6904
rect -3581 -6928 -3517 -6924
rect -3581 -6984 -3577 -6928
rect -3577 -6984 -3521 -6928
rect -3521 -6984 -3517 -6928
rect -3581 -6988 -3517 -6984
rect -3581 -7008 -3517 -7004
rect -3581 -7064 -3577 -7008
rect -3577 -7064 -3521 -7008
rect -3521 -7064 -3517 -7008
rect -3581 -7068 -3517 -7064
rect -3581 -7088 -3517 -7084
rect -3581 -7144 -3577 -7088
rect -3577 -7144 -3521 -7088
rect -3521 -7144 -3517 -7088
rect -3581 -7148 -3517 -7144
rect -3581 -7168 -3517 -7164
rect -3581 -7224 -3577 -7168
rect -3577 -7224 -3521 -7168
rect -3521 -7224 -3517 -7168
rect -3581 -7228 -3517 -7224
rect -3581 -7248 -3517 -7244
rect -3581 -7304 -3577 -7248
rect -3577 -7304 -3521 -7248
rect -3521 -7304 -3517 -7248
rect -3581 -7308 -3517 -7304
rect -3581 -7328 -3517 -7324
rect -3581 -7384 -3577 -7328
rect -3577 -7384 -3521 -7328
rect -3521 -7384 -3517 -7328
rect -3581 -7388 -3517 -7384
rect -3581 -7408 -3517 -7404
rect -3581 -7464 -3577 -7408
rect -3577 -7464 -3521 -7408
rect -3521 -7464 -3517 -7408
rect -3581 -7468 -3517 -7464
rect -3581 -7488 -3517 -7484
rect -3581 -7544 -3577 -7488
rect -3577 -7544 -3521 -7488
rect -3521 -7544 -3517 -7488
rect -3581 -7548 -3517 -7544
rect -3581 -7568 -3517 -7564
rect -3581 -7624 -3577 -7568
rect -3577 -7624 -3521 -7568
rect -3521 -7624 -3517 -7568
rect -3581 -7628 -3517 -7624
rect -3581 -7648 -3517 -7644
rect -3581 -7704 -3577 -7648
rect -3577 -7704 -3521 -7648
rect -3521 -7704 -3517 -7648
rect -3581 -7708 -3517 -7704
rect -3581 -7728 -3517 -7724
rect -3581 -7784 -3577 -7728
rect -3577 -7784 -3521 -7728
rect -3521 -7784 -3517 -7728
rect -3581 -7788 -3517 -7784
rect -3581 -7808 -3517 -7804
rect -3581 -7864 -3577 -7808
rect -3577 -7864 -3521 -7808
rect -3521 -7864 -3517 -7808
rect -3581 -7868 -3517 -7864
rect -3581 -7888 -3517 -7884
rect -3581 -7944 -3577 -7888
rect -3577 -7944 -3521 -7888
rect -3521 -7944 -3517 -7888
rect -3581 -7948 -3517 -7944
rect -3581 -7968 -3517 -7964
rect -3581 -8024 -3577 -7968
rect -3577 -8024 -3521 -7968
rect -3521 -8024 -3517 -7968
rect -3581 -8028 -3517 -8024
rect -3581 -8048 -3517 -8044
rect -3581 -8104 -3577 -8048
rect -3577 -8104 -3521 -8048
rect -3521 -8104 -3517 -8048
rect -3581 -8108 -3517 -8104
rect -3581 -8128 -3517 -8124
rect -3581 -8184 -3577 -8128
rect -3577 -8184 -3521 -8128
rect -3521 -8184 -3517 -8128
rect -3581 -8188 -3517 -8184
rect -3581 -8208 -3517 -8204
rect -3581 -8264 -3577 -8208
rect -3577 -8264 -3521 -8208
rect -3521 -8264 -3517 -8208
rect -3581 -8268 -3517 -8264
rect -3581 -8288 -3517 -8284
rect -3581 -8344 -3577 -8288
rect -3577 -8344 -3521 -8288
rect -3521 -8344 -3517 -8288
rect -3581 -8348 -3517 -8344
rect -3581 -8368 -3517 -8364
rect -3581 -8424 -3577 -8368
rect -3577 -8424 -3521 -8368
rect -3521 -8424 -3517 -8368
rect -3581 -8428 -3517 -8424
rect -3581 -8448 -3517 -8444
rect -3581 -8504 -3577 -8448
rect -3577 -8504 -3521 -8448
rect -3521 -8504 -3517 -8448
rect -3581 -8508 -3517 -8504
rect -3581 -8528 -3517 -8524
rect -3581 -8584 -3577 -8528
rect -3577 -8584 -3521 -8528
rect -3521 -8584 -3517 -8528
rect -3581 -8588 -3517 -8584
rect -3581 -8608 -3517 -8604
rect -3581 -8664 -3577 -8608
rect -3577 -8664 -3521 -8608
rect -3521 -8664 -3517 -8608
rect -3581 -8668 -3517 -8664
rect -3581 -8688 -3517 -8684
rect -3581 -8744 -3577 -8688
rect -3577 -8744 -3521 -8688
rect -3521 -8744 -3517 -8688
rect -3581 -8748 -3517 -8744
rect -3581 -8768 -3517 -8764
rect -3581 -8824 -3577 -8768
rect -3577 -8824 -3521 -8768
rect -3521 -8824 -3517 -8768
rect -3581 -8828 -3517 -8824
rect -3581 -8848 -3517 -8844
rect -3581 -8904 -3577 -8848
rect -3577 -8904 -3521 -8848
rect -3521 -8904 -3517 -8848
rect -3581 -8908 -3517 -8904
rect -3581 -8928 -3517 -8924
rect -3581 -8984 -3577 -8928
rect -3577 -8984 -3521 -8928
rect -3521 -8984 -3517 -8928
rect -3581 -8988 -3517 -8984
rect -3581 -9008 -3517 -9004
rect -3581 -9064 -3577 -9008
rect -3577 -9064 -3521 -9008
rect -3521 -9064 -3517 -9008
rect -3581 -9068 -3517 -9064
rect -3581 -9088 -3517 -9084
rect -3581 -9144 -3577 -9088
rect -3577 -9144 -3521 -9088
rect -3521 -9144 -3517 -9088
rect -3581 -9148 -3517 -9144
rect -3581 -9168 -3517 -9164
rect -3581 -9224 -3577 -9168
rect -3577 -9224 -3521 -9168
rect -3521 -9224 -3517 -9168
rect -3581 -9228 -3517 -9224
rect -3581 -9248 -3517 -9244
rect -3581 -9304 -3577 -9248
rect -3577 -9304 -3521 -9248
rect -3521 -9304 -3517 -9248
rect -3581 -9308 -3517 -9304
rect -3581 -9328 -3517 -9324
rect -3581 -9384 -3577 -9328
rect -3577 -9384 -3521 -9328
rect -3521 -9384 -3517 -9328
rect -3581 -9388 -3517 -9384
rect -3581 -9408 -3517 -9404
rect -3581 -9464 -3577 -9408
rect -3577 -9464 -3521 -9408
rect -3521 -9464 -3517 -9408
rect -3581 -9468 -3517 -9464
rect -3581 -9488 -3517 -9484
rect -3581 -9544 -3577 -9488
rect -3577 -9544 -3521 -9488
rect -3521 -9544 -3517 -9488
rect -3581 -9548 -3517 -9544
rect -3581 -9568 -3517 -9564
rect -3581 -9624 -3577 -9568
rect -3577 -9624 -3521 -9568
rect -3521 -9624 -3517 -9568
rect -3581 -9628 -3517 -9624
rect -3581 -9648 -3517 -9644
rect -3581 -9704 -3577 -9648
rect -3577 -9704 -3521 -9648
rect -3521 -9704 -3517 -9648
rect -3581 -9708 -3517 -9704
rect -3581 -9728 -3517 -9724
rect -3581 -9784 -3577 -9728
rect -3577 -9784 -3521 -9728
rect -3521 -9784 -3517 -9728
rect -3581 -9788 -3517 -9784
rect -3581 -9808 -3517 -9804
rect -3581 -9864 -3577 -9808
rect -3577 -9864 -3521 -9808
rect -3521 -9864 -3517 -9808
rect -3581 -9868 -3517 -9864
rect -3581 -9888 -3517 -9884
rect -3581 -9944 -3577 -9888
rect -3577 -9944 -3521 -9888
rect -3521 -9944 -3517 -9888
rect -3581 -9948 -3517 -9944
rect -3581 -9968 -3517 -9964
rect -3581 -10024 -3577 -9968
rect -3577 -10024 -3521 -9968
rect -3521 -10024 -3517 -9968
rect -3581 -10028 -3517 -10024
rect -3581 -10048 -3517 -10044
rect -3581 -10104 -3577 -10048
rect -3577 -10104 -3521 -10048
rect -3521 -10104 -3517 -10048
rect -3581 -10108 -3517 -10104
rect -575 -6855 -511 -6851
rect -575 -6911 -571 -6855
rect -571 -6911 -515 -6855
rect -515 -6911 -511 -6855
rect -575 -6915 -511 -6911
rect -575 -6935 -511 -6931
rect -575 -6991 -571 -6935
rect -571 -6991 -515 -6935
rect -515 -6991 -511 -6935
rect -575 -6995 -511 -6991
rect -575 -7015 -511 -7011
rect -575 -7071 -571 -7015
rect -571 -7071 -515 -7015
rect -515 -7071 -511 -7015
rect -575 -7075 -511 -7071
rect -575 -7095 -511 -7091
rect -575 -7151 -571 -7095
rect -571 -7151 -515 -7095
rect -515 -7151 -511 -7095
rect -575 -7155 -511 -7151
rect -575 -7175 -511 -7171
rect -575 -7231 -571 -7175
rect -571 -7231 -515 -7175
rect -515 -7231 -511 -7175
rect -575 -7235 -511 -7231
rect -575 -7255 -511 -7251
rect -575 -7311 -571 -7255
rect -571 -7311 -515 -7255
rect -515 -7311 -511 -7255
rect -575 -7315 -511 -7311
rect -575 -7335 -511 -7331
rect -575 -7391 -571 -7335
rect -571 -7391 -515 -7335
rect -515 -7391 -511 -7335
rect -575 -7395 -511 -7391
rect -575 -7415 -511 -7411
rect -575 -7471 -571 -7415
rect -571 -7471 -515 -7415
rect -515 -7471 -511 -7415
rect -575 -7475 -511 -7471
rect -575 -7495 -511 -7491
rect -575 -7551 -571 -7495
rect -571 -7551 -515 -7495
rect -515 -7551 -511 -7495
rect -575 -7555 -511 -7551
rect -575 -7575 -511 -7571
rect -575 -7631 -571 -7575
rect -571 -7631 -515 -7575
rect -515 -7631 -511 -7575
rect -575 -7635 -511 -7631
rect -575 -7655 -511 -7651
rect -575 -7711 -571 -7655
rect -571 -7711 -515 -7655
rect -515 -7711 -511 -7655
rect -575 -7715 -511 -7711
rect -575 -7735 -511 -7731
rect -575 -7791 -571 -7735
rect -571 -7791 -515 -7735
rect -515 -7791 -511 -7735
rect -575 -7795 -511 -7791
rect -575 -7815 -511 -7811
rect -575 -7871 -571 -7815
rect -571 -7871 -515 -7815
rect -515 -7871 -511 -7815
rect -575 -7875 -511 -7871
rect -575 -7895 -511 -7891
rect -575 -7951 -571 -7895
rect -571 -7951 -515 -7895
rect -515 -7951 -511 -7895
rect -575 -7955 -511 -7951
rect -575 -7975 -511 -7971
rect -575 -8031 -571 -7975
rect -571 -8031 -515 -7975
rect -515 -8031 -511 -7975
rect -575 -8035 -511 -8031
rect -575 -8055 -511 -8051
rect -575 -8111 -571 -8055
rect -571 -8111 -515 -8055
rect -515 -8111 -511 -8055
rect -575 -8115 -511 -8111
rect -575 -8135 -511 -8131
rect -575 -8191 -571 -8135
rect -571 -8191 -515 -8135
rect -515 -8191 -511 -8135
rect -575 -8195 -511 -8191
rect -575 -8215 -511 -8211
rect -575 -8271 -571 -8215
rect -571 -8271 -515 -8215
rect -515 -8271 -511 -8215
rect -575 -8275 -511 -8271
rect -575 -8295 -511 -8291
rect -575 -8351 -571 -8295
rect -571 -8351 -515 -8295
rect -515 -8351 -511 -8295
rect -575 -8355 -511 -8351
rect -575 -8375 -511 -8371
rect -575 -8431 -571 -8375
rect -571 -8431 -515 -8375
rect -515 -8431 -511 -8375
rect -575 -8435 -511 -8431
rect -575 -8455 -511 -8451
rect -575 -8511 -571 -8455
rect -571 -8511 -515 -8455
rect -515 -8511 -511 -8455
rect -575 -8515 -511 -8511
rect -575 -8535 -511 -8531
rect -575 -8591 -571 -8535
rect -571 -8591 -515 -8535
rect -515 -8591 -511 -8535
rect -575 -8595 -511 -8591
rect -575 -8615 -511 -8611
rect -575 -8671 -571 -8615
rect -571 -8671 -515 -8615
rect -515 -8671 -511 -8615
rect -575 -8675 -511 -8671
rect -575 -8695 -511 -8691
rect -575 -8751 -571 -8695
rect -571 -8751 -515 -8695
rect -515 -8751 -511 -8695
rect -575 -8755 -511 -8751
rect -575 -8775 -511 -8771
rect -575 -8831 -571 -8775
rect -571 -8831 -515 -8775
rect -515 -8831 -511 -8775
rect -575 -8835 -511 -8831
rect -575 -8855 -511 -8851
rect -575 -8911 -571 -8855
rect -571 -8911 -515 -8855
rect -515 -8911 -511 -8855
rect -575 -8915 -511 -8911
rect -575 -8935 -511 -8931
rect -575 -8991 -571 -8935
rect -571 -8991 -515 -8935
rect -515 -8991 -511 -8935
rect -575 -8995 -511 -8991
rect -575 -9015 -511 -9011
rect -575 -9071 -571 -9015
rect -571 -9071 -515 -9015
rect -515 -9071 -511 -9015
rect -575 -9075 -511 -9071
rect -575 -9095 -511 -9091
rect -575 -9151 -571 -9095
rect -571 -9151 -515 -9095
rect -515 -9151 -511 -9095
rect -575 -9155 -511 -9151
rect -575 -9175 -511 -9171
rect -575 -9231 -571 -9175
rect -571 -9231 -515 -9175
rect -515 -9231 -511 -9175
rect -575 -9235 -511 -9231
rect -575 -9255 -511 -9251
rect -575 -9311 -571 -9255
rect -571 -9311 -515 -9255
rect -515 -9311 -511 -9255
rect -575 -9315 -511 -9311
rect -575 -9335 -511 -9331
rect -575 -9391 -571 -9335
rect -571 -9391 -515 -9335
rect -515 -9391 -511 -9335
rect -575 -9395 -511 -9391
rect -575 -9415 -511 -9411
rect -575 -9471 -571 -9415
rect -571 -9471 -515 -9415
rect -515 -9471 -511 -9415
rect -575 -9475 -511 -9471
rect -575 -9495 -511 -9491
rect -575 -9551 -571 -9495
rect -571 -9551 -515 -9495
rect -515 -9551 -511 -9495
rect -575 -9555 -511 -9551
rect -575 -9575 -511 -9571
rect -575 -9631 -571 -9575
rect -571 -9631 -515 -9575
rect -515 -9631 -511 -9575
rect -575 -9635 -511 -9631
rect -575 -9655 -511 -9651
rect -575 -9711 -571 -9655
rect -571 -9711 -515 -9655
rect -515 -9711 -511 -9655
rect -575 -9715 -511 -9711
rect -575 -9735 -511 -9731
rect -575 -9791 -571 -9735
rect -571 -9791 -515 -9735
rect -515 -9791 -511 -9735
rect -575 -9795 -511 -9791
rect -575 -9815 -511 -9811
rect -575 -9871 -571 -9815
rect -571 -9871 -515 -9815
rect -515 -9871 -511 -9815
rect -575 -9875 -511 -9871
rect -575 -9895 -511 -9891
rect -575 -9951 -571 -9895
rect -571 -9951 -515 -9895
rect -515 -9951 -511 -9895
rect -575 -9955 -511 -9951
rect -575 -9975 -511 -9971
rect -575 -10031 -571 -9975
rect -571 -10031 -515 -9975
rect -515 -10031 -511 -9975
rect -575 -10035 -511 -10031
rect -575 -10055 -511 -10051
rect -575 -10111 -571 -10055
rect -571 -10111 -515 -10055
rect -515 -10111 -511 -10055
rect -575 -10115 -511 -10111
<< metal4 >>
rect -57093 88360 62907 88442
rect -57093 86524 -55011 88360
rect -53175 86524 -43253 88360
rect -42697 86524 -35253 88360
rect -34697 86524 -27253 88360
rect -26697 86524 -19253 88360
rect -18697 86524 -11253 88360
rect -10697 86524 -3253 88360
rect -2697 86524 4747 88360
rect 5303 86524 12747 88360
rect 13303 86524 20747 88360
rect 21303 86524 28747 88360
rect 29303 86524 36747 88360
rect 37303 86524 44747 88360
rect 45303 86524 54989 88360
rect 56825 86524 62907 88360
rect -57093 86442 62907 86524
rect -57093 84360 62907 84442
rect -57093 82524 -51011 84360
rect -49175 82524 -39253 84360
rect -38697 82524 -31253 84360
rect -30697 82524 -23253 84360
rect -22697 82524 -15253 84360
rect -14697 82524 -7253 84360
rect -6697 82524 747 84360
rect 1303 82524 8747 84360
rect 9303 82524 16747 84360
rect 17303 82524 24747 84360
rect 25303 82524 32747 84360
rect 33303 82524 40747 84360
rect 41303 82524 48747 84360
rect 49303 82524 58989 84360
rect 60825 82524 62907 84360
rect -57093 82442 62907 82524
rect -16930 76692 -16690 76806
rect -16930 76628 -16831 76692
rect -16767 76628 -16690 76692
rect -16930 76612 -16690 76628
rect -16930 76548 -16831 76612
rect -16767 76548 -16690 76612
rect -16930 76532 -16690 76548
rect -16930 76468 -16831 76532
rect -16767 76468 -16690 76532
rect -16930 76452 -16690 76468
rect -16930 76388 -16831 76452
rect -16767 76388 -16690 76452
rect -16930 76372 -16690 76388
rect -16930 76308 -16831 76372
rect -16767 76308 -16690 76372
rect -16930 76292 -16690 76308
rect -16930 76228 -16831 76292
rect -16767 76228 -16690 76292
rect -16930 76212 -16690 76228
rect -16930 76148 -16831 76212
rect -16767 76148 -16690 76212
rect -16930 76132 -16690 76148
rect -16930 76068 -16831 76132
rect -16767 76068 -16690 76132
rect -16930 76052 -16690 76068
rect -16930 75988 -16831 76052
rect -16767 75988 -16690 76052
rect -16930 75972 -16690 75988
rect -16930 75908 -16831 75972
rect -16767 75908 -16690 75972
rect -16930 75892 -16690 75908
rect -16930 75828 -16831 75892
rect -16767 75828 -16690 75892
rect -16930 75812 -16690 75828
rect -16930 75748 -16831 75812
rect -16767 75748 -16690 75812
rect -16930 75732 -16690 75748
rect -16930 75668 -16831 75732
rect -16767 75668 -16690 75732
rect -16930 75652 -16690 75668
rect -16930 75588 -16831 75652
rect -16767 75588 -16690 75652
rect -16930 75572 -16690 75588
rect -16930 75508 -16831 75572
rect -16767 75508 -16690 75572
rect -16930 75492 -16690 75508
rect -16930 75428 -16831 75492
rect -16767 75428 -16690 75492
rect -16930 75412 -16690 75428
rect -16930 75348 -16831 75412
rect -16767 75348 -16690 75412
rect -16930 75332 -16690 75348
rect -16930 75268 -16831 75332
rect -16767 75268 -16690 75332
rect -16930 75252 -16690 75268
rect -13914 76698 -13674 76891
rect -13914 76634 -13830 76698
rect -13766 76634 -13674 76698
rect -13914 76618 -13674 76634
rect -13914 76554 -13830 76618
rect -13766 76554 -13674 76618
rect -13914 76538 -13674 76554
rect -13914 76474 -13830 76538
rect -13766 76474 -13674 76538
rect -13914 76458 -13674 76474
rect -13914 76394 -13830 76458
rect -13766 76394 -13674 76458
rect -13914 76378 -13674 76394
rect -13914 76314 -13830 76378
rect -13766 76314 -13674 76378
rect -13914 76298 -13674 76314
rect -13914 76234 -13830 76298
rect -13766 76234 -13674 76298
rect -13914 76218 -13674 76234
rect -13914 76154 -13830 76218
rect -13766 76154 -13674 76218
rect -13914 76138 -13674 76154
rect -13914 76074 -13830 76138
rect -13766 76074 -13674 76138
rect -13914 76058 -13674 76074
rect -13914 75994 -13830 76058
rect -13766 75994 -13674 76058
rect -13914 75978 -13674 75994
rect -13914 75914 -13830 75978
rect -13766 75914 -13674 75978
rect -13914 75898 -13674 75914
rect -13914 75834 -13830 75898
rect -13766 75834 -13674 75898
rect -13914 75818 -13674 75834
rect -13914 75754 -13830 75818
rect -13766 75754 -13674 75818
rect -13914 75738 -13674 75754
rect -13914 75674 -13830 75738
rect -13766 75674 -13674 75738
rect -13914 75658 -13674 75674
rect -13914 75594 -13830 75658
rect -13766 75594 -13674 75658
rect -13914 75578 -13674 75594
rect -13914 75514 -13830 75578
rect -13766 75514 -13674 75578
rect -13914 75498 -13674 75514
rect -13914 75434 -13830 75498
rect -13766 75434 -13674 75498
rect -13914 75418 -13674 75434
rect -13914 75354 -13830 75418
rect -13766 75354 -13674 75418
rect -13914 75338 -13674 75354
rect -13914 75274 -13830 75338
rect -13766 75274 -13674 75338
rect -13914 75258 -13674 75274
rect -13914 75253 -13830 75258
rect -16930 75188 -16831 75252
rect -16767 75188 -16690 75252
rect -16930 75172 -16690 75188
rect -16930 75108 -16831 75172
rect -16767 75108 -16690 75172
rect -16930 75092 -16690 75108
rect -16930 75068 -16831 75092
rect -19241 75066 -16831 75068
rect -19241 74830 -19094 75066
rect -18858 75028 -16831 75066
rect -16767 75028 -16690 75092
rect -18858 75012 -16690 75028
rect -15243 75251 -13830 75253
rect -15243 75015 -15096 75251
rect -14860 75194 -13830 75251
rect -13766 75194 -13674 75258
rect -14860 75178 -13674 75194
rect -14860 75114 -13830 75178
rect -13766 75114 -13674 75178
rect 11083 76694 11323 76878
rect 11083 76630 11175 76694
rect 11239 76630 11323 76694
rect 11083 76614 11323 76630
rect 11083 76550 11175 76614
rect 11239 76550 11323 76614
rect 11083 76534 11323 76550
rect 11083 76470 11175 76534
rect 11239 76470 11323 76534
rect 11083 76454 11323 76470
rect 11083 76390 11175 76454
rect 11239 76390 11323 76454
rect 11083 76374 11323 76390
rect 11083 76310 11175 76374
rect 11239 76310 11323 76374
rect 11083 76294 11323 76310
rect 11083 76230 11175 76294
rect 11239 76230 11323 76294
rect 11083 76214 11323 76230
rect 11083 76150 11175 76214
rect 11239 76150 11323 76214
rect 11083 76134 11323 76150
rect 11083 76070 11175 76134
rect 11239 76070 11323 76134
rect 11083 76054 11323 76070
rect 11083 75990 11175 76054
rect 11239 75990 11323 76054
rect 11083 75974 11323 75990
rect 11083 75910 11175 75974
rect 11239 75910 11323 75974
rect 11083 75894 11323 75910
rect 11083 75830 11175 75894
rect 11239 75830 11323 75894
rect 11083 75814 11323 75830
rect 11083 75750 11175 75814
rect 11239 75750 11323 75814
rect 11083 75734 11323 75750
rect 11083 75670 11175 75734
rect 11239 75670 11323 75734
rect 11083 75654 11323 75670
rect 11083 75590 11175 75654
rect 11239 75590 11323 75654
rect 11083 75574 11323 75590
rect 11083 75510 11175 75574
rect 11239 75510 11323 75574
rect 11083 75494 11323 75510
rect 11083 75430 11175 75494
rect 11239 75430 11323 75494
rect 11083 75414 11323 75430
rect 11083 75350 11175 75414
rect 11239 75350 11323 75414
rect 11083 75334 11323 75350
rect 11083 75270 11175 75334
rect 11239 75270 11323 75334
rect 11083 75254 11323 75270
rect 11083 75190 11175 75254
rect 11239 75190 11323 75254
rect 11083 75174 11323 75190
rect 11083 75172 11175 75174
rect -14860 75098 -13674 75114
rect -14860 75034 -13830 75098
rect -13766 75034 -13674 75098
rect -14860 75018 -13674 75034
rect -14860 75015 -13830 75018
rect -15243 75013 -13830 75015
rect -18858 74948 -16831 75012
rect -16767 74948 -16690 75012
rect -18858 74932 -16690 74948
rect -18858 74868 -16831 74932
rect -16767 74868 -16690 74932
rect -18858 74852 -16690 74868
rect -18858 74830 -16831 74852
rect -19241 74828 -16831 74830
rect -16930 74788 -16831 74828
rect -16767 74788 -16690 74852
rect -16930 74772 -16690 74788
rect -16930 74708 -16831 74772
rect -16767 74708 -16690 74772
rect -16930 74692 -16690 74708
rect -16930 74628 -16831 74692
rect -16767 74628 -16690 74692
rect -16930 74612 -16690 74628
rect -16930 74548 -16831 74612
rect -16767 74548 -16690 74612
rect -16930 74532 -16690 74548
rect -16930 74468 -16831 74532
rect -16767 74468 -16690 74532
rect -16930 74452 -16690 74468
rect -16930 74388 -16831 74452
rect -16767 74388 -16690 74452
rect -16930 74372 -16690 74388
rect -16930 74308 -16831 74372
rect -16767 74308 -16690 74372
rect -16930 74292 -16690 74308
rect -16930 74228 -16831 74292
rect -16767 74228 -16690 74292
rect -16930 74212 -16690 74228
rect -16930 74148 -16831 74212
rect -16767 74148 -16690 74212
rect -16930 74132 -16690 74148
rect -16930 74068 -16831 74132
rect -16767 74068 -16690 74132
rect -16930 74052 -16690 74068
rect -16930 73988 -16831 74052
rect -16767 73988 -16690 74052
rect -16930 73972 -16690 73988
rect -16930 73908 -16831 73972
rect -16767 73908 -16690 73972
rect -16930 73892 -16690 73908
rect -16930 73828 -16831 73892
rect -16767 73828 -16690 73892
rect -16930 73812 -16690 73828
rect -16930 73748 -16831 73812
rect -16767 73748 -16690 73812
rect -16930 73732 -16690 73748
rect -16930 73668 -16831 73732
rect -16767 73668 -16690 73732
rect -16930 73652 -16690 73668
rect -16930 73588 -16831 73652
rect -16767 73588 -16690 73652
rect -16930 73572 -16690 73588
rect -16930 73508 -16831 73572
rect -16767 73508 -16690 73572
rect -16930 73492 -16690 73508
rect -16930 73428 -16831 73492
rect -16767 73428 -16690 73492
rect -16930 72559 -16690 73428
rect -13914 74954 -13830 75013
rect -13766 74954 -13674 75018
rect -13914 74938 -13674 74954
rect -13914 74874 -13830 74938
rect -13766 74874 -13674 74938
rect 11082 75110 11175 75172
rect 11239 75172 11323 75174
rect 14083 76707 14323 76876
rect 14083 76643 14176 76707
rect 14240 76643 14323 76707
rect 14083 76627 14323 76643
rect 14083 76563 14176 76627
rect 14240 76563 14323 76627
rect 14083 76547 14323 76563
rect 14083 76483 14176 76547
rect 14240 76483 14323 76547
rect 14083 76467 14323 76483
rect 14083 76403 14176 76467
rect 14240 76403 14323 76467
rect 14083 76387 14323 76403
rect 14083 76323 14176 76387
rect 14240 76323 14323 76387
rect 14083 76307 14323 76323
rect 14083 76243 14176 76307
rect 14240 76243 14323 76307
rect 14083 76227 14323 76243
rect 14083 76163 14176 76227
rect 14240 76163 14323 76227
rect 14083 76147 14323 76163
rect 14083 76083 14176 76147
rect 14240 76083 14323 76147
rect 14083 76067 14323 76083
rect 14083 76003 14176 76067
rect 14240 76003 14323 76067
rect 14083 75987 14323 76003
rect 14083 75923 14176 75987
rect 14240 75923 14323 75987
rect 14083 75907 14323 75923
rect 14083 75843 14176 75907
rect 14240 75843 14323 75907
rect 14083 75827 14323 75843
rect 14083 75763 14176 75827
rect 14240 75763 14323 75827
rect 14083 75747 14323 75763
rect 14083 75683 14176 75747
rect 14240 75683 14323 75747
rect 14083 75667 14323 75683
rect 14083 75603 14176 75667
rect 14240 75603 14323 75667
rect 14083 75587 14323 75603
rect 14083 75523 14176 75587
rect 14240 75523 14323 75587
rect 14083 75507 14323 75523
rect 14083 75443 14176 75507
rect 14240 75443 14323 75507
rect 14083 75427 14323 75443
rect 14083 75363 14176 75427
rect 14240 75363 14323 75427
rect 14083 75347 14323 75363
rect 14083 75283 14176 75347
rect 14240 75283 14323 75347
rect 14083 75267 14323 75283
rect 14083 75203 14176 75267
rect 14240 75203 14323 75267
rect 14083 75187 14323 75203
rect 11239 75170 13288 75172
rect 11239 75110 12905 75170
rect 11082 75094 12905 75110
rect 11082 75030 11175 75094
rect 11239 75030 12905 75094
rect 11082 75014 12905 75030
rect 11082 74950 11175 75014
rect 11239 74950 12905 75014
rect 11082 74934 12905 74950
rect 13141 74934 13288 75170
rect 11082 74932 11175 74934
rect -13914 74858 -13674 74874
rect -13914 74794 -13830 74858
rect -13766 74794 -13674 74858
rect -13914 74778 -13674 74794
rect -13914 74714 -13830 74778
rect -13766 74714 -13674 74778
rect -13914 74698 -13674 74714
rect -13914 74634 -13830 74698
rect -13766 74634 -13674 74698
rect -13914 74618 -13674 74634
rect -13914 74554 -13830 74618
rect -13766 74554 -13674 74618
rect -13914 74538 -13674 74554
rect -13914 74474 -13830 74538
rect -13766 74474 -13674 74538
rect -13914 74458 -13674 74474
rect -13914 74394 -13830 74458
rect -13766 74394 -13674 74458
rect -13914 74378 -13674 74394
rect -13914 74314 -13830 74378
rect -13766 74314 -13674 74378
rect -13914 74298 -13674 74314
rect -13914 74234 -13830 74298
rect -13766 74234 -13674 74298
rect -13914 74218 -13674 74234
rect -13914 74154 -13830 74218
rect -13766 74154 -13674 74218
rect -13914 74138 -13674 74154
rect -13914 74074 -13830 74138
rect -13766 74074 -13674 74138
rect -13914 74058 -13674 74074
rect -13914 73994 -13830 74058
rect -13766 73994 -13674 74058
rect -13914 73978 -13674 73994
rect -13914 73914 -13830 73978
rect -13766 73914 -13674 73978
rect -13914 73898 -13674 73914
rect -13914 73834 -13830 73898
rect -13766 73834 -13674 73898
rect -13914 73818 -13674 73834
rect -13914 73754 -13830 73818
rect -13766 73754 -13674 73818
rect -13914 73738 -13674 73754
rect -13914 73674 -13830 73738
rect -13766 73674 -13674 73738
rect -13914 73658 -13674 73674
rect -13914 73594 -13830 73658
rect -13766 73594 -13674 73658
rect -13914 73578 -13674 73594
rect -13914 73514 -13830 73578
rect -13766 73514 -13674 73578
rect -13914 73498 -13674 73514
rect -13914 73434 -13830 73498
rect -13766 73434 -13674 73498
rect -13914 73242 -13674 73434
rect 11083 74870 11175 74932
rect 11239 74932 13288 74934
rect 14083 75123 14176 75187
rect 14240 75164 14323 75187
rect 14240 75162 17287 75164
rect 14240 75123 16904 75162
rect 14083 75107 16904 75123
rect 14083 75043 14176 75107
rect 14240 75043 16904 75107
rect 14083 75027 16904 75043
rect 14083 74963 14176 75027
rect 14240 74963 16904 75027
rect 14083 74947 16904 74963
rect 11239 74870 11323 74932
rect 11083 74854 11323 74870
rect 11083 74790 11175 74854
rect 11239 74790 11323 74854
rect 11083 74774 11323 74790
rect 11083 74710 11175 74774
rect 11239 74710 11323 74774
rect 11083 74694 11323 74710
rect 11083 74630 11175 74694
rect 11239 74630 11323 74694
rect 11083 74614 11323 74630
rect 11083 74550 11175 74614
rect 11239 74550 11323 74614
rect 11083 74534 11323 74550
rect 11083 74470 11175 74534
rect 11239 74470 11323 74534
rect 11083 74454 11323 74470
rect 11083 74390 11175 74454
rect 11239 74390 11323 74454
rect 11083 74374 11323 74390
rect 11083 74310 11175 74374
rect 11239 74310 11323 74374
rect 11083 74294 11323 74310
rect 11083 74230 11175 74294
rect 11239 74230 11323 74294
rect 11083 74214 11323 74230
rect 11083 74150 11175 74214
rect 11239 74150 11323 74214
rect 11083 74134 11323 74150
rect 11083 74070 11175 74134
rect 11239 74070 11323 74134
rect 11083 74054 11323 74070
rect 11083 73990 11175 74054
rect 11239 73990 11323 74054
rect 11083 73974 11323 73990
rect 11083 73910 11175 73974
rect 11239 73910 11323 73974
rect 11083 73894 11323 73910
rect 11083 73830 11175 73894
rect 11239 73830 11323 73894
rect 11083 73814 11323 73830
rect 11083 73750 11175 73814
rect 11239 73750 11323 73814
rect 11083 73734 11323 73750
rect 11083 73670 11175 73734
rect 11239 73670 11323 73734
rect 11083 73654 11323 73670
rect 11083 73590 11175 73654
rect 11239 73590 11323 73654
rect 11083 73574 11323 73590
rect 11083 73510 11175 73574
rect 11239 73510 11323 73574
rect 11083 73494 11323 73510
rect 11083 73430 11175 73494
rect 11239 73430 11323 73494
rect 11083 73244 11323 73430
rect 14083 74883 14176 74947
rect 14240 74926 16904 74947
rect 17140 74926 17287 75162
rect 14240 74924 17287 74926
rect 14240 74883 14323 74924
rect 14083 74867 14323 74883
rect 14083 74803 14176 74867
rect 14240 74803 14323 74867
rect 14083 74787 14323 74803
rect 14083 74723 14176 74787
rect 14240 74723 14323 74787
rect 14083 74707 14323 74723
rect 14083 74643 14176 74707
rect 14240 74643 14323 74707
rect 14083 74627 14323 74643
rect 14083 74563 14176 74627
rect 14240 74563 14323 74627
rect 14083 74547 14323 74563
rect 14083 74483 14176 74547
rect 14240 74483 14323 74547
rect 14083 74467 14323 74483
rect 14083 74403 14176 74467
rect 14240 74403 14323 74467
rect 14083 74387 14323 74403
rect 14083 74323 14176 74387
rect 14240 74323 14323 74387
rect 14083 74307 14323 74323
rect 14083 74243 14176 74307
rect 14240 74243 14323 74307
rect 14083 74227 14323 74243
rect 14083 74163 14176 74227
rect 14240 74163 14323 74227
rect 14083 74147 14323 74163
rect 14083 74083 14176 74147
rect 14240 74083 14323 74147
rect 14083 74067 14323 74083
rect 14083 74003 14176 74067
rect 14240 74003 14323 74067
rect 14083 73987 14323 74003
rect 14083 73923 14176 73987
rect 14240 73923 14323 73987
rect 14083 73907 14323 73923
rect 14083 73843 14176 73907
rect 14240 73843 14323 73907
rect 14083 73827 14323 73843
rect 14083 73763 14176 73827
rect 14240 73763 14323 73827
rect 14083 73747 14323 73763
rect 14083 73683 14176 73747
rect 14240 73683 14323 73747
rect 14083 73667 14323 73683
rect 14083 73603 14176 73667
rect 14240 73603 14323 73667
rect 14083 73587 14323 73603
rect 14083 73523 14176 73587
rect 14240 73523 14323 73587
rect 14083 73507 14323 73523
rect 14083 73443 14176 73507
rect 14240 73443 14323 73507
rect 14083 73232 14323 73443
rect -16930 72495 -14071 72559
rect -16665 71802 -16599 71803
rect -16665 71738 -16664 71802
rect -16600 71738 -16599 71802
rect -15486 71799 -15422 72495
rect -15270 71805 -15204 71806
rect -16665 71737 -16599 71738
rect -15487 71798 -15421 71799
rect -16664 70898 -16600 71737
rect -15487 71734 -15486 71798
rect -15422 71734 -15421 71798
rect -15270 71741 -15269 71805
rect -15205 71741 -15204 71805
rect -14135 71803 -14071 72495
rect -15270 71740 -15204 71741
rect -14136 71802 -14070 71803
rect -15487 71733 -15421 71734
rect -15269 70994 -15205 71740
rect -14136 71738 -14135 71802
rect -14071 71738 -14070 71802
rect -14136 71737 -14070 71738
rect -15269 70992 -14712 70994
rect -15269 70898 -15095 70992
rect -16664 70834 -15095 70898
rect -16664 70303 -16600 70834
rect -15242 70756 -15095 70834
rect -14859 70756 -14712 70992
rect -15242 70754 -14712 70756
rect -16664 70298 -16489 70303
rect -19241 70235 -18665 70237
rect -19241 69999 -19094 70235
rect -18858 70143 -18665 70235
rect -16664 70234 -16554 70298
rect -16490 70234 -16489 70298
rect -15227 70286 -15163 70754
rect -15228 70285 -15162 70286
rect -16555 70233 -16489 70234
rect -15441 70284 -15375 70285
rect -15441 70220 -15440 70284
rect -15376 70220 -15375 70284
rect -15228 70221 -15227 70285
rect -15163 70221 -15162 70285
rect -15228 70220 -15162 70221
rect -14064 70285 -13998 70286
rect -14064 70221 -14063 70285
rect -13999 70221 -13998 70285
rect -14064 70220 -13998 70221
rect -15441 70219 -15375 70220
rect -15440 70143 -15376 70219
rect -14063 70143 -13999 70220
rect -18858 70079 -13999 70143
rect -18858 69999 -18665 70079
rect -19241 69997 -18665 69999
rect 36630 69334 36696 69335
rect 36630 69270 36631 69334
rect 36695 69270 36696 69334
rect 36630 69258 36696 69270
rect -15239 68913 -14709 68915
rect -15239 68807 -15092 68913
rect -16577 68743 -15092 68807
rect -16577 67614 -16513 68743
rect -15962 68262 -15898 68743
rect -15239 68677 -15092 68743
rect -14856 68807 -14709 68913
rect -14856 68743 -14240 68807
rect -14856 68677 -14709 68743
rect -15239 68675 -14709 68677
rect -15422 68516 -15358 68542
rect -15423 68492 -15357 68516
rect -15423 68428 -15422 68492
rect -15358 68428 -15357 68492
rect -15423 68412 -15357 68428
rect -15423 68348 -15422 68412
rect -15358 68348 -15357 68412
rect -15423 68332 -15357 68348
rect -15423 68268 -15422 68332
rect -15358 68268 -15357 68332
rect -15964 68255 -15889 68262
rect -15964 68191 -15959 68255
rect -15895 68191 -15889 68255
rect -15964 68175 -15889 68191
rect -15964 68111 -15959 68175
rect -15895 68111 -15889 68175
rect -15423 68252 -15357 68268
rect -14874 68265 -14810 68675
rect -15423 68188 -15422 68252
rect -15358 68188 -15357 68252
rect -15423 68165 -15357 68188
rect -14880 68258 -14805 68265
rect -14880 68194 -14875 68258
rect -14811 68194 -14805 68258
rect -14880 68178 -14805 68194
rect -15964 68104 -15889 68111
rect -16578 67613 -16512 67614
rect -16578 67549 -16577 67613
rect -16513 67549 -16512 67613
rect -15422 67608 -15358 68165
rect -14880 68114 -14875 68178
rect -14811 68114 -14805 68178
rect -14880 68107 -14805 68114
rect -14304 67619 -14240 68743
rect 36064 68741 36132 68743
rect 36064 68677 36066 68741
rect 36130 68677 36132 68741
rect 36064 68675 36132 68677
rect 36065 68638 36131 68675
rect 35475 68081 35543 68083
rect 35475 68017 35477 68081
rect 35541 68017 35543 68081
rect 35475 68015 35543 68017
rect -14305 67618 -14239 67619
rect -16578 67548 -16512 67549
rect -15423 67607 -15357 67608
rect -15423 67543 -15422 67607
rect -15358 67543 -15357 67607
rect -14305 67554 -14304 67618
rect -14240 67554 -14239 67618
rect -14305 67553 -14239 67554
rect -15423 67542 -15357 67543
rect -19245 67120 -18715 67122
rect -19245 66884 -19098 67120
rect -18862 67030 -18715 67120
rect -15422 67030 -15358 67542
rect -18862 66966 -15358 67030
rect -18862 66884 -18715 66966
rect -19245 66882 -18715 66884
rect -13096 66770 -13032 66772
rect -13097 66769 -13031 66770
rect -13097 66705 -13096 66769
rect -13032 66705 -13031 66769
rect -13097 66704 -13031 66705
rect -8074 66769 -8008 66770
rect -8074 66705 -8073 66769
rect -8009 66705 -8008 66769
rect -8074 66704 -8008 66705
rect -13096 59581 -13032 66704
rect -12316 66446 -12250 66447
rect -12316 66382 -12315 66446
rect -12251 66382 -12250 66446
rect -12316 66381 -12250 66382
rect -12315 59581 -12251 66381
rect -11305 66014 -11241 66018
rect -11306 66013 -11240 66014
rect -11306 65949 -11305 66013
rect -11241 65949 -11240 66013
rect -11306 65948 -11240 65949
rect -11305 59581 -11241 65948
rect -10536 65761 -10472 65768
rect -10537 65760 -10471 65761
rect -10537 65696 -10536 65760
rect -10472 65696 -10471 65760
rect -10537 65695 -10471 65696
rect -11072 63533 -10736 63558
rect -11072 63229 -11056 63533
rect -10752 63229 -10736 63533
rect -11072 63204 -10736 63229
rect -10536 59581 -10472 65695
rect -8073 65330 -8009 66704
rect -7267 66446 -7201 66447
rect -7267 66382 -7266 66446
rect -7202 66382 -7201 66446
rect -7267 66381 -7201 66382
rect -8074 65329 -8008 65330
rect -8074 65265 -8073 65329
rect -8009 65265 -8008 65329
rect -8074 65264 -8008 65265
rect -7266 65077 -7202 66381
rect -2674 66013 -2608 66014
rect -2674 65949 -2673 66013
rect -2609 65949 -2608 66013
rect -2674 65948 -2608 65949
rect -2673 65330 -2609 65948
rect -1867 65760 -1801 65761
rect -1867 65696 -1866 65760
rect -1802 65696 -1801 65760
rect -1867 65695 -1801 65696
rect -2674 65329 -2608 65330
rect -2674 65265 -2673 65329
rect -2609 65265 -2599 65329
rect -2674 65264 -2608 65265
rect -1866 65077 -1802 65695
rect -7267 65076 -7201 65077
rect -7267 65012 -7266 65076
rect -7202 65012 -7201 65076
rect -7267 65011 -7201 65012
rect -1867 65076 -1801 65077
rect -1867 65012 -1866 65076
rect -1802 65012 -1791 65076
rect -1867 65011 -1801 65012
rect 16717 64728 33332 64767
rect 16717 64664 17431 64728
rect 17495 64664 23959 64728
rect 24023 64664 31575 64728
rect 31639 64664 33332 64728
rect 16717 64648 33332 64664
rect 16717 64584 17431 64648
rect 17495 64584 23959 64648
rect 24023 64584 31575 64648
rect 31639 64584 33332 64648
rect 16717 64579 33332 64584
rect 16717 64573 28901 64579
rect 16717 64568 20907 64573
rect 16717 64504 17431 64568
rect 17495 64504 20907 64568
rect 16717 64488 20907 64504
rect 16717 64424 17431 64488
rect 17495 64424 20907 64488
rect 16717 64408 20907 64424
rect 16717 64344 17431 64408
rect 17495 64344 20907 64408
rect 16717 64337 20907 64344
rect 21143 64568 28901 64573
rect 21143 64504 23959 64568
rect 24023 64504 28901 64568
rect 21143 64488 28901 64504
rect 21143 64424 23959 64488
rect 24023 64424 28901 64488
rect 21143 64408 28901 64424
rect 21143 64344 23959 64408
rect 24023 64344 28901 64408
rect 21143 64343 28901 64344
rect 29137 64568 33332 64579
rect 29137 64504 31575 64568
rect 31639 64504 33332 64568
rect 29137 64488 33332 64504
rect 29137 64424 31575 64488
rect 31639 64424 33332 64488
rect 29137 64408 33332 64424
rect 29137 64344 31575 64408
rect 31639 64344 33332 64408
rect 29137 64343 33332 64344
rect 21143 64337 33332 64343
rect 16717 64328 33332 64337
rect 16717 64264 17431 64328
rect 17495 64264 23959 64328
rect 24023 64264 31575 64328
rect 31639 64264 33332 64328
rect 16717 64248 33332 64264
rect 16717 64184 17431 64248
rect 17495 64184 23959 64248
rect 24023 64184 31575 64248
rect 31639 64184 33332 64248
rect 16717 64147 33332 64184
rect -3241 63409 -2711 63411
rect -8074 63404 -7630 63405
rect -10188 63402 -10122 63403
rect -9885 63402 -9441 63403
rect -8074 63402 -8044 63404
rect -10188 63338 -10187 63402
rect -10123 63338 -9855 63402
rect -9791 63338 -9775 63402
rect -9711 63338 -9695 63402
rect -9631 63338 -9615 63402
rect -9551 63338 -9535 63402
rect -9471 63340 -8044 63402
rect -7980 63340 -7964 63404
rect -7900 63340 -7884 63404
rect -7820 63340 -7804 63404
rect -7740 63340 -7724 63404
rect -7660 63402 -7630 63404
rect -3241 63402 -3094 63409
rect -7660 63400 -3094 63402
rect -7660 63340 -6249 63400
rect -9471 63338 -6249 63340
rect -10188 63337 -10122 63338
rect -9885 63337 -9441 63338
rect -6279 63336 -6249 63338
rect -6185 63336 -6169 63400
rect -6105 63336 -6089 63400
rect -6025 63336 -6009 63400
rect -5945 63336 -5929 63400
rect -5865 63398 -3094 63400
rect -5865 63338 -4450 63398
rect -5865 63336 -5835 63338
rect -6279 63335 -5835 63336
rect -4480 63334 -4450 63338
rect -4386 63334 -4370 63398
rect -4306 63334 -4290 63398
rect -4226 63334 -4210 63398
rect -4146 63334 -4130 63398
rect -4066 63338 -3094 63398
rect -4066 63334 -4036 63338
rect -4480 63333 -4036 63334
rect -6940 63204 -6698 63207
rect -6940 62968 -6937 63204
rect -6701 62968 -6698 63204
rect -3241 63173 -3094 63338
rect -2858 63403 -2711 63409
rect -2858 63402 -2245 63403
rect -2858 63338 -2659 63402
rect -2595 63338 -2579 63402
rect -2515 63338 -2499 63402
rect -2435 63338 -2419 63402
rect -2355 63338 -2339 63402
rect -2275 63398 243 63402
rect -2275 63338 -857 63398
rect -2858 63337 -2245 63338
rect -2858 63173 -2711 63337
rect -887 63334 -857 63338
rect -793 63334 -777 63398
rect -713 63334 -697 63398
rect -633 63334 -617 63398
rect -553 63334 -537 63398
rect -473 63338 243 63398
rect -473 63334 -443 63338
rect -887 63333 -443 63334
rect -3241 63171 -2711 63173
rect 756 63230 1288 63233
rect 756 63224 904 63230
rect 1140 63224 1288 63230
rect 756 63000 790 63224
rect 1254 63000 1288 63224
rect 756 62994 904 63000
rect 1140 62994 1288 63000
rect 756 62991 1288 62994
rect -6940 62965 -6698 62968
rect 16715 62725 33227 62767
rect 16715 62661 17976 62725
rect 18040 62661 19064 62725
rect 19128 62661 21240 62725
rect 21304 62661 22328 62725
rect 22392 62661 23416 62725
rect 23480 62661 24504 62725
rect 24568 62661 25592 62725
rect 25656 62661 26680 62725
rect 26744 62661 28856 62725
rect 28920 62661 29944 62725
rect 30008 62661 31032 62725
rect 31096 62717 33227 62725
rect 31096 62661 33290 62717
rect 16715 62645 33290 62661
rect 16715 62582 17976 62645
rect 16715 62346 16910 62582
rect 17146 62581 17976 62582
rect 18040 62581 19064 62645
rect 19128 62581 21240 62645
rect 21304 62581 22328 62645
rect 22392 62581 23416 62645
rect 23480 62581 24504 62645
rect 24568 62581 25592 62645
rect 25656 62581 26680 62645
rect 26744 62581 28856 62645
rect 28920 62581 29944 62645
rect 30008 62581 31032 62645
rect 31096 62581 33290 62645
rect 17146 62575 33290 62581
rect 17146 62565 24906 62575
rect 17146 62501 17976 62565
rect 18040 62501 19064 62565
rect 19128 62501 21240 62565
rect 21304 62501 22328 62565
rect 22392 62501 23416 62565
rect 23480 62501 24504 62565
rect 24568 62501 24906 62565
rect 17146 62485 24906 62501
rect 17146 62421 17976 62485
rect 18040 62421 19064 62485
rect 19128 62421 21240 62485
rect 21304 62421 22328 62485
rect 22392 62421 23416 62485
rect 23480 62421 24504 62485
rect 24568 62421 24906 62485
rect 17146 62405 24906 62421
rect 17146 62346 17976 62405
rect 16715 62341 17976 62346
rect 18040 62341 19064 62405
rect 19128 62341 21240 62405
rect 21304 62341 22328 62405
rect 22392 62341 23416 62405
rect 23480 62341 24504 62405
rect 24568 62341 24906 62405
rect 16715 62339 24906 62341
rect 25142 62571 33290 62575
rect 25142 62565 32909 62571
rect 25142 62501 25592 62565
rect 25656 62501 26680 62565
rect 26744 62501 28856 62565
rect 28920 62501 29944 62565
rect 30008 62501 31032 62565
rect 31096 62501 32909 62565
rect 25142 62485 32909 62501
rect 25142 62421 25592 62485
rect 25656 62421 26680 62485
rect 26744 62421 28856 62485
rect 28920 62421 29944 62485
rect 30008 62421 31032 62485
rect 31096 62421 32909 62485
rect 25142 62405 32909 62421
rect 25142 62341 25592 62405
rect 25656 62341 26680 62405
rect 26744 62341 28856 62405
rect 28920 62341 29944 62405
rect 30008 62341 31032 62405
rect 31096 62341 32909 62405
rect 25142 62339 32909 62341
rect 16715 62335 32909 62339
rect 33145 62335 33290 62571
rect 16715 62325 33290 62335
rect 16715 62261 17976 62325
rect 18040 62261 19064 62325
rect 19128 62261 21240 62325
rect 21304 62261 22328 62325
rect 22392 62261 23416 62325
rect 23480 62261 24504 62325
rect 24568 62261 25592 62325
rect 25656 62261 26680 62325
rect 26744 62261 28856 62325
rect 28920 62261 29944 62325
rect 30008 62261 31032 62325
rect 31096 62261 33290 62325
rect 16715 62245 33290 62261
rect 16715 62181 17976 62245
rect 18040 62181 19064 62245
rect 19128 62181 21240 62245
rect 21304 62181 22328 62245
rect 22392 62181 23416 62245
rect 23480 62181 24504 62245
rect 24568 62181 25592 62245
rect 25656 62181 26680 62245
rect 26744 62181 28856 62245
rect 28920 62181 29944 62245
rect 30008 62181 31032 62245
rect 31096 62189 33290 62245
rect 31096 62181 33227 62189
rect 16715 62147 33227 62181
rect -13469 59517 -13032 59581
rect -19238 50688 -18708 50690
rect -19238 50452 -19091 50688
rect -18855 50452 -18708 50688
rect -19238 50450 -18708 50452
rect -27236 49824 -26706 49826
rect -27236 49588 -27089 49824
rect -26853 49720 -26706 49824
rect -26826 49656 -26810 49720
rect -26746 49656 -26706 49720
rect -26853 49588 -26706 49656
rect -27236 49586 -26706 49588
rect -26125 49221 -22704 49223
rect -26125 49178 -23087 49221
rect -26125 49114 -25964 49178
rect -25900 49114 -25884 49178
rect -25820 49114 -25804 49178
rect -25740 49114 -25724 49178
rect -25660 49114 -23087 49178
rect -26125 48985 -23087 49114
rect -22851 48985 -22704 49221
rect -26125 48983 -22704 48985
rect -27162 43278 -26922 43373
rect -27162 43214 -27071 43278
rect -27007 43214 -26922 43278
rect -27162 43198 -26922 43214
rect -27162 43134 -27071 43198
rect -27007 43156 -26922 43198
rect -27007 43154 -26709 43156
rect -27162 43118 -27054 43134
rect -27162 43054 -27071 43118
rect -27162 43038 -27054 43054
rect -27162 42974 -27071 43038
rect -27162 42958 -27054 42974
rect -27162 42894 -27071 42958
rect -26818 42918 -26709 43154
rect -13469 43062 -13405 59517
rect -13096 52391 -13032 59517
rect -12693 59517 -12251 59581
rect -13097 52390 -13031 52391
rect -13097 52326 -13096 52390
rect -13032 52326 -13031 52390
rect -13097 52325 -13031 52326
rect -13470 43061 -13404 43062
rect -13470 42997 -13469 43061
rect -13405 42997 -13404 43061
rect -13470 42996 -13404 42997
rect -13469 42992 -13405 42996
rect -27007 42916 -26709 42918
rect -27007 42894 -26922 42916
rect -27162 42878 -26922 42894
rect -27162 42814 -27071 42878
rect -27007 42814 -26922 42878
rect -27162 42137 -26922 42814
rect -12693 42399 -12629 59517
rect -12315 52714 -12251 59517
rect -11713 59517 -11241 59581
rect -12316 52713 -12250 52714
rect -12316 52649 -12315 52713
rect -12251 52649 -12250 52713
rect -12316 52648 -12250 52649
rect -11713 44606 -11649 59517
rect -11305 53147 -11241 59517
rect -10905 59517 -10472 59581
rect -11306 53146 -11240 53147
rect -11306 53082 -11305 53146
rect -11241 53082 -11240 53146
rect -11306 53081 -11240 53082
rect -11362 47256 -11296 47257
rect -11362 47192 -11361 47256
rect -11297 47192 -11296 47256
rect -11362 47191 -11296 47192
rect -11361 44606 -11297 47191
rect -11713 44542 -11297 44606
rect -10905 44619 -10841 59517
rect -10536 53403 -10472 59517
rect 344 60806 640 60887
rect -6978 55329 -6706 55397
rect -6978 55093 -6960 55329
rect -6724 55093 -6706 55329
rect -6978 55009 -6706 55093
rect -6978 54773 -6960 55009
rect -6724 54773 -6706 55009
rect -6978 54706 -6706 54773
rect -6865 54597 -6801 54706
rect -6867 54596 -6801 54597
rect -8558 54595 -8492 54596
rect -6867 54595 -6866 54596
rect -8558 54531 -8557 54595
rect -8493 54532 -6866 54595
rect -6802 54595 -6801 54596
rect -5162 54595 -5096 54596
rect -3366 54595 -3300 54596
rect -1537 54595 -1471 54596
rect -6802 54532 -5161 54595
rect -8493 54531 -5161 54532
rect -5097 54531 -3365 54595
rect -3301 54531 -1536 54595
rect -1472 54531 240 54595
rect -8558 54530 -8492 54531
rect -5162 54530 -5096 54531
rect -3366 54530 -3300 54531
rect -1537 54530 -1471 54531
rect -3237 54420 -2707 54422
rect -6110 54404 -5866 54405
rect -9705 54403 -9461 54404
rect -6110 54403 -6100 54404
rect -9731 54339 -9695 54403
rect -9631 54339 -9615 54403
rect -9551 54339 -9535 54403
rect -9471 54402 -6100 54403
rect -9471 54339 -7900 54402
rect -9705 54338 -9461 54339
rect -7910 54338 -7900 54339
rect -7836 54338 -7820 54402
rect -7756 54338 -7740 54402
rect -7676 54340 -6100 54402
rect -6036 54340 -6020 54404
rect -5956 54340 -5940 54404
rect -5876 54403 -5866 54404
rect -4312 54403 -4068 54404
rect -3237 54403 -3090 54420
rect -5876 54340 -4302 54403
rect -7676 54339 -4302 54340
rect -4238 54339 -4222 54403
rect -4158 54339 -4142 54403
rect -4078 54339 -3090 54403
rect -7676 54338 -7666 54339
rect -4312 54338 -4068 54339
rect -7910 54337 -7666 54338
rect -3237 54184 -3090 54339
rect -2854 54403 -2707 54420
rect 176 54405 240 54531
rect -2514 54404 -2270 54405
rect 175 54404 241 54405
rect -2514 54403 -2504 54404
rect -2854 54340 -2504 54403
rect -2440 54340 -2424 54404
rect -2360 54340 -2344 54404
rect -2280 54403 -2270 54404
rect -711 54403 -467 54404
rect -2280 54340 -701 54403
rect -2854 54339 -701 54340
rect -637 54339 -621 54403
rect -557 54339 -541 54403
rect -477 54339 -467 54403
rect 175 54340 176 54404
rect 240 54340 241 54404
rect 175 54339 241 54340
rect -2854 54184 -2707 54339
rect -711 54338 -467 54339
rect -3237 54182 -2707 54184
rect -7266 54083 -7200 54084
rect -7266 54019 -7265 54083
rect -7201 54019 -7200 54083
rect -7266 54018 -7200 54019
rect -1866 54083 -1800 54084
rect -1866 54019 -1865 54083
rect -1801 54019 -1791 54083
rect -1866 54018 -1800 54019
rect -8074 53830 -8008 53831
rect -8074 53766 -8073 53830
rect -8009 53766 -8008 53830
rect -8074 53765 -8008 53766
rect -10537 53402 -10471 53403
rect -10537 53338 -10536 53402
rect -10472 53338 -10471 53402
rect -10537 53337 -10471 53338
rect -8073 52391 -8009 53765
rect -7265 52714 -7201 54018
rect -2674 53830 -2608 53831
rect -2674 53766 -2673 53830
rect -2609 53766 -2599 53830
rect -2674 53765 -2608 53766
rect -2673 53147 -2609 53765
rect -1865 53403 -1801 54018
rect -1866 53402 -1800 53403
rect -1866 53338 -1865 53402
rect -1801 53338 -1800 53402
rect 344 53400 361 60806
rect -1866 53337 -1800 53338
rect -2674 53146 -2608 53147
rect -2674 53082 -2673 53146
rect -2609 53082 -2608 53146
rect 338 53142 361 53400
rect 505 60125 640 60806
rect 10176 60818 10552 60837
rect 505 60124 768 60125
rect 505 60122 1286 60124
rect 505 59886 903 60122
rect 1139 59886 1286 60122
rect 10176 60113 10212 60818
rect 505 59884 1286 59886
rect 8761 60111 10212 60113
rect 505 57511 640 59884
rect 8761 59875 8908 60111
rect 9144 59875 10212 60111
rect 8761 59873 10212 59875
rect 505 57271 757 57511
rect 505 56750 640 57271
rect 505 56749 668 56750
rect 505 56747 1286 56749
rect 505 56511 903 56747
rect 1139 56511 1286 56747
rect 10176 56738 10212 59873
rect 505 56509 1286 56511
rect 8760 56736 10212 56738
rect 505 56508 668 56509
rect 505 53400 640 56508
rect 8760 56500 8907 56736
rect 9143 56500 10212 56736
rect 8760 56498 10212 56500
rect 505 53399 671 53400
rect 505 53372 1315 53399
rect 505 53142 903 53372
rect 338 53136 903 53142
rect 1139 53345 1315 53372
rect 10176 53363 10212 56498
rect 8760 53361 10212 53363
rect 1139 53167 1344 53345
rect 1139 53136 1315 53167
rect 338 53104 1315 53136
rect 8760 53125 8907 53361
rect 9143 53125 10212 53361
rect 8760 53123 10212 53125
rect -2674 53081 -2608 53082
rect -7266 52713 -7200 52714
rect -7266 52649 -7265 52713
rect -7201 52649 -7200 52713
rect -7266 52648 -7200 52649
rect -8074 52390 -8008 52391
rect -8074 52326 -8073 52390
rect -8009 52326 -8008 52390
rect -8074 52325 -8008 52326
rect 10176 52033 10212 53123
rect 10069 51855 10212 52033
rect -9010 51699 -6707 51701
rect -9010 51463 -7090 51699
rect -6854 51463 -6707 51699
rect -9010 51461 -6707 51463
rect -9010 51250 -8770 51461
rect -9010 51243 -8769 51250
rect -9010 51179 -8844 51243
rect -8780 51179 -8769 51243
rect -7723 51247 -7657 51248
rect -7723 51183 -7722 51247
rect -7658 51183 -7657 51247
rect -7723 51182 -7657 51183
rect -9010 51163 -8769 51179
rect -9010 51099 -8844 51163
rect -8780 51099 -8769 51163
rect -9010 51083 -8769 51099
rect -9010 51019 -8844 51083
rect -8780 51019 -8769 51083
rect -9010 51014 -8769 51019
rect -8855 51013 -8769 51014
rect -8875 50776 -8777 50792
rect -8875 50712 -8859 50776
rect -8795 50712 -8777 50776
rect -8875 50696 -8777 50712
rect -8875 50632 -8859 50696
rect -8795 50632 -8777 50696
rect -8875 50616 -8777 50632
rect -8875 50552 -8859 50616
rect -8795 50552 -8777 50616
rect -8875 50536 -8777 50552
rect -8875 50472 -8859 50536
rect -8795 50472 -8777 50536
rect -8875 50456 -8777 50472
rect -8875 50392 -8859 50456
rect -8795 50392 -8777 50456
rect -8875 50377 -8777 50392
rect -8481 50441 -8415 50442
rect -8481 50377 -8480 50441
rect -8416 50377 -8415 50441
rect -8481 50376 -8415 50377
rect -8480 50073 -8416 50376
rect -8481 50072 -8415 50073
rect -8481 50008 -8480 50072
rect -8416 50008 -8415 50072
rect -8481 50007 -8415 50008
rect -10488 46633 -10422 46634
rect -10488 46569 -10487 46633
rect -10423 46569 -10422 46633
rect -10488 46568 -10422 46569
rect -10487 44619 -10423 46568
rect -10905 44555 -10423 44619
rect -12694 42398 -12628 42399
rect -12694 42334 -12693 42398
rect -12629 42334 -12628 42398
rect -12694 42333 -12628 42334
rect -12693 42328 -12629 42333
rect -27162 42073 -27071 42137
rect -27007 42073 -26922 42137
rect -21476 42163 -21410 42164
rect -21476 42099 -21475 42163
rect -21411 42099 -17680 42163
rect -21476 42098 -21410 42099
rect -27162 42057 -26922 42073
rect -27162 41993 -27071 42057
rect -27007 41993 -26922 42057
rect -27162 41977 -26922 41993
rect -27162 41913 -27071 41977
rect -27007 41913 -26922 41977
rect -27162 41897 -26922 41913
rect -27162 41833 -27071 41897
rect -27007 41833 -26922 41897
rect -27162 41817 -26922 41833
rect -27162 41753 -27071 41817
rect -27007 41753 -26922 41817
rect -27162 41737 -26922 41753
rect -27162 41673 -27071 41737
rect -27007 41673 -26922 41737
rect -27162 41657 -26922 41673
rect -27162 41593 -27071 41657
rect -27007 41593 -26922 41657
rect -27162 41577 -26922 41593
rect -27162 41513 -27071 41577
rect -27007 41513 -26922 41577
rect -27162 41497 -26922 41513
rect -27162 41433 -27071 41497
rect -27007 41433 -26922 41497
rect -27162 41417 -26922 41433
rect -27162 41353 -27071 41417
rect -27007 41353 -26922 41417
rect -27162 41337 -26922 41353
rect -27162 41273 -27071 41337
rect -27007 41273 -26922 41337
rect -27162 41257 -26922 41273
rect -27162 41193 -27071 41257
rect -27007 41193 -26922 41257
rect -27162 41177 -26922 41193
rect -27162 41113 -27071 41177
rect -27007 41113 -26922 41177
rect -27162 41097 -26922 41113
rect -27162 41033 -27071 41097
rect -27007 41033 -26922 41097
rect -27162 40611 -26922 41033
rect -27162 40547 -27066 40611
rect -27002 40547 -26922 40611
rect -27162 40531 -26922 40547
rect -27162 40467 -27066 40531
rect -27002 40467 -26922 40531
rect -27162 40451 -26922 40467
rect -27162 40387 -27066 40451
rect -27002 40387 -26922 40451
rect -27162 40371 -26922 40387
rect -27162 40307 -27066 40371
rect -27002 40307 -26922 40371
rect -27162 40291 -26922 40307
rect -27162 40227 -27066 40291
rect -27002 40227 -26922 40291
rect -27162 40211 -26922 40227
rect -27162 40147 -27066 40211
rect -27002 40147 -26922 40211
rect -27162 40131 -26922 40147
rect -27162 40067 -27066 40131
rect -27002 40067 -26922 40131
rect -27162 40051 -26922 40067
rect -27162 39987 -27066 40051
rect -27002 39987 -26922 40051
rect -27162 39971 -26922 39987
rect -27162 39907 -27066 39971
rect -27002 39950 -26922 39971
rect -27002 39948 -26699 39950
rect -27162 39891 -27049 39907
rect -27162 39827 -27066 39891
rect -27162 39811 -27049 39827
rect -27162 39747 -27066 39811
rect -27162 39731 -27049 39747
rect -27162 39667 -27066 39731
rect -26813 39712 -26699 39948
rect -17744 39824 -17680 42099
rect -17744 39760 -17097 39824
rect -27002 39710 -26699 39712
rect -27002 39667 -26922 39710
rect -27162 39651 -26922 39667
rect -27162 39587 -27066 39651
rect -27002 39587 -26922 39651
rect -27162 39571 -26922 39587
rect -27162 39507 -27066 39571
rect -27002 39507 -26922 39571
rect -31813 39148 -31747 39167
rect -31813 39084 -31812 39148
rect -31748 39084 -31747 39148
rect -31813 39068 -31747 39084
rect -31813 39004 -31812 39068
rect -31748 39023 -31747 39068
rect -27162 39108 -26922 39507
rect -27162 39044 -27072 39108
rect -27008 39044 -26922 39108
rect -27162 39028 -26922 39044
rect -31748 39004 -30945 39023
rect -31813 38988 -30945 39004
rect -31813 38924 -31812 38988
rect -31748 38959 -30945 38988
rect -31748 38924 -31747 38959
rect -31813 38908 -31747 38924
rect -31813 38844 -31812 38908
rect -31748 38844 -31747 38908
rect -31813 38826 -31747 38844
rect -31812 38609 -31746 38614
rect -31812 38545 -31811 38609
rect -31747 38545 -31746 38609
rect -31812 38529 -31746 38545
rect -35218 38496 -34755 38498
rect -35218 38260 -35105 38496
rect -34869 38415 -34755 38496
rect -31812 38465 -31811 38529
rect -31747 38465 -31746 38529
rect -31009 38509 -30945 38959
rect -27162 38964 -27072 39028
rect -27008 38964 -26922 39028
rect -27162 38948 -26922 38964
rect -27162 38884 -27072 38948
rect -27008 38884 -26922 38948
rect -27162 38868 -26922 38884
rect -27162 38804 -27072 38868
rect -27008 38804 -26922 38868
rect -27162 38788 -26922 38804
rect -27162 38724 -27072 38788
rect -27008 38724 -26922 38788
rect -27162 38708 -26922 38724
rect -27162 38644 -27072 38708
rect -27008 38644 -26922 38708
rect -27162 38628 -26922 38644
rect -27162 38564 -27072 38628
rect -27008 38564 -26922 38628
rect -27162 38548 -26922 38564
rect -31812 38449 -31746 38465
rect -31812 38415 -31811 38449
rect -34869 38385 -31811 38415
rect -31747 38385 -31746 38449
rect -34869 38369 -31746 38385
rect -34869 38351 -31811 38369
rect -34869 38260 -34755 38351
rect -35218 38258 -34755 38260
rect -31812 38305 -31811 38351
rect -31747 38305 -31746 38369
rect -31812 38289 -31746 38305
rect -31812 38225 -31811 38289
rect -31747 38225 -31746 38289
rect -31206 38507 -30743 38509
rect -31206 38271 -31093 38507
rect -30857 38413 -30743 38507
rect -27162 38484 -27072 38548
rect -27008 38484 -26922 38548
rect -27162 38468 -26922 38484
rect -29615 38413 -29149 38414
rect -30857 38349 -29614 38413
rect -29550 38349 -29534 38413
rect -29470 38349 -29454 38413
rect -29390 38349 -29374 38413
rect -29310 38349 -29294 38413
rect -29230 38349 -29214 38413
rect -29150 38349 -29149 38413
rect -30857 38271 -30743 38349
rect -29615 38348 -29149 38349
rect -27162 38404 -27072 38468
rect -27008 38404 -26922 38468
rect -27162 38388 -26922 38404
rect -31206 38269 -30743 38271
rect -27162 38324 -27072 38388
rect -27008 38324 -26922 38388
rect -27162 38308 -26922 38324
rect -31812 38209 -31746 38225
rect -31812 38145 -31811 38209
rect -31747 38145 -31746 38209
rect -31812 38140 -31746 38145
rect -27162 38244 -27072 38308
rect -27008 38244 -26922 38308
rect -31218 37409 -30755 37411
rect -31218 37173 -31105 37409
rect -30869 37323 -30755 37409
rect -27162 37341 -26922 38244
rect -18956 39502 -18716 39689
rect -18956 39438 -18877 39502
rect -18813 39438 -18716 39502
rect -18956 39422 -18716 39438
rect -18956 39358 -18877 39422
rect -18813 39358 -18716 39422
rect -18956 39342 -18716 39358
rect -18956 39278 -18877 39342
rect -18813 39278 -18716 39342
rect -18956 39262 -18716 39278
rect -18956 39198 -18877 39262
rect -18813 39198 -18716 39262
rect -18956 39182 -18716 39198
rect -18956 39118 -18877 39182
rect -18813 39118 -18716 39182
rect -18956 39102 -18716 39118
rect -18956 39038 -18877 39102
rect -18813 39038 -18716 39102
rect -18956 39022 -18716 39038
rect -18956 38958 -18877 39022
rect -18813 38958 -18716 39022
rect -18956 38942 -18716 38958
rect -18956 38878 -18877 38942
rect -18813 38878 -18716 38942
rect -18956 38862 -18716 38878
rect -18956 38798 -18877 38862
rect -18813 38798 -18716 38862
rect -18956 38782 -18716 38798
rect -11713 38791 -11649 44542
rect -11714 38790 -11648 38791
rect -13395 38783 -13331 38784
rect -18956 38718 -18877 38782
rect -18813 38718 -18716 38782
rect -14898 38719 -13331 38783
rect -11714 38726 -11713 38790
rect -11649 38726 -11648 38790
rect -11714 38725 -11648 38726
rect -11713 38724 -11649 38725
rect -18956 38702 -18716 38718
rect -18956 38638 -18877 38702
rect -18813 38638 -18716 38702
rect -18956 38622 -18716 38638
rect -18956 38558 -18877 38622
rect -18813 38558 -18716 38622
rect -18956 38542 -18716 38558
rect -18956 38478 -18877 38542
rect -18813 38478 -18716 38542
rect -18956 38462 -18716 38478
rect -18956 38398 -18877 38462
rect -18813 38398 -18716 38462
rect -18956 38382 -18716 38398
rect -18956 38318 -18877 38382
rect -18813 38318 -18716 38382
rect -18956 38302 -18716 38318
rect -18956 38238 -18877 38302
rect -18813 38238 -18716 38302
rect -18956 38222 -18716 38238
rect -18956 38158 -18877 38222
rect -18813 38158 -18716 38222
rect -18956 38142 -18716 38158
rect -18956 38078 -18877 38142
rect -18813 38078 -18716 38142
rect -18956 38062 -18716 38078
rect -23192 37904 -22729 38013
rect -18956 37998 -18877 38062
rect -18813 37998 -18716 38062
rect -18956 37982 -18716 37998
rect -18956 37918 -18877 37982
rect -18813 37918 -18716 37982
rect -18956 37904 -18716 37918
rect -23192 37902 -18716 37904
rect -23192 37894 -18877 37902
rect -23192 37658 -23079 37894
rect -22843 37838 -18877 37894
rect -18813 37838 -18716 37902
rect -22843 37822 -18716 37838
rect -22843 37758 -18877 37822
rect -18813 37758 -18716 37822
rect -15217 38281 -14731 38300
rect -15217 37817 -15206 38281
rect -14742 37817 -14731 38281
rect -15217 37798 -14731 37817
rect -22843 37742 -18716 37758
rect -22843 37678 -18877 37742
rect -18813 37678 -18716 37742
rect -22843 37664 -18716 37678
rect -22843 37658 -22729 37664
rect -23192 37540 -22729 37658
rect -18956 37662 -18716 37664
rect -18956 37598 -18877 37662
rect -18813 37598 -18716 37662
rect -18956 37582 -18716 37598
rect -29653 37323 -29142 37324
rect -30869 37259 -29630 37323
rect -29566 37259 -29550 37323
rect -29486 37259 -29470 37323
rect -29406 37259 -29390 37323
rect -29326 37259 -29310 37323
rect -29246 37259 -29230 37323
rect -29166 37259 -29142 37323
rect -30869 37173 -30755 37259
rect -29653 37258 -29142 37259
rect -27162 37277 -27069 37341
rect -27005 37277 -26922 37341
rect -27162 37261 -26922 37277
rect -31218 37171 -30755 37173
rect -27162 37197 -27069 37261
rect -27005 37197 -26922 37261
rect -27162 37181 -26922 37197
rect -27162 37117 -27069 37181
rect -27005 37117 -26922 37181
rect -27162 37101 -26922 37117
rect -27162 37037 -27069 37101
rect -27005 37037 -26922 37101
rect -27162 37021 -26922 37037
rect -27162 36957 -27069 37021
rect -27005 36957 -26922 37021
rect -27162 36941 -26922 36957
rect -27162 36877 -27069 36941
rect -27005 36877 -26922 36941
rect -27162 36861 -26922 36877
rect -27162 36797 -27069 36861
rect -27005 36797 -26922 36861
rect -27162 36781 -26922 36797
rect -27162 36717 -27069 36781
rect -27005 36717 -26922 36781
rect -27162 36701 -26922 36717
rect -27162 36637 -27069 36701
rect -27005 36637 -26922 36701
rect -27162 36621 -26922 36637
rect -27162 36557 -27069 36621
rect -27005 36557 -26922 36621
rect -27162 36541 -26922 36557
rect -27162 36477 -27069 36541
rect -27005 36477 -26922 36541
rect -27162 36124 -26922 36477
rect -27162 36060 -27069 36124
rect -27005 36060 -26922 36124
rect -27162 36044 -26922 36060
rect -27162 35980 -27069 36044
rect -27005 35980 -26922 36044
rect -27162 35964 -26922 35980
rect -27162 35900 -27069 35964
rect -27005 35900 -26922 35964
rect -18956 37518 -18877 37582
rect -18813 37518 -18716 37582
rect -18956 37502 -18716 37518
rect -18956 37438 -18877 37502
rect -18813 37438 -18716 37502
rect -18956 37422 -18716 37438
rect -18956 37358 -18877 37422
rect -18813 37358 -18716 37422
rect -18956 37342 -18716 37358
rect -18956 37278 -18877 37342
rect -18813 37278 -18716 37342
rect -18956 37262 -18716 37278
rect -18956 37198 -18877 37262
rect -18813 37198 -18716 37262
rect -18956 37182 -18716 37198
rect -18956 37118 -18877 37182
rect -18813 37118 -18716 37182
rect -18956 37102 -18716 37118
rect -18956 37038 -18877 37102
rect -18813 37038 -18716 37102
rect -18956 37022 -18716 37038
rect -18956 36958 -18877 37022
rect -18813 36958 -18716 37022
rect -18956 36942 -18716 36958
rect -18956 36878 -18877 36942
rect -18813 36878 -18716 36942
rect -18956 36862 -18716 36878
rect -18956 36798 -18877 36862
rect -18813 36798 -18716 36862
rect -18956 36782 -18716 36798
rect -18956 36718 -18877 36782
rect -18813 36718 -18716 36782
rect -18956 36702 -18716 36718
rect -18956 36638 -18877 36702
rect -18813 36638 -18716 36702
rect -18956 36622 -18716 36638
rect -18956 36558 -18877 36622
rect -18813 36558 -18716 36622
rect -18956 36542 -18716 36558
rect -18956 36478 -18877 36542
rect -18813 36478 -18716 36542
rect -18956 36462 -18716 36478
rect -18956 36398 -18877 36462
rect -18813 36398 -18716 36462
rect -18956 36382 -18716 36398
rect -18956 36318 -18877 36382
rect -18813 36318 -18716 36382
rect -18956 36302 -18716 36318
rect -18956 36238 -18877 36302
rect -18813 36238 -18716 36302
rect -18956 36222 -18716 36238
rect -18956 36158 -18877 36222
rect -18813 36158 -18716 36222
rect -18956 35957 -18716 36158
rect -17743 36329 -17006 36393
rect -27162 35884 -26922 35900
rect -27162 35820 -27069 35884
rect -27005 35881 -26922 35884
rect -27005 35879 -26699 35881
rect -27162 35804 -27049 35820
rect -27162 35740 -27069 35804
rect -27162 35724 -27049 35740
rect -27162 35660 -27069 35724
rect -27162 35644 -27049 35660
rect -27162 35580 -27069 35644
rect -26813 35643 -26699 35879
rect -27005 35641 -26699 35643
rect -27005 35580 -26922 35641
rect -27162 35564 -26922 35580
rect -27162 35500 -27069 35564
rect -27005 35500 -26922 35564
rect -27162 35484 -26922 35500
rect -27162 35420 -27069 35484
rect -27005 35420 -26922 35484
rect -27162 35404 -26922 35420
rect -27162 35340 -27069 35404
rect -27005 35340 -26922 35404
rect -27162 35324 -26922 35340
rect -27162 35260 -27069 35324
rect -27005 35260 -26922 35324
rect -27162 35244 -26922 35260
rect -27162 35180 -27069 35244
rect -27005 35180 -26922 35244
rect -27162 35164 -26922 35180
rect -27162 35100 -27069 35164
rect -27005 35100 -26922 35164
rect -27162 35084 -26922 35100
rect -27162 35020 -27069 35084
rect -27005 35020 -26922 35084
rect -27162 34686 -26922 35020
rect -27162 34622 -27072 34686
rect -27008 34622 -26922 34686
rect -27162 34606 -26922 34622
rect -27162 34542 -27072 34606
rect -27008 34542 -26922 34606
rect -27162 34526 -26922 34542
rect -27162 34462 -27072 34526
rect -27008 34462 -26922 34526
rect -27162 34446 -26922 34462
rect -27162 34382 -27072 34446
rect -27008 34382 -26922 34446
rect -27162 34366 -26922 34382
rect -27162 34302 -27072 34366
rect -27008 34302 -26922 34366
rect -27162 34286 -26922 34302
rect -27162 34222 -27072 34286
rect -27008 34222 -26922 34286
rect -27162 34206 -26922 34222
rect -27162 34142 -27072 34206
rect -27008 34142 -26922 34206
rect -27162 34126 -26922 34142
rect -27162 34062 -27072 34126
rect -27008 34062 -26922 34126
rect -27162 34046 -26922 34062
rect -27162 33982 -27072 34046
rect -27008 33982 -26922 34046
rect -27162 33966 -26922 33982
rect -27162 33902 -27072 33966
rect -27008 33902 -26922 33966
rect -27162 33886 -26922 33902
rect -27162 33822 -27072 33886
rect -27008 33822 -26922 33886
rect -27162 33806 -26922 33822
rect -27162 33742 -27072 33806
rect -27008 33742 -26922 33806
rect -27162 33726 -26922 33742
rect -27162 33662 -27072 33726
rect -27008 33662 -26922 33726
rect -27162 33646 -26922 33662
rect -27162 33582 -27072 33646
rect -27008 33582 -26922 33646
rect -27162 33566 -26922 33582
rect -27162 33502 -27072 33566
rect -27008 33502 -26922 33566
rect -27162 32864 -26922 33502
rect -21519 33551 -21453 33552
rect -17743 33551 -17679 36329
rect -21519 33487 -21518 33551
rect -21454 33487 -17679 33551
rect -21519 33486 -21453 33487
rect -15139 33180 -15075 35346
rect -13395 34677 -13331 38719
rect -10905 38448 -10841 44555
rect -9209 43061 -9143 43062
rect -9209 42997 -9208 43061
rect -9144 42997 -9143 43061
rect -9209 42996 -9143 42997
rect -10070 42398 -10004 42399
rect -10070 42334 -10069 42398
rect -10005 42334 -10004 42398
rect -10070 42333 -10004 42334
rect -10906 38447 -10840 38448
rect -10906 38383 -10905 38447
rect -10841 38383 -10840 38447
rect -10906 38382 -10840 38383
rect -10905 38376 -10841 38382
rect -10069 35352 -10005 42333
rect -9208 35942 -9144 42996
rect -8480 37372 -8416 50007
rect -7722 49425 -7658 51182
rect -5972 51121 -5695 51124
rect -5972 51099 139 51121
rect -5972 51057 -3084 51099
rect -2848 51057 139 51099
rect -5972 51046 -3341 51057
rect -5972 50902 -5660 51046
rect -3916 50913 -3341 51046
rect -2557 51047 139 51057
rect -2557 50913 -1642 51047
rect -3916 50902 -3084 50913
rect -5972 50863 -3084 50902
rect -2848 50903 -1642 50913
rect -778 50903 139 51047
rect -2848 50863 139 50903
rect -5972 50845 139 50863
rect -5972 50720 -5695 50845
rect -7723 49424 -7657 49425
rect -7723 49360 -7722 49424
rect -7658 49360 -7657 49424
rect -7723 49359 -7657 49360
rect -7722 37900 -7658 49359
rect -5972 47776 -5912 50720
rect -5768 48791 -5695 50720
rect -138 50735 139 50845
rect -138 48791 -51 50735
rect -5768 48771 -51 48791
rect -5768 48535 -3090 48771
rect -2854 48535 -51 48771
rect -5768 48514 -51 48535
rect -5768 47776 -5695 48514
rect -5972 47688 -5695 47776
rect -138 47791 -51 48514
rect 93 47791 139 50735
rect 600 49997 1298 50017
rect 600 49761 903 49997
rect 1139 49761 1298 49997
rect 10176 49988 10212 51855
rect 600 49722 1298 49761
rect 8760 49986 10212 49988
rect 8760 49750 8907 49986
rect 9143 49750 10212 49986
rect 8760 49748 10212 49750
rect -138 47715 139 47791
rect 10176 47634 10212 49748
rect 10516 47634 10552 60818
rect 16717 60728 33332 60767
rect 16717 60664 17431 60728
rect 17495 60664 18519 60728
rect 18583 60664 19607 60728
rect 19671 60664 20695 60728
rect 20759 60664 21783 60728
rect 21847 60664 22871 60728
rect 22935 60664 23959 60728
rect 24023 60664 25047 60728
rect 25111 60664 26135 60728
rect 26199 60664 27223 60728
rect 27287 60664 28311 60728
rect 28375 60664 29399 60728
rect 29463 60664 30487 60728
rect 30551 60664 31575 60728
rect 31639 60664 33332 60728
rect 16717 60648 33332 60664
rect 16717 60584 17431 60648
rect 17495 60584 18519 60648
rect 18583 60584 19607 60648
rect 19671 60584 20695 60648
rect 20759 60584 21783 60648
rect 21847 60584 22871 60648
rect 22935 60584 23959 60648
rect 24023 60584 25047 60648
rect 25111 60584 26135 60648
rect 26199 60584 27223 60648
rect 27287 60584 28311 60648
rect 28375 60584 29399 60648
rect 29463 60584 30487 60648
rect 30551 60584 31575 60648
rect 31639 60584 33332 60648
rect 16717 60579 33332 60584
rect 16717 60573 28901 60579
rect 16717 60568 20907 60573
rect 16717 60504 17431 60568
rect 17495 60504 18519 60568
rect 18583 60504 19607 60568
rect 19671 60504 20695 60568
rect 20759 60504 20907 60568
rect 16717 60488 20907 60504
rect 16717 60424 17431 60488
rect 17495 60424 18519 60488
rect 18583 60424 19607 60488
rect 19671 60424 20695 60488
rect 20759 60424 20907 60488
rect 16717 60408 20907 60424
rect 16717 60344 17431 60408
rect 17495 60344 18519 60408
rect 18583 60344 19607 60408
rect 19671 60344 20695 60408
rect 20759 60344 20907 60408
rect 16717 60337 20907 60344
rect 21143 60568 28901 60573
rect 21143 60504 21783 60568
rect 21847 60504 22871 60568
rect 22935 60504 23959 60568
rect 24023 60504 25047 60568
rect 25111 60504 26135 60568
rect 26199 60504 27223 60568
rect 27287 60504 28311 60568
rect 28375 60504 28901 60568
rect 21143 60488 28901 60504
rect 21143 60424 21783 60488
rect 21847 60424 22871 60488
rect 22935 60424 23959 60488
rect 24023 60424 25047 60488
rect 25111 60424 26135 60488
rect 26199 60424 27223 60488
rect 27287 60424 28311 60488
rect 28375 60424 28901 60488
rect 21143 60408 28901 60424
rect 21143 60344 21783 60408
rect 21847 60344 22871 60408
rect 22935 60344 23959 60408
rect 24023 60344 25047 60408
rect 25111 60344 26135 60408
rect 26199 60344 27223 60408
rect 27287 60344 28311 60408
rect 28375 60344 28901 60408
rect 21143 60343 28901 60344
rect 29137 60568 33332 60579
rect 29137 60504 29399 60568
rect 29463 60504 30487 60568
rect 30551 60504 31575 60568
rect 31639 60504 33332 60568
rect 29137 60488 33332 60504
rect 29137 60424 29399 60488
rect 29463 60424 30487 60488
rect 30551 60424 31575 60488
rect 31639 60424 33332 60488
rect 29137 60408 33332 60424
rect 29137 60344 29399 60408
rect 29463 60344 30487 60408
rect 30551 60344 31575 60408
rect 31639 60344 33332 60408
rect 29137 60343 33332 60344
rect 21143 60337 33332 60343
rect 16717 60328 33332 60337
rect 16717 60264 17431 60328
rect 17495 60264 18519 60328
rect 18583 60264 19607 60328
rect 19671 60264 20695 60328
rect 20759 60264 21783 60328
rect 21847 60264 22871 60328
rect 22935 60264 23959 60328
rect 24023 60264 25047 60328
rect 25111 60264 26135 60328
rect 26199 60264 27223 60328
rect 27287 60264 28311 60328
rect 28375 60264 29399 60328
rect 29463 60264 30487 60328
rect 30551 60264 31575 60328
rect 31639 60264 33332 60328
rect 16717 60248 33332 60264
rect 16717 60184 17431 60248
rect 17495 60184 18519 60248
rect 18583 60184 19607 60248
rect 19671 60184 20695 60248
rect 20759 60184 21783 60248
rect 21847 60184 22871 60248
rect 22935 60184 23959 60248
rect 24023 60184 25047 60248
rect 25111 60184 26135 60248
rect 26199 60184 27223 60248
rect 27287 60184 28311 60248
rect 28375 60184 29399 60248
rect 29463 60184 30487 60248
rect 30551 60184 31575 60248
rect 31639 60184 33332 60248
rect 16717 60147 33332 60184
rect 16715 58725 33227 58767
rect 16715 58661 17976 58725
rect 18040 58661 19064 58725
rect 19128 58661 20152 58725
rect 20216 58661 21240 58725
rect 21304 58661 22328 58725
rect 22392 58661 23416 58725
rect 23480 58661 24504 58725
rect 24568 58661 25592 58725
rect 25656 58661 26680 58725
rect 26744 58661 27768 58725
rect 27832 58661 28856 58725
rect 28920 58661 29944 58725
rect 30008 58661 31032 58725
rect 31096 58717 33227 58725
rect 31096 58661 33290 58717
rect 16715 58645 33290 58661
rect 16715 58582 17976 58645
rect 16715 58346 16910 58582
rect 17146 58581 17976 58582
rect 18040 58581 19064 58645
rect 19128 58581 20152 58645
rect 20216 58581 21240 58645
rect 21304 58581 22328 58645
rect 22392 58581 23416 58645
rect 23480 58581 24504 58645
rect 24568 58581 25592 58645
rect 25656 58581 26680 58645
rect 26744 58581 27768 58645
rect 27832 58581 28856 58645
rect 28920 58581 29944 58645
rect 30008 58581 31032 58645
rect 31096 58581 33290 58645
rect 17146 58575 33290 58581
rect 17146 58565 24906 58575
rect 17146 58501 17976 58565
rect 18040 58501 19064 58565
rect 19128 58501 20152 58565
rect 20216 58501 21240 58565
rect 21304 58501 22328 58565
rect 22392 58501 23416 58565
rect 23480 58501 24504 58565
rect 24568 58501 24906 58565
rect 17146 58485 24906 58501
rect 17146 58421 17976 58485
rect 18040 58421 19064 58485
rect 19128 58421 20152 58485
rect 20216 58421 21240 58485
rect 21304 58421 22328 58485
rect 22392 58421 23416 58485
rect 23480 58421 24504 58485
rect 24568 58421 24906 58485
rect 17146 58405 24906 58421
rect 17146 58346 17976 58405
rect 16715 58341 17976 58346
rect 18040 58341 19064 58405
rect 19128 58341 20152 58405
rect 20216 58341 21240 58405
rect 21304 58341 22328 58405
rect 22392 58341 23416 58405
rect 23480 58341 24504 58405
rect 24568 58341 24906 58405
rect 16715 58339 24906 58341
rect 25142 58571 33290 58575
rect 25142 58565 32909 58571
rect 25142 58501 25592 58565
rect 25656 58501 26680 58565
rect 26744 58501 27768 58565
rect 27832 58501 28856 58565
rect 28920 58501 29944 58565
rect 30008 58501 31032 58565
rect 31096 58501 32909 58565
rect 25142 58485 32909 58501
rect 25142 58421 25592 58485
rect 25656 58421 26680 58485
rect 26744 58421 27768 58485
rect 27832 58421 28856 58485
rect 28920 58421 29944 58485
rect 30008 58421 31032 58485
rect 31096 58421 32909 58485
rect 25142 58405 32909 58421
rect 25142 58341 25592 58405
rect 25656 58341 26680 58405
rect 26744 58341 27768 58405
rect 27832 58341 28856 58405
rect 28920 58341 29944 58405
rect 30008 58341 31032 58405
rect 31096 58341 32909 58405
rect 25142 58339 32909 58341
rect 16715 58335 32909 58339
rect 33145 58335 33290 58571
rect 16715 58325 33290 58335
rect 16715 58261 17976 58325
rect 18040 58261 19064 58325
rect 19128 58261 20152 58325
rect 20216 58261 21240 58325
rect 21304 58261 22328 58325
rect 22392 58261 23416 58325
rect 23480 58261 24504 58325
rect 24568 58261 25592 58325
rect 25656 58261 26680 58325
rect 26744 58261 27768 58325
rect 27832 58261 28856 58325
rect 28920 58261 29944 58325
rect 30008 58261 31032 58325
rect 31096 58261 33290 58325
rect 16715 58245 33290 58261
rect 16715 58181 17976 58245
rect 18040 58181 19064 58245
rect 19128 58181 20152 58245
rect 20216 58181 21240 58245
rect 21304 58181 22328 58245
rect 22392 58181 23416 58245
rect 23480 58181 24504 58245
rect 24568 58181 25592 58245
rect 25656 58181 26680 58245
rect 26744 58181 27768 58245
rect 27832 58181 28856 58245
rect 28920 58181 29944 58245
rect 30008 58181 31032 58245
rect 31096 58189 33290 58245
rect 31096 58181 33227 58189
rect 16715 58147 33227 58181
rect 16717 56728 33332 56767
rect 16717 56664 17431 56728
rect 17495 56664 18519 56728
rect 18583 56664 19607 56728
rect 19671 56664 20695 56728
rect 20759 56664 21783 56728
rect 21847 56664 22871 56728
rect 22935 56664 23959 56728
rect 24023 56664 25047 56728
rect 25111 56664 26135 56728
rect 26199 56664 27223 56728
rect 27287 56664 28311 56728
rect 28375 56664 29399 56728
rect 29463 56664 30487 56728
rect 30551 56664 31575 56728
rect 31639 56664 33332 56728
rect 16717 56648 33332 56664
rect 16717 56584 17431 56648
rect 17495 56584 18519 56648
rect 18583 56584 19607 56648
rect 19671 56584 20695 56648
rect 20759 56584 21783 56648
rect 21847 56584 22871 56648
rect 22935 56584 23959 56648
rect 24023 56584 25047 56648
rect 25111 56584 26135 56648
rect 26199 56584 27223 56648
rect 27287 56584 28311 56648
rect 28375 56584 29399 56648
rect 29463 56584 30487 56648
rect 30551 56584 31575 56648
rect 31639 56584 33332 56648
rect 16717 56579 33332 56584
rect 16717 56573 28901 56579
rect 16717 56568 20907 56573
rect 16717 56504 17431 56568
rect 17495 56504 18519 56568
rect 18583 56504 19607 56568
rect 19671 56504 20695 56568
rect 20759 56504 20907 56568
rect 16717 56488 20907 56504
rect 16717 56424 17431 56488
rect 17495 56424 18519 56488
rect 18583 56424 19607 56488
rect 19671 56424 20695 56488
rect 20759 56424 20907 56488
rect 16717 56408 20907 56424
rect 16717 56344 17431 56408
rect 17495 56344 18519 56408
rect 18583 56344 19607 56408
rect 19671 56344 20695 56408
rect 20759 56344 20907 56408
rect 16717 56337 20907 56344
rect 21143 56568 28901 56573
rect 21143 56504 21783 56568
rect 21847 56504 22871 56568
rect 22935 56504 23959 56568
rect 24023 56504 25047 56568
rect 25111 56504 26135 56568
rect 26199 56504 27223 56568
rect 27287 56504 28311 56568
rect 28375 56504 28901 56568
rect 21143 56488 28901 56504
rect 21143 56424 21783 56488
rect 21847 56424 22871 56488
rect 22935 56424 23959 56488
rect 24023 56424 25047 56488
rect 25111 56424 26135 56488
rect 26199 56424 27223 56488
rect 27287 56424 28311 56488
rect 28375 56424 28901 56488
rect 21143 56408 28901 56424
rect 21143 56344 21783 56408
rect 21847 56344 22871 56408
rect 22935 56344 23959 56408
rect 24023 56344 25047 56408
rect 25111 56344 26135 56408
rect 26199 56344 27223 56408
rect 27287 56344 28311 56408
rect 28375 56344 28901 56408
rect 21143 56343 28901 56344
rect 29137 56568 33332 56579
rect 29137 56504 29399 56568
rect 29463 56504 30487 56568
rect 30551 56504 31575 56568
rect 31639 56504 33332 56568
rect 29137 56488 33332 56504
rect 29137 56424 29399 56488
rect 29463 56424 30487 56488
rect 30551 56424 31575 56488
rect 31639 56424 33332 56488
rect 29137 56408 33332 56424
rect 29137 56344 29399 56408
rect 29463 56344 30487 56408
rect 30551 56344 31575 56408
rect 31639 56344 33332 56408
rect 29137 56343 33332 56344
rect 21143 56337 33332 56343
rect 16717 56328 33332 56337
rect 16717 56264 17431 56328
rect 17495 56264 18519 56328
rect 18583 56264 19607 56328
rect 19671 56264 20695 56328
rect 20759 56264 21783 56328
rect 21847 56264 22871 56328
rect 22935 56264 23959 56328
rect 24023 56264 25047 56328
rect 25111 56264 26135 56328
rect 26199 56264 27223 56328
rect 27287 56264 28311 56328
rect 28375 56264 29399 56328
rect 29463 56264 30487 56328
rect 30551 56264 31575 56328
rect 31639 56264 33332 56328
rect 16717 56248 33332 56264
rect 16717 56184 17431 56248
rect 17495 56184 18519 56248
rect 18583 56184 19607 56248
rect 19671 56184 20695 56248
rect 20759 56184 21783 56248
rect 21847 56184 22871 56248
rect 22935 56184 23959 56248
rect 24023 56184 25047 56248
rect 25111 56184 26135 56248
rect 26199 56184 27223 56248
rect 27287 56184 28311 56248
rect 28375 56184 29399 56248
rect 29463 56184 30487 56248
rect 30551 56184 31575 56248
rect 31639 56184 33332 56248
rect 16717 56147 33332 56184
rect 16715 54725 33227 54767
rect 16715 54661 17976 54725
rect 18040 54661 19064 54725
rect 19128 54661 20152 54725
rect 20216 54661 21240 54725
rect 21304 54661 22328 54725
rect 22392 54661 23416 54725
rect 23480 54661 24504 54725
rect 24568 54661 25592 54725
rect 25656 54661 26680 54725
rect 26744 54661 27768 54725
rect 27832 54661 28856 54725
rect 28920 54661 29944 54725
rect 30008 54661 31032 54725
rect 31096 54717 33227 54725
rect 31096 54661 33290 54717
rect 16715 54645 33290 54661
rect 16715 54582 17976 54645
rect 16715 54346 16910 54582
rect 17146 54581 17976 54582
rect 18040 54581 19064 54645
rect 19128 54581 20152 54645
rect 20216 54581 21240 54645
rect 21304 54581 22328 54645
rect 22392 54581 23416 54645
rect 23480 54581 24504 54645
rect 24568 54581 25592 54645
rect 25656 54581 26680 54645
rect 26744 54581 27768 54645
rect 27832 54581 28856 54645
rect 28920 54581 29944 54645
rect 30008 54581 31032 54645
rect 31096 54581 33290 54645
rect 17146 54575 33290 54581
rect 17146 54565 24906 54575
rect 17146 54501 17976 54565
rect 18040 54501 19064 54565
rect 19128 54501 20152 54565
rect 20216 54501 21240 54565
rect 21304 54501 22328 54565
rect 22392 54501 23416 54565
rect 23480 54501 24504 54565
rect 24568 54501 24906 54565
rect 17146 54485 24906 54501
rect 17146 54421 17976 54485
rect 18040 54421 19064 54485
rect 19128 54421 20152 54485
rect 20216 54421 21240 54485
rect 21304 54421 22328 54485
rect 22392 54421 23416 54485
rect 23480 54421 24504 54485
rect 24568 54421 24906 54485
rect 17146 54405 24906 54421
rect 17146 54346 17976 54405
rect 16715 54341 17976 54346
rect 18040 54341 19064 54405
rect 19128 54341 20152 54405
rect 20216 54341 21240 54405
rect 21304 54341 22328 54405
rect 22392 54341 23416 54405
rect 23480 54341 24504 54405
rect 24568 54341 24906 54405
rect 16715 54339 24906 54341
rect 25142 54571 33290 54575
rect 25142 54565 32909 54571
rect 25142 54501 25592 54565
rect 25656 54501 26680 54565
rect 26744 54501 27768 54565
rect 27832 54501 28856 54565
rect 28920 54501 29944 54565
rect 30008 54501 31032 54565
rect 31096 54501 32909 54565
rect 25142 54485 32909 54501
rect 25142 54421 25592 54485
rect 25656 54421 26680 54485
rect 26744 54421 27768 54485
rect 27832 54421 28856 54485
rect 28920 54421 29944 54485
rect 30008 54421 31032 54485
rect 31096 54421 32909 54485
rect 25142 54405 32909 54421
rect 25142 54341 25592 54405
rect 25656 54341 26680 54405
rect 26744 54341 27768 54405
rect 27832 54341 28856 54405
rect 28920 54341 29944 54405
rect 30008 54341 31032 54405
rect 31096 54341 32909 54405
rect 25142 54339 32909 54341
rect 16715 54335 32909 54339
rect 33145 54335 33290 54571
rect 16715 54325 33290 54335
rect 16715 54261 17976 54325
rect 18040 54261 19064 54325
rect 19128 54261 20152 54325
rect 20216 54261 21240 54325
rect 21304 54261 22328 54325
rect 22392 54261 23416 54325
rect 23480 54261 24504 54325
rect 24568 54261 25592 54325
rect 25656 54261 26680 54325
rect 26744 54261 27768 54325
rect 27832 54261 28856 54325
rect 28920 54261 29944 54325
rect 30008 54261 31032 54325
rect 31096 54261 33290 54325
rect 16715 54245 33290 54261
rect 16715 54181 17976 54245
rect 18040 54181 19064 54245
rect 19128 54181 20152 54245
rect 20216 54181 21240 54245
rect 21304 54181 22328 54245
rect 22392 54181 23416 54245
rect 23480 54181 24504 54245
rect 24568 54181 25592 54245
rect 25656 54181 26680 54245
rect 26744 54181 27768 54245
rect 27832 54181 28856 54245
rect 28920 54181 29944 54245
rect 30008 54181 31032 54245
rect 31096 54189 33290 54245
rect 31096 54181 33227 54189
rect 16715 54147 33227 54181
rect 16717 52728 33332 52767
rect 16717 52664 17431 52728
rect 17495 52664 18519 52728
rect 18583 52664 19607 52728
rect 19671 52664 20695 52728
rect 20759 52664 21783 52728
rect 21847 52664 22871 52728
rect 22935 52664 23959 52728
rect 24023 52664 25047 52728
rect 25111 52664 26135 52728
rect 26199 52664 27223 52728
rect 27287 52664 28311 52728
rect 28375 52664 29399 52728
rect 29463 52664 30487 52728
rect 30551 52664 31575 52728
rect 31639 52664 33332 52728
rect 16717 52648 33332 52664
rect 16717 52584 17431 52648
rect 17495 52584 18519 52648
rect 18583 52584 19607 52648
rect 19671 52584 20695 52648
rect 20759 52584 21783 52648
rect 21847 52584 22871 52648
rect 22935 52584 23959 52648
rect 24023 52584 25047 52648
rect 25111 52584 26135 52648
rect 26199 52584 27223 52648
rect 27287 52584 28311 52648
rect 28375 52584 29399 52648
rect 29463 52584 30487 52648
rect 30551 52584 31575 52648
rect 31639 52584 33332 52648
rect 16717 52579 33332 52584
rect 16717 52573 28901 52579
rect 16717 52568 20907 52573
rect 16717 52504 17431 52568
rect 17495 52504 18519 52568
rect 18583 52504 19607 52568
rect 19671 52504 20695 52568
rect 20759 52504 20907 52568
rect 16717 52488 20907 52504
rect 16717 52424 17431 52488
rect 17495 52424 18519 52488
rect 18583 52424 19607 52488
rect 19671 52424 20695 52488
rect 20759 52424 20907 52488
rect 16717 52408 20907 52424
rect 16717 52344 17431 52408
rect 17495 52344 18519 52408
rect 18583 52344 19607 52408
rect 19671 52344 20695 52408
rect 20759 52344 20907 52408
rect 16717 52337 20907 52344
rect 21143 52568 28901 52573
rect 21143 52504 21783 52568
rect 21847 52504 22871 52568
rect 22935 52504 23959 52568
rect 24023 52504 25047 52568
rect 25111 52504 26135 52568
rect 26199 52504 27223 52568
rect 27287 52504 28311 52568
rect 28375 52504 28901 52568
rect 21143 52488 28901 52504
rect 21143 52424 21783 52488
rect 21847 52424 22871 52488
rect 22935 52424 23959 52488
rect 24023 52424 25047 52488
rect 25111 52424 26135 52488
rect 26199 52424 27223 52488
rect 27287 52424 28311 52488
rect 28375 52424 28901 52488
rect 21143 52408 28901 52424
rect 21143 52344 21783 52408
rect 21847 52344 22871 52408
rect 22935 52344 23959 52408
rect 24023 52344 25047 52408
rect 25111 52344 26135 52408
rect 26199 52344 27223 52408
rect 27287 52344 28311 52408
rect 28375 52344 28901 52408
rect 21143 52343 28901 52344
rect 29137 52568 33332 52579
rect 29137 52504 29399 52568
rect 29463 52504 30487 52568
rect 30551 52504 31575 52568
rect 31639 52504 33332 52568
rect 29137 52488 33332 52504
rect 29137 52424 29399 52488
rect 29463 52424 30487 52488
rect 30551 52424 31575 52488
rect 31639 52424 33332 52488
rect 29137 52408 33332 52424
rect 29137 52344 29399 52408
rect 29463 52344 30487 52408
rect 30551 52344 31575 52408
rect 31639 52344 33332 52408
rect 29137 52343 33332 52344
rect 21143 52337 33332 52343
rect 16717 52328 33332 52337
rect 16717 52264 17431 52328
rect 17495 52264 18519 52328
rect 18583 52264 19607 52328
rect 19671 52264 20695 52328
rect 20759 52264 21783 52328
rect 21847 52264 22871 52328
rect 22935 52264 23959 52328
rect 24023 52264 25047 52328
rect 25111 52264 26135 52328
rect 26199 52264 27223 52328
rect 27287 52264 28311 52328
rect 28375 52264 29399 52328
rect 29463 52264 30487 52328
rect 30551 52264 31575 52328
rect 31639 52264 33332 52328
rect 16717 52248 33332 52264
rect 16717 52184 17431 52248
rect 17495 52184 18519 52248
rect 18583 52184 19607 52248
rect 19671 52184 20695 52248
rect 20759 52184 21783 52248
rect 21847 52184 22871 52248
rect 22935 52184 23959 52248
rect 24023 52184 25047 52248
rect 25111 52184 26135 52248
rect 26199 52184 27223 52248
rect 27287 52184 28311 52248
rect 28375 52184 29399 52248
rect 29463 52184 30487 52248
rect 30551 52184 31575 52248
rect 31639 52184 33332 52248
rect 16717 52147 33332 52184
rect 16715 50725 33227 50767
rect 16715 50661 17976 50725
rect 18040 50661 20152 50725
rect 20216 50661 21240 50725
rect 21304 50661 23416 50725
rect 23480 50661 24504 50725
rect 24568 50661 25592 50725
rect 25656 50661 27768 50725
rect 27832 50661 28856 50725
rect 28920 50661 31032 50725
rect 31096 50717 33227 50725
rect 31096 50661 33290 50717
rect 16715 50645 33290 50661
rect 16715 50582 17976 50645
rect 16715 50346 16910 50582
rect 17146 50581 17976 50582
rect 18040 50581 20152 50645
rect 20216 50581 21240 50645
rect 21304 50581 23416 50645
rect 23480 50581 24504 50645
rect 24568 50581 25592 50645
rect 25656 50581 27768 50645
rect 27832 50581 28856 50645
rect 28920 50581 31032 50645
rect 31096 50581 33290 50645
rect 17146 50575 33290 50581
rect 17146 50565 24906 50575
rect 17146 50501 17976 50565
rect 18040 50501 20152 50565
rect 20216 50501 21240 50565
rect 21304 50501 23416 50565
rect 23480 50501 24504 50565
rect 24568 50501 24906 50565
rect 17146 50485 24906 50501
rect 17146 50421 17976 50485
rect 18040 50421 20152 50485
rect 20216 50421 21240 50485
rect 21304 50421 23416 50485
rect 23480 50421 24504 50485
rect 24568 50421 24906 50485
rect 17146 50405 24906 50421
rect 17146 50346 17976 50405
rect 16715 50341 17976 50346
rect 18040 50341 20152 50405
rect 20216 50341 21240 50405
rect 21304 50341 23416 50405
rect 23480 50341 24504 50405
rect 24568 50341 24906 50405
rect 16715 50339 24906 50341
rect 25142 50571 33290 50575
rect 25142 50565 32909 50571
rect 25142 50501 25592 50565
rect 25656 50501 27768 50565
rect 27832 50501 28856 50565
rect 28920 50501 31032 50565
rect 31096 50501 32909 50565
rect 25142 50485 32909 50501
rect 25142 50421 25592 50485
rect 25656 50421 27768 50485
rect 27832 50421 28856 50485
rect 28920 50421 31032 50485
rect 31096 50421 32909 50485
rect 25142 50405 32909 50421
rect 25142 50341 25592 50405
rect 25656 50341 27768 50405
rect 27832 50341 28856 50405
rect 28920 50341 31032 50405
rect 31096 50341 32909 50405
rect 25142 50339 32909 50341
rect 16715 50335 32909 50339
rect 33145 50335 33290 50571
rect 16715 50325 33290 50335
rect 16715 50261 17976 50325
rect 18040 50261 20152 50325
rect 20216 50261 21240 50325
rect 21304 50261 23416 50325
rect 23480 50261 24504 50325
rect 24568 50261 25592 50325
rect 25656 50261 27768 50325
rect 27832 50261 28856 50325
rect 28920 50261 31032 50325
rect 31096 50261 33290 50325
rect 16715 50245 33290 50261
rect 16715 50181 17976 50245
rect 18040 50181 20152 50245
rect 20216 50181 21240 50245
rect 21304 50181 23416 50245
rect 23480 50181 24504 50245
rect 24568 50181 25592 50245
rect 25656 50181 27768 50245
rect 27832 50181 28856 50245
rect 28920 50181 31032 50245
rect 31096 50189 33290 50245
rect 31096 50181 33227 50189
rect 16715 50147 33227 50181
rect 16717 48728 33332 48767
rect 16717 48664 17431 48728
rect 17495 48664 18519 48728
rect 18583 48664 19607 48728
rect 19671 48664 20695 48728
rect 20759 48664 21783 48728
rect 21847 48664 22871 48728
rect 22935 48664 23959 48728
rect 24023 48664 29399 48728
rect 29463 48664 30487 48728
rect 30551 48664 31575 48728
rect 31639 48664 33332 48728
rect 16717 48648 33332 48664
rect 16717 48584 17431 48648
rect 17495 48584 18519 48648
rect 18583 48584 19607 48648
rect 19671 48584 20695 48648
rect 20759 48584 21783 48648
rect 21847 48584 22871 48648
rect 22935 48584 23959 48648
rect 24023 48584 29399 48648
rect 29463 48584 30487 48648
rect 30551 48584 31575 48648
rect 31639 48584 33332 48648
rect 16717 48579 33332 48584
rect 16717 48573 28901 48579
rect 16717 48568 20907 48573
rect 16717 48504 17431 48568
rect 17495 48504 18519 48568
rect 18583 48504 19607 48568
rect 19671 48504 20695 48568
rect 20759 48504 20907 48568
rect 16717 48488 20907 48504
rect 16717 48424 17431 48488
rect 17495 48424 18519 48488
rect 18583 48424 19607 48488
rect 19671 48424 20695 48488
rect 20759 48424 20907 48488
rect 16717 48408 20907 48424
rect 16717 48344 17431 48408
rect 17495 48344 18519 48408
rect 18583 48344 19607 48408
rect 19671 48344 20695 48408
rect 20759 48344 20907 48408
rect 16717 48337 20907 48344
rect 21143 48568 28901 48573
rect 21143 48504 21783 48568
rect 21847 48504 22871 48568
rect 22935 48504 23959 48568
rect 24023 48504 28901 48568
rect 21143 48488 28901 48504
rect 21143 48424 21783 48488
rect 21847 48424 22871 48488
rect 22935 48424 23959 48488
rect 24023 48424 28901 48488
rect 21143 48408 28901 48424
rect 21143 48344 21783 48408
rect 21847 48344 22871 48408
rect 22935 48344 23959 48408
rect 24023 48344 28901 48408
rect 21143 48343 28901 48344
rect 29137 48568 33332 48579
rect 29137 48504 29399 48568
rect 29463 48504 30487 48568
rect 30551 48504 31575 48568
rect 31639 48504 33332 48568
rect 29137 48488 33332 48504
rect 29137 48424 29399 48488
rect 29463 48424 30487 48488
rect 30551 48424 31575 48488
rect 31639 48424 33332 48488
rect 29137 48408 33332 48424
rect 29137 48344 29399 48408
rect 29463 48344 30487 48408
rect 30551 48344 31575 48408
rect 31639 48344 33332 48408
rect 29137 48343 33332 48344
rect 21143 48337 33332 48343
rect 16717 48328 33332 48337
rect 16717 48264 17431 48328
rect 17495 48264 18519 48328
rect 18583 48264 19607 48328
rect 19671 48264 20695 48328
rect 20759 48264 21783 48328
rect 21847 48264 22871 48328
rect 22935 48264 23959 48328
rect 24023 48264 29399 48328
rect 29463 48264 30487 48328
rect 30551 48264 31575 48328
rect 31639 48264 33332 48328
rect 16717 48248 33332 48264
rect 16717 48184 17431 48248
rect 17495 48184 18519 48248
rect 18583 48184 19607 48248
rect 19671 48184 20695 48248
rect 20759 48184 21783 48248
rect 21847 48184 22871 48248
rect 22935 48184 23959 48248
rect 24023 48184 29399 48248
rect 29463 48184 30487 48248
rect 30551 48184 31575 48248
rect 31639 48184 33332 48248
rect 16717 48147 33332 48184
rect 10176 47616 10552 47634
rect -6412 47256 -6346 47257
rect -6412 47192 -6411 47256
rect -6347 47192 12030 47256
rect -6412 47191 -6346 47192
rect -6412 46633 -6346 46634
rect -6412 46569 -6411 46633
rect -6347 46569 11411 46633
rect -6412 46568 -6346 46569
rect -5972 46238 -5674 46319
rect -5972 39854 -5895 46238
rect -5751 45377 -5674 46238
rect 10179 46109 10552 46129
rect 330 45833 619 45964
rect -5751 45079 -5652 45377
rect -5751 44658 -5674 45079
rect -5751 44601 -2659 44658
rect -5751 44365 -3094 44601
rect -2858 44365 -2659 44601
rect -5751 44318 -2659 44365
rect 330 44329 379 45833
rect 523 44544 619 45833
rect 10179 44544 10213 46109
rect 523 44512 1372 44544
rect 523 44329 899 44512
rect -5751 39891 -5674 44318
rect 330 44276 899 44329
rect 1135 44276 1372 44512
rect 330 44255 1372 44276
rect 10087 44255 10213 44544
rect 10179 43238 10213 44255
rect 8760 43236 10213 43238
rect 8760 43000 8907 43236
rect 9143 43000 10213 43236
rect 8760 42998 10213 43000
rect 325 41371 565 41411
rect -5751 39884 -135 39891
rect -5751 39854 -3086 39884
rect -5972 39828 -3086 39854
rect -2850 39828 -135 39884
rect -5972 39748 -5668 39828
rect -5713 39684 -5668 39748
rect -164 39684 -135 39828
rect 325 39867 360 41371
rect 504 40868 565 41371
rect 762 40868 1292 40869
rect 504 40867 1292 40868
rect 504 40631 909 40867
rect 1145 40631 1292 40867
rect 504 40629 1292 40631
rect 504 40628 928 40629
rect 504 39867 565 40628
rect 325 39810 565 39867
rect 10179 39885 10213 42998
rect 10517 39885 10552 46109
rect 10179 39866 10552 39885
rect -5713 39648 -3086 39684
rect -2850 39648 -135 39684
rect -5713 39636 -135 39648
rect 756 39438 1286 39440
rect 756 39202 903 39438
rect 1139 39350 1286 39438
rect 1139 39286 2638 39350
rect 1139 39202 1286 39286
rect 756 39200 1286 39202
rect 2512 38873 2638 39286
rect 2512 38809 2522 38873
rect 2586 38809 2638 38873
rect 2512 38793 2638 38809
rect -4714 38790 -4648 38791
rect -4714 38726 -4713 38790
rect -4649 38726 -4648 38790
rect -4714 38725 -4648 38726
rect 2512 38729 2522 38793
rect 2586 38729 2638 38793
rect -7723 37899 -7657 37900
rect -7723 37835 -7722 37899
rect -7658 37835 -7657 37899
rect -7723 37834 -7657 37835
rect -8481 37371 -8415 37372
rect -8481 37307 -8480 37371
rect -8416 37307 -8415 37371
rect -8481 37306 -8415 37307
rect -9209 35941 -9143 35942
rect -9209 35877 -9208 35941
rect -9144 35877 -9143 35941
rect -9209 35876 -9143 35877
rect -10070 35351 -10004 35352
rect -10070 35287 -10069 35351
rect -10005 35287 -10004 35351
rect -10070 35286 -10004 35287
rect -13396 34676 -13330 34677
rect -13396 34612 -13395 34676
rect -13331 34612 -13330 34676
rect -13396 34611 -13330 34612
rect -4713 34196 -4649 38725
rect 2512 38713 2638 38729
rect 2512 38649 2522 38713
rect 2586 38649 2638 38713
rect 2512 38632 2638 38649
rect -4124 38447 -4058 38448
rect -4124 38383 -4123 38447
rect -4059 38383 -4058 38447
rect -4124 38382 -4058 38383
rect 2514 38400 2640 38422
rect -4714 34195 -4648 34196
rect -4714 34131 -4713 34195
rect -4649 34131 -4648 34195
rect -4714 34130 -4648 34131
rect -4123 33851 -4059 38382
rect 2514 38336 2532 38400
rect 2596 38336 2640 38400
rect 2514 38320 2640 38336
rect 2514 38256 2532 38320
rect 2596 38256 2640 38320
rect 2514 38240 2640 38256
rect 2514 38176 2532 38240
rect 2596 38176 2640 38240
rect 2514 38160 2640 38176
rect 2514 38096 2532 38160
rect 2596 38096 2640 38160
rect 2514 38080 2640 38096
rect 2514 38016 2532 38080
rect 2596 38016 2640 38080
rect 2514 37971 2640 38016
rect 4761 38051 5291 38053
rect 4761 37971 4908 38051
rect 2514 37907 4908 37971
rect -2398 37900 -2334 37901
rect -2399 37899 -2333 37900
rect -761 37899 -695 37900
rect 1472 37899 1538 37900
rect -2399 37835 -2398 37899
rect -2334 37835 -2333 37899
rect -777 37835 -760 37899
rect -696 37835 1473 37899
rect 1537 37835 1569 37899
rect 2514 37875 2614 37907
rect -2399 37834 -2333 37835
rect -761 37834 -695 37835
rect 1472 37834 1538 37835
rect -2815 37372 -2751 37375
rect -2816 37371 -2750 37372
rect -2816 37307 -2815 37371
rect -2751 37307 -2750 37371
rect -2816 37306 -2750 37307
rect -4124 33850 -4058 33851
rect -4124 33786 -4123 33850
rect -4059 33786 -4058 33850
rect -4124 33785 -4058 33786
rect -15140 33179 -15074 33180
rect -15140 33115 -15139 33179
rect -15075 33115 -15074 33179
rect -15140 33114 -15074 33115
rect -27162 32800 -27077 32864
rect -27013 32800 -26922 32864
rect -27162 32784 -26922 32800
rect -27162 32720 -27077 32784
rect -27013 32767 -26922 32784
rect -27013 32765 -26704 32767
rect -27162 32704 -27051 32720
rect -27162 32640 -27077 32704
rect -27162 32624 -27051 32640
rect -27162 32560 -27077 32624
rect -27162 32544 -27051 32560
rect -27162 32480 -27077 32544
rect -26815 32529 -26704 32765
rect -27013 32527 -26704 32529
rect -27013 32480 -26922 32527
rect -27162 32464 -26922 32480
rect -27162 32400 -27077 32464
rect -27013 32400 -26922 32464
rect -27162 32329 -26922 32400
rect -3919 29752 -3853 29753
rect -3919 29688 -3918 29752
rect -3854 29688 -3853 29752
rect -3919 29687 -3853 29688
rect -5279 29330 -5215 29332
rect -5280 29329 -5214 29330
rect -5280 29265 -5279 29329
rect -5215 29265 -5214 29329
rect -5280 29264 -5214 29265
rect -15741 28708 -15500 28709
rect -19238 28706 -15500 28708
rect -19238 28470 -19091 28706
rect -18855 28470 -15500 28706
rect -19238 28468 -15500 28470
rect -17700 27612 -17460 28468
rect -15741 28063 -15500 28468
rect -15741 27999 -15695 28063
rect -15631 27999 -15500 28063
rect -15741 27983 -15500 27999
rect -15741 27919 -15695 27983
rect -15631 27919 -15500 27983
rect -15741 27903 -15500 27919
rect -15741 27839 -15695 27903
rect -15631 27839 -15500 27903
rect -15741 27823 -15500 27839
rect -15741 27759 -15695 27823
rect -15631 27759 -15500 27823
rect -15741 27743 -15500 27759
rect -15741 27679 -15695 27743
rect -15631 27679 -15500 27743
rect -15741 27619 -15500 27679
rect -12394 28065 -12266 28089
rect -12394 28001 -12385 28065
rect -12321 28003 -12266 28065
rect -11237 28053 -10707 28055
rect -11237 28003 -11090 28053
rect -12321 28001 -11090 28003
rect -12394 27985 -11090 28001
rect -12394 27921 -12385 27985
rect -12321 27921 -11090 27985
rect -12394 27905 -11090 27921
rect -12394 27841 -12385 27905
rect -12321 27875 -11090 27905
rect -12321 27841 -12266 27875
rect -12394 27825 -12266 27841
rect -12394 27761 -12385 27825
rect -12321 27761 -12266 27825
rect -12394 27745 -12266 27761
rect -12394 27681 -12385 27745
rect -12321 27681 -12266 27745
rect -12394 27658 -12266 27681
rect -17700 27548 -17603 27612
rect -17539 27548 -17460 27612
rect -17700 27461 -17460 27548
rect -15234 27441 -14704 27443
rect -15234 27205 -15087 27441
rect -14851 27388 -14704 27441
rect -12386 27428 -12258 27461
rect -12395 27424 -12258 27428
rect -12395 27388 -12378 27424
rect -14851 27360 -12378 27388
rect -12314 27388 -12258 27424
rect -12314 27360 -12247 27388
rect -14851 27344 -12247 27360
rect -14851 27280 -12378 27344
rect -12314 27280 -12247 27344
rect -14851 27264 -12247 27280
rect -14851 27260 -12378 27264
rect -14851 27205 -14704 27260
rect -15234 27203 -14704 27205
rect -12395 27200 -12378 27260
rect -12314 27260 -12247 27264
rect -12314 27200 -12258 27260
rect -12395 27197 -12258 27200
rect -12386 27188 -12258 27197
rect -35224 26906 -34761 26908
rect -35224 26670 -35111 26906
rect -34875 26670 -34761 26906
rect -35224 26612 -34761 26670
rect -38191 26594 -34761 26612
rect -38191 26530 -38155 26594
rect -38091 26530 -38075 26594
rect -38011 26530 -37995 26594
rect -37931 26530 -37915 26594
rect -37851 26530 -37835 26594
rect -37771 26530 -37755 26594
rect -37691 26530 -37675 26594
rect -37611 26530 -37595 26594
rect -37531 26530 -37515 26594
rect -37451 26530 -37435 26594
rect -37371 26530 -37355 26594
rect -37291 26530 -37275 26594
rect -37211 26530 -37195 26594
rect -37131 26530 -37115 26594
rect -37051 26530 -37035 26594
rect -36971 26530 -36955 26594
rect -36891 26530 -36875 26594
rect -36811 26530 -36795 26594
rect -36731 26530 -36715 26594
rect -36651 26530 -36635 26594
rect -36571 26530 -36555 26594
rect -36491 26530 -36475 26594
rect -36411 26530 -36395 26594
rect -36331 26530 -36315 26594
rect -36251 26530 -36235 26594
rect -36171 26530 -36155 26594
rect -36091 26530 -36075 26594
rect -36011 26530 -35995 26594
rect -35931 26530 -35915 26594
rect -35851 26530 -35835 26594
rect -35771 26530 -35755 26594
rect -35691 26530 -35675 26594
rect -35611 26530 -35595 26594
rect -35531 26530 -35515 26594
rect -35451 26530 -35435 26594
rect -35371 26530 -35355 26594
rect -35291 26530 -35275 26594
rect -35211 26530 -35195 26594
rect -35131 26530 -35115 26594
rect -35051 26530 -35035 26594
rect -34971 26530 -34955 26594
rect -34891 26530 -34761 26594
rect -38191 26514 -34761 26530
rect -38191 26513 -34855 26514
rect -12422 26463 -12294 26493
rect -17691 26383 -17458 26461
rect -17691 26319 -17603 26383
rect -17539 26319 -17458 26383
rect -12422 26399 -12381 26463
rect -12317 26399 -12294 26463
rect -12422 26383 -12294 26399
rect -17691 25810 -17458 26319
rect -15742 26274 -15509 26354
rect -15742 26210 -15713 26274
rect -15649 26210 -15509 26274
rect -15742 26194 -15509 26210
rect -15742 26130 -15713 26194
rect -15649 26130 -15509 26194
rect -15742 26114 -15509 26130
rect -15742 26050 -15713 26114
rect -15649 26050 -15509 26114
rect -12422 26319 -12381 26383
rect -12317 26330 -12294 26383
rect -11717 26330 -11589 27875
rect -11237 27817 -11090 27875
rect -10854 27817 -10707 28053
rect -11237 27815 -10707 27817
rect -5279 27533 -5215 29264
rect -5280 27532 -5214 27533
rect -5280 27468 -5279 27532
rect -5215 27468 -5214 27532
rect -5280 27467 -5214 27468
rect -12317 26319 -11589 26330
rect -12422 26303 -11589 26319
rect -12422 26239 -12381 26303
rect -12317 26239 -11589 26303
rect -12422 26223 -11589 26239
rect -12422 26159 -12381 26223
rect -12317 26202 -11589 26223
rect -12317 26159 -12294 26202
rect -12422 26143 -12294 26159
rect -12422 26079 -12381 26143
rect -12317 26079 -12294 26143
rect -12422 26053 -12294 26079
rect -15742 25810 -15509 26050
rect -15238 25816 -14708 25818
rect -15238 25810 -15091 25816
rect -19246 25808 -18716 25810
rect -19246 25572 -19099 25808
rect -18863 25799 -18716 25808
rect -18860 25575 -18716 25799
rect -18863 25572 -18716 25575
rect -19246 25570 -18716 25572
rect -17691 25580 -15091 25810
rect -14855 25765 -14708 25816
rect -12383 25765 -12255 25856
rect -14855 25637 -12255 25765
rect -14855 25580 -14708 25637
rect -12383 25595 -12255 25637
rect -17691 25578 -14708 25580
rect -17691 25577 -14847 25578
rect -27228 25512 -26698 25514
rect -27228 25276 -27081 25512
rect -26845 25433 -26698 25512
rect -25450 25480 -25368 25483
rect -25450 25433 -25441 25480
rect -26845 25416 -25441 25433
rect -25377 25433 -25368 25480
rect -25377 25416 -25316 25433
rect -26845 25400 -25316 25416
rect -26845 25336 -25441 25400
rect -25377 25336 -25316 25400
rect -26845 25320 -25316 25336
rect -26845 25305 -25441 25320
rect -26845 25276 -26698 25305
rect -27228 25274 -26698 25276
rect -25450 25256 -25441 25305
rect -25377 25305 -25316 25320
rect -25377 25256 -25368 25305
rect -25450 25240 -25368 25256
rect -25450 25176 -25441 25240
rect -25377 25176 -25368 25240
rect -25450 25174 -25368 25176
rect -17691 24970 -17458 25577
rect -11717 25313 -11589 26202
rect -11324 25665 -11260 25666
rect -11325 25664 -11259 25665
rect -11325 25600 -11324 25664
rect -11260 25600 -11259 25664
rect -11325 25599 -11259 25600
rect -25453 24941 -25364 24946
rect -25453 24877 -25441 24941
rect -25377 24893 -25364 24941
rect -23236 24915 -22706 24917
rect -23236 24893 -23089 24915
rect -25377 24877 -23089 24893
rect -25453 24861 -23089 24877
rect -25453 24797 -25441 24861
rect -25377 24797 -23089 24861
rect -25453 24781 -23089 24797
rect -25453 24717 -25441 24781
rect -25377 24765 -23089 24781
rect -25377 24717 -25364 24765
rect -25453 24713 -25364 24717
rect -23236 24679 -23089 24765
rect -22853 24679 -22706 24915
rect -17691 24906 -17603 24970
rect -17539 24906 -17458 24970
rect -17691 24811 -17458 24906
rect -12398 25185 -11589 25313
rect -23236 24677 -22706 24679
rect -12398 24697 -12270 25185
rect -11978 24872 -11912 24873
rect -11978 24808 -11977 24872
rect -11913 24808 -11912 24872
rect -11978 24807 -11912 24808
rect -12398 24633 -12393 24697
rect -12329 24633 -12270 24697
rect -12398 24617 -12270 24633
rect -12398 24553 -12393 24617
rect -12329 24553 -12270 24617
rect -12398 24537 -12270 24553
rect -12398 24473 -12393 24537
rect -12329 24473 -12270 24537
rect -12398 24441 -12270 24473
rect -12434 24233 -12306 24264
rect -12434 24169 -12389 24233
rect -12325 24169 -12306 24233
rect -12434 24153 -12306 24169
rect -12434 24089 -12389 24153
rect -12325 24089 -12306 24153
rect -12434 24073 -12306 24089
rect -12434 24009 -12389 24073
rect -12325 24009 -12306 24073
rect -17692 23741 -17452 23854
rect -17692 23731 -17603 23741
rect -18811 23730 -17603 23731
rect -19239 23728 -17603 23730
rect -39205 23712 -38742 23714
rect -39205 23476 -39092 23712
rect -38856 23710 -38742 23712
rect -38856 23586 -34770 23710
rect -38856 23522 -38149 23586
rect -38085 23522 -38069 23586
rect -38005 23522 -37989 23586
rect -37925 23522 -37909 23586
rect -37845 23522 -37829 23586
rect -37765 23522 -37749 23586
rect -37685 23522 -37669 23586
rect -37605 23522 -37589 23586
rect -37525 23522 -37509 23586
rect -37445 23522 -37429 23586
rect -37365 23522 -37349 23586
rect -37285 23522 -37269 23586
rect -37205 23522 -37189 23586
rect -37125 23522 -37109 23586
rect -37045 23522 -37029 23586
rect -36965 23522 -36949 23586
rect -36885 23522 -36869 23586
rect -36805 23522 -36789 23586
rect -36725 23522 -36709 23586
rect -36645 23522 -36629 23586
rect -36565 23522 -36549 23586
rect -36485 23522 -36469 23586
rect -36405 23522 -36389 23586
rect -36325 23522 -36309 23586
rect -36245 23522 -36229 23586
rect -36165 23522 -36149 23586
rect -36085 23522 -36069 23586
rect -36005 23522 -35989 23586
rect -35925 23522 -35909 23586
rect -35845 23522 -35829 23586
rect -35765 23522 -35749 23586
rect -35685 23522 -35669 23586
rect -35605 23522 -35589 23586
rect -35525 23522 -35509 23586
rect -35445 23522 -35429 23586
rect -35365 23522 -35349 23586
rect -35285 23522 -35269 23586
rect -35205 23522 -35189 23586
rect -35125 23522 -35109 23586
rect -35045 23522 -35029 23586
rect -34965 23522 -34949 23586
rect -34885 23522 -34770 23586
rect -38856 23476 -34770 23522
rect -19239 23492 -19092 23728
rect -18856 23677 -17603 23728
rect -17539 23677 -17452 23741
rect -18856 23492 -17452 23677
rect -19239 23491 -17452 23492
rect -15726 23637 -15493 23639
rect -15237 23637 -14707 23639
rect -15726 23633 -15090 23637
rect -15726 23569 -15724 23633
rect -15660 23569 -15090 23633
rect -15726 23553 -15090 23569
rect -19239 23490 -18709 23491
rect -39205 23474 -34770 23476
rect -15726 23489 -15724 23553
rect -15660 23489 -15090 23553
rect -15726 23473 -15090 23489
rect -15726 23409 -15724 23473
rect -15660 23409 -15090 23473
rect -15726 23404 -15090 23409
rect -15237 23401 -15090 23404
rect -14854 23592 -14707 23637
rect -12434 23592 -12306 24009
rect -14854 23464 -12306 23592
rect -11977 23519 -11913 24807
rect -11324 23888 -11260 25599
rect -11325 23887 -11259 23888
rect -11325 23823 -11324 23887
rect -11260 23823 -11259 23887
rect -11325 23822 -11259 23823
rect -11978 23518 -11912 23519
rect -14854 23401 -14707 23464
rect -15237 23399 -14707 23401
rect -16600 22724 -16534 22725
rect -16600 22660 -16599 22724
rect -16535 22660 -16534 22724
rect -16600 22659 -16534 22660
rect -16599 20652 -16535 22659
rect -13885 22584 -13757 23464
rect -11978 23454 -11977 23518
rect -11913 23454 -11912 23518
rect -11978 23453 -11912 23454
rect -11977 23442 -11913 23453
rect -12390 23277 -12318 23278
rect -12390 23259 -12258 23277
rect -12390 23195 -12386 23259
rect -12322 23195 -12258 23259
rect -12390 23179 -12258 23195
rect -12390 23115 -12386 23179
rect -12322 23115 -12258 23179
rect -12390 23108 -12258 23115
rect -11246 23152 -10716 23154
rect -11246 23108 -11099 23152
rect -12390 23099 -11099 23108
rect -12390 23035 -12386 23099
rect -12322 23035 -11099 23099
rect -12390 23019 -11099 23035
rect -12390 22955 -12386 23019
rect -12322 22980 -11099 23019
rect -12322 22955 -12258 22980
rect -12390 22939 -12258 22955
rect -12390 22875 -12386 22939
rect -12322 22875 -12258 22939
rect -11246 22916 -11099 22980
rect -10863 22916 -10716 23152
rect -11246 22914 -10716 22916
rect -12390 22856 -12258 22875
rect -12386 22837 -12258 22856
rect -12400 22623 -12272 22651
rect -12400 22584 -12389 22623
rect -13885 22559 -12389 22584
rect -12325 22559 -12272 22623
rect -13885 22543 -12272 22559
rect -13885 22479 -12389 22543
rect -12325 22479 -12272 22543
rect -13885 22463 -12272 22479
rect -13885 22456 -12389 22463
rect -12400 22399 -12389 22456
rect -12325 22399 -12272 22463
rect -12400 22350 -12272 22399
rect -16600 20651 -16534 20652
rect -16600 20587 -16599 20651
rect -16535 20587 -16534 20651
rect -16600 20586 -16534 20587
rect -35218 19231 -34755 19233
rect -35218 19066 -35105 19231
rect -38169 19058 -35105 19066
rect -38169 18994 -38147 19058
rect -38083 18994 -38067 19058
rect -38003 18994 -37987 19058
rect -37923 18994 -37907 19058
rect -37843 18994 -37827 19058
rect -37763 18994 -37747 19058
rect -37683 18994 -37667 19058
rect -37603 18994 -37587 19058
rect -37523 18994 -37507 19058
rect -37443 18994 -37427 19058
rect -37363 18994 -37347 19058
rect -37283 18994 -37267 19058
rect -37203 18994 -37187 19058
rect -37123 18994 -37107 19058
rect -37043 18994 -37027 19058
rect -36963 18994 -36947 19058
rect -36883 18994 -36867 19058
rect -36803 18994 -36787 19058
rect -36723 18994 -36707 19058
rect -36643 18994 -36627 19058
rect -36563 18994 -36547 19058
rect -36483 18994 -36467 19058
rect -36403 18994 -36387 19058
rect -36323 18994 -36307 19058
rect -36243 18994 -36227 19058
rect -36163 18994 -36147 19058
rect -36083 18994 -36067 19058
rect -36003 18994 -35987 19058
rect -35923 18994 -35907 19058
rect -35843 18994 -35827 19058
rect -35763 18994 -35747 19058
rect -35683 18994 -35667 19058
rect -35603 18994 -35587 19058
rect -35523 18994 -35507 19058
rect -35443 18994 -35427 19058
rect -35363 18994 -35347 19058
rect -35283 18994 -35267 19058
rect -35203 18994 -35187 19058
rect -35123 18994 -35107 19058
rect -34869 18995 -34755 19231
rect -5279 19044 -5215 27467
rect -3918 26856 -3854 29687
rect -3919 26855 -3853 26856
rect -3919 26791 -3918 26855
rect -3854 26791 -3853 26855
rect -3919 26790 -3853 26791
rect -3918 19044 -3854 26790
rect -2815 19514 -2751 37306
rect -2816 19513 -2750 19514
rect -2816 19449 -2815 19513
rect -2751 19449 -2750 19513
rect -2816 19448 -2750 19449
rect -2398 19213 -2334 37834
rect 4761 37815 4908 37907
rect 5144 37815 5291 38051
rect 4761 37813 5291 37815
rect -761 37370 -695 37371
rect 1995 37370 2061 37371
rect -761 37306 -760 37370
rect -696 37306 1996 37370
rect 2060 37306 2094 37370
rect -761 37305 -695 37306
rect 1995 37305 2061 37306
rect 2167 37135 2233 37150
rect 757 37093 1287 37095
rect 757 36857 904 37093
rect 1140 36996 1287 37093
rect 2167 37071 2168 37135
rect 2232 37071 2233 37135
rect 2167 37055 2233 37071
rect 2167 36996 2168 37055
rect 1140 36991 2168 36996
rect 2232 36991 2233 37055
rect 1140 36975 2233 36991
rect 1140 36932 2168 36975
rect 1140 36857 1287 36932
rect 2167 36911 2168 36932
rect 2232 36911 2233 36975
rect 2167 36897 2233 36911
rect 757 36855 1287 36857
rect 2169 36669 2233 36680
rect 2168 36651 2234 36669
rect 2168 36587 2169 36651
rect 2233 36587 2234 36651
rect 2168 36571 2234 36587
rect 2168 36507 2169 36571
rect 2233 36567 2234 36571
rect 4768 36658 5298 36660
rect 4768 36567 4915 36658
rect 2233 36507 4915 36567
rect 2168 36503 4915 36507
rect 2168 36491 2234 36503
rect 2168 36427 2169 36491
rect 2233 36427 2234 36491
rect 2168 36411 2234 36427
rect 4768 36422 4915 36503
rect 5151 36422 5298 36658
rect 4768 36420 5298 36422
rect 2168 36347 2169 36411
rect 2233 36347 2234 36411
rect 2168 36331 2234 36347
rect 2168 36267 2169 36331
rect 2233 36267 2234 36331
rect 2168 36249 2234 36267
rect 3664 36095 3783 36115
rect 5179 36105 5243 36420
rect 3581 36094 3812 36095
rect 3581 36030 3584 36094
rect 3648 36030 3664 36094
rect 3728 36030 3744 36094
rect 3808 36030 3812 36094
rect 3581 36029 3812 36030
rect 5054 36093 5352 36105
rect 5629 36098 5748 36115
rect 5054 36029 5091 36093
rect 5155 36029 5171 36093
rect 5235 36029 5251 36093
rect 5315 36029 5352 36093
rect 774 36014 1304 36016
rect 774 35778 921 36014
rect 1157 35957 1304 36014
rect 3664 35957 3783 36029
rect 5054 36017 5352 36029
rect 5573 36094 5802 36098
rect 5573 36030 5575 36094
rect 5639 36030 5655 36094
rect 5719 36030 5735 36094
rect 5799 36030 5802 36094
rect 6981 36090 7100 36125
rect 9645 36092 9764 36100
rect 5573 36026 5802 36030
rect 6935 36086 7158 36090
rect 5629 35957 5748 36026
rect 6935 36022 6974 36086
rect 7038 36022 7054 36086
rect 7118 36022 7158 36086
rect 9574 36089 9803 36092
rect 6935 36019 7158 36022
rect 8758 36026 9288 36028
rect 6981 35957 7100 36019
rect 8758 35957 8905 36026
rect 1157 35838 8905 35957
rect 1157 35778 1304 35838
rect 8758 35790 8905 35838
rect 9141 35957 9288 36026
rect 9574 36025 9576 36089
rect 9640 36025 9656 36089
rect 9720 36025 9736 36089
rect 9800 36025 9803 36089
rect 9574 36022 9803 36025
rect 9645 35957 9764 36022
rect 9141 35838 9764 35957
rect 9141 35790 9288 35838
rect 8758 35788 9288 35790
rect 774 35776 1304 35778
rect 3120 35644 3241 35673
rect 3120 35580 3148 35644
rect 3212 35580 3241 35644
rect 3120 35552 3241 35580
rect 7502 35613 7623 35642
rect 3121 35418 3240 35552
rect 7502 35549 7530 35613
rect 7594 35549 7623 35613
rect 7502 35521 7623 35549
rect 9069 35622 9190 35651
rect 9069 35558 9097 35622
rect 9161 35558 9190 35622
rect 9069 35530 9190 35558
rect 4774 35480 5304 35482
rect 4774 35418 4921 35480
rect 3046 35299 4921 35418
rect 4774 35244 4921 35299
rect 5157 35418 5304 35480
rect 7503 35418 7622 35521
rect 9070 35418 9189 35530
rect 5157 35299 9189 35418
rect 5157 35244 5304 35299
rect 4774 35242 5304 35244
rect 4701 31450 4765 32172
rect 7965 31812 8029 32172
rect 7964 31811 8030 31812
rect 7964 31747 7965 31811
rect 8029 31747 8030 31811
rect 7964 31746 8030 31747
rect 3944 31386 4765 31450
rect 4941 31390 5739 31454
rect 6991 31390 7789 31454
rect 7965 31450 8029 31746
rect 4701 31372 4765 31386
rect 7965 31386 8786 31450
rect 11347 31392 11411 46569
rect 11346 31391 11412 31392
rect 7965 31372 8029 31386
rect 11346 31327 11347 31391
rect 11411 31327 11412 31391
rect 11346 31326 11412 31327
rect 3698 30389 3762 31187
rect 4353 30432 4419 30433
rect 4353 30368 4354 30432
rect 4418 30368 4705 30432
rect 5965 30394 6029 31192
rect 6701 30394 6765 31192
rect 8327 30437 8393 30438
rect 8028 30373 8328 30437
rect 8392 30373 8393 30437
rect 8968 30389 9032 31187
rect 8327 30372 8393 30373
rect 4353 30367 4419 30368
rect 3325 30305 3391 30306
rect 3325 30241 3326 30305
rect 3390 30241 3743 30305
rect 3325 30240 3391 30241
rect 3698 29389 3762 30187
rect 4701 29396 4765 30194
rect 5965 29394 6029 30192
rect 6701 29394 6765 30192
rect 7965 29396 8029 30194
rect 8968 29389 9032 30187
rect 3698 28389 3762 29167
rect 4967 28378 5031 29176
rect 5965 28394 6029 29192
rect 6701 28394 6765 29192
rect 7699 28378 7763 29176
rect 8968 28389 9032 29187
rect 10632 28804 10698 28805
rect 10632 28740 10633 28804
rect 10697 28740 10698 28804
rect 10632 28739 10698 28740
rect 3698 27389 3762 28187
rect 5965 27394 6029 28192
rect 6701 27394 6765 28192
rect 8968 27389 9032 28187
rect 4703 27188 4767 27200
rect 7963 27188 8027 27200
rect 3966 27124 4767 27188
rect 4966 27124 5764 27188
rect 6966 27124 7764 27188
rect 7963 27124 8764 27188
rect 4703 26402 4767 27124
rect 7963 26402 8027 27124
rect 7600 24848 7666 24849
rect 7600 24784 7601 24848
rect 7665 24784 7666 24848
rect 7600 24783 7666 24784
rect 5718 24595 5782 24717
rect 5714 24582 5784 24595
rect 5714 24518 5717 24582
rect 5781 24518 5784 24582
rect 7265 24593 7331 24594
rect 7265 24529 7266 24593
rect 7330 24529 7331 24593
rect 7265 24528 7331 24529
rect 5714 24502 5784 24518
rect 5714 24438 5717 24502
rect 5781 24438 5784 24502
rect 5714 24422 5784 24438
rect 5714 24358 5717 24422
rect 5781 24358 5784 24422
rect 5714 24342 5784 24358
rect 5714 24278 5717 24342
rect 5781 24278 5784 24342
rect 5714 24262 5784 24278
rect 5714 24198 5717 24262
rect 5781 24198 5784 24262
rect 5714 24185 5784 24198
rect 4779 23157 5244 23160
rect 4779 23151 4893 23157
rect 5129 23151 5244 23157
rect 4779 22927 4819 23151
rect 5203 22927 5244 23151
rect 5718 23064 5782 24185
rect 7266 23888 7330 24528
rect 7265 23887 7331 23888
rect 7265 23823 7266 23887
rect 7330 23823 7331 23887
rect 7265 23822 7331 23823
rect 5717 23063 5783 23064
rect 5717 22999 5718 23063
rect 5782 22999 5783 23063
rect 5717 22998 5783 22999
rect 4779 22921 4893 22927
rect 5129 22921 5244 22927
rect 4779 22918 5244 22921
rect 7601 22274 7665 24783
rect 8128 24530 8194 24531
rect 8128 24466 8129 24530
rect 8193 24466 8194 24530
rect 8128 24465 8194 24466
rect 8129 22725 8193 24465
rect 8774 23493 9237 23495
rect 8774 23333 8887 23493
rect 8774 23269 8793 23333
rect 8857 23269 8873 23333
rect 8774 23257 8887 23269
rect 9123 23257 9237 23493
rect 8774 23255 9237 23257
rect 8786 23245 8944 23255
rect 8128 22724 8194 22725
rect 8128 22660 8129 22724
rect 8193 22660 8194 22724
rect 8128 22659 8194 22660
rect 8129 22651 8193 22659
rect 7600 22273 7666 22274
rect 7600 22209 7601 22273
rect 7665 22209 7666 22273
rect 7600 22208 7666 22209
rect 10633 20950 10697 28739
rect 11347 26351 11411 31326
rect 11966 30773 12030 47192
rect 16715 46725 33227 46767
rect 16715 46661 17976 46725
rect 18040 46661 19064 46725
rect 19128 46661 20152 46725
rect 20216 46661 21240 46725
rect 21304 46661 22328 46725
rect 22392 46661 24504 46725
rect 24568 46661 25592 46725
rect 25656 46661 26680 46725
rect 26744 46661 27768 46725
rect 27832 46661 28856 46725
rect 28920 46661 29944 46725
rect 30008 46661 31032 46725
rect 31096 46717 33227 46725
rect 31096 46661 33290 46717
rect 16715 46645 33290 46661
rect 16715 46582 17976 46645
rect 16715 46346 16910 46582
rect 17146 46581 17976 46582
rect 18040 46581 19064 46645
rect 19128 46581 20152 46645
rect 20216 46581 21240 46645
rect 21304 46581 22328 46645
rect 22392 46581 24504 46645
rect 24568 46581 25592 46645
rect 25656 46581 26680 46645
rect 26744 46581 27768 46645
rect 27832 46581 28856 46645
rect 28920 46581 29944 46645
rect 30008 46581 31032 46645
rect 31096 46581 33290 46645
rect 17146 46575 33290 46581
rect 17146 46565 24906 46575
rect 17146 46501 17976 46565
rect 18040 46501 19064 46565
rect 19128 46501 20152 46565
rect 20216 46501 21240 46565
rect 21304 46501 22328 46565
rect 22392 46501 24504 46565
rect 24568 46501 24906 46565
rect 17146 46485 24906 46501
rect 17146 46421 17976 46485
rect 18040 46421 19064 46485
rect 19128 46421 20152 46485
rect 20216 46421 21240 46485
rect 21304 46421 22328 46485
rect 22392 46421 24504 46485
rect 24568 46421 24906 46485
rect 17146 46405 24906 46421
rect 17146 46346 17976 46405
rect 16715 46341 17976 46346
rect 18040 46341 19064 46405
rect 19128 46341 20152 46405
rect 20216 46341 21240 46405
rect 21304 46341 22328 46405
rect 22392 46341 24504 46405
rect 24568 46341 24906 46405
rect 16715 46339 24906 46341
rect 25142 46571 33290 46575
rect 25142 46565 32909 46571
rect 25142 46501 25592 46565
rect 25656 46501 26680 46565
rect 26744 46501 27768 46565
rect 27832 46501 28856 46565
rect 28920 46501 29944 46565
rect 30008 46501 31032 46565
rect 31096 46501 32909 46565
rect 25142 46485 32909 46501
rect 25142 46421 25592 46485
rect 25656 46421 26680 46485
rect 26744 46421 27768 46485
rect 27832 46421 28856 46485
rect 28920 46421 29944 46485
rect 30008 46421 31032 46485
rect 31096 46421 32909 46485
rect 25142 46405 32909 46421
rect 25142 46341 25592 46405
rect 25656 46341 26680 46405
rect 26744 46341 27768 46405
rect 27832 46341 28856 46405
rect 28920 46341 29944 46405
rect 30008 46341 31032 46405
rect 31096 46341 32909 46405
rect 25142 46339 32909 46341
rect 16715 46335 32909 46339
rect 33145 46335 33290 46571
rect 16715 46325 33290 46335
rect 16715 46261 17976 46325
rect 18040 46261 19064 46325
rect 19128 46261 20152 46325
rect 20216 46261 21240 46325
rect 21304 46261 22328 46325
rect 22392 46261 24504 46325
rect 24568 46261 25592 46325
rect 25656 46261 26680 46325
rect 26744 46261 27768 46325
rect 27832 46261 28856 46325
rect 28920 46261 29944 46325
rect 30008 46261 31032 46325
rect 31096 46261 33290 46325
rect 16715 46245 33290 46261
rect 16715 46181 17976 46245
rect 18040 46181 19064 46245
rect 19128 46181 20152 46245
rect 20216 46181 21240 46245
rect 21304 46181 22328 46245
rect 22392 46181 24504 46245
rect 24568 46181 25592 46245
rect 25656 46181 26680 46245
rect 26744 46181 27768 46245
rect 27832 46181 28856 46245
rect 28920 46181 29944 46245
rect 30008 46181 31032 46245
rect 31096 46189 33290 46245
rect 31096 46181 33227 46189
rect 16715 46147 33227 46181
rect 18244 45748 18310 45749
rect 18244 45684 18245 45748
rect 18309 45684 18310 45748
rect 18244 45683 18310 45684
rect 18790 45748 18856 45749
rect 18790 45684 18791 45748
rect 18855 45684 18856 45748
rect 26405 45742 26471 45743
rect 18790 45683 18856 45684
rect 19336 45739 19402 45740
rect 18245 44702 18309 45683
rect 18791 45073 18855 45683
rect 19336 45675 19337 45739
rect 19401 45675 19402 45739
rect 19336 45674 19402 45675
rect 19881 45738 19947 45739
rect 19881 45674 19882 45738
rect 19946 45674 19947 45738
rect 25862 45738 25928 45739
rect 23144 45727 23210 45728
rect 18790 45072 18856 45073
rect 18790 45008 18791 45072
rect 18855 45008 18856 45072
rect 18790 45007 18856 45008
rect 18244 44701 18310 44702
rect 18244 44637 18245 44701
rect 18309 44637 18310 44701
rect 18244 44636 18310 44637
rect 18245 38437 18309 44636
rect 13830 38436 13896 38437
rect 13830 38372 13831 38436
rect 13895 38372 13896 38436
rect 13830 38371 13896 38372
rect 18244 38436 18310 38437
rect 18244 38372 18245 38436
rect 18309 38372 18310 38436
rect 18244 38371 18310 38372
rect 13831 31392 13895 38371
rect 18791 37862 18855 45007
rect 19337 41012 19401 45674
rect 19881 45673 19947 45674
rect 21512 45726 21578 45727
rect 19882 41383 19946 45673
rect 21512 45662 21513 45726
rect 21577 45662 21578 45726
rect 21512 45661 21578 45662
rect 22055 45723 22121 45724
rect 19881 41382 19947 41383
rect 19881 41318 19882 41382
rect 19946 41318 19947 41382
rect 19881 41317 19947 41318
rect 19336 41011 19402 41012
rect 19336 40947 19337 41011
rect 19401 40947 19402 41011
rect 19336 40946 19402 40947
rect 14585 37861 14651 37862
rect 14585 37797 14586 37861
rect 14650 37797 14651 37861
rect 14585 37796 14651 37797
rect 18790 37861 18856 37862
rect 18790 37797 18791 37861
rect 18855 37797 18856 37861
rect 18790 37796 18856 37797
rect 13830 31391 13896 31392
rect 13830 31327 13831 31391
rect 13895 31327 13896 31391
rect 13830 31326 13896 31327
rect 14586 30773 14650 37796
rect 19337 37311 19401 40946
rect 15229 37310 15295 37311
rect 15229 37246 15230 37310
rect 15294 37246 15295 37310
rect 15229 37245 15295 37246
rect 19336 37310 19402 37311
rect 19336 37246 19337 37310
rect 19401 37246 19402 37310
rect 19336 37245 19402 37246
rect 11965 30772 12031 30773
rect 11965 30708 11966 30772
rect 12030 30708 12031 30772
rect 11965 30707 12031 30708
rect 14585 30772 14651 30773
rect 14585 30708 14586 30772
rect 14650 30708 14651 30772
rect 14585 30707 14651 30708
rect 11966 28805 12030 30707
rect 11965 28804 12031 28805
rect 11965 28740 11966 28804
rect 12030 28740 12031 28804
rect 11965 28739 12031 28740
rect 11966 28734 12030 28739
rect 11346 26350 11412 26351
rect 11346 26286 11347 26350
rect 11411 26286 11412 26350
rect 11346 26285 11412 26286
rect 11836 26350 11902 26351
rect 11836 26286 11837 26350
rect 11901 26286 11902 26350
rect 11836 26285 11902 26286
rect 11347 26280 11411 26285
rect 11080 24203 11144 24209
rect 11079 24202 11145 24203
rect 11079 24138 11080 24202
rect 11144 24138 11145 24202
rect 11079 24137 11145 24138
rect 10632 20886 10698 20950
rect 11080 20886 11144 24137
rect 11837 22917 11901 26285
rect 13849 26009 13915 26010
rect 13849 25945 13850 26009
rect 13914 25945 13915 26009
rect 13849 25944 13915 25945
rect 13265 25598 13331 25599
rect 13265 25534 13266 25598
rect 13330 25534 13331 25598
rect 13265 25533 13331 25534
rect 12588 23211 12652 23220
rect 12587 23210 12653 23211
rect 12587 23146 12588 23210
rect 12652 23146 12653 23210
rect 12587 23145 12653 23146
rect 11836 22916 11902 22917
rect 11475 22915 11541 22916
rect 11475 22851 11476 22915
rect 11540 22851 11541 22915
rect 11836 22852 11837 22916
rect 11901 22852 11902 22916
rect 11836 22851 11902 22852
rect 11475 22850 11541 22851
rect 10632 20820 11144 20886
rect 11080 20335 11144 20820
rect 11079 20334 11145 20335
rect 11079 20270 11080 20334
rect 11144 20270 11145 20334
rect 11079 20269 11145 20270
rect 11476 19804 11540 22850
rect 12072 21656 12136 21664
rect 12071 21655 12137 21656
rect 12071 21591 12072 21655
rect 12136 21591 12137 21655
rect 12071 21590 12137 21591
rect 11475 19803 11541 19804
rect 11475 19739 11476 19803
rect 11540 19739 11541 19803
rect 11475 19738 11541 19739
rect 4797 19231 5260 19233
rect -2399 19212 -2333 19213
rect -2399 19148 -2398 19212
rect -2334 19148 -2333 19212
rect -2399 19147 -2333 19148
rect 4797 19172 4910 19231
rect 5146 19172 5260 19231
rect -35043 18994 -35027 18995
rect -34963 18994 -34947 18995
rect -34883 18994 -34755 18995
rect -38169 18993 -34755 18994
rect -5280 19043 -5214 19044
rect -38169 18986 -34860 18993
rect -5280 18979 -5279 19043
rect -5215 18979 -5214 19043
rect -5280 18978 -5214 18979
rect -3919 19043 -3853 19044
rect -3919 18979 -3918 19043
rect -3854 18979 -3853 19043
rect -3919 18978 -3853 18979
rect -27238 17961 -26708 17963
rect -27238 17725 -27091 17961
rect -26855 17913 -26708 17961
rect -25453 17913 -25386 17923
rect -26855 17886 -25378 17913
rect -26855 17822 -25452 17886
rect -25388 17822 -25378 17886
rect -26855 17806 -25378 17822
rect -26855 17785 -25452 17806
rect -26855 17725 -26708 17785
rect -27238 17723 -26708 17725
rect -25453 17742 -25452 17785
rect -25388 17785 -25378 17806
rect -3212 17862 -2747 17865
rect -3212 17856 -3098 17862
rect -2862 17856 -2747 17862
rect -25388 17742 -25386 17785
rect -25453 17726 -25386 17742
rect -25453 17662 -25452 17726
rect -25388 17662 -25386 17726
rect -25453 17626 -25386 17662
rect -3212 17632 -3172 17856
rect -2788 17632 -2747 17856
rect -3212 17626 -3098 17632
rect -2862 17626 -2747 17632
rect -3212 17623 -2747 17626
rect -25451 17398 -25377 17405
rect -25451 17336 -25446 17398
rect -25454 17334 -25446 17336
rect -25382 17336 -25377 17398
rect -25382 17334 -24738 17336
rect -25454 17318 -24738 17334
rect -25454 17254 -25446 17318
rect -25382 17254 -24738 17318
rect -25454 17238 -24738 17254
rect -25454 17208 -25446 17238
rect -25451 17174 -25446 17208
rect -25382 17208 -24738 17238
rect -25382 17174 -25377 17208
rect -25451 17168 -25377 17174
rect -39204 16198 -38741 16200
rect -39204 15962 -39091 16198
rect -38855 16078 -38741 16198
rect -38855 16076 -34857 16078
rect -38855 16063 -34851 16076
rect -38855 15999 -38145 16063
rect -38081 15999 -38065 16063
rect -38001 15999 -37985 16063
rect -37921 15999 -37905 16063
rect -37841 15999 -37825 16063
rect -37761 15999 -37745 16063
rect -37681 15999 -37665 16063
rect -37601 15999 -37585 16063
rect -37521 15999 -37505 16063
rect -37441 15999 -37425 16063
rect -37361 15999 -37345 16063
rect -37281 15999 -37265 16063
rect -37201 15999 -37185 16063
rect -37121 15999 -37105 16063
rect -37041 15999 -37025 16063
rect -36961 15999 -36945 16063
rect -36881 15999 -36865 16063
rect -36801 15999 -36785 16063
rect -36721 15999 -36705 16063
rect -36641 15999 -36625 16063
rect -36561 15999 -36545 16063
rect -36481 15999 -36465 16063
rect -36401 15999 -36385 16063
rect -36321 15999 -36305 16063
rect -36241 15999 -36225 16063
rect -36161 15999 -36145 16063
rect -36081 15999 -36065 16063
rect -36001 15999 -35985 16063
rect -35921 15999 -35905 16063
rect -35841 15999 -35825 16063
rect -35761 15999 -35745 16063
rect -35681 15999 -35665 16063
rect -35601 15999 -35585 16063
rect -35521 15999 -35505 16063
rect -35441 15999 -35425 16063
rect -35361 15999 -35345 16063
rect -35281 15999 -35265 16063
rect -35201 15999 -35185 16063
rect -35121 15999 -35105 16063
rect -35041 15999 -35025 16063
rect -34961 15999 -34945 16063
rect -34881 15999 -34851 16063
rect -38855 15986 -34851 15999
rect -38855 15984 -34857 15986
rect -38855 15962 -38741 15984
rect -39204 15960 -38741 15962
rect -24866 15445 -24738 17208
rect -18719 17145 -17699 17209
rect -16119 17145 -15099 17209
rect -13519 17145 -12499 17209
rect -10417 17157 -10351 17158
rect -10912 17093 -10416 17157
rect -10352 17093 -10351 17157
rect -10417 17092 -10351 17093
rect -2398 16989 -2334 19147
rect 4797 19028 4873 19172
rect 5177 19028 5260 19172
rect 4797 18995 4910 19028
rect 5146 18995 5260 19028
rect 4797 18993 5260 18995
rect 10231 19058 10297 19059
rect 10231 18994 10232 19058
rect 10296 18994 10297 19058
rect 10231 18993 10297 18994
rect -1505 18910 -1439 18911
rect -1505 18846 -1504 18910
rect -1440 18846 -1439 18910
rect -1505 18845 -1439 18846
rect -3928 16925 -2334 16989
rect -23253 15488 -22723 15490
rect -23253 15445 -23106 15488
rect -24866 15317 -23106 15445
rect -27231 14475 -26701 14477
rect -27231 14239 -27084 14475
rect -26848 14425 -26701 14475
rect -25518 14425 -25443 14447
rect -26848 14413 -25414 14425
rect -26848 14349 -25513 14413
rect -25449 14349 -25414 14413
rect -26848 14333 -25414 14349
rect -26848 14297 -25513 14333
rect -26848 14239 -26701 14297
rect -27231 14237 -26701 14239
rect -25518 14269 -25513 14297
rect -25449 14297 -25414 14333
rect -25449 14269 -25443 14297
rect -25518 14253 -25443 14269
rect -25518 14189 -25513 14253
rect -25449 14189 -25443 14253
rect -25518 14156 -25443 14189
rect -25519 13919 -25445 13926
rect -25519 13874 -25514 13919
rect -25520 13855 -25514 13874
rect -25450 13874 -25445 13919
rect -24866 13874 -24738 15317
rect -23253 15252 -23106 15317
rect -22870 15252 -22723 15488
rect -23253 15250 -22723 15252
rect -20013 14880 -19949 15900
rect -14185 15370 -14055 15403
rect -14185 15306 -14152 15370
rect -14088 15306 -14055 15370
rect -14185 15273 -14055 15306
rect -14184 14892 -14056 15273
rect -11255 14873 -11191 15893
rect -7218 15810 -6755 15812
rect -7218 15574 -7105 15810
rect -6869 15708 -6755 15810
rect -5787 15708 -5721 15709
rect -6869 15644 -5786 15708
rect -5722 15644 -5721 15708
rect -6869 15574 -6755 15644
rect -5787 15643 -5721 15644
rect -7218 15572 -6755 15574
rect -3928 15455 -3864 16925
rect -3201 16448 -2738 16450
rect -3201 16212 -3088 16448
rect -2852 16212 -2738 16448
rect -3201 16210 -2738 16212
rect -3510 16205 -3444 16206
rect -3510 16141 -3509 16205
rect -3445 16141 -3444 16205
rect -3510 16140 -3444 16141
rect -3929 15454 -3863 15455
rect -3929 15390 -3928 15454
rect -3864 15390 -3863 15454
rect -3929 15389 -3863 15390
rect -7221 14450 -6758 14452
rect -7221 14214 -7108 14450
rect -6872 14345 -6758 14450
rect -4903 14413 -4831 14447
rect -4903 14349 -4899 14413
rect -4835 14349 -4831 14413
rect -4903 14345 -4831 14349
rect -6872 14333 -4828 14345
rect -6872 14281 -4899 14333
rect -6872 14214 -6758 14281
rect -4903 14269 -4899 14281
rect -4835 14281 -4828 14333
rect -4835 14269 -4831 14281
rect -4903 14235 -4831 14269
rect -7221 14212 -6758 14214
rect -18224 14073 -18158 14074
rect -18224 14009 -18223 14073
rect -18159 14009 -17732 14073
rect -18224 14008 -18158 14009
rect -25450 13855 -24738 13874
rect -25520 13839 -24738 13855
rect -25520 13775 -25514 13839
rect -25450 13775 -24738 13839
rect -25520 13759 -24738 13775
rect -25520 13746 -25514 13759
rect -25519 13695 -25514 13746
rect -25450 13746 -24738 13759
rect -25450 13695 -25445 13746
rect -25519 13689 -25445 13695
rect -16124 13625 -15104 13689
rect -20013 12280 -19949 13300
rect -11255 12273 -11191 13293
rect -18722 10995 -17702 11059
rect -16122 10995 -15102 11059
rect -13522 10995 -12502 11059
rect -7221 10910 -6758 10912
rect -7221 10674 -7108 10910
rect -6872 10832 -6758 10910
rect -6163 10832 -5936 10834
rect -6872 10827 -5929 10832
rect -6872 10768 -6162 10827
rect -6872 10674 -6758 10768
rect -6163 10763 -6162 10768
rect -6098 10763 -6082 10827
rect -6018 10763 -6002 10827
rect -5938 10768 -5929 10827
rect -5938 10763 -5936 10768
rect -6163 10757 -5936 10763
rect -7221 10672 -6758 10674
rect -10971 10223 -10905 10224
rect -10971 10159 -10970 10223
rect -10906 10159 -10905 10223
rect -10971 10158 -10905 10159
rect -10970 9696 -10906 10158
rect -7211 9660 -6748 9662
rect -7211 9424 -7098 9660
rect -6862 9572 -6748 9660
rect -6168 9584 -5928 9593
rect -6168 9572 -6160 9584
rect -6862 9520 -6160 9572
rect -6096 9520 -6080 9584
rect -6016 9520 -6000 9584
rect -5936 9572 -5928 9584
rect -5936 9520 -5909 9572
rect -6862 9508 -5909 9520
rect -6862 9424 -6748 9508
rect -7211 9422 -6748 9424
rect -18719 9345 -17699 9409
rect -16119 9345 -15099 9409
rect -13519 9345 -12499 9409
rect -20013 7080 -19949 8100
rect -16782 7607 -16652 7640
rect -16782 7543 -16749 7607
rect -16685 7543 -16652 7607
rect -16782 7510 -16652 7543
rect -16781 7040 -16653 7510
rect -11255 7073 -11191 8093
rect -7215 7241 -6750 7244
rect -7215 7235 -7101 7241
rect -6865 7235 -6750 7241
rect -7215 7011 -7175 7235
rect -6791 7011 -6750 7235
rect -7215 7005 -7101 7011
rect -6865 7005 -6750 7011
rect -7215 7002 -6750 7005
rect -27239 6708 -26709 6710
rect -27239 6472 -27092 6708
rect -26856 6646 -26709 6708
rect -25522 6650 -25445 6670
rect -25522 6646 -25516 6650
rect -26856 6586 -25516 6646
rect -25452 6646 -25445 6650
rect -25452 6586 -25404 6646
rect -26856 6570 -25404 6586
rect -26856 6518 -25516 6570
rect -26856 6472 -26709 6518
rect -27239 6470 -26709 6472
rect -25522 6506 -25516 6518
rect -25452 6518 -25404 6570
rect -25452 6506 -25445 6518
rect -25522 6490 -25445 6506
rect -25522 6426 -25516 6490
rect -25452 6426 -25445 6490
rect -25522 6407 -25445 6426
rect -18252 6303 -18186 6304
rect -18252 6239 -18251 6303
rect -18187 6239 -17700 6303
rect -18252 6238 -18186 6239
rect -25523 6163 -25446 6175
rect -25523 6099 -25517 6163
rect -25453 6141 -25446 6163
rect -4911 6164 -4847 6176
rect -25453 6099 -25388 6141
rect -25523 6083 -25388 6099
rect -25523 6019 -25517 6083
rect -25453 6019 -25388 6083
rect -25523 6003 -25388 6019
rect -25523 5939 -25517 6003
rect -25453 5939 -25388 6003
rect -25523 5928 -25388 5939
rect -25516 4984 -25388 5928
rect -4911 6128 -4840 6164
rect -4911 6064 -4906 6128
rect -4842 6064 -4840 6128
rect -4911 6048 -4840 6064
rect -4911 5984 -4906 6048
rect -4842 5984 -4840 6048
rect -3928 6043 -3864 15389
rect -3509 14645 -3445 16140
rect -3134 14999 -3070 15001
rect -3145 14970 -3060 14999
rect -3145 14906 -3135 14970
rect -3071 14906 -3060 14970
rect -3145 14890 -3060 14906
rect -3145 14826 -3135 14890
rect -3071 14826 -3060 14890
rect -3145 14810 -3060 14826
rect -3145 14746 -3135 14810
rect -3071 14746 -3060 14810
rect -3145 14718 -3060 14746
rect -3510 14644 -3444 14645
rect -3510 14580 -3509 14644
rect -3445 14580 -3444 14644
rect -3510 14579 -3444 14580
rect -4911 5949 -4840 5984
rect -3929 6042 -3863 6043
rect -3929 5978 -3928 6042
rect -3864 5978 -3863 6042
rect -3929 5977 -3863 5978
rect -3928 5973 -3864 5977
rect -16124 5825 -15104 5889
rect -7211 5762 -6748 5764
rect -7211 5526 -7098 5762
rect -6862 5670 -6748 5762
rect -4911 5670 -4847 5949
rect -6862 5606 -4847 5670
rect -6862 5526 -6748 5606
rect -7211 5524 -6748 5526
rect -23232 5042 -22702 5044
rect -23232 4984 -23085 5042
rect -25516 4856 -23085 4984
rect -23232 4806 -23085 4856
rect -22849 4806 -22702 5042
rect -23232 4804 -22702 4806
rect -20013 4480 -19949 5500
rect -11255 4473 -11191 5493
rect -3509 5234 -3445 14579
rect -3134 14048 -3070 14718
rect -3199 14046 -2736 14048
rect -3199 13810 -3086 14046
rect -2850 13942 -2736 14046
rect -2850 13878 -2305 13942
rect -2850 13810 -2736 13878
rect -3199 13808 -2736 13810
rect -2369 12955 -2305 13878
rect -1809 13121 -1724 13134
rect -1809 13057 -1799 13121
rect -1735 13057 -1724 13121
rect -1809 13041 -1724 13057
rect -1809 12977 -1799 13041
rect -1735 12977 -1724 13041
rect -1809 12961 -1724 12977
rect -1809 12955 -1799 12961
rect -2369 12897 -1799 12955
rect -1735 12897 -1724 12961
rect -2369 12891 -1724 12897
rect -2369 11390 -2305 12891
rect -1809 12881 -1724 12891
rect -1809 12817 -1799 12881
rect -1735 12817 -1724 12881
rect -1809 12801 -1724 12817
rect -1809 12737 -1799 12801
rect -1735 12737 -1724 12801
rect -1809 12725 -1724 12737
rect -1760 11526 -1692 11530
rect -1760 11462 -1758 11526
rect -1694 11462 -1692 11526
rect -1760 11446 -1692 11462
rect -1760 11390 -1758 11446
rect -2369 11382 -1758 11390
rect -1694 11382 -1692 11446
rect -2369 11366 -1692 11382
rect -2369 11326 -1758 11366
rect -1760 11302 -1758 11326
rect -1694 11302 -1692 11366
rect -1760 11286 -1692 11302
rect -1760 11222 -1758 11286
rect -1694 11222 -1692 11286
rect -1760 11206 -1692 11222
rect -1760 11142 -1758 11206
rect -1694 11142 -1692 11206
rect -1760 11139 -1692 11142
rect -1760 9923 -1694 9931
rect -1760 9859 -1759 9923
rect -1695 9859 -1694 9923
rect -1760 9843 -1694 9859
rect -1760 9779 -1759 9843
rect -1695 9779 -1694 9843
rect -1760 9775 -1694 9779
rect -2390 9763 -1694 9775
rect -2390 9711 -1759 9763
rect -3201 8800 -2738 8802
rect -3201 8707 -3088 8800
rect -3201 8643 -3185 8707
rect -3121 8643 -3088 8707
rect -3201 8564 -3088 8643
rect -2852 8710 -2738 8800
rect -2390 8710 -2326 9711
rect -1760 9699 -1759 9711
rect -1695 9699 -1694 9763
rect -1760 9683 -1694 9699
rect -1760 9619 -1759 9683
rect -1695 9619 -1694 9683
rect -1760 9603 -1694 9619
rect -1760 9539 -1759 9603
rect -1695 9539 -1694 9603
rect -1760 9531 -1694 9539
rect -2852 8646 -2326 8710
rect -2852 8564 -2738 8646
rect -3201 8562 -2738 8564
rect -2390 8179 -2326 8646
rect -1759 8322 -1689 8331
rect -1759 8258 -1756 8322
rect -1692 8258 -1689 8322
rect -1759 8242 -1689 8258
rect -1759 8179 -1756 8242
rect -2390 8178 -1756 8179
rect -1692 8178 -1689 8242
rect -2390 8162 -1689 8178
rect -2390 8115 -1756 8162
rect -1759 8098 -1756 8115
rect -1692 8098 -1689 8162
rect -1759 8082 -1689 8098
rect -1759 8018 -1756 8082
rect -1692 8018 -1689 8082
rect -1759 8002 -1689 8018
rect -1759 7938 -1756 8002
rect -1692 7938 -1689 8002
rect -1759 7929 -1689 7938
rect -3199 6741 -2736 6743
rect -3199 6649 -3086 6741
rect -3199 6585 -3184 6649
rect -3120 6585 -3086 6649
rect -3199 6505 -3086 6585
rect -2850 6651 -2736 6741
rect -2850 6587 -2335 6651
rect -2850 6505 -2736 6587
rect -3199 6503 -2736 6505
rect -3194 5548 -3109 5578
rect -3194 5484 -3184 5548
rect -3120 5484 -3109 5548
rect -3194 5468 -3109 5484
rect -3194 5411 -3184 5468
rect -3201 5404 -3184 5411
rect -3120 5411 -3109 5468
rect -2399 5411 -2335 6587
rect -3120 5404 -2335 5411
rect -3201 5388 -2335 5404
rect -3201 5347 -3184 5388
rect -3194 5324 -3184 5347
rect -3120 5347 -2335 5388
rect -3120 5324 -3109 5347
rect -3194 5295 -3109 5324
rect -3510 5233 -3444 5234
rect -3510 5169 -3509 5233
rect -3445 5169 -3444 5233
rect -3510 5168 -3444 5169
rect -18722 3195 -17702 3259
rect -16122 3195 -15102 3259
rect -13522 3195 -12502 3259
rect -1504 -3060 -1440 18845
rect 8279 18718 8345 18719
rect 8279 18654 8280 18718
rect 8344 18654 8345 18718
rect 8279 18653 8345 18654
rect -1134 18651 -1068 18652
rect -1134 18587 -1133 18651
rect -1069 18587 -1068 18651
rect -1134 18586 -1068 18587
rect -1133 -2703 -1069 18586
rect -681 18312 -615 18313
rect -681 18248 -680 18312
rect -616 18248 -615 18312
rect -681 18247 -615 18248
rect -680 -2288 -616 18247
rect -285 18031 -219 18032
rect -285 17967 -284 18031
rect -220 17967 -219 18031
rect -285 17966 -219 17967
rect -284 -1862 -220 17966
rect 789 17616 1252 17618
rect 789 17380 902 17616
rect 1138 17380 1252 17616
rect 789 17378 1252 17380
rect 4294 17289 4360 17290
rect 6226 17289 6292 17290
rect 8280 17289 8344 18653
rect 8789 17401 9252 17403
rect 8789 17289 8902 17401
rect 4294 17225 4295 17289
rect 4359 17225 6227 17289
rect 6291 17225 8902 17289
rect 4294 17224 4360 17225
rect 6226 17224 6292 17225
rect 8789 17165 8902 17225
rect 9138 17289 9252 17401
rect 10232 17289 10296 18993
rect 9138 17225 10296 17289
rect 9138 17165 9252 17225
rect 8789 17163 9252 17165
rect 4794 16593 5256 16746
rect 4794 16447 4907 16593
rect 250 16414 4907 16447
rect 5143 16447 5256 16593
rect 5143 16414 11140 16447
rect 250 16270 263 16414
rect 11127 16270 11140 16414
rect 250 16237 4907 16270
rect 4792 16190 4907 16237
rect 4794 16037 4907 16190
rect 5143 16237 11140 16270
rect 5143 16037 5256 16237
rect 4794 15884 5256 16037
rect 12072 12363 12136 21590
rect 12588 13171 12652 23145
rect 12861 21094 13103 21097
rect 12861 20858 12864 21094
rect 13100 20858 13103 21094
rect 12861 20855 13103 20858
rect 12849 18793 13091 18796
rect 12849 18557 12852 18793
rect 13088 18557 13091 18793
rect 12849 18554 13091 18557
rect 13266 17763 13330 25533
rect 13850 18571 13914 25944
rect 15230 24849 15294 37245
rect 19882 36729 19946 41317
rect 21513 40113 21577 45661
rect 22055 45659 22056 45723
rect 22120 45659 22121 45723
rect 22055 45658 22121 45659
rect 21512 40112 21578 40113
rect 21512 40048 21513 40112
rect 21577 40048 21578 40112
rect 21512 40047 21578 40048
rect 15989 36728 16055 36729
rect 15989 36664 15990 36728
rect 16054 36664 16055 36728
rect 15989 36663 16055 36664
rect 19881 36728 19947 36729
rect 19881 36664 19882 36728
rect 19946 36664 19947 36728
rect 19881 36663 19947 36664
rect 15229 24848 15295 24849
rect 15229 24784 15230 24848
rect 15294 24784 15295 24848
rect 15229 24783 15295 24784
rect 15990 24531 16054 36663
rect 16720 36050 16786 36051
rect 16720 35986 16721 36050
rect 16785 35986 16786 36050
rect 16720 35985 16786 35986
rect 16721 29753 16785 35985
rect 17411 35343 17477 35344
rect 17411 35279 17412 35343
rect 17476 35279 17477 35343
rect 17411 35278 17477 35279
rect 16720 29752 16786 29753
rect 16720 29688 16721 29752
rect 16785 29688 16786 29752
rect 16720 29687 16786 29688
rect 17412 29330 17476 35278
rect 18251 34583 18317 34584
rect 18251 34519 18252 34583
rect 18316 34519 18317 34583
rect 18251 34518 18317 34519
rect 17411 29329 17477 29330
rect 17411 29265 17412 29329
rect 17476 29265 17477 29329
rect 17411 29264 17477 29265
rect 17412 29261 17476 29264
rect 15989 24530 16055 24531
rect 15989 24466 15990 24530
rect 16054 24466 16055 24530
rect 15989 24465 16055 24466
rect 18252 23519 18316 34518
rect 21513 33747 21577 40047
rect 22057 39742 22121 45658
rect 22597 45722 22663 45723
rect 22597 45658 22598 45722
rect 22662 45658 22663 45722
rect 23144 45663 23145 45727
rect 23209 45663 23210 45727
rect 25862 45674 25863 45738
rect 25927 45674 25928 45738
rect 26405 45678 26406 45742
rect 26470 45678 26471 45742
rect 29128 45738 29194 45739
rect 26405 45677 26471 45678
rect 26947 45736 27013 45737
rect 25862 45673 25928 45674
rect 23144 45662 23210 45663
rect 22597 45657 22663 45658
rect 22598 43923 22662 45657
rect 22596 43922 22662 43923
rect 22596 43858 22597 43922
rect 22661 43858 22662 43922
rect 22596 43857 22662 43858
rect 22056 39741 22122 39742
rect 22056 39677 22057 39741
rect 22121 39677 22122 39741
rect 22056 39676 22122 39677
rect 22057 34584 22121 39676
rect 22598 35344 22662 43857
rect 23145 43552 23209 45662
rect 25863 44892 25927 45673
rect 25862 44891 25928 44892
rect 25862 44827 25863 44891
rect 25927 44827 25928 44891
rect 25862 44826 25928 44827
rect 23144 43551 23210 43552
rect 23144 43487 23145 43551
rect 23209 43487 23210 43551
rect 23144 43486 23210 43487
rect 23145 36051 23209 43486
rect 25863 38419 25927 44826
rect 26406 44527 26470 45677
rect 26947 45672 26948 45736
rect 27012 45672 27013 45736
rect 26947 45671 27013 45672
rect 27504 45727 27570 45728
rect 26405 44526 26471 44527
rect 26405 44462 26406 44526
rect 26470 44462 26471 44526
rect 26405 44461 26471 44462
rect 25862 38418 25928 38419
rect 25862 38354 25863 38418
rect 25927 38354 25928 38418
rect 25862 38353 25928 38354
rect 26406 37839 26470 44461
rect 26948 41202 27012 45671
rect 27504 45663 27505 45727
rect 27569 45663 27570 45727
rect 29128 45674 29129 45738
rect 29193 45674 29194 45738
rect 30222 45735 30288 45736
rect 29128 45673 29194 45674
rect 29672 45731 29738 45732
rect 27504 45662 27570 45663
rect 26947 41201 27013 41202
rect 26947 41137 26948 41201
rect 27012 41137 27013 41201
rect 26947 41136 27013 41137
rect 26405 37838 26471 37839
rect 26405 37774 26406 37838
rect 26470 37774 26471 37838
rect 26405 37773 26471 37774
rect 23144 36050 23210 36051
rect 23144 35986 23145 36050
rect 23209 35986 23210 36050
rect 23144 35985 23210 35986
rect 22597 35343 22663 35344
rect 22597 35279 22598 35343
rect 22662 35279 22663 35343
rect 22597 35278 22663 35279
rect 22598 35258 22662 35278
rect 22055 34583 22121 34584
rect 22055 34519 22056 34583
rect 22120 34519 22121 34583
rect 26948 34523 27012 41136
rect 27505 40837 27569 45662
rect 27504 40836 27570 40837
rect 27504 40772 27505 40836
rect 27569 40772 27570 40836
rect 27504 40771 27570 40772
rect 22055 34518 22121 34519
rect 26947 34522 27013 34523
rect 26947 34458 26948 34522
rect 27012 34458 27013 34522
rect 26947 34457 27013 34458
rect 27505 33814 27569 40771
rect 29129 39567 29193 45673
rect 29672 45667 29673 45731
rect 29737 45667 29738 45731
rect 29672 45666 29738 45667
rect 30222 45671 30223 45735
rect 30287 45671 30288 45735
rect 30222 45670 30288 45671
rect 30755 45735 30821 45736
rect 30755 45671 30756 45735
rect 30820 45671 30821 45735
rect 30755 45670 30821 45671
rect 29673 39932 29737 45666
rect 30222 43376 30286 45670
rect 30756 43742 30820 45670
rect 30755 43741 30821 43742
rect 30755 43677 30756 43741
rect 30820 43677 30821 43741
rect 30755 43676 30821 43677
rect 30221 43375 30287 43376
rect 30221 43311 30222 43375
rect 30286 43311 30287 43375
rect 30221 43310 30287 43311
rect 29672 39931 29738 39932
rect 29672 39867 29673 39931
rect 29737 39867 29738 39931
rect 29672 39866 29738 39867
rect 29128 39566 29194 39567
rect 29128 39502 29129 39566
rect 29193 39502 29194 39566
rect 29128 39501 29194 39502
rect 29129 35259 29193 39501
rect 29673 35971 29737 39866
rect 30222 36594 30286 43310
rect 30756 37230 30820 43676
rect 32413 38418 32479 38419
rect 32413 38354 32414 38418
rect 32478 38354 32479 38418
rect 32413 38353 32479 38354
rect 31823 37838 31889 37839
rect 31823 37774 31824 37838
rect 31888 37774 31889 37838
rect 31823 37773 31889 37774
rect 30755 37229 30821 37230
rect 30755 37165 30756 37229
rect 30820 37165 30821 37229
rect 30755 37164 30821 37165
rect 31230 37229 31296 37230
rect 31230 37165 31231 37229
rect 31295 37165 31296 37229
rect 31230 37164 31296 37165
rect 30221 36593 30287 36594
rect 30221 36529 30222 36593
rect 30286 36529 30287 36593
rect 30221 36528 30287 36529
rect 30583 36593 30649 36594
rect 30583 36529 30584 36593
rect 30648 36529 30649 36593
rect 30583 36528 30649 36529
rect 29672 35970 29738 35971
rect 29672 35906 29673 35970
rect 29737 35906 29738 35970
rect 29672 35905 29738 35906
rect 29989 35970 30055 35971
rect 29989 35906 29990 35970
rect 30054 35906 30055 35970
rect 29989 35905 30055 35906
rect 29128 35258 29194 35259
rect 29128 35194 29129 35258
rect 29193 35194 29194 35258
rect 29128 35193 29194 35194
rect 29406 35258 29472 35259
rect 29406 35194 29407 35258
rect 29471 35194 29472 35258
rect 29406 35193 29472 35194
rect 28827 34522 28893 34523
rect 28827 34458 28828 34522
rect 28892 34458 28893 34522
rect 28827 34457 28893 34458
rect 27504 33813 27570 33814
rect 27504 33749 27505 33813
rect 27569 33749 27570 33813
rect 27504 33748 27570 33749
rect 28314 33813 28380 33814
rect 28314 33749 28315 33813
rect 28379 33749 28380 33813
rect 28314 33748 28380 33749
rect 19254 33746 19320 33747
rect 19254 33682 19255 33746
rect 19319 33682 19320 33746
rect 19254 33681 19320 33682
rect 21512 33746 21579 33747
rect 21512 33682 21513 33746
rect 21577 33682 21579 33746
rect 21512 33681 21579 33682
rect 19255 23888 19319 33681
rect 25878 26009 25944 26010
rect 25878 25945 25879 26009
rect 25943 25945 25944 26009
rect 25878 25944 25944 25945
rect 19254 23887 19320 23888
rect 19254 23823 19255 23887
rect 19319 23823 19320 23887
rect 19254 23822 19320 23823
rect 18251 23518 18317 23519
rect 18251 23454 18252 23518
rect 18316 23454 18317 23518
rect 18251 23453 18317 23454
rect 23688 19382 23754 19383
rect 14686 19328 14750 19332
rect 14686 19327 14752 19328
rect 14686 19263 14687 19327
rect 14751 19263 14752 19327
rect 23688 19318 23689 19382
rect 23753 19318 23754 19382
rect 23688 19317 23754 19318
rect 14686 19262 14752 19263
rect 14686 19095 14750 19262
rect 16889 19185 17131 19188
rect 14686 19094 14753 19095
rect 16889 19094 16892 19185
rect 14686 19030 16892 19094
rect 14114 18571 14180 18572
rect 13850 18507 14115 18571
rect 14179 18507 14180 18571
rect 14114 18506 14180 18507
rect 14367 17763 14433 17764
rect 13266 17699 14368 17763
rect 14432 17699 14433 17763
rect 14367 17698 14433 17699
rect 14689 17543 14753 19030
rect 16889 18949 16892 19030
rect 17128 18949 17131 19185
rect 16889 18946 17131 18949
rect 20893 19158 21135 19161
rect 20893 18922 20896 19158
rect 21132 18922 21135 19158
rect 20893 18919 21135 18922
rect 23689 19083 23753 19317
rect 24903 19153 25145 19156
rect 24903 19083 24906 19153
rect 23689 19019 24906 19083
rect 23689 17553 23753 19019
rect 24903 18917 24906 19019
rect 25142 18917 25145 19153
rect 24903 18914 25145 18917
rect 25613 18571 25679 18572
rect 25879 18571 25943 25944
rect 26462 25598 26528 25599
rect 26462 25534 26463 25598
rect 26527 25534 26528 25598
rect 26462 25533 26528 25534
rect 25613 18507 25614 18571
rect 25678 18507 25943 18571
rect 25613 18506 25679 18507
rect 25360 17764 25426 17765
rect 26463 17764 26527 25533
rect 27111 23211 27175 23222
rect 27110 23210 27176 23211
rect 27110 23146 27111 23210
rect 27175 23146 27176 23210
rect 27110 23145 27176 23146
rect 25360 17700 25361 17764
rect 25425 17700 26527 17764
rect 25360 17699 25426 17700
rect 23688 17552 23754 17553
rect 14688 17542 14754 17543
rect 14688 17478 14689 17542
rect 14753 17478 14754 17542
rect 23688 17488 23689 17552
rect 23753 17488 23754 17552
rect 23688 17487 23754 17488
rect 14688 17477 14754 17478
rect 12843 17188 13085 17191
rect 12843 16952 12846 17188
rect 13082 16952 13085 17188
rect 12843 16949 13085 16952
rect 23685 15788 23751 15789
rect 14685 15734 14824 15769
rect 14664 15711 14824 15734
rect 23685 15724 23686 15788
rect 23750 15724 23751 15788
rect 23685 15723 23751 15724
rect 14664 15647 14686 15711
rect 14750 15647 14824 15711
rect 14664 15625 14824 15647
rect 14685 15524 14824 15625
rect 16797 15592 17039 15595
rect 16797 15524 16800 15592
rect 14685 15423 16800 15524
rect 12862 15317 13104 15320
rect 12862 15081 12865 15317
rect 13101 15081 13104 15317
rect 12862 15078 13104 15081
rect 14685 13966 14824 15423
rect 16797 15356 16800 15423
rect 17036 15356 17039 15592
rect 16797 15353 17039 15356
rect 20836 15587 21078 15590
rect 20836 15351 20839 15587
rect 21075 15351 21078 15587
rect 20836 15348 21078 15351
rect 23686 15473 23750 15723
rect 24905 15560 25147 15563
rect 24905 15473 24908 15560
rect 23686 15409 24908 15473
rect 23686 13998 23750 15409
rect 24905 15324 24908 15409
rect 25144 15324 25147 15560
rect 24905 15321 25147 15324
rect 14684 13965 14824 13966
rect 14684 13901 14685 13965
rect 14749 13901 14824 13965
rect 23685 13997 23751 13998
rect 23685 13933 23686 13997
rect 23750 13933 23751 13997
rect 23685 13932 23751 13933
rect 14684 13900 14824 13901
rect 12884 13616 13126 13619
rect 12884 13380 12887 13616
rect 13123 13380 13126 13616
rect 12884 13377 13126 13380
rect 14114 13171 14180 13172
rect 12588 13107 14115 13171
rect 14179 13107 14180 13171
rect 14114 13106 14180 13107
rect 14367 12363 14433 12364
rect 12072 12299 14368 12363
rect 14432 12299 14433 12363
rect 14367 12298 14433 12299
rect 14685 12180 14824 13900
rect 27111 13171 27175 23145
rect 27657 21656 27721 21665
rect 27656 21655 27722 21656
rect 27656 21591 27657 21655
rect 27721 21591 27722 21655
rect 27656 21590 27722 21591
rect 25678 13107 27175 13171
rect 27657 12364 27721 21590
rect 25425 12300 27721 12364
rect 14685 12116 14702 12180
rect 14766 12116 14824 12180
rect 23690 12190 23756 12191
rect 23690 12126 23691 12190
rect 23755 12126 23756 12190
rect 23690 12125 23756 12126
rect 12897 11761 13139 11764
rect 12897 11525 12900 11761
rect 13136 11525 13139 11761
rect 12897 11522 13139 11525
rect 12783 10651 13246 10653
rect 12783 10617 12896 10651
rect 10804 10538 12896 10617
rect 6482 10518 12896 10538
rect 6482 10374 6498 10518
rect 11202 10439 12896 10518
rect 11202 10374 11338 10439
rect 12783 10415 12896 10439
rect 13132 10617 13246 10651
rect 13132 10439 13289 10617
rect 13132 10415 13246 10439
rect 12783 10413 13246 10415
rect 6482 10355 11338 10374
rect 10804 10326 11338 10355
rect 14685 10383 14824 12116
rect 20890 11999 21132 12002
rect 20890 11763 20893 11999
rect 21129 11763 21132 11999
rect 20890 11760 21132 11763
rect 23691 11890 23755 12125
rect 24893 11969 25135 11972
rect 24893 11890 24896 11969
rect 23691 11826 24896 11890
rect 14685 10350 14691 10383
rect 14690 10319 14691 10350
rect 14755 10350 14824 10383
rect 23691 10381 23755 11826
rect 24893 11733 24896 11826
rect 25132 11733 25135 11969
rect 24893 11730 25135 11733
rect 23690 10380 23756 10381
rect 14755 10319 14756 10350
rect 14690 10318 14756 10319
rect 23690 10316 23691 10380
rect 23755 10316 23756 10380
rect 23690 10315 23756 10316
rect 8814 335 9277 337
rect 794 323 1257 325
rect 794 233 907 323
rect 321 221 907 233
rect 1143 233 1257 323
rect 4603 233 4917 290
rect 8814 233 8927 335
rect 1143 221 8927 233
rect 9163 233 9277 335
rect 12169 233 12420 334
rect 16791 323 17254 325
rect 16791 233 16904 323
rect 9163 221 16904 233
rect 17140 233 17254 323
rect 17140 221 21108 233
rect 321 77 322 221
rect 21106 77 21108 221
rect 321 66 21108 77
rect 28315 -1862 28379 33748
rect -284 -1926 28379 -1862
rect 28828 -2288 28892 34457
rect -680 -2352 28892 -2288
rect 29407 -2703 29471 35193
rect -1133 -2767 29471 -2703
rect 29990 -3060 30054 35905
rect -1504 -3124 30054 -3060
rect 21201 -3509 21267 -3508
rect 30584 -3509 30648 36528
rect 21201 -3573 21202 -3509
rect 21266 -3573 30648 -3509
rect 21201 -3574 21267 -3573
rect 21201 -3981 21267 -3980
rect 31231 -3981 31295 37164
rect 21201 -4045 21202 -3981
rect 21266 -4045 31295 -3981
rect 21201 -4046 21267 -4045
rect 21201 -4516 21267 -4515
rect 31824 -4516 31888 37773
rect 21201 -4580 21202 -4516
rect 21266 -4580 31888 -4516
rect 21201 -4581 21267 -4580
rect 21201 -4979 21267 -4978
rect 32414 -4979 32478 38353
rect 32791 24132 33254 24134
rect 32791 23896 32904 24132
rect 33140 24048 33254 24132
rect 33140 23984 35216 24048
rect 33140 23896 33254 23984
rect 32791 23894 33254 23896
rect 35152 23867 35216 23984
rect 35151 23866 35217 23867
rect 35151 23802 35152 23866
rect 35216 23802 35217 23866
rect 35151 23801 35217 23802
rect 32790 21672 33253 21674
rect 32790 21436 32903 21672
rect 33139 21585 33253 21672
rect 35151 21585 35217 21586
rect 33139 21521 35152 21585
rect 35216 21521 35217 21585
rect 33139 21436 33253 21521
rect 35151 21520 35217 21521
rect 32790 21434 33253 21436
rect 35477 21380 35541 68015
rect 36066 24019 36130 68638
rect 36065 24018 36131 24019
rect 36065 23954 36066 24018
rect 36130 23954 36131 24018
rect 36065 23953 36131 23954
rect 35476 21379 35542 21380
rect 35476 21315 35477 21379
rect 35541 21315 35542 21379
rect 35476 21314 35542 21315
rect 35477 8532 35541 21314
rect 36066 9155 36130 23953
rect 36065 9154 36131 9155
rect 36065 9090 36066 9154
rect 36130 9090 36131 9154
rect 36065 9089 36131 9090
rect 35477 8531 35554 8532
rect 35477 8467 35489 8531
rect 35553 8467 35554 8531
rect 35477 8466 35554 8467
rect 32793 7291 33256 7293
rect 32793 7055 32906 7291
rect 33142 7223 33256 7291
rect 35027 7223 35093 7224
rect 33142 7159 35028 7223
rect 35092 7159 35093 7223
rect 33142 7055 33256 7159
rect 35027 7158 35093 7159
rect 32793 7053 33256 7055
rect 32784 5991 33247 5993
rect 32784 5755 32897 5991
rect 33133 5885 33247 5991
rect 35026 5885 35092 5886
rect 33133 5821 35027 5885
rect 35091 5821 35092 5885
rect 33133 5755 33247 5821
rect 35026 5820 35092 5821
rect 32784 5753 33247 5755
rect 32790 4576 33253 4578
rect 32790 4340 32903 4576
rect 33139 4492 33253 4576
rect 35034 4492 35100 4493
rect 33139 4428 35035 4492
rect 35099 4428 35100 4492
rect 33139 4340 33253 4428
rect 35034 4427 35100 4428
rect 32790 4338 33253 4340
rect 32786 3203 33249 3205
rect 32786 2967 32899 3203
rect 33135 3122 33249 3203
rect 35030 3122 35096 3123
rect 33135 3058 35031 3122
rect 35095 3058 35096 3122
rect 33135 2967 33249 3058
rect 35030 3057 35096 3058
rect 32786 2965 33249 2967
rect 35477 1592 35541 8466
rect 36066 2215 36130 9089
rect 36631 8470 36695 69258
rect 44736 45172 45324 45179
rect 44736 45072 44908 45172
rect 45144 45072 45324 45172
rect 44736 45008 44758 45072
rect 44822 45008 44838 45072
rect 44902 45008 44908 45072
rect 45144 45008 45158 45072
rect 45222 45008 45238 45072
rect 45302 45008 45324 45072
rect 44736 44936 44908 45008
rect 45144 44936 45324 45008
rect 44736 44931 45324 44936
rect 41587 44528 41827 44551
rect 41515 44526 41875 44528
rect 41515 44462 41543 44526
rect 41607 44462 41623 44526
rect 41687 44462 41703 44526
rect 41767 44462 41783 44526
rect 41847 44462 41875 44526
rect 41515 44461 41875 44462
rect 41587 44304 41827 44461
rect 40800 44302 41827 44304
rect 40800 44066 40913 44302
rect 41149 44066 41827 44302
rect 40800 44064 41827 44066
rect 41587 43378 41827 44064
rect 44795 44011 45258 44013
rect 44795 43926 44908 44011
rect 44765 43921 44908 43926
rect 45144 43926 45258 44011
rect 45144 43921 45294 43926
rect 44765 43857 44797 43921
rect 44861 43857 44877 43921
rect 45181 43857 45197 43921
rect 45261 43857 45294 43921
rect 44765 43853 44908 43857
rect 44795 43775 44908 43853
rect 45144 43853 45294 43857
rect 45144 43775 45258 43853
rect 44795 43773 45258 43775
rect 41513 43376 41873 43378
rect 41513 43312 41541 43376
rect 41605 43312 41621 43376
rect 41685 43312 41701 43376
rect 41765 43312 41781 43376
rect 41845 43312 41873 43376
rect 41513 43311 41873 43312
rect 41587 43295 41827 43311
rect 44779 41502 45242 41504
rect 44779 41384 44892 41502
rect 44755 41379 44892 41384
rect 45128 41384 45242 41502
rect 45128 41379 45284 41384
rect 44755 41315 44787 41379
rect 44851 41315 44867 41379
rect 45171 41315 45187 41379
rect 45251 41315 45284 41379
rect 44755 41311 44892 41315
rect 44779 41266 44892 41311
rect 45128 41311 45284 41315
rect 45128 41266 45242 41311
rect 44779 41264 45242 41266
rect 41494 40837 41734 40855
rect 41431 40835 41791 40837
rect 41431 40771 41459 40835
rect 41523 40771 41539 40835
rect 41603 40771 41619 40835
rect 41683 40771 41699 40835
rect 41763 40771 41791 40835
rect 41431 40770 41791 40771
rect 41494 40559 41734 40770
rect 40808 40557 41734 40559
rect 40808 40321 40921 40557
rect 41157 40321 41734 40557
rect 40808 40319 41734 40321
rect 41494 39568 41734 40319
rect 44772 40191 45235 40193
rect 44772 40114 44885 40191
rect 44755 40109 44885 40114
rect 45121 40114 45235 40191
rect 45121 40109 45284 40114
rect 44755 40045 44787 40109
rect 44851 40045 44867 40109
rect 45171 40045 45187 40109
rect 45251 40045 45284 40109
rect 44755 40041 44885 40045
rect 44772 39955 44885 40041
rect 45121 40041 45284 40045
rect 45121 39955 45235 40041
rect 44772 39953 45235 39955
rect 41429 39566 41789 39568
rect 41429 39502 41457 39566
rect 41521 39502 41537 39566
rect 41601 39502 41617 39566
rect 41681 39502 41697 39566
rect 41761 39502 41789 39566
rect 41429 39501 41789 39502
rect 41494 39483 41734 39501
rect 42785 24250 46299 24252
rect 42785 24151 44914 24250
rect 45150 24151 46299 24250
rect 42785 24087 42891 24151
rect 42955 24087 42971 24151
rect 43035 24087 43051 24151
rect 43115 24087 43131 24151
rect 43195 24087 43211 24151
rect 43275 24087 43291 24151
rect 43355 24087 43371 24151
rect 43435 24087 43451 24151
rect 43515 24087 43531 24151
rect 43595 24087 43611 24151
rect 43675 24087 43691 24151
rect 43755 24087 43771 24151
rect 43835 24087 43851 24151
rect 43915 24087 43931 24151
rect 43995 24087 44011 24151
rect 44075 24087 44091 24151
rect 44155 24087 44171 24151
rect 44235 24087 44251 24151
rect 44315 24087 44331 24151
rect 44395 24087 44411 24151
rect 44475 24087 44491 24151
rect 44555 24087 44571 24151
rect 44635 24087 44651 24151
rect 44715 24087 44731 24151
rect 44795 24087 44811 24151
rect 44875 24087 44891 24151
rect 45195 24087 45211 24151
rect 45275 24087 45291 24151
rect 45355 24087 45371 24151
rect 45435 24087 45451 24151
rect 45515 24087 45531 24151
rect 45595 24087 45611 24151
rect 45675 24087 45691 24151
rect 45755 24087 45771 24151
rect 45835 24087 45851 24151
rect 45915 24087 45931 24151
rect 45995 24087 46011 24151
rect 46075 24087 46091 24151
rect 46155 24087 46299 24151
rect 42785 24014 44914 24087
rect 45150 24014 46299 24087
rect 42785 24012 46299 24014
rect 37661 23675 40175 23728
rect 37661 23611 39351 23675
rect 39415 23611 40175 23675
rect 37661 23595 40175 23611
rect 37661 23583 39351 23595
rect 37661 23519 37823 23583
rect 37887 23531 39351 23583
rect 39415 23531 40175 23595
rect 37887 23519 40175 23531
rect 37661 23488 40175 23519
rect 37818 23190 37906 23195
rect 39334 23190 39422 23201
rect 37274 23188 39497 23190
rect 37274 23182 39346 23188
rect 37274 23118 37830 23182
rect 37894 23124 39346 23182
rect 39410 23124 39497 23188
rect 37894 23118 39497 23124
rect 37274 23108 39497 23118
rect 37274 23102 39346 23108
rect 37274 23038 37830 23102
rect 37894 23044 39346 23102
rect 39410 23044 39497 23108
rect 37894 23038 39497 23044
rect 37274 23028 39497 23038
rect 37274 23022 39346 23028
rect 37274 22958 37830 23022
rect 37894 22964 39346 23022
rect 39410 22964 39497 23028
rect 37894 22958 39497 22964
rect 37274 22954 39497 22958
rect 37274 22816 37510 22954
rect 37818 22945 37906 22954
rect 39334 22951 39422 22954
rect 36913 22815 37510 22816
rect 36913 22579 36917 22815
rect 37153 22580 37510 22815
rect 37153 22579 37157 22580
rect 36913 22578 37157 22579
rect 37274 21827 37510 22580
rect 39935 22732 40175 23488
rect 39935 22730 41264 22732
rect 39935 22494 40914 22730
rect 41150 22494 41264 22730
rect 39935 22492 41264 22494
rect 39935 22402 40175 22492
rect 37732 22349 40175 22402
rect 37732 22285 39351 22349
rect 39415 22285 40175 22349
rect 37732 22269 40175 22285
rect 37732 22247 39351 22269
rect 37732 22183 37829 22247
rect 37893 22205 39351 22247
rect 39415 22205 40175 22269
rect 37893 22183 40175 22205
rect 37732 22162 40175 22183
rect 37825 22150 37897 22162
rect 39340 21827 39428 21835
rect 37274 21822 39497 21827
rect 37274 21794 39352 21822
rect 37274 21730 37824 21794
rect 37888 21758 39352 21794
rect 39416 21758 39497 21822
rect 37888 21742 39497 21758
rect 37888 21730 39352 21742
rect 37274 21714 39352 21730
rect 37274 21650 37824 21714
rect 37888 21678 39352 21714
rect 39416 21678 39497 21742
rect 37888 21662 39497 21678
rect 37888 21650 39352 21662
rect 37274 21598 39352 21650
rect 39416 21598 39497 21662
rect 37274 21591 39497 21598
rect 39340 21585 39428 21591
rect 48791 21244 49254 21245
rect 42729 21243 49254 21244
rect 42729 21155 48904 21243
rect 42729 21091 42889 21155
rect 42953 21091 42969 21155
rect 43033 21091 43049 21155
rect 43113 21091 43129 21155
rect 43193 21091 43209 21155
rect 43273 21091 43289 21155
rect 43353 21091 43369 21155
rect 43433 21091 43449 21155
rect 43513 21091 43529 21155
rect 43593 21091 43609 21155
rect 43673 21091 43689 21155
rect 43753 21091 43769 21155
rect 43833 21091 43849 21155
rect 43913 21091 43929 21155
rect 43993 21091 44009 21155
rect 44073 21091 44089 21155
rect 44153 21091 44169 21155
rect 44233 21091 44249 21155
rect 44313 21091 44329 21155
rect 44393 21091 44409 21155
rect 44473 21091 44489 21155
rect 44553 21091 44569 21155
rect 44633 21091 44649 21155
rect 44713 21091 44729 21155
rect 44793 21091 44809 21155
rect 44873 21091 44889 21155
rect 44953 21091 44969 21155
rect 45033 21091 45049 21155
rect 45113 21091 45129 21155
rect 45193 21091 45209 21155
rect 45273 21091 45289 21155
rect 45353 21091 45369 21155
rect 45433 21091 45449 21155
rect 45513 21091 45529 21155
rect 45593 21091 45609 21155
rect 45673 21091 45689 21155
rect 45753 21091 45769 21155
rect 45833 21091 45849 21155
rect 45913 21091 45929 21155
rect 45993 21091 46009 21155
rect 46073 21091 46089 21155
rect 46153 21091 48904 21155
rect 42729 21007 48904 21091
rect 49140 21007 49254 21243
rect 42729 21005 49254 21007
rect 42729 21004 49031 21005
rect 36881 8791 37155 8810
rect 36881 8555 36900 8791
rect 37136 8555 37155 8791
rect 36881 8537 37155 8555
rect 36630 8469 36696 8470
rect 36630 8405 36631 8469
rect 36695 8405 36696 8469
rect 36630 8404 36696 8405
rect 36065 2214 36131 2215
rect 36065 2150 36066 2214
rect 36130 2150 36131 2214
rect 36065 2149 36131 2150
rect 36066 2136 36130 2149
rect 35477 1591 35554 1592
rect 35477 1527 35489 1591
rect 35553 1527 35554 1591
rect 36631 1530 36695 8404
rect 36971 7350 37067 8537
rect 37895 7593 38131 8554
rect 37895 7541 38667 7593
rect 37895 7477 38576 7541
rect 38640 7477 38667 7541
rect 37895 7461 38667 7477
rect 37895 7397 38576 7461
rect 38640 7397 38667 7461
rect 37895 7357 38667 7397
rect 39402 7590 39638 8553
rect 39402 7554 40189 7590
rect 39402 7490 40095 7554
rect 40159 7490 40189 7554
rect 39402 7474 40189 7490
rect 39402 7410 40095 7474
rect 40159 7410 40189 7474
rect 36970 7333 37068 7350
rect 36970 7269 36987 7333
rect 37051 7269 37068 7333
rect 36970 7252 37068 7269
rect 36971 6525 37067 7252
rect 37895 7138 38131 7357
rect 37894 6902 38131 7138
rect 37895 6525 38131 6902
rect 39402 7354 40189 7410
rect 44796 7444 45259 7446
rect 39402 6525 39638 7354
rect 44796 7233 44909 7444
rect 42601 7219 44909 7233
rect 45145 7233 45259 7444
rect 45145 7219 45924 7233
rect 40800 7168 41265 7171
rect 40800 7162 40914 7168
rect 41150 7162 41265 7168
rect 40800 6938 40840 7162
rect 41224 6938 41265 7162
rect 42601 7155 42630 7219
rect 42694 7155 42710 7219
rect 42774 7155 42790 7219
rect 42854 7155 42870 7219
rect 42934 7155 42950 7219
rect 43014 7155 43030 7219
rect 43094 7155 43110 7219
rect 43174 7155 43190 7219
rect 43254 7155 43270 7219
rect 43334 7155 43350 7219
rect 43414 7155 43430 7219
rect 43494 7155 43510 7219
rect 43574 7155 43590 7219
rect 43654 7155 43670 7219
rect 43734 7155 43750 7219
rect 43814 7155 43830 7219
rect 43894 7155 43910 7219
rect 43974 7155 43990 7219
rect 44054 7155 44070 7219
rect 44134 7155 44150 7219
rect 44214 7155 44230 7219
rect 44294 7155 44310 7219
rect 44374 7155 44390 7219
rect 44454 7155 44470 7219
rect 44534 7155 44550 7219
rect 44614 7155 44630 7219
rect 44694 7155 44710 7219
rect 44774 7155 44790 7219
rect 44854 7155 44870 7219
rect 44934 7155 44950 7208
rect 45014 7155 45030 7208
rect 45094 7155 45110 7208
rect 45174 7155 45190 7219
rect 45254 7155 45270 7219
rect 45334 7155 45350 7219
rect 45414 7155 45430 7219
rect 45494 7155 45510 7219
rect 45574 7155 45590 7219
rect 45654 7155 45670 7219
rect 45734 7155 45750 7219
rect 45814 7155 45830 7219
rect 45894 7155 45924 7219
rect 42601 7142 45924 7155
rect 40800 6932 40914 6938
rect 41150 6932 41265 6938
rect 40800 6929 41265 6932
rect 36938 6289 36941 6525
rect 37177 6289 39638 6525
rect 36970 6249 37068 6289
rect 36970 6185 36987 6249
rect 37051 6185 37068 6249
rect 36970 6168 37068 6185
rect 36971 5178 37067 6168
rect 36970 5161 37068 5178
rect 36970 5109 36987 5161
rect 37051 5109 37068 5161
rect 37895 5109 38131 6289
rect 38562 6210 38646 6289
rect 38562 6146 38571 6210
rect 38635 6205 38646 6210
rect 39402 6275 39638 6289
rect 39402 6207 40175 6275
rect 38635 6146 38645 6205
rect 38562 6130 38645 6146
rect 38562 6066 38571 6130
rect 38635 6066 38645 6130
rect 38562 6043 38645 6066
rect 39402 6143 40100 6207
rect 40164 6143 40175 6207
rect 39402 6127 40175 6143
rect 39402 6063 40100 6127
rect 40164 6063 40175 6127
rect 39402 6039 40175 6063
rect 39402 5109 39638 6039
rect 36899 4873 36902 5109
rect 37138 4873 39638 5109
rect 36971 4090 37067 4873
rect 36971 4073 37069 4090
rect 36971 4009 36988 4073
rect 37052 4009 37069 4073
rect 36971 3992 37069 4009
rect 36971 2832 37067 3992
rect 37895 3500 38131 4873
rect 38561 4857 38644 4873
rect 38561 4793 38570 4857
rect 38634 4793 38644 4857
rect 38561 4777 38644 4793
rect 38561 4713 38570 4777
rect 38634 4713 38644 4777
rect 38561 4690 38644 4713
rect 39402 4835 40189 4873
rect 39402 4771 40100 4835
rect 40164 4771 40189 4835
rect 39402 4755 40189 4771
rect 39402 4691 40100 4755
rect 40164 4691 40189 4755
rect 39402 4637 40189 4691
rect 39402 3503 39638 4637
rect 40798 4267 41263 4268
rect 40798 4265 46002 4267
rect 40798 4259 40912 4265
rect 41148 4259 46002 4265
rect 40798 4035 40838 4259
rect 41222 4220 46002 4259
rect 41222 4156 42607 4220
rect 42671 4156 42687 4220
rect 42751 4156 42767 4220
rect 42831 4156 42847 4220
rect 42911 4156 42927 4220
rect 42991 4156 43007 4220
rect 43071 4156 43087 4220
rect 43151 4156 43167 4220
rect 43231 4156 43247 4220
rect 43311 4156 43327 4220
rect 43391 4156 43407 4220
rect 43471 4156 43487 4220
rect 43551 4156 43567 4220
rect 43631 4156 43647 4220
rect 43711 4156 43727 4220
rect 43791 4156 43807 4220
rect 43871 4156 43887 4220
rect 43951 4156 43967 4220
rect 44031 4156 44047 4220
rect 44111 4156 44127 4220
rect 44191 4156 44207 4220
rect 44271 4156 44287 4220
rect 44351 4156 44367 4220
rect 44431 4156 44447 4220
rect 44511 4156 44527 4220
rect 44591 4156 44607 4220
rect 44671 4156 44687 4220
rect 44751 4156 44767 4220
rect 44831 4156 44847 4220
rect 44911 4156 44927 4220
rect 44991 4156 45007 4220
rect 45071 4156 45087 4220
rect 45151 4156 45167 4220
rect 45231 4156 45247 4220
rect 45311 4156 45327 4220
rect 45391 4156 45407 4220
rect 45471 4156 45487 4220
rect 45551 4156 45567 4220
rect 45631 4156 45647 4220
rect 45711 4156 45727 4220
rect 45791 4156 45807 4220
rect 45871 4156 45887 4220
rect 45951 4156 46002 4220
rect 41222 4035 46002 4156
rect 40798 4029 40912 4035
rect 41148 4029 46002 4035
rect 40798 4027 46002 4029
rect 40798 4026 41263 4027
rect 37895 3480 38646 3500
rect 37895 3457 38647 3480
rect 37895 3393 38573 3457
rect 38637 3393 38647 3457
rect 37895 3377 38647 3393
rect 37895 3313 38573 3377
rect 38637 3313 38647 3377
rect 37895 3290 38647 3313
rect 39402 3451 40187 3503
rect 39402 3387 40097 3451
rect 40161 3387 40187 3451
rect 39402 3371 40187 3387
rect 39402 3307 40097 3371
rect 40161 3307 40187 3371
rect 37895 3264 38646 3290
rect 39402 3267 40187 3307
rect 36889 2813 37163 2832
rect 36889 2577 36908 2813
rect 37144 2577 37163 2813
rect 37895 2750 38131 3264
rect 39402 2820 39638 3267
rect 36889 2559 37163 2577
rect 36881 1851 37155 1870
rect 36881 1615 36900 1851
rect 37136 1615 37155 1851
rect 36881 1597 37155 1615
rect 35477 1526 35554 1527
rect 36630 1529 36696 1530
rect 35477 1493 35541 1526
rect 36630 1465 36631 1529
rect 36695 1465 36696 1529
rect 36630 1464 36696 1465
rect 36631 1436 36695 1464
rect 36971 410 37067 1597
rect 37895 653 38131 1614
rect 37895 601 38667 653
rect 37895 537 38576 601
rect 38640 537 38667 601
rect 37895 521 38667 537
rect 37895 457 38576 521
rect 38640 457 38667 521
rect 37895 417 38667 457
rect 39402 650 39638 1613
rect 39402 614 40189 650
rect 39402 550 40095 614
rect 40159 550 40189 614
rect 39402 534 40189 550
rect 39402 470 40095 534
rect 40159 470 40189 534
rect 36970 393 37068 410
rect 32793 351 33256 353
rect 32793 115 32906 351
rect 33142 283 33256 351
rect 36970 329 36987 393
rect 37051 329 37068 393
rect 36970 312 37068 329
rect 35027 283 35093 284
rect 33142 219 35028 283
rect 35092 219 35093 283
rect 33142 115 33256 219
rect 35027 218 35093 219
rect 32793 113 33256 115
rect 36971 -415 37067 312
rect 37895 198 38131 417
rect 37894 -38 38131 198
rect 37895 -415 38131 -38
rect 39402 414 40189 470
rect 44799 519 45262 521
rect 39402 -415 39638 414
rect 44799 310 44912 519
rect 42598 286 44912 310
rect 45148 310 45262 519
rect 45148 286 45931 310
rect 40800 228 41265 231
rect 40800 222 40914 228
rect 41150 222 41265 228
rect 40800 -2 40840 222
rect 41224 -2 41265 222
rect 42598 222 42632 286
rect 42696 222 42712 286
rect 42776 222 42792 286
rect 42856 222 42872 286
rect 42936 222 42952 286
rect 43016 222 43032 286
rect 43096 222 43112 286
rect 43176 222 43192 286
rect 43256 222 43272 286
rect 43336 222 43352 286
rect 43416 222 43432 286
rect 43496 222 43512 286
rect 43576 222 43592 286
rect 43656 222 43672 286
rect 43736 222 43752 286
rect 43816 222 43832 286
rect 43896 222 43912 286
rect 43976 222 43992 286
rect 44056 222 44072 286
rect 44136 222 44152 286
rect 44216 222 44232 286
rect 44296 222 44312 286
rect 44376 222 44392 286
rect 44456 222 44472 286
rect 44536 222 44552 286
rect 44616 222 44632 286
rect 44696 222 44712 286
rect 44776 222 44792 286
rect 44856 222 44872 286
rect 44936 222 44952 283
rect 45016 222 45032 283
rect 45096 222 45112 283
rect 45176 222 45192 286
rect 45256 222 45272 286
rect 45336 222 45352 286
rect 45416 222 45432 286
rect 45496 222 45512 286
rect 45576 222 45592 286
rect 45656 222 45672 286
rect 45736 222 45752 286
rect 45816 222 45832 286
rect 45896 222 45931 286
rect 42598 198 45931 222
rect 40800 -8 40914 -2
rect 41150 -8 41265 -2
rect 40800 -11 41265 -8
rect 36938 -651 36941 -415
rect 37177 -651 39638 -415
rect 36970 -691 37068 -651
rect 36970 -755 36987 -691
rect 37051 -755 37068 -691
rect 36970 -772 37068 -755
rect 32784 -949 33247 -947
rect 32784 -1185 32897 -949
rect 33133 -1055 33247 -949
rect 35026 -1055 35092 -1054
rect 33133 -1119 35027 -1055
rect 35091 -1119 35092 -1055
rect 33133 -1185 33247 -1119
rect 35026 -1120 35092 -1119
rect 32784 -1187 33247 -1185
rect 36971 -1762 37067 -772
rect 36970 -1779 37068 -1762
rect 36970 -1831 36987 -1779
rect 37051 -1831 37068 -1779
rect 37895 -1831 38131 -651
rect 38562 -730 38646 -651
rect 38562 -794 38571 -730
rect 38635 -735 38646 -730
rect 39402 -665 39638 -651
rect 39402 -733 40175 -665
rect 38635 -794 38645 -735
rect 38562 -810 38645 -794
rect 38562 -874 38571 -810
rect 38635 -874 38645 -810
rect 38562 -897 38645 -874
rect 39402 -797 40100 -733
rect 40164 -797 40175 -733
rect 39402 -813 40175 -797
rect 39402 -877 40100 -813
rect 40164 -877 40175 -813
rect 39402 -901 40175 -877
rect 39402 -1831 39638 -901
rect 36899 -2067 36902 -1831
rect 37138 -2067 39638 -1831
rect 32790 -2364 33253 -2362
rect 32790 -2600 32903 -2364
rect 33139 -2448 33253 -2364
rect 35034 -2448 35100 -2447
rect 33139 -2512 35035 -2448
rect 35099 -2512 35100 -2448
rect 33139 -2600 33253 -2512
rect 35034 -2513 35100 -2512
rect 32790 -2602 33253 -2600
rect 36971 -2850 37067 -2067
rect 36971 -2867 37069 -2850
rect 36971 -2931 36988 -2867
rect 37052 -2931 37069 -2867
rect 36971 -2948 37069 -2931
rect 32786 -3737 33249 -3735
rect 32786 -3973 32899 -3737
rect 33135 -3818 33249 -3737
rect 35030 -3818 35096 -3817
rect 33135 -3882 35031 -3818
rect 35095 -3882 35096 -3818
rect 33135 -3973 33249 -3882
rect 35030 -3883 35096 -3882
rect 32786 -3975 33249 -3973
rect 36971 -4108 37067 -2948
rect 37895 -3440 38131 -2067
rect 38561 -2083 38644 -2067
rect 38561 -2147 38570 -2083
rect 38634 -2147 38644 -2083
rect 38561 -2163 38644 -2147
rect 38561 -2227 38570 -2163
rect 38634 -2227 38644 -2163
rect 38561 -2250 38644 -2227
rect 39402 -2105 40189 -2067
rect 39402 -2169 40100 -2105
rect 40164 -2169 40189 -2105
rect 39402 -2185 40189 -2169
rect 39402 -2249 40100 -2185
rect 40164 -2249 40189 -2185
rect 39402 -2303 40189 -2249
rect 39402 -3437 39638 -2303
rect 40798 -2673 41263 -2672
rect 40798 -2679 41517 -2673
rect 40798 -2680 40905 -2679
rect 40785 -2681 40905 -2680
rect 41141 -2680 41517 -2679
rect 41141 -2681 46063 -2680
rect 40785 -2905 40838 -2681
rect 41222 -2720 46063 -2681
rect 41222 -2784 42588 -2720
rect 42652 -2784 42668 -2720
rect 42732 -2784 42748 -2720
rect 42812 -2784 42828 -2720
rect 42892 -2784 42908 -2720
rect 42972 -2784 42988 -2720
rect 43052 -2784 43068 -2720
rect 43132 -2784 43148 -2720
rect 43212 -2784 43228 -2720
rect 43292 -2784 43308 -2720
rect 43372 -2784 43388 -2720
rect 43452 -2784 43468 -2720
rect 43532 -2784 43548 -2720
rect 43612 -2784 43628 -2720
rect 43692 -2784 43708 -2720
rect 43772 -2784 43788 -2720
rect 43852 -2784 43868 -2720
rect 43932 -2784 43948 -2720
rect 44012 -2784 44028 -2720
rect 44092 -2784 44108 -2720
rect 44172 -2784 44188 -2720
rect 44252 -2784 44268 -2720
rect 44332 -2784 44348 -2720
rect 44412 -2784 44428 -2720
rect 44492 -2784 44508 -2720
rect 44572 -2784 44588 -2720
rect 44652 -2784 44668 -2720
rect 44732 -2784 44748 -2720
rect 44812 -2784 44828 -2720
rect 44892 -2784 44908 -2720
rect 44972 -2784 44988 -2720
rect 45052 -2784 45068 -2720
rect 45132 -2784 45148 -2720
rect 45212 -2784 45228 -2720
rect 45292 -2784 45308 -2720
rect 45372 -2784 45388 -2720
rect 45452 -2784 45468 -2720
rect 45532 -2784 45548 -2720
rect 45612 -2784 45628 -2720
rect 45692 -2784 45708 -2720
rect 45772 -2784 45788 -2720
rect 45852 -2784 45868 -2720
rect 45932 -2784 46063 -2720
rect 41222 -2905 46063 -2784
rect 40785 -2915 40905 -2905
rect 41141 -2915 46063 -2905
rect 40785 -2920 46063 -2915
rect 37895 -3460 38646 -3440
rect 37895 -3483 38647 -3460
rect 37895 -3547 38573 -3483
rect 38637 -3547 38647 -3483
rect 37895 -3563 38647 -3547
rect 37895 -3627 38573 -3563
rect 38637 -3627 38647 -3563
rect 37895 -3650 38647 -3627
rect 39402 -3489 40187 -3437
rect 39402 -3553 40097 -3489
rect 40161 -3553 40187 -3489
rect 39402 -3569 40187 -3553
rect 39402 -3633 40097 -3569
rect 40161 -3633 40187 -3569
rect 37895 -3676 38646 -3650
rect 39402 -3673 40187 -3633
rect 36889 -4127 37163 -4108
rect 36889 -4363 36908 -4127
rect 37144 -4363 37163 -4127
rect 37895 -4190 38131 -3676
rect 39402 -4120 39638 -3673
rect 36889 -4381 37163 -4363
rect 21201 -5043 21202 -4979
rect 21266 -5043 32478 -4979
rect 21201 -5044 21267 -5043
rect -3198 -6175 -487 -6173
rect -3198 -6411 -3085 -6175
rect -2849 -6411 -487 -6175
rect -3198 -6413 -487 -6411
rect -3596 -6844 -3502 -6821
rect -600 -6824 -487 -6413
rect -3596 -6908 -3581 -6844
rect -3517 -6908 -3502 -6844
rect -3596 -6924 -3502 -6908
rect -3596 -6988 -3581 -6924
rect -3517 -6988 -3502 -6924
rect -3596 -7004 -3502 -6988
rect -3596 -7068 -3581 -7004
rect -3517 -7068 -3502 -7004
rect -3596 -7084 -3502 -7068
rect -3596 -7148 -3581 -7084
rect -3517 -7148 -3502 -7084
rect -3596 -7164 -3502 -7148
rect -3596 -7228 -3581 -7164
rect -3517 -7228 -3502 -7164
rect -3596 -7244 -3502 -7228
rect -3596 -7308 -3581 -7244
rect -3517 -7308 -3502 -7244
rect -3596 -7324 -3502 -7308
rect -3596 -7388 -3581 -7324
rect -3517 -7388 -3502 -7324
rect -3596 -7404 -3502 -7388
rect -3596 -7468 -3581 -7404
rect -3517 -7468 -3502 -7404
rect -3596 -7484 -3502 -7468
rect -3596 -7548 -3581 -7484
rect -3517 -7548 -3502 -7484
rect -3596 -7564 -3502 -7548
rect -3596 -7628 -3581 -7564
rect -3517 -7628 -3502 -7564
rect -3596 -7644 -3502 -7628
rect -3596 -7708 -3581 -7644
rect -3517 -7708 -3502 -7644
rect -3596 -7724 -3502 -7708
rect -3596 -7788 -3581 -7724
rect -3517 -7788 -3502 -7724
rect -3596 -7804 -3502 -7788
rect -3596 -7868 -3581 -7804
rect -3517 -7868 -3502 -7804
rect -3596 -7884 -3502 -7868
rect -3596 -7948 -3581 -7884
rect -3517 -7948 -3502 -7884
rect -3596 -7964 -3502 -7948
rect -3596 -8028 -3581 -7964
rect -3517 -8028 -3502 -7964
rect -3596 -8044 -3502 -8028
rect -3596 -8108 -3581 -8044
rect -3517 -8108 -3502 -8044
rect -3596 -8124 -3502 -8108
rect -3596 -8188 -3581 -8124
rect -3517 -8188 -3502 -8124
rect -3596 -8204 -3502 -8188
rect -3596 -8268 -3581 -8204
rect -3517 -8268 -3502 -8204
rect -3596 -8276 -3502 -8268
rect -601 -6851 -485 -6824
rect -601 -6915 -575 -6851
rect -511 -6915 -485 -6851
rect -601 -6931 -485 -6915
rect -601 -6995 -575 -6931
rect -511 -6995 -485 -6931
rect -601 -7011 -485 -6995
rect -601 -7075 -575 -7011
rect -511 -7075 -485 -7011
rect -601 -7091 -485 -7075
rect -601 -7155 -575 -7091
rect -511 -7155 -485 -7091
rect -601 -7171 -485 -7155
rect -601 -7235 -575 -7171
rect -511 -7235 -485 -7171
rect -601 -7251 -485 -7235
rect -601 -7315 -575 -7251
rect -511 -7315 -485 -7251
rect -601 -7331 -485 -7315
rect -601 -7395 -575 -7331
rect -511 -7395 -485 -7331
rect -601 -7411 -485 -7395
rect -601 -7475 -575 -7411
rect -511 -7475 -485 -7411
rect -601 -7491 -485 -7475
rect -601 -7555 -575 -7491
rect -511 -7555 -485 -7491
rect -601 -7571 -485 -7555
rect -601 -7635 -575 -7571
rect -511 -7635 -485 -7571
rect -601 -7651 -485 -7635
rect -601 -7715 -575 -7651
rect -511 -7715 -485 -7651
rect -601 -7731 -485 -7715
rect -601 -7795 -575 -7731
rect -511 -7795 -485 -7731
rect -601 -7811 -485 -7795
rect -601 -7875 -575 -7811
rect -511 -7875 -485 -7811
rect -601 -7891 -485 -7875
rect -601 -7955 -575 -7891
rect -511 -7955 -485 -7891
rect -601 -7971 -485 -7955
rect -601 -8035 -575 -7971
rect -511 -8035 -485 -7971
rect -601 -8051 -485 -8035
rect -601 -8115 -575 -8051
rect -511 -8115 -485 -8051
rect -601 -8131 -485 -8115
rect -601 -8195 -575 -8131
rect -511 -8195 -485 -8131
rect -601 -8211 -485 -8195
rect -601 -8275 -575 -8211
rect -511 -8275 -485 -8211
rect -7204 -8278 -3494 -8276
rect -7204 -8514 -7091 -8278
rect -6855 -8284 -3494 -8278
rect -6855 -8348 -3581 -8284
rect -3517 -8348 -3494 -8284
rect -6855 -8364 -3494 -8348
rect -6855 -8428 -3581 -8364
rect -3517 -8428 -3494 -8364
rect -6855 -8444 -3494 -8428
rect -6855 -8508 -3581 -8444
rect -3517 -8508 -3494 -8444
rect -6855 -8514 -3494 -8508
rect -7204 -8516 -3494 -8514
rect -601 -8291 -485 -8275
rect -601 -8355 -575 -8291
rect -511 -8355 -485 -8291
rect -601 -8371 -485 -8355
rect -601 -8435 -575 -8371
rect -511 -8435 -485 -8371
rect -601 -8451 -485 -8435
rect -601 -8515 -575 -8451
rect -511 -8515 -485 -8451
rect -3596 -8524 -3502 -8516
rect -3596 -8588 -3581 -8524
rect -3517 -8588 -3502 -8524
rect -3596 -8604 -3502 -8588
rect -3596 -8668 -3581 -8604
rect -3517 -8668 -3502 -8604
rect -3596 -8684 -3502 -8668
rect -3596 -8748 -3581 -8684
rect -3517 -8748 -3502 -8684
rect -3596 -8764 -3502 -8748
rect -3596 -8828 -3581 -8764
rect -3517 -8828 -3502 -8764
rect -3596 -8844 -3502 -8828
rect -3596 -8908 -3581 -8844
rect -3517 -8908 -3502 -8844
rect -3596 -8924 -3502 -8908
rect -3596 -8988 -3581 -8924
rect -3517 -8988 -3502 -8924
rect -3596 -9004 -3502 -8988
rect -3596 -9068 -3581 -9004
rect -3517 -9068 -3502 -9004
rect -3596 -9084 -3502 -9068
rect -3596 -9148 -3581 -9084
rect -3517 -9148 -3502 -9084
rect -3596 -9164 -3502 -9148
rect -3596 -9228 -3581 -9164
rect -3517 -9228 -3502 -9164
rect -3596 -9244 -3502 -9228
rect -3596 -9308 -3581 -9244
rect -3517 -9308 -3502 -9244
rect -3596 -9324 -3502 -9308
rect -3596 -9388 -3581 -9324
rect -3517 -9388 -3502 -9324
rect -3596 -9404 -3502 -9388
rect -3596 -9468 -3581 -9404
rect -3517 -9468 -3502 -9404
rect -3596 -9484 -3502 -9468
rect -3596 -9548 -3581 -9484
rect -3517 -9548 -3502 -9484
rect -3596 -9564 -3502 -9548
rect -3596 -9628 -3581 -9564
rect -3517 -9628 -3502 -9564
rect -3596 -9644 -3502 -9628
rect -3596 -9708 -3581 -9644
rect -3517 -9708 -3502 -9644
rect -3596 -9724 -3502 -9708
rect -3596 -9788 -3581 -9724
rect -3517 -9788 -3502 -9724
rect -3596 -9804 -3502 -9788
rect -3596 -9868 -3581 -9804
rect -3517 -9868 -3502 -9804
rect -3596 -9884 -3502 -9868
rect -3596 -9948 -3581 -9884
rect -3517 -9948 -3502 -9884
rect -3596 -9964 -3502 -9948
rect -3596 -10028 -3581 -9964
rect -3517 -10028 -3502 -9964
rect -3596 -10044 -3502 -10028
rect -3596 -10108 -3581 -10044
rect -3517 -10108 -3502 -10044
rect -3596 -10131 -3502 -10108
rect -601 -8531 -485 -8515
rect -601 -8595 -575 -8531
rect -511 -8595 -485 -8531
rect -601 -8611 -485 -8595
rect -601 -8675 -575 -8611
rect -511 -8675 -485 -8611
rect -601 -8691 -485 -8675
rect -601 -8755 -575 -8691
rect -511 -8755 -485 -8691
rect -601 -8771 -485 -8755
rect -601 -8835 -575 -8771
rect -511 -8835 -485 -8771
rect -601 -8851 -485 -8835
rect -601 -8915 -575 -8851
rect -511 -8915 -485 -8851
rect -601 -8931 -485 -8915
rect -601 -8995 -575 -8931
rect -511 -8995 -485 -8931
rect -601 -9011 -485 -8995
rect -601 -9075 -575 -9011
rect -511 -9075 -485 -9011
rect -601 -9091 -485 -9075
rect -601 -9155 -575 -9091
rect -511 -9155 -485 -9091
rect -601 -9171 -485 -9155
rect -601 -9235 -575 -9171
rect -511 -9235 -485 -9171
rect -601 -9251 -485 -9235
rect -601 -9315 -575 -9251
rect -511 -9315 -485 -9251
rect -601 -9331 -485 -9315
rect -601 -9395 -575 -9331
rect -511 -9395 -485 -9331
rect -601 -9411 -485 -9395
rect -601 -9475 -575 -9411
rect -511 -9475 -485 -9411
rect -601 -9491 -485 -9475
rect -601 -9555 -575 -9491
rect -511 -9555 -485 -9491
rect -601 -9571 -485 -9555
rect -601 -9635 -575 -9571
rect -511 -9635 -485 -9571
rect -601 -9651 -485 -9635
rect -601 -9715 -575 -9651
rect -511 -9715 -485 -9651
rect -601 -9731 -485 -9715
rect -601 -9795 -575 -9731
rect -511 -9795 -485 -9731
rect -601 -9811 -485 -9795
rect -601 -9875 -575 -9811
rect -511 -9875 -485 -9811
rect -601 -9891 -485 -9875
rect -601 -9955 -575 -9891
rect -511 -9955 -485 -9891
rect -601 -9971 -485 -9955
rect -601 -10035 -575 -9971
rect -511 -10035 -485 -9971
rect -601 -10051 -485 -10035
rect -601 -10115 -575 -10051
rect -511 -10115 -485 -10051
rect -601 -10141 -485 -10115
rect -57093 -16103 62907 -16021
rect -57093 -17939 -55011 -16103
rect -53175 -17939 -43253 -16103
rect -42697 -17939 -35253 -16103
rect -34697 -17939 -27253 -16103
rect -26697 -17939 -19253 -16103
rect -18697 -17939 -11253 -16103
rect -10697 -17939 -3253 -16103
rect -2697 -17939 4747 -16103
rect 5303 -17939 12747 -16103
rect 13303 -17939 20747 -16103
rect 21303 -17939 28747 -16103
rect 29303 -17939 36747 -16103
rect 37303 -17939 44747 -16103
rect 45303 -17939 54989 -16103
rect 56825 -17939 62907 -16103
rect -57093 -18021 62907 -17939
rect -57093 -20103 62907 -20021
rect -57093 -21939 -51011 -20103
rect -49175 -21939 -39253 -20103
rect -38697 -21939 -31253 -20103
rect -30697 -21939 -23253 -20103
rect -22697 -21939 -15253 -20103
rect -14697 -21939 -7253 -20103
rect -6697 -21939 747 -20103
rect 1303 -21939 8747 -20103
rect 9303 -21939 16747 -20103
rect 17303 -21939 24747 -20103
rect 25303 -21939 32747 -20103
rect 33303 -21939 40747 -20103
rect 41303 -21939 48747 -20103
rect 49303 -21939 58989 -20103
rect 60825 -21939 62907 -20103
rect -57093 -22021 62907 -21939
<< via4 >>
rect -55011 86524 -53175 88360
rect -43253 86524 -42697 88360
rect -35253 86524 -34697 88360
rect -27253 86524 -26697 88360
rect -19253 86524 -18697 88360
rect -11253 86524 -10697 88360
rect -3253 86524 -2697 88360
rect 4747 86524 5303 88360
rect 12747 86524 13303 88360
rect 20747 86524 21303 88360
rect 28747 86524 29303 88360
rect 36747 86524 37303 88360
rect 44747 86524 45303 88360
rect 54989 86524 56825 88360
rect -51011 82524 -49175 84360
rect -39253 82524 -38697 84360
rect -31253 82524 -30697 84360
rect -23253 82524 -22697 84360
rect -15253 82524 -14697 84360
rect -7253 82524 -6697 84360
rect 747 82524 1303 84360
rect 8747 82524 9303 84360
rect 16747 82524 17303 84360
rect 24747 82524 25303 84360
rect 32747 82524 33303 84360
rect 40747 82524 41303 84360
rect 48747 82524 49303 84360
rect 58989 82524 60825 84360
rect -19094 74830 -18858 75066
rect -15096 75015 -14860 75251
rect 12905 74934 13141 75170
rect 16904 74926 17140 75162
rect -15095 70756 -14859 70992
rect -19094 69999 -18858 70235
rect -15092 68677 -14856 68913
rect -19098 66884 -18862 67120
rect -11022 63263 -10786 63499
rect 20907 64337 21143 64573
rect 28901 64343 29137 64579
rect -6937 63198 -6701 63204
rect -6937 62974 -6931 63198
rect -6931 62974 -6707 63198
rect -6707 62974 -6701 63198
rect -6937 62968 -6701 62974
rect -3094 63173 -2858 63409
rect 904 63224 1140 63230
rect 904 63000 1140 63224
rect 904 62994 1140 63000
rect 16910 62346 17146 62582
rect 24906 62339 25142 62575
rect 32909 62335 33145 62571
rect -19091 50596 -18855 50688
rect -19091 50532 -19005 50596
rect -19005 50532 -18941 50596
rect -18941 50532 -18855 50596
rect -19091 50452 -18855 50532
rect -27089 49720 -26853 49824
rect -27089 49656 -27050 49720
rect -27050 49656 -26986 49720
rect -26986 49656 -26970 49720
rect -26970 49656 -26906 49720
rect -26906 49656 -26890 49720
rect -26890 49656 -26853 49720
rect -27089 49588 -26853 49656
rect -23087 48985 -22851 49221
rect -27054 43134 -27007 43154
rect -27007 43134 -26818 43154
rect -27054 43118 -26818 43134
rect -27054 43054 -27007 43118
rect -27007 43054 -26818 43118
rect -27054 43038 -26818 43054
rect -27054 42974 -27007 43038
rect -27007 42974 -26818 43038
rect -27054 42958 -26818 42974
rect -27054 42918 -27007 42958
rect -27007 42918 -26818 42958
rect -6960 55093 -6724 55329
rect -6960 54773 -6724 55009
rect -3090 54184 -2854 54420
rect 903 59886 1139 60122
rect 8908 59875 9144 60111
rect 903 56511 1139 56747
rect 8907 56500 9143 56736
rect 903 53136 1139 53372
rect 8907 53125 9143 53361
rect -7090 51463 -6854 51699
rect -27049 39907 -27002 39948
rect -27002 39907 -26813 39948
rect -27049 39891 -26813 39907
rect -27049 39827 -27002 39891
rect -27002 39827 -26813 39891
rect -27049 39811 -26813 39827
rect -27049 39747 -27002 39811
rect -27002 39747 -26813 39811
rect -27049 39731 -26813 39747
rect -27049 39712 -27002 39731
rect -27002 39712 -26813 39731
rect -35105 38260 -34869 38496
rect -31093 38271 -30857 38507
rect -31105 37173 -30869 37409
rect -23079 37658 -22843 37894
rect -15092 37931 -14856 38167
rect -27049 35820 -27005 35879
rect -27005 35820 -26813 35879
rect -27049 35804 -26813 35820
rect -27049 35740 -27005 35804
rect -27005 35740 -26813 35804
rect -27049 35724 -26813 35740
rect -27049 35660 -27005 35724
rect -27005 35660 -26813 35724
rect -27049 35644 -26813 35660
rect -27049 35643 -27005 35644
rect -27005 35643 -26813 35644
rect -3084 51057 -2848 51099
rect -3084 50913 -2848 51057
rect -3084 50863 -2848 50913
rect -3090 48535 -2854 48771
rect 903 49761 1139 49997
rect 8907 49750 9143 49986
rect 20907 60337 21143 60573
rect 28901 60343 29137 60579
rect 16910 58346 17146 58582
rect 24906 58339 25142 58575
rect 32909 58335 33145 58571
rect 20907 56337 21143 56573
rect 28901 56343 29137 56579
rect 16910 54346 17146 54582
rect 24906 54339 25142 54575
rect 32909 54335 33145 54571
rect 20907 52337 21143 52573
rect 28901 52343 29137 52579
rect 16910 50346 17146 50582
rect 24906 50339 25142 50575
rect 32909 50335 33145 50571
rect 20907 48337 21143 48573
rect 28901 48343 29137 48579
rect -3094 44365 -2858 44601
rect 899 44276 1135 44512
rect 8907 43000 9143 43236
rect -3086 39828 -2850 39884
rect -3086 39684 -2850 39828
rect 909 40631 1145 40867
rect -3086 39648 -2850 39684
rect 903 39202 1139 39438
rect -27051 32720 -27013 32765
rect -27013 32720 -26815 32765
rect -27051 32704 -26815 32720
rect -27051 32640 -27013 32704
rect -27013 32640 -26815 32704
rect -27051 32624 -26815 32640
rect -27051 32560 -27013 32624
rect -27013 32560 -26815 32624
rect -27051 32544 -26815 32560
rect -27051 32529 -27013 32544
rect -27013 32529 -26815 32544
rect -19091 28470 -18855 28706
rect -15087 27205 -14851 27441
rect -35111 26670 -34875 26906
rect -11090 27817 -10854 28053
rect -19099 25799 -18863 25808
rect -19099 25575 -19084 25799
rect -19084 25575 -18863 25799
rect -19099 25572 -18863 25575
rect -15091 25580 -14855 25816
rect -27081 25276 -26845 25512
rect -23089 24679 -22853 24915
rect -39092 23476 -38856 23712
rect -19092 23492 -18856 23728
rect -15090 23401 -14854 23637
rect -11099 22916 -10863 23152
rect -35105 19058 -34869 19231
rect -35105 18995 -35043 19058
rect -35043 18995 -35027 19058
rect -35027 18995 -34963 19058
rect -34963 18995 -34947 19058
rect -34947 18995 -34883 19058
rect -34883 18995 -34869 19058
rect 4908 37815 5144 38051
rect 904 36857 1140 37093
rect 4915 36422 5151 36658
rect 921 35778 1157 36014
rect 8905 35790 9141 36026
rect 4921 35244 5157 35480
rect 4893 23151 5129 23157
rect 4893 22927 5129 23151
rect 4893 22921 5129 22927
rect 8887 23333 9123 23493
rect 8887 23269 8937 23333
rect 8937 23269 9123 23333
rect 8887 23257 9123 23269
rect 16910 46346 17146 46582
rect 24906 46339 25142 46575
rect 32909 46335 33145 46571
rect 4910 19172 5146 19231
rect -27091 17725 -26855 17961
rect -3098 17856 -2862 17862
rect -3098 17632 -2862 17856
rect -3098 17626 -2862 17632
rect -39091 15962 -38855 16198
rect 4910 19028 5146 19172
rect 4910 18995 5146 19028
rect -27084 14239 -26848 14475
rect -23106 15252 -22870 15488
rect -7105 15574 -6869 15810
rect -3088 16212 -2852 16448
rect -7108 14214 -6872 14450
rect -7108 10674 -6872 10910
rect -7098 9424 -6862 9660
rect -7101 7235 -6865 7241
rect -7101 7011 -6865 7235
rect -7101 7005 -6865 7011
rect -27092 6472 -26856 6708
rect -7098 5526 -6862 5762
rect -23085 4806 -22849 5042
rect -3086 13810 -2850 14046
rect -3088 8564 -2852 8800
rect -3086 6505 -2850 6741
rect 902 17525 1138 17616
rect 902 17461 981 17525
rect 981 17461 1045 17525
rect 1045 17461 1138 17525
rect 902 17380 1138 17461
rect 8902 17165 9138 17401
rect 4907 16414 5143 16593
rect 4907 16357 5143 16414
rect 4907 16270 5143 16273
rect 4907 16037 5143 16270
rect 12864 21027 13100 21094
rect 12864 20963 12936 21027
rect 12936 20963 13000 21027
rect 13000 20963 13100 21027
rect 12864 20858 13100 20963
rect 12852 18688 13088 18793
rect 12852 18624 12930 18688
rect 12930 18624 12994 18688
rect 12994 18624 13088 18688
rect 12852 18557 13088 18624
rect 16892 18949 17128 19185
rect 20896 19062 21132 19158
rect 20896 18998 20971 19062
rect 20971 18998 21035 19062
rect 21035 18998 21132 19062
rect 20896 18922 21132 18998
rect 24906 18917 25142 19153
rect 12846 17083 13082 17188
rect 12846 17019 12956 17083
rect 12956 17019 13020 17083
rect 13020 17019 13082 17083
rect 12846 16952 13082 17019
rect 12865 15228 13101 15317
rect 12865 15164 12973 15228
rect 12973 15164 13037 15228
rect 13037 15164 13101 15228
rect 12865 15081 13101 15164
rect 16800 15356 17036 15592
rect 20839 15496 21075 15587
rect 20839 15432 20928 15496
rect 20928 15432 20992 15496
rect 20992 15432 21075 15496
rect 20839 15351 21075 15432
rect 24908 15324 25144 15560
rect 12887 13528 13123 13616
rect 12887 13464 13003 13528
rect 13003 13464 13067 13528
rect 13067 13464 13123 13528
rect 12887 13380 13123 13464
rect 12900 11676 13136 11761
rect 12900 11612 13001 11676
rect 13001 11612 13065 11676
rect 13065 11612 13136 11676
rect 12900 11525 13136 11612
rect 12896 10415 13132 10651
rect 20893 11906 21129 11999
rect 20893 11842 20985 11906
rect 20985 11842 21049 11906
rect 21049 11842 21129 11906
rect 20893 11763 21129 11842
rect 24896 11733 25132 11969
rect 907 221 1143 323
rect 8927 221 9163 335
rect 16904 221 17140 323
rect 907 87 1143 221
rect 8927 99 9163 221
rect 16904 87 17140 221
rect 32904 23896 33140 24132
rect 32903 21436 33139 21672
rect 32906 7055 33142 7291
rect 32897 5755 33133 5991
rect 32903 4340 33139 4576
rect 32899 2967 33135 3203
rect 44908 45072 45144 45172
rect 44908 45008 44918 45072
rect 44918 45008 44982 45072
rect 44982 45008 44998 45072
rect 44998 45008 45062 45072
rect 45062 45008 45078 45072
rect 45078 45008 45142 45072
rect 45142 45008 45144 45072
rect 44908 44936 45144 45008
rect 40913 44066 41149 44302
rect 44908 43921 45144 44011
rect 44908 43857 44941 43921
rect 44941 43857 44957 43921
rect 44957 43857 45021 43921
rect 45021 43857 45037 43921
rect 45037 43857 45101 43921
rect 45101 43857 45117 43921
rect 45117 43857 45144 43921
rect 44908 43775 45144 43857
rect 44892 41379 45128 41502
rect 44892 41315 44931 41379
rect 44931 41315 44947 41379
rect 44947 41315 45011 41379
rect 45011 41315 45027 41379
rect 45027 41315 45091 41379
rect 45091 41315 45107 41379
rect 45107 41315 45128 41379
rect 44892 41266 45128 41315
rect 40921 40321 41157 40557
rect 44885 40109 45121 40191
rect 44885 40045 44931 40109
rect 44931 40045 44947 40109
rect 44947 40045 45011 40109
rect 45011 40045 45027 40109
rect 45027 40045 45091 40109
rect 45091 40045 45107 40109
rect 45107 40045 45121 40109
rect 44885 39955 45121 40045
rect 44914 24151 45150 24250
rect 44914 24087 44955 24151
rect 44955 24087 44971 24151
rect 44971 24087 45035 24151
rect 45035 24087 45051 24151
rect 45051 24087 45115 24151
rect 45115 24087 45131 24151
rect 45131 24087 45150 24151
rect 44914 24014 45150 24087
rect 36917 22809 37153 22815
rect 36917 22585 36923 22809
rect 36923 22585 37147 22809
rect 37147 22585 37153 22809
rect 36917 22579 37153 22585
rect 40914 22494 41150 22730
rect 48904 21007 49140 21243
rect 36900 8786 37136 8791
rect 36900 8562 36907 8786
rect 36907 8562 37131 8786
rect 37131 8562 37136 8786
rect 36900 8555 37136 8562
rect 44909 7219 45145 7444
rect 40914 7162 41150 7168
rect 40914 6938 41150 7162
rect 44909 7208 44934 7219
rect 44934 7208 44950 7219
rect 44950 7208 45014 7219
rect 45014 7208 45030 7219
rect 45030 7208 45094 7219
rect 45094 7208 45110 7219
rect 45110 7208 45145 7219
rect 40914 6932 41150 6938
rect 36941 6289 37177 6525
rect 36902 5097 36987 5109
rect 36987 5097 37051 5109
rect 37051 5097 37138 5109
rect 36902 4873 37138 5097
rect 40912 4259 41148 4265
rect 40912 4035 41148 4259
rect 40912 4029 41148 4035
rect 36908 2577 37144 2813
rect 36900 1846 37136 1851
rect 36900 1622 36907 1846
rect 36907 1622 37131 1846
rect 37131 1622 37136 1846
rect 36900 1615 37136 1622
rect 32906 115 33142 351
rect 44912 286 45148 519
rect 40914 222 41150 228
rect 40914 -2 41150 222
rect 44912 283 44936 286
rect 44936 283 44952 286
rect 44952 283 45016 286
rect 45016 283 45032 286
rect 45032 283 45096 286
rect 45096 283 45112 286
rect 45112 283 45148 286
rect 40914 -8 41150 -2
rect 36941 -651 37177 -415
rect 32897 -1185 33133 -949
rect 36902 -1843 36987 -1831
rect 36987 -1843 37051 -1831
rect 37051 -1843 37138 -1831
rect 36902 -2067 37138 -1843
rect 32903 -2600 33139 -2364
rect 32899 -3973 33135 -3737
rect 40905 -2681 41141 -2679
rect 40905 -2905 41141 -2681
rect 40905 -2915 41141 -2905
rect 36908 -4363 37144 -4127
rect -3085 -6411 -2849 -6175
rect -7091 -8514 -6855 -8278
rect -55011 -17939 -53175 -16103
rect -43253 -17939 -42697 -16103
rect -35253 -17939 -34697 -16103
rect -27253 -17939 -26697 -16103
rect -19253 -17939 -18697 -16103
rect -11253 -17939 -10697 -16103
rect -3253 -17939 -2697 -16103
rect 4747 -17939 5303 -16103
rect 12747 -17939 13303 -16103
rect 20747 -17939 21303 -16103
rect 28747 -17939 29303 -16103
rect 36747 -17939 37303 -16103
rect 44747 -17939 45303 -16103
rect 54989 -17939 56825 -16103
rect -51011 -21939 -49175 -20103
rect -39253 -21939 -38697 -20103
rect -31253 -21939 -30697 -20103
rect -23253 -21939 -22697 -20103
rect -15253 -21939 -14697 -20103
rect -7253 -21939 -6697 -20103
rect 747 -21939 1303 -20103
rect 8747 -21939 9303 -20103
rect 16747 -21939 17303 -20103
rect 24747 -21939 25303 -20103
rect 32747 -21939 33303 -20103
rect 40747 -21939 41303 -20103
rect 48747 -21939 49303 -20103
rect 58989 -21939 60825 -20103
<< metal5 >>
rect -55093 88466 -53093 90442
rect -55117 88360 -53069 88466
rect -55117 86524 -55011 88360
rect -53175 86524 -53069 88360
rect -55117 86418 -53069 86524
rect -55093 -15997 -53093 86418
rect -51093 84466 -49093 90441
rect 54907 88466 56907 90441
rect -43309 88360 -42641 88466
rect -43309 86524 -43253 88360
rect -42697 86524 -42641 88360
rect -43309 86418 -42641 86524
rect -51117 84360 -49069 84466
rect -51117 82524 -51011 84360
rect -49175 82524 -49069 84360
rect -51117 82418 -49069 82524
rect -55117 -16103 -53069 -15997
rect -55117 -17939 -55011 -16103
rect -53175 -17939 -53069 -16103
rect -55117 -18045 -53069 -17939
rect -55093 -24021 -53093 -18045
rect -51093 -19997 -49093 82418
rect -43285 -15997 -42665 86418
rect -39285 84466 -38665 88466
rect -35309 88360 -34641 88466
rect -35309 86524 -35253 88360
rect -34697 86524 -34641 88360
rect -35309 86418 -34641 86524
rect -39309 84360 -38641 84466
rect -39309 82524 -39253 84360
rect -38697 82524 -38641 84360
rect -39309 82418 -38641 82524
rect -39285 23712 -38665 82418
rect -39285 23476 -39092 23712
rect -38856 23476 -38665 23712
rect -39285 16198 -38665 23476
rect -39285 15962 -39091 16198
rect -38855 15962 -38665 16198
rect -43309 -16103 -42641 -15997
rect -43309 -17939 -43253 -16103
rect -42697 -17939 -42641 -16103
rect -43309 -18045 -42641 -17939
rect -51117 -20103 -49069 -19997
rect -51117 -21939 -51011 -20103
rect -49175 -21939 -49069 -20103
rect -51117 -22045 -49069 -21939
rect -43285 -22045 -42665 -18045
rect -39285 -19997 -38665 15962
rect -35285 38496 -34665 86418
rect -31285 84466 -30665 88466
rect -27309 88360 -26641 88466
rect -27309 86524 -27253 88360
rect -26697 86524 -26641 88360
rect -27309 86418 -26641 86524
rect -31309 84360 -30641 84466
rect -31309 82524 -31253 84360
rect -30697 82524 -30641 84360
rect -31309 82418 -30641 82524
rect -35285 38260 -35105 38496
rect -34869 38260 -34665 38496
rect -35285 26906 -34665 38260
rect -35285 26670 -35111 26906
rect -34875 26670 -34665 26906
rect -35285 19231 -34665 26670
rect -35285 18995 -35105 19231
rect -34869 18995 -34665 19231
rect -35285 -15997 -34665 18995
rect -31285 38507 -30665 82418
rect -31285 38271 -31093 38507
rect -30857 38271 -30665 38507
rect -31285 37409 -30665 38271
rect -31285 37173 -31105 37409
rect -30869 37173 -30665 37409
rect -35309 -16103 -34641 -15997
rect -35309 -17939 -35253 -16103
rect -34697 -17939 -34641 -16103
rect -35309 -18045 -34641 -17939
rect -39309 -20103 -38641 -19997
rect -39309 -21939 -39253 -20103
rect -38697 -21939 -38641 -20103
rect -39309 -22045 -38641 -21939
rect -35285 -22045 -34665 -18045
rect -31285 -19997 -30665 37173
rect -27285 49824 -26665 86418
rect -23285 84466 -22665 88466
rect -19309 88360 -18641 88466
rect -19309 86524 -19253 88360
rect -18697 86524 -18641 88360
rect -19309 86418 -18641 86524
rect -23309 84360 -22641 84466
rect -23309 82524 -23253 84360
rect -22697 82524 -22641 84360
rect -23309 82418 -22641 82524
rect -27285 49588 -27089 49824
rect -26853 49588 -26665 49824
rect -27285 43154 -26665 49588
rect -27285 42918 -27054 43154
rect -26818 42918 -26665 43154
rect -27285 39948 -26665 42918
rect -27285 39712 -27049 39948
rect -26813 39712 -26665 39948
rect -27285 35879 -26665 39712
rect -27285 35643 -27049 35879
rect -26813 35643 -26665 35879
rect -27285 32765 -26665 35643
rect -27285 32529 -27051 32765
rect -26815 32529 -26665 32765
rect -27285 25512 -26665 32529
rect -27285 25276 -27081 25512
rect -26845 25276 -26665 25512
rect -27285 17961 -26665 25276
rect -27285 17725 -27091 17961
rect -26855 17725 -26665 17961
rect -27285 14475 -26665 17725
rect -27285 14239 -27084 14475
rect -26848 14239 -26665 14475
rect -27285 6708 -26665 14239
rect -27285 6472 -27092 6708
rect -26856 6472 -26665 6708
rect -27285 -15997 -26665 6472
rect -23285 49221 -22665 82418
rect -23285 48985 -23087 49221
rect -22851 48985 -22665 49221
rect -23285 37894 -22665 48985
rect -23285 37658 -23079 37894
rect -22843 37658 -22665 37894
rect -23285 24915 -22665 37658
rect -23285 24679 -23089 24915
rect -22853 24679 -22665 24915
rect -23285 15488 -22665 24679
rect -23285 15252 -23106 15488
rect -22870 15252 -22665 15488
rect -23285 5042 -22665 15252
rect -23285 4806 -23085 5042
rect -22849 4806 -22665 5042
rect -27309 -16103 -26641 -15997
rect -27309 -17939 -27253 -16103
rect -26697 -17939 -26641 -16103
rect -27309 -18045 -26641 -17939
rect -31309 -20103 -30641 -19997
rect -31309 -21939 -31253 -20103
rect -30697 -21939 -30641 -20103
rect -31309 -22045 -30641 -21939
rect -27285 -22045 -26665 -18045
rect -23285 -19997 -22665 4806
rect -19285 75066 -18665 86418
rect -15285 84466 -14665 88466
rect -11309 88360 -10641 88466
rect -11309 86524 -11253 88360
rect -10697 86524 -10641 88360
rect -11309 86418 -10641 86524
rect -15309 84360 -14641 84466
rect -15309 82524 -15253 84360
rect -14697 82524 -14641 84360
rect -15309 82418 -14641 82524
rect -19285 74830 -19094 75066
rect -18858 74830 -18665 75066
rect -19285 70235 -18665 74830
rect -19285 69999 -19094 70235
rect -18858 69999 -18665 70235
rect -19285 67120 -18665 69999
rect -19285 66884 -19098 67120
rect -18862 66884 -18665 67120
rect -19285 50688 -18665 66884
rect -19285 50452 -19091 50688
rect -18855 50452 -18665 50688
rect -19285 28706 -18665 50452
rect -19285 28470 -19091 28706
rect -18855 28470 -18665 28706
rect -19285 25808 -18665 28470
rect -19285 25572 -19099 25808
rect -18863 25572 -18665 25808
rect -19285 23728 -18665 25572
rect -19285 23492 -19092 23728
rect -18856 23492 -18665 23728
rect -19285 -15997 -18665 23492
rect -15285 75251 -14665 82418
rect -15285 75015 -15096 75251
rect -14860 75015 -14665 75251
rect -15285 70992 -14665 75015
rect -15285 70756 -15095 70992
rect -14859 70756 -14665 70992
rect -15285 68913 -14665 70756
rect -15285 68677 -15092 68913
rect -14856 68677 -14665 68913
rect -15285 38167 -14665 68677
rect -15285 37931 -15092 38167
rect -14856 37931 -14665 38167
rect -15285 27441 -14665 37931
rect -15285 27205 -15087 27441
rect -14851 27205 -14665 27441
rect -15285 25816 -14665 27205
rect -15285 25580 -15091 25816
rect -14855 25580 -14665 25816
rect -15285 23637 -14665 25580
rect -15285 23401 -15090 23637
rect -14854 23401 -14665 23637
rect -19309 -16103 -18641 -15997
rect -19309 -17939 -19253 -16103
rect -18697 -17939 -18641 -16103
rect -19309 -18045 -18641 -17939
rect -23309 -20103 -22641 -19997
rect -23309 -21939 -23253 -20103
rect -22697 -21939 -22641 -20103
rect -23309 -22045 -22641 -21939
rect -19285 -22045 -18665 -18045
rect -15285 -19997 -14665 23401
rect -11285 63499 -10665 86418
rect -7285 84466 -6665 88466
rect -3309 88360 -2641 88466
rect -3309 86524 -3253 88360
rect -2697 86524 -2641 88360
rect -3309 86418 -2641 86524
rect -7309 84360 -6641 84466
rect -7309 82524 -7253 84360
rect -6697 82524 -6641 84360
rect -7309 82418 -6641 82524
rect -11285 63263 -11022 63499
rect -10786 63263 -10665 63499
rect -11285 28053 -10665 63263
rect -11285 27817 -11090 28053
rect -10854 27817 -10665 28053
rect -11285 23152 -10665 27817
rect -11285 22916 -11099 23152
rect -10863 22916 -10665 23152
rect -11285 -15997 -10665 22916
rect -7285 63204 -6665 82418
rect -7285 62968 -6937 63204
rect -6701 62968 -6665 63204
rect -7285 55329 -6665 62968
rect -7285 55093 -6960 55329
rect -6724 55093 -6665 55329
rect -7285 55009 -6665 55093
rect -7285 54773 -6960 55009
rect -6724 54773 -6665 55009
rect -7285 51699 -6665 54773
rect -7285 51463 -7090 51699
rect -6854 51463 -6665 51699
rect -7285 15810 -6665 51463
rect -7285 15574 -7105 15810
rect -6869 15574 -6665 15810
rect -7285 14450 -6665 15574
rect -7285 14214 -7108 14450
rect -6872 14214 -6665 14450
rect -7285 10910 -6665 14214
rect -7285 10674 -7108 10910
rect -6872 10674 -6665 10910
rect -7285 9660 -6665 10674
rect -7285 9424 -7098 9660
rect -6862 9424 -6665 9660
rect -7285 7241 -6665 9424
rect -7285 7005 -7101 7241
rect -6865 7005 -6665 7241
rect -7285 5762 -6665 7005
rect -7285 5526 -7098 5762
rect -6862 5526 -6665 5762
rect -7285 -8278 -6665 5526
rect -7285 -8514 -7091 -8278
rect -6855 -8514 -6665 -8278
rect -11309 -16103 -10641 -15997
rect -11309 -17939 -11253 -16103
rect -10697 -17939 -10641 -16103
rect -11309 -18045 -10641 -17939
rect -15309 -20103 -14641 -19997
rect -15309 -21939 -15253 -20103
rect -14697 -21939 -14641 -20103
rect -15309 -22045 -14641 -21939
rect -11285 -22045 -10665 -18045
rect -7285 -19997 -6665 -8514
rect -3285 63409 -2665 86418
rect 715 84466 1335 88466
rect 4691 88360 5359 88466
rect 4691 86524 4747 88360
rect 5303 86524 5359 88360
rect 4691 86418 5359 86524
rect 691 84360 1359 84466
rect 691 82524 747 84360
rect 1303 82524 1359 84360
rect 691 82418 1359 82524
rect -3285 63173 -3094 63409
rect -2858 63173 -2665 63409
rect -3285 54420 -2665 63173
rect -3285 54184 -3090 54420
rect -2854 54184 -2665 54420
rect -3285 51099 -2665 54184
rect -3285 50863 -3084 51099
rect -2848 50863 -2665 51099
rect -3285 48771 -2665 50863
rect -3285 48535 -3090 48771
rect -2854 48535 -2665 48771
rect -3285 44601 -2665 48535
rect -3285 44365 -3094 44601
rect -2858 44365 -2665 44601
rect -3285 39884 -2665 44365
rect -3285 39648 -3086 39884
rect -2850 39648 -2665 39884
rect -3285 17862 -2665 39648
rect -3285 17626 -3098 17862
rect -2862 17626 -2665 17862
rect -3285 16448 -2665 17626
rect -3285 16212 -3088 16448
rect -2852 16212 -2665 16448
rect -3285 14046 -2665 16212
rect -3285 13810 -3086 14046
rect -2850 13810 -2665 14046
rect -3285 8800 -2665 13810
rect -3285 8564 -3088 8800
rect -2852 8564 -2665 8800
rect -3285 6741 -2665 8564
rect -3285 6505 -3086 6741
rect -2850 6505 -2665 6741
rect -3285 -6175 -2665 6505
rect -3285 -6411 -3085 -6175
rect -2849 -6411 -2665 -6175
rect -3285 -15997 -2665 -6411
rect 715 63230 1335 82418
rect 715 62994 904 63230
rect 1140 62994 1335 63230
rect 715 60122 1335 62994
rect 715 59886 903 60122
rect 1139 59886 1335 60122
rect 715 56747 1335 59886
rect 715 56511 903 56747
rect 1139 56511 1335 56747
rect 715 53372 1335 56511
rect 715 53136 903 53372
rect 1139 53136 1335 53372
rect 715 49997 1335 53136
rect 715 49761 903 49997
rect 1139 49761 1335 49997
rect 715 44512 1335 49761
rect 715 44276 899 44512
rect 1135 44276 1335 44512
rect 715 40867 1335 44276
rect 715 40631 909 40867
rect 1145 40631 1335 40867
rect 715 39438 1335 40631
rect 715 39202 903 39438
rect 1139 39202 1335 39438
rect 715 37093 1335 39202
rect 715 36857 904 37093
rect 1140 36857 1335 37093
rect 715 36014 1335 36857
rect 715 35778 921 36014
rect 1157 35778 1335 36014
rect 715 17616 1335 35778
rect 715 17380 902 17616
rect 1138 17380 1335 17616
rect 715 323 1335 17380
rect 715 87 907 323
rect 1143 87 1335 323
rect -3309 -16103 -2641 -15997
rect -3309 -17939 -3253 -16103
rect -2697 -17939 -2641 -16103
rect -3309 -18045 -2641 -17939
rect -7309 -20103 -6641 -19997
rect -7309 -21939 -7253 -20103
rect -6697 -21939 -6641 -20103
rect -7309 -22045 -6641 -21939
rect -3285 -22045 -2665 -18045
rect 715 -19997 1335 87
rect 4715 38051 5335 86418
rect 8715 84466 9335 88466
rect 12691 88360 13359 88466
rect 12691 86524 12747 88360
rect 13303 86524 13359 88360
rect 12691 86418 13359 86524
rect 8691 84360 9359 84466
rect 8691 82524 8747 84360
rect 9303 82524 9359 84360
rect 8691 82418 9359 82524
rect 4715 37815 4908 38051
rect 5144 37815 5335 38051
rect 4715 36658 5335 37815
rect 4715 36422 4915 36658
rect 5151 36422 5335 36658
rect 4715 35480 5335 36422
rect 4715 35244 4921 35480
rect 5157 35244 5335 35480
rect 4715 23157 5335 35244
rect 4715 22921 4893 23157
rect 5129 22921 5335 23157
rect 4715 19231 5335 22921
rect 4715 18995 4910 19231
rect 5146 18995 5335 19231
rect 4715 16593 5335 18995
rect 4715 16357 4907 16593
rect 5143 16357 5335 16593
rect 4715 16273 5335 16357
rect 4715 16037 4907 16273
rect 5143 16037 5335 16273
rect 4715 -15997 5335 16037
rect 8715 60111 9335 82418
rect 8715 59875 8908 60111
rect 9144 59875 9335 60111
rect 8715 56736 9335 59875
rect 8715 56500 8907 56736
rect 9143 56500 9335 56736
rect 8715 53361 9335 56500
rect 8715 53125 8907 53361
rect 9143 53125 9335 53361
rect 8715 49986 9335 53125
rect 8715 49750 8907 49986
rect 9143 49750 9335 49986
rect 8715 43236 9335 49750
rect 8715 43000 8907 43236
rect 9143 43000 9335 43236
rect 8715 36026 9335 43000
rect 8715 35790 8905 36026
rect 9141 35790 9335 36026
rect 8715 23493 9335 35790
rect 8715 23257 8887 23493
rect 9123 23257 9335 23493
rect 8715 17401 9335 23257
rect 8715 17165 8902 17401
rect 9138 17165 9335 17401
rect 8715 335 9335 17165
rect 8715 99 8927 335
rect 9163 99 9335 335
rect 4691 -16103 5359 -15997
rect 4691 -17939 4747 -16103
rect 5303 -17939 5359 -16103
rect 4691 -18045 5359 -17939
rect 691 -20103 1359 -19997
rect 691 -21939 747 -20103
rect 1303 -21939 1359 -20103
rect 691 -22045 1359 -21939
rect 4715 -22045 5335 -18045
rect 8715 -19997 9335 99
rect 12715 75170 13335 86418
rect 16715 84466 17335 88466
rect 20691 88360 21359 88466
rect 20691 86524 20747 88360
rect 21303 86524 21359 88360
rect 20691 86418 21359 86524
rect 16691 84360 17359 84466
rect 16691 82524 16747 84360
rect 17303 82524 17359 84360
rect 16691 82418 17359 82524
rect 12715 74934 12905 75170
rect 13141 74934 13335 75170
rect 12715 21094 13335 74934
rect 12715 20858 12864 21094
rect 13100 20858 13335 21094
rect 12715 18793 13335 20858
rect 12715 18557 12852 18793
rect 13088 18557 13335 18793
rect 12715 17188 13335 18557
rect 12715 16952 12846 17188
rect 13082 16952 13335 17188
rect 12715 15317 13335 16952
rect 12715 15081 12865 15317
rect 13101 15081 13335 15317
rect 12715 13616 13335 15081
rect 12715 13380 12887 13616
rect 13123 13380 13335 13616
rect 12715 11761 13335 13380
rect 12715 11525 12900 11761
rect 13136 11525 13335 11761
rect 12715 10651 13335 11525
rect 12715 10415 12896 10651
rect 13132 10415 13335 10651
rect 12715 -15997 13335 10415
rect 16715 75162 17335 82418
rect 16715 74926 16904 75162
rect 17140 74926 17335 75162
rect 16715 62582 17335 74926
rect 16715 62346 16910 62582
rect 17146 62346 17335 62582
rect 16715 58582 17335 62346
rect 16715 58346 16910 58582
rect 17146 58346 17335 58582
rect 16715 54582 17335 58346
rect 16715 54346 16910 54582
rect 17146 54346 17335 54582
rect 16715 50582 17335 54346
rect 16715 50346 16910 50582
rect 17146 50346 17335 50582
rect 16715 46582 17335 50346
rect 16715 46346 16910 46582
rect 17146 46346 17335 46582
rect 16715 19185 17335 46346
rect 16715 18949 16892 19185
rect 17128 18949 17335 19185
rect 16715 15592 17335 18949
rect 16715 15356 16800 15592
rect 17036 15356 17335 15592
rect 16715 323 17335 15356
rect 16715 87 16904 323
rect 17140 87 17335 323
rect 12691 -16103 13359 -15997
rect 12691 -17939 12747 -16103
rect 13303 -17939 13359 -16103
rect 12691 -18045 13359 -17939
rect 8691 -20103 9359 -19997
rect 8691 -21939 8747 -20103
rect 9303 -21939 9359 -20103
rect 8691 -22045 9359 -21939
rect 12715 -22045 13335 -18045
rect 16715 -19997 17335 87
rect 20715 64573 21335 86418
rect 24715 84466 25335 88466
rect 28691 88360 29359 88466
rect 28691 86524 28747 88360
rect 29303 86524 29359 88360
rect 28691 86418 29359 86524
rect 24691 84360 25359 84466
rect 24691 82524 24747 84360
rect 25303 82524 25359 84360
rect 24691 82418 25359 82524
rect 20715 64337 20907 64573
rect 21143 64337 21335 64573
rect 20715 60573 21335 64337
rect 20715 60337 20907 60573
rect 21143 60337 21335 60573
rect 20715 56573 21335 60337
rect 20715 56337 20907 56573
rect 21143 56337 21335 56573
rect 20715 52573 21335 56337
rect 20715 52337 20907 52573
rect 21143 52337 21335 52573
rect 20715 48573 21335 52337
rect 20715 48337 20907 48573
rect 21143 48337 21335 48573
rect 20715 19158 21335 48337
rect 20715 18922 20896 19158
rect 21132 18922 21335 19158
rect 20715 15587 21335 18922
rect 20715 15351 20839 15587
rect 21075 15351 21335 15587
rect 20715 11999 21335 15351
rect 20715 11763 20893 11999
rect 21129 11763 21335 11999
rect 20715 -15997 21335 11763
rect 24715 62575 25335 82418
rect 24715 62339 24906 62575
rect 25142 62339 25335 62575
rect 24715 58575 25335 62339
rect 24715 58339 24906 58575
rect 25142 58339 25335 58575
rect 24715 54575 25335 58339
rect 24715 54339 24906 54575
rect 25142 54339 25335 54575
rect 24715 50575 25335 54339
rect 24715 50339 24906 50575
rect 25142 50339 25335 50575
rect 24715 46575 25335 50339
rect 24715 46339 24906 46575
rect 25142 46339 25335 46575
rect 24715 19153 25335 46339
rect 24715 18917 24906 19153
rect 25142 18917 25335 19153
rect 24715 15560 25335 18917
rect 24715 15324 24908 15560
rect 25144 15324 25335 15560
rect 24715 11969 25335 15324
rect 24715 11733 24896 11969
rect 25132 11733 25335 11969
rect 20691 -16103 21359 -15997
rect 20691 -17939 20747 -16103
rect 21303 -17939 21359 -16103
rect 20691 -18045 21359 -17939
rect 16691 -20103 17359 -19997
rect 16691 -21939 16747 -20103
rect 17303 -21939 17359 -20103
rect 16691 -22045 17359 -21939
rect 20715 -22045 21335 -18045
rect 24715 -19997 25335 11733
rect 28715 64579 29335 86418
rect 32715 84466 33335 88466
rect 36691 88360 37359 88466
rect 36691 86524 36747 88360
rect 37303 86524 37359 88360
rect 36691 86418 37359 86524
rect 32691 84360 33359 84466
rect 32691 82524 32747 84360
rect 33303 82524 33359 84360
rect 32691 82418 33359 82524
rect 28715 64343 28901 64579
rect 29137 64343 29335 64579
rect 28715 60579 29335 64343
rect 28715 60343 28901 60579
rect 29137 60343 29335 60579
rect 28715 56579 29335 60343
rect 28715 56343 28901 56579
rect 29137 56343 29335 56579
rect 28715 52579 29335 56343
rect 28715 52343 28901 52579
rect 29137 52343 29335 52579
rect 28715 48579 29335 52343
rect 28715 48343 28901 48579
rect 29137 48343 29335 48579
rect 28715 -15997 29335 48343
rect 32715 62571 33335 82418
rect 32715 62335 32909 62571
rect 33145 62335 33335 62571
rect 32715 58571 33335 62335
rect 32715 58335 32909 58571
rect 33145 58335 33335 58571
rect 32715 54571 33335 58335
rect 32715 54335 32909 54571
rect 33145 54335 33335 54571
rect 32715 50571 33335 54335
rect 32715 50335 32909 50571
rect 33145 50335 33335 50571
rect 32715 46571 33335 50335
rect 32715 46335 32909 46571
rect 33145 46335 33335 46571
rect 32715 24132 33335 46335
rect 32715 23896 32904 24132
rect 33140 23896 33335 24132
rect 32715 21672 33335 23896
rect 32715 21436 32903 21672
rect 33139 21436 33335 21672
rect 32715 7291 33335 21436
rect 32715 7055 32906 7291
rect 33142 7055 33335 7291
rect 32715 5991 33335 7055
rect 32715 5755 32897 5991
rect 33133 5755 33335 5991
rect 32715 4576 33335 5755
rect 32715 4340 32903 4576
rect 33139 4340 33335 4576
rect 32715 3203 33335 4340
rect 32715 2967 32899 3203
rect 33135 2967 33335 3203
rect 32715 351 33335 2967
rect 32715 115 32906 351
rect 33142 115 33335 351
rect 32715 -949 33335 115
rect 32715 -1185 32897 -949
rect 33133 -1185 33335 -949
rect 32715 -2364 33335 -1185
rect 32715 -2600 32903 -2364
rect 33139 -2600 33335 -2364
rect 32715 -3737 33335 -2600
rect 32715 -3973 32899 -3737
rect 33135 -3973 33335 -3737
rect 28691 -16103 29359 -15997
rect 28691 -17939 28747 -16103
rect 29303 -17939 29359 -16103
rect 28691 -18045 29359 -17939
rect 24691 -20103 25359 -19997
rect 24691 -21939 24747 -20103
rect 25303 -21939 25359 -20103
rect 24691 -22045 25359 -21939
rect 28715 -22045 29335 -18045
rect 32715 -19997 33335 -3973
rect 36715 22815 37335 86418
rect 40715 84466 41335 88466
rect 44691 88360 45359 88466
rect 44691 86524 44747 88360
rect 45303 86524 45359 88360
rect 44691 86418 45359 86524
rect 40691 84360 41359 84466
rect 40691 82524 40747 84360
rect 41303 82524 41359 84360
rect 40691 82418 41359 82524
rect 36715 22579 36917 22815
rect 37153 22579 37335 22815
rect 36715 8791 37335 22579
rect 36715 8555 36900 8791
rect 37136 8555 37335 8791
rect 36715 6525 37335 8555
rect 36715 6289 36941 6525
rect 37177 6289 37335 6525
rect 36715 5109 37335 6289
rect 36715 4873 36902 5109
rect 37138 4873 37335 5109
rect 36715 2813 37335 4873
rect 36715 2577 36908 2813
rect 37144 2577 37335 2813
rect 36715 1851 37335 2577
rect 36715 1615 36900 1851
rect 37136 1615 37335 1851
rect 36715 -415 37335 1615
rect 36715 -651 36941 -415
rect 37177 -651 37335 -415
rect 36715 -1831 37335 -651
rect 36715 -2067 36902 -1831
rect 37138 -2067 37335 -1831
rect 36715 -4127 37335 -2067
rect 36715 -4363 36908 -4127
rect 37144 -4363 37335 -4127
rect 36715 -15997 37335 -4363
rect 40715 44302 41335 82418
rect 40715 44066 40913 44302
rect 41149 44066 41335 44302
rect 40715 40557 41335 44066
rect 40715 40321 40921 40557
rect 41157 40321 41335 40557
rect 40715 22730 41335 40321
rect 40715 22494 40914 22730
rect 41150 22494 41335 22730
rect 40715 7168 41335 22494
rect 40715 6932 40914 7168
rect 41150 6932 41335 7168
rect 40715 4265 41335 6932
rect 40715 4029 40912 4265
rect 41148 4029 41335 4265
rect 40715 228 41335 4029
rect 40715 -8 40914 228
rect 41150 -8 41335 228
rect 40715 -2679 41335 -8
rect 40715 -2915 40905 -2679
rect 41141 -2915 41335 -2679
rect 36691 -16103 37359 -15997
rect 36691 -17939 36747 -16103
rect 37303 -17939 37359 -16103
rect 36691 -18045 37359 -17939
rect 32691 -20103 33359 -19997
rect 32691 -21939 32747 -20103
rect 33303 -21939 33359 -20103
rect 32691 -22045 33359 -21939
rect 36715 -22045 37335 -18045
rect 40715 -19997 41335 -2915
rect 44715 45172 45335 86418
rect 48715 84466 49335 88466
rect 54883 88360 56931 88466
rect 54883 86524 54989 88360
rect 56825 86524 56931 88360
rect 54883 86418 56931 86524
rect 48691 84360 49359 84466
rect 48691 82524 48747 84360
rect 49303 82524 49359 84360
rect 48691 82418 49359 82524
rect 44715 44936 44908 45172
rect 45144 44936 45335 45172
rect 44715 44011 45335 44936
rect 44715 43775 44908 44011
rect 45144 43775 45335 44011
rect 44715 41502 45335 43775
rect 44715 41266 44892 41502
rect 45128 41266 45335 41502
rect 44715 40191 45335 41266
rect 44715 39955 44885 40191
rect 45121 39955 45335 40191
rect 44715 24250 45335 39955
rect 44715 24014 44914 24250
rect 45150 24014 45335 24250
rect 44715 7444 45335 24014
rect 44715 7208 44909 7444
rect 45145 7208 45335 7444
rect 44715 519 45335 7208
rect 44715 283 44912 519
rect 45148 283 45335 519
rect 44715 -15997 45335 283
rect 48715 21243 49335 82418
rect 48715 21007 48904 21243
rect 49140 21007 49335 21243
rect 44691 -16103 45359 -15997
rect 44691 -17939 44747 -16103
rect 45303 -17939 45359 -16103
rect 44691 -18045 45359 -17939
rect 40691 -20103 41359 -19997
rect 40691 -21939 40747 -20103
rect 41303 -21939 41359 -20103
rect 40691 -22045 41359 -21939
rect 44715 -22045 45335 -18045
rect 48715 -19997 49335 21007
rect 54907 -15997 56907 86418
rect 58907 84466 60907 90441
rect 58883 84360 60931 84466
rect 58883 82524 58989 84360
rect 60825 82524 60931 84360
rect 58883 82418 60931 82524
rect 54883 -16103 56931 -15997
rect 54883 -17939 54989 -16103
rect 56825 -17939 56931 -16103
rect 54883 -18045 56931 -17939
rect 48691 -20103 49359 -19997
rect 48691 -21939 48747 -20103
rect 49303 -21939 49359 -20103
rect 48691 -22045 49359 -21939
rect -51093 -24021 -49093 -22045
rect 54907 -24021 56907 -18045
rect 58907 -19997 60907 82418
rect 58883 -20103 60931 -19997
rect 58883 -21939 58989 -20103
rect 60825 -21939 60931 -20103
rect 58883 -22045 60931 -21939
rect 58907 -24021 60907 -22045
use a_mux2_en  a_mux2_en_0
timestamp 1654583406
transform 0 -1 -16584 1 0 68726
box -2638 -2585 3429 115
use a_mux2_en  a_mux2_en_1
timestamp 1654583406
transform 1 0 36330 0 1 23897
box -2638 -2585 3429 115
use a_mux4_en  a_mux4_en_0
timestamp 1654583406
transform 1 0 37083 0 1 8326
box -3690 -5314 3456 148
use a_mux4_en  a_mux4_en_1
timestamp 1654583406
transform 1 0 37083 0 1 1386
box -3690 -5314 3456 148
use clock_v2  clock_v2_0
timestamp 1654583406
transform 0 1 31620 -1 0 62637
box -3621 -14204 17033 36
use comparator_v2  comparator_v2_0
timestamp 1654583406
transform 0 -1 -18981 -1 0 39564
box -3788 -193 7250 10729
use esd_cell  esd_cell_0
timestamp 1654583101
transform 0 -1 14206 1 0 73319
box -65 -55 3553 3095
use esd_cell  esd_cell_1
timestamp 1654583101
transform 0 -1 -13798 1 0 73319
box -65 -55 3553 3095
use esd_cell  esd_cell_2
timestamp 1654583101
transform 1 0 42777 0 1 21122
box -65 -55 3553 3095
use esd_cell  esd_cell_3
timestamp 1654583101
transform 1 0 -38260 0 1 16027
box -65 -55 3553 3095
use esd_cell  esd_cell_4
timestamp 1654583101
transform 1 0 -38260 0 1 23557
box -65 -55 3553 3095
use esd_cell  esd_cell_5
timestamp 1654583101
transform 1 0 42522 0 1 4189
box -65 -55 3553 3095
use esd_cell  esd_cell_6
timestamp 1654583101
transform 1 0 42522 0 1 -2751
box -65 -55 3553 3095
use esd_cell  esd_cell_7
timestamp 1654583101
transform 0 1 -3548 -1 0 -6736
box -65 -55 3553 3095
use onebit_dac  onebit_dac_0
timestamp 1654583101
transform 1 0 -17091 0 1 24436
box -313 -1154 1895 1114
use onebit_dac  onebit_dac_1
timestamp 1654583101
transform 1 0 -17086 0 1 27078
box -313 -1154 1895 1114
use ota  ota_0
timestamp 1654583101
transform 0 -1 -7145 1 0 47315
box -7664 -17587 18520 2944
use ota_w_test  ota_w_test_0
timestamp 1654583101
transform 1 0 7664 0 1 17642
box -7664 -17587 18520 2944
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_0
timestamp 1654583101
transform 0 1 9865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_1
timestamp 1654583101
transform 0 1 9865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_2
timestamp 1654583101
transform 0 1 7865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_3
timestamp 1654583101
transform 0 1 7865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_4
timestamp 1654583101
transform 0 1 8865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_5
timestamp 1654583101
transform 0 1 8865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_6
timestamp 1654583101
transform 0 -1 4865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_7
timestamp 1654583101
transform 0 -1 5865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_8
timestamp 1654583101
transform 0 -1 4865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_9
timestamp 1654583101
transform 0 -1 5865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_10
timestamp 1654583101
transform 0 1 6865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_11
timestamp 1654583101
transform 0 1 6865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_12
timestamp 1654583101
transform 0 -1 2865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_13
timestamp 1654583101
transform 0 -1 3865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_14
timestamp 1654583101
transform 0 -1 2865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_15
timestamp 1654583101
transform 0 -1 3865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_16
timestamp 1654583101
transform 0 1 9865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_17
timestamp 1654583101
transform 0 1 9865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_18
timestamp 1654583101
transform 0 1 9865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_19
timestamp 1654583101
transform 0 1 7865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_20
timestamp 1654583101
transform 0 1 7865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_21
timestamp 1654583101
transform 0 1 7865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_22
timestamp 1654583101
transform 0 1 8865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_23
timestamp 1654583101
transform 0 1 8865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_24
timestamp 1654583101
transform 0 1 8865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_25
timestamp 1654583101
transform 0 -1 4865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_26
timestamp 1654583101
transform 0 -1 5865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_27
timestamp 1654583101
transform 0 -1 4865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_28
timestamp 1654583101
transform 0 -1 4865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_29
timestamp 1654583101
transform 0 -1 5865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_30
timestamp 1654583101
transform 0 -1 5865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_31
timestamp 1654583101
transform 0 1 6865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_32
timestamp 1654583101
transform 0 1 6865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_33
timestamp 1654583101
transform 0 1 6865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_34
timestamp 1654583101
transform 0 -1 2865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_35
timestamp 1654583101
transform 0 -1 3865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_36
timestamp 1654583101
transform 0 -1 2865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_37
timestamp 1654583101
transform 0 -1 2865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_38
timestamp 1654583101
transform 0 -1 3865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_39
timestamp 1654583101
transform 0 -1 3865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_40
timestamp 1654583101
transform 0 1 8865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_41
timestamp 1654583101
transform 0 1 9865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_42
timestamp 1654583101
transform 0 -1 5865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_43
timestamp 1654583101
transform 0 1 6865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_44
timestamp 1654583101
transform 0 1 7865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_45
timestamp 1654583101
transform 0 -1 4865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_46
timestamp 1654583101
transform 0 -1 2865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_47
timestamp 1654583101
transform 0 -1 3865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_48
timestamp 1654583101
transform 0 1 9865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_49
timestamp 1654583101
transform 0 1 8865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_50
timestamp 1654583101
transform 0 1 8865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_51
timestamp 1654583101
transform 0 1 8865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_52
timestamp 1654583101
transform 0 1 9865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_53
timestamp 1654583101
transform 0 1 9865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_54
timestamp 1654583101
transform 0 -1 5865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_55
timestamp 1654583101
transform 0 -1 5865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_56
timestamp 1654583101
transform 0 -1 5865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_57
timestamp 1654583101
transform 0 1 6865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_58
timestamp 1654583101
transform 0 1 6865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_59
timestamp 1654583101
transform 0 1 6865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_60
timestamp 1654583101
transform 0 1 7865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_61
timestamp 1654583101
transform 0 1 7865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_62
timestamp 1654583101
transform 0 1 7865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_63
timestamp 1654583101
transform 0 -1 4865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_64
timestamp 1654583101
transform 0 -1 4865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_65
timestamp 1654583101
transform 0 -1 4865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_66
timestamp 1654583101
transform 0 -1 2865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_67
timestamp 1654583101
transform 0 -1 3865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_68
timestamp 1654583101
transform 0 -1 2865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_69
timestamp 1654583101
transform 0 -1 2865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_70
timestamp 1654583101
transform 0 -1 3865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_71
timestamp 1654583101
transform 0 -1 3865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_0
timestamp 1654583101
transform 1 0 -9068 0 1 19276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_1
timestamp 1654583101
transform 1 0 -11668 0 1 19276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_2
timestamp 1654583101
transform 1 0 -14268 0 1 19276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_3
timestamp 1654583101
transform 1 0 -16868 0 1 19276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_4
timestamp 1654583101
transform 1 0 -19468 0 1 19276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_5
timestamp 1654583101
transform 1 0 -22068 0 1 19276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_6
timestamp 1654583101
transform 1 0 -9068 0 1 14076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_7
timestamp 1654583101
transform 1 0 -9068 0 1 16676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_8
timestamp 1654583101
transform 1 0 -9068 0 1 8876
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_9
timestamp 1654583101
transform 1 0 -9068 0 1 11476
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_10
timestamp 1654583101
transform 1 0 -9068 0 1 6276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_11
timestamp 1654583101
transform 1 0 -9068 0 1 3676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_12
timestamp 1654583101
transform 1 0 -9068 0 1 1076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_13
timestamp 1654583101
transform 1 0 -11668 0 1 16676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_14
timestamp 1654583101
transform 1 0 -14268 0 1 16676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_15
timestamp 1654583101
transform 1 0 -16868 0 1 16676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_16
timestamp 1654583101
transform 1 0 -19468 0 1 16676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_17
timestamp 1654583101
transform 1 0 -22068 0 1 16676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_18
timestamp 1654583101
transform 1 0 -11668 0 1 14076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_19
timestamp 1654583101
transform 1 0 -14268 0 1 14076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_20
timestamp 1654583101
transform 1 0 -16868 0 1 14076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_21
timestamp 1654583101
transform 1 0 -19468 0 1 14076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_22
timestamp 1654583101
transform 1 0 -22068 0 1 14076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_23
timestamp 1654583101
transform 1 0 -11668 0 1 11476
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_24
timestamp 1654583101
transform 1 0 -14268 0 1 11476
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_25
timestamp 1654583101
transform 1 0 -11668 0 1 8876
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_26
timestamp 1654583101
transform 1 0 -14268 0 1 8876
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_27
timestamp 1654583101
transform 1 0 -16868 0 1 11476
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_28
timestamp 1654583101
transform 1 0 -19468 0 1 11476
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_29
timestamp 1654583101
transform 1 0 -16868 0 1 8876
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_30
timestamp 1654583101
transform 1 0 -19468 0 1 8876
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_31
timestamp 1654583101
transform 1 0 -22068 0 1 8876
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_32
timestamp 1654583101
transform 1 0 -22068 0 1 11476
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_33
timestamp 1654583101
transform 1 0 -11668 0 1 3676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_34
timestamp 1654583101
transform 1 0 -14268 0 1 3676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_35
timestamp 1654583101
transform 1 0 -11668 0 1 6276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_36
timestamp 1654583101
transform 1 0 -14268 0 1 6276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_37
timestamp 1654583101
transform 1 0 -19468 0 1 3676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_38
timestamp 1654583101
transform 1 0 -16868 0 1 3676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_39
timestamp 1654583101
transform 1 0 -16868 0 1 6276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_40
timestamp 1654583101
transform 1 0 -19468 0 1 6276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_41
timestamp 1654583101
transform 1 0 -22068 0 1 6276
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_42
timestamp 1654583101
transform 1 0 -22068 0 1 3676
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_43
timestamp 1654583101
transform 1 0 -14268 0 1 1076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_44
timestamp 1654583101
transform 1 0 -11668 0 1 1076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_45
timestamp 1654583101
transform 1 0 -19468 0 1 1076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_46
timestamp 1654583101
transform 1 0 -16868 0 1 1076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_47
timestamp 1654583101
transform 1 0 -22068 0 1 1076
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_0
timestamp 1654583101
transform 1 0 -15946 0 -1 39777
box -1310 -1260 1210 1260
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_1
timestamp 1654583101
transform 1 0 -15946 0 -1 36367
box -1310 -1260 1210 1260
use sky130_fd_pr__nfet_01v8_CFEPS5  sky130_fd_pr__nfet_01v8_CFEPS5_0
timestamp 1654583101
transform 1 0 -31520 0 -1 38989
box -301 -264 301 266
use sky130_fd_pr__pfet_01v8_hvt_XAYTAL  sky130_fd_pr__pfet_01v8_hvt_XAYTAL_0
timestamp 1654583101
transform 1 0 -31520 0 1 38390
box -311 -319 311 319
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0
timestamp 1654583406
transform 1 0 42422 0 1 44495
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1654583406
transform 1 0 42422 0 1 43345
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1654583406
transform 1 0 -26628 0 1 49146
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1654583406
transform 1 0 42422 0 1 40805
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_4
timestamp 1654583406
transform 1 0 42422 0 1 39535
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0
timestamp 1654583406
transform 1 0 43158 0 1 44495
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1654583406
transform 1 0 43158 0 1 43345
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1654583406
transform 1 0 43158 0 1 40805
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1654583406
transform 1 0 43158 0 1 39535
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1654583406
transform 1 0 45458 0 1 44495
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1654583406
transform 1 0 45458 0 1 43345
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1654583406
transform 1 0 41962 0 1 44495
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1654583406
transform 1 0 41962 0 1 43345
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1654583406
transform 1 0 -25892 0 1 49146
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1654583406
transform 1 0 -27088 0 1 49146
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1654583406
transform 1 0 45458 0 1 40805
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1654583406
transform 1 0 41962 0 1 40805
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1654583406
transform 1 0 45458 0 1 39535
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1654583406
transform 1 0 41962 0 1 39535
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0
timestamp 1654583101
transform 1 0 39938 0 1 44495
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_1
timestamp 1654583101
transform 1 0 39938 0 1 43345
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_2
timestamp 1654583101
transform 1 0 39938 0 1 40805
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_3
timestamp 1654583101
transform 1 0 39938 0 1 39535
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1654583406
transform 1 0 45366 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654583406
transform 1 0 45366 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1654583406
transform 1 0 42330 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1654583406
transform 1 0 43066 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1654583406
transform 1 0 42330 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1654583406
transform 1 0 43066 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1654583406
transform 1 0 41870 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1654583406
transform 1 0 41870 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1654583406
transform 1 0 39846 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1654583406
transform 1 0 39846 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1654583406
transform 1 0 -26720 0 1 49146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1654583406
transform 1 0 -25984 0 1 49146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1654583406
transform 1 0 45366 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1654583406
transform 1 0 42330 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1654583406
transform 1 0 43066 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1654583406
transform 1 0 41870 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1654583406
transform 1 0 45366 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1654583406
transform 1 0 42330 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1654583406
transform 1 0 43066 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1654583406
transform 1 0 41870 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1654583406
transform 1 0 39846 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1654583406
transform 1 0 39846 0 1 39535
box -38 -48 130 592
use transmission_gate  transmission_gate_0
timestamp 1654583101
transform -1 0 -7618 0 -1 51315
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1654583101
transform 1 0 1359 0 -1 38947
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1654583101
transform 0 -1 9873 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1654583101
transform 0 1 6861 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1654583101
transform 0 -1 5873 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1654583101
transform 0 -1 3873 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1654583101
transform 1 0 1007 0 -1 37197
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1654583101
transform 0 1 9022 1 0 22174
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1654583101
transform -1 0 6948 0 1 23654
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1654583101
transform 0 -1 3845 1 0 22174
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1654583101
transform 0 -1 9839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1654583101
transform 0 -1 7839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_12
timestamp 1654583101
transform 0 -1 5839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_13
timestamp 1654583101
transform 0 -1 3839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_14
timestamp 1654583101
transform 0 1 -826 -1 0 18922
box -216 -51 1283 1063
use transmission_gate  transmission_gate_15
timestamp 1654583101
transform 1 0 -13548 0 1 27131
box -216 -51 1283 1063
use transmission_gate  transmission_gate_16
timestamp 1654583101
transform 1 0 -13548 0 1 25531
box -216 -51 1283 1063
use transmission_gate  transmission_gate_17
timestamp 1654583101
transform 1 0 -13548 0 1 23931
box -216 -51 1283 1063
use transmission_gate  transmission_gate_18
timestamp 1654583101
transform 1 0 -13548 0 1 22331
box -216 -51 1283 1063
use transmission_gate  transmission_gate_19
timestamp 1654583101
transform 1 0 -26607 0 1 24644
box -216 -51 1283 1063
use transmission_gate  transmission_gate_20
timestamp 1654583101
transform 1 0 -26607 0 1 17101
box -216 -51 1283 1063
use transmission_gate  transmission_gate_21
timestamp 1654583101
transform -1 0 -1901 0 -1 15522
box -216 -51 1283 1063
use transmission_gate  transmission_gate_22
timestamp 1654583101
transform 1 0 -6071 0 -1 14526
box -216 -51 1283 1063
use transmission_gate  transmission_gate_23
timestamp 1654583101
transform 0 1 -6231 1 0 8354
box -216 -51 1283 1063
use transmission_gate  transmission_gate_24
timestamp 1654583101
transform 0 1 -6231 -1 0 11991
box -216 -51 1283 1063
use transmission_gate  transmission_gate_25
timestamp 1654583101
transform 1 0 -2967 0 1 8995
box -216 -51 1283 1063
use transmission_gate  transmission_gate_26
timestamp 1654583101
transform 1 0 -2967 0 1 10595
box -216 -51 1283 1063
use transmission_gate  transmission_gate_27
timestamp 1654583101
transform 1 0 -2967 0 1 12195
box -216 -51 1283 1063
use transmission_gate  transmission_gate_28
timestamp 1654583101
transform -1 0 -1903 0 -1 6110
box -216 -51 1283 1063
use transmission_gate  transmission_gate_29
timestamp 1654583101
transform 1 0 -6071 0 1 5869
box -216 -51 1283 1063
use transmission_gate  transmission_gate_30
timestamp 1654583101
transform 1 0 -2967 0 1 7395
box -216 -51 1283 1063
use transmission_gate  transmission_gate_31
timestamp 1654583101
transform 1 0 -26675 0 1 13627
box -216 -51 1283 1063
use transmission_gate  transmission_gate_32
timestamp 1654583101
transform 1 0 -26675 0 1 5859
box -216 -51 1283 1063
<< labels >>
flabel metal3 s -56975 25027 -56975 25027 1 FreeSans 20000 0 0 0 ip
port 1 nsew
flabel metal3 s -57006 17492 -57006 17492 1 FreeSans 20000 0 0 0 in
port 2 nsew
flabel metal3 s -56866 37447 -56866 37447 1 FreeSans 20000 0 0 0 op
port 3 nsew
flabel metal3 s -56957 50045 -56957 50045 1 FreeSans 20000 0 0 0 rst_n
port 4 nsew
flabel metal3 s -16863 90254 -16863 90254 1 FreeSans 20000 0 0 0 a_probe_1
port 5 nsew
flabel metal3 s 11101 90277 11101 90277 1 FreeSans 20000 0 0 0 i_bias_2
port 6 nsew
flabel metal3 s 23035 90264 23035 90264 1 FreeSans 20000 0 0 0 clk
port 7 nsew
flabel metal3 s 62718 76068 62718 76068 1 FreeSans 20000 0 0 0 a_mod_grp_ctrl_1
port 8 nsew
flabel metal3 s 62776 68706 62776 68706 1 FreeSans 20000 0 0 0 a_mod_grp_ctrl_0
port 9 nsew
flabel metal3 s 62776 61266 62776 61266 1 FreeSans 20000 0 0 0 debug
port 10 nsew
flabel metal3 s 62793 55222 62793 55222 1 FreeSans 20000 0 0 0 d_clk_grp_1_ctrl_0
port 11 nsew
flabel metal3 s 62783 50992 62783 50992 1 FreeSans 20000 0 0 0 d_clk_grp_1_ctrl_1
port 12 nsew
flabel metal3 s 62738 47250 62738 47250 1 FreeSans 20000 0 0 0 d_probe_0
port 13 nsew
flabel metal3 s 62730 43660 62730 43660 1 FreeSans 20000 0 0 0 d_probe_1
port 14 nsew
flabel metal3 s 62755 33541 62755 33541 1 FreeSans 20000 0 0 0 d_probe_2
port 15 nsew
flabel metal3 s 62821 30323 62821 30323 1 FreeSans 20000 0 0 0 d_probe_3
port 16 nsew
flabel metal3 s 62686 40251 62686 40251 1 FreeSans 20000 0 0 0 d_clk_grp_2_ctrl_0
port 17 nsew
flabel metal3 s 62811 36995 62811 36995 1 FreeSans 20000 0 0 0 d_clk_grp_2_ctrl_1
port 18 nsew
flabel metal3 s 62769 22636 62769 22636 1 FreeSans 20000 0 0 0 a_probe_0
port 19 nsew
flabel metal3 s 62810 5693 62810 5693 1 FreeSans 20000 0 0 0 a_probe_2
port 20 nsew
flabel metal3 s 62725 -1241 62725 -1241 1 FreeSans 20000 0 0 0 a_probe_3
port 21 nsew
flabel metal3 s -998 -23902 -998 -23902 1 FreeSans 20000 0 0 0 i_bias_1
port 22 nsew
flabel metal5 s -54092 90092 -54092 90092 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s -50052 90052 -50052 90052 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
flabel metal5 s 55900 90138 55900 90138 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s 59914 90094 59914 90094 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
flabel metal5 s -54102 -23638 -54102 -23638 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s -50108 -23638 -50108 -23638 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
flabel metal5 s 55928 -23634 55928 -23634 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s 59912 -23508 59912 -23508 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
<< end >>
