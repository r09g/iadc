magic
tech sky130A
magscale 1 2
timestamp 1653390068
<< metal1 >>
rect 1558 6112 1568 6176
rect 1632 6112 1642 6176
rect 1568 3846 1632 6112
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 3157 5084 3221 5494
rect 3147 5020 3157 5084
rect 3221 5020 3231 5084
rect 4221 4928 6166 4932
rect 4148 4864 4158 4928
rect 4222 4868 6166 4928
rect 6230 4868 6240 4932
rect 4222 4864 4232 4868
rect 3298 4328 3308 4392
rect 3372 4328 3382 4392
rect 3308 4265 3372 4328
rect 4874 4326 5207 4390
rect 5271 4326 5281 4390
rect 1568 3782 1866 3846
rect 323 3419 333 3483
rect 397 3419 1571 3483
rect 1635 3419 1645 3483
rect 1802 3154 1866 3782
rect 323 3090 333 3154
rect 397 3090 1866 3154
rect 3308 2223 3371 4265
rect 4874 3642 4938 4326
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 3298 2159 3308 2223
rect 3372 2159 3382 2223
rect 3962 1582 3972 1646
rect 4036 1582 6152 1646
rect 6216 1582 6226 1646
rect 290 1307 300 1371
rect 364 1307 4326 1371
rect 4390 1307 4400 1371
<< via1 >>
rect 1568 6112 1632 6176
rect 3157 5494 3221 5558
rect 3157 5020 3221 5084
rect 4158 4864 4222 4928
rect 6166 4868 6230 4932
rect 3308 4328 3372 4392
rect 5207 4326 5271 4390
rect 333 3419 397 3483
rect 1571 3419 1635 3483
rect 333 3090 397 3154
rect 4874 3578 4938 3642
rect 3308 2159 3372 2223
rect 3972 1582 4036 1646
rect 6152 1582 6216 1646
rect 300 1307 364 1371
rect 4326 1307 4390 1371
<< metal2 >>
rect 1568 6176 1632 6186
rect 1568 6102 1632 6112
rect 3410 5781 3474 5791
rect 1570 5763 1634 5773
rect 1570 3843 1634 5699
rect 3157 5558 3221 5568
rect 3157 5484 3221 5494
rect 3410 5169 3474 5717
rect 3410 5095 3474 5105
rect 3157 5084 3221 5094
rect 3157 5010 3221 5020
rect 4158 4928 4222 4938
rect 4158 4854 4222 4864
rect 4704 4928 4768 4938
rect 5706 4928 5770 4938
rect 4768 4864 5706 4928
rect 4704 4854 4768 4864
rect 5706 4854 5770 4864
rect 6166 4932 6230 4942
rect 6166 4858 6230 4868
rect 3308 4392 3372 4402
rect 3308 4318 3372 4328
rect 5207 4390 5271 4400
rect 5207 4316 5271 4326
rect 3306 4042 3370 4052
rect 1570 3779 1866 3843
rect 333 3483 397 3493
rect 333 3409 397 3419
rect 765 3483 829 3493
rect 1378 3483 1442 3493
rect 829 3419 1378 3483
rect 765 3409 829 3419
rect 1378 3409 1442 3419
rect 1571 3483 1635 3493
rect 1571 3409 1635 3419
rect 333 3154 397 3164
rect 333 3080 397 3090
rect 764 3153 828 3163
rect 1802 3153 1866 3779
rect 828 3089 1866 3153
rect 764 3079 828 3089
rect 3306 2623 3370 3978
rect 4876 3980 4940 3990
rect 5206 3980 5270 3990
rect 4940 3916 5206 3980
rect 4876 3906 4940 3916
rect 5206 3906 5270 3916
rect 4874 3642 4938 3652
rect 4874 3568 4938 3578
rect 3306 2549 3370 2559
rect 3308 2223 3372 2233
rect 3308 2149 3372 2159
rect 3972 1646 4036 1656
rect 3972 1572 4036 1582
rect 4264 1642 4328 1652
rect 5736 1642 5800 1652
rect 4328 1578 5736 1642
rect 4264 1568 4328 1578
rect 5736 1568 5800 1578
rect 6152 1646 6216 1656
rect 6152 1572 6216 1582
rect 300 1371 364 1381
rect 300 1297 364 1307
rect 730 1371 794 1381
rect 3943 1371 4007 1381
rect 794 1307 3943 1371
rect 730 1297 794 1307
rect 3943 1297 4007 1307
rect 4326 1371 4390 1381
rect 4326 1297 4390 1307
<< via2 >>
rect 1568 6112 1632 6176
rect 1570 5699 1634 5763
rect 3410 5717 3474 5781
rect 3157 5494 3221 5558
rect 3410 5105 3474 5169
rect 3157 5020 3221 5084
rect 4158 4864 4222 4928
rect 4704 4864 4768 4928
rect 5706 4864 5770 4928
rect 6166 4868 6230 4932
rect 3308 4328 3372 4392
rect 5207 4326 5271 4390
rect 3306 3978 3370 4042
rect 333 3419 397 3483
rect 765 3419 829 3483
rect 1378 3419 1442 3483
rect 1571 3419 1635 3483
rect 333 3090 397 3154
rect 764 3089 828 3153
rect 4876 3916 4940 3980
rect 5206 3916 5270 3980
rect 4874 3578 4938 3642
rect 3306 2559 3370 2623
rect 3308 2159 3372 2223
rect 3972 1582 4036 1646
rect 4264 1578 4328 1642
rect 5736 1578 5800 1642
rect 6152 1582 6216 1646
rect 300 1307 364 1371
rect 730 1307 794 1371
rect 3943 1307 4007 1371
rect 4326 1307 4390 1371
<< metal3 >>
rect 1558 6176 1642 6181
rect 1558 6112 1568 6176
rect 1632 6112 1896 6176
rect 3157 6133 3698 6197
rect 1558 6107 1642 6112
rect 1556 5763 1648 5796
rect 1556 5699 1570 5763
rect 1634 5699 1648 5763
rect 1556 5674 1648 5699
rect 3157 5563 3221 6133
rect 3400 5781 3484 5810
rect 3400 5717 3410 5781
rect 3474 5717 3484 5781
rect 3400 5693 3484 5717
rect 3147 5558 3231 5563
rect 544 5311 608 5551
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 3147 5489 3231 5494
rect 544 5247 5105 5311
rect 3379 5169 3508 5177
rect 3379 5105 3410 5169
rect 3474 5105 3508 5169
rect 3379 5097 3508 5105
rect 3147 5084 3231 5089
rect 754 5020 3157 5084
rect 3221 5020 3231 5084
rect 754 4663 818 5020
rect 3147 5015 3231 5020
rect 4148 4928 4232 4933
rect 1241 4864 4158 4928
rect 4222 4864 4232 4928
rect 333 3488 397 3761
rect 323 3483 407 3488
rect 323 3419 333 3483
rect 397 3419 407 3483
rect 323 3414 407 3419
rect 743 3483 849 3501
rect 743 3419 765 3483
rect 829 3419 849 3483
rect 743 3404 849 3419
rect 323 3154 407 3159
rect 323 3090 333 3154
rect 397 3090 407 3154
rect 323 3085 407 3090
rect 745 3158 837 3183
rect 745 3153 838 3158
rect 745 3089 764 3153
rect 828 3089 838 3153
rect 333 2812 397 3085
rect 745 3084 838 3089
rect 745 3061 837 3084
rect 300 1376 364 1946
rect 290 1371 374 1376
rect 290 1307 300 1371
rect 364 1307 374 1371
rect 290 1302 374 1307
rect 710 1371 811 1387
rect 710 1307 730 1371
rect 794 1307 811 1371
rect 710 1289 811 1307
rect 1241 354 1305 4864
rect 4148 4859 4232 4864
rect 4681 4928 4791 4944
rect 4681 4864 4704 4928
rect 4768 4864 4791 4928
rect 4681 4850 4791 4864
rect 3298 4392 3382 4397
rect 3298 4328 3308 4392
rect 3372 4328 3698 4392
rect 3298 4323 3382 4328
rect 3283 4042 3389 4065
rect 3283 3978 3306 4042
rect 3370 3978 3389 4042
rect 3283 3958 3389 3978
rect 4862 3980 4953 4019
rect 4862 3916 4876 3980
rect 4940 3916 4953 3980
rect 4862 3879 4953 3916
rect 1367 3483 1454 3517
rect 1367 3419 1378 3483
rect 1442 3419 1454 3483
rect 1367 3388 1454 3419
rect 1561 3483 1645 3488
rect 1561 3419 1571 3483
rect 1635 3419 1645 3483
rect 1561 3414 1645 3419
rect 2348 3432 2412 3740
rect 4864 3642 4948 3647
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 4864 3573 4948 3578
rect 999 290 1305 354
rect 1571 365 1635 3414
rect 2348 3368 4212 3432
rect 4148 2819 4212 3368
rect 3284 2623 3390 2645
rect 3284 2559 3306 2623
rect 3370 2559 3390 2623
rect 3284 2538 3390 2559
rect 3298 2223 3382 2228
rect 2887 2159 3308 2223
rect 3372 2159 3382 2223
rect 3298 2154 3382 2159
rect 3962 1646 4046 1651
rect 3083 1582 3972 1646
rect 4036 1582 4046 1646
rect 1571 301 1897 365
rect 3083 363 3147 1582
rect 3962 1577 4046 1582
rect 4243 1642 4348 1666
rect 4243 1578 4264 1642
rect 4328 1578 4348 1642
rect 4243 1557 4348 1578
rect 3923 1371 4024 1390
rect 3923 1307 3943 1371
rect 4007 1307 4024 1371
rect 3923 1292 4024 1307
rect 4316 1371 4400 1376
rect 4316 1307 4326 1371
rect 4390 1307 4400 1371
rect 4316 1302 4400 1307
rect 4326 1060 4390 1302
rect 4874 448 4938 3573
rect 5041 616 5105 5247
rect 5683 4928 5793 4943
rect 6166 4937 6230 5491
rect 5683 4864 5706 4928
rect 5770 4864 5793 4928
rect 5683 4849 5793 4864
rect 6156 4932 6240 4937
rect 6156 4868 6166 4932
rect 6230 4868 6240 4932
rect 6156 4863 6240 4868
rect 5197 4390 5281 4395
rect 5197 4326 5207 4390
rect 5271 4326 5495 4390
rect 5197 4321 5281 4326
rect 5193 3980 5284 4018
rect 5193 3916 5206 3980
rect 5270 3916 5284 3980
rect 5193 3878 5284 3916
rect 5715 1642 5820 1664
rect 6152 1651 6216 1903
rect 5715 1578 5736 1642
rect 5800 1578 5820 1642
rect 5715 1555 5820 1578
rect 6142 1646 6226 1651
rect 6142 1582 6152 1646
rect 6216 1582 6226 1646
rect 6142 1577 6226 1582
rect 5041 552 5566 616
rect 4610 384 4941 448
rect 2812 299 3147 363
<< via3 >>
rect 1570 5699 1634 5763
rect 3410 5717 3474 5781
rect 3410 5105 3474 5169
rect 765 3419 829 3483
rect 764 3089 828 3153
rect 730 1307 794 1371
rect 4704 4864 4768 4928
rect 3306 3978 3370 4042
rect 4876 3916 4940 3980
rect 1378 3419 1442 3483
rect 3306 2559 3370 2623
rect 4264 1578 4328 1642
rect 3943 1307 4007 1371
rect 5706 4864 5770 4928
rect 5206 3916 5270 3980
rect 5736 1578 5800 1642
<< metal4 >>
rect 3409 5781 3475 5782
rect 1569 5763 1635 5764
rect 1569 5699 1570 5763
rect 1634 5699 1949 5763
rect 3409 5717 3410 5781
rect 3474 5717 3744 5781
rect 3409 5716 3475 5717
rect 1569 5698 1635 5699
rect 544 5311 608 5551
rect 544 5247 5105 5311
rect 3409 5169 3475 5170
rect 320 5105 3410 5169
rect 3474 5105 3475 5169
rect 320 4612 384 5105
rect 3409 5104 3475 5105
rect 4703 4928 4769 4929
rect 1242 4864 4704 4928
rect 4768 4864 4770 4928
rect 765 3484 829 3761
rect 764 3483 830 3484
rect 764 3419 765 3483
rect 829 3419 830 3483
rect 764 3418 830 3419
rect 763 3153 829 3154
rect 763 3089 764 3153
rect 828 3089 829 3153
rect 763 3088 829 3089
rect 764 2811 828 3088
rect 730 1372 794 1946
rect 729 1371 795 1372
rect 729 1307 730 1371
rect 794 1307 795 1371
rect 729 1306 795 1307
rect 1242 859 1306 4864
rect 4703 4863 4769 4864
rect 3305 4042 3371 4043
rect 3305 3978 3306 4042
rect 3370 3978 3746 4042
rect 4875 3980 4941 3981
rect 3305 3977 3371 3978
rect 4875 3916 4876 3980
rect 4940 3916 4941 3980
rect 4875 3915 4941 3916
rect 1377 3483 1443 3484
rect 1377 3419 1378 3483
rect 1442 3419 1443 3483
rect 1377 3418 1443 3419
rect 2348 3432 2412 3740
rect 998 795 1306 859
rect 1378 813 1442 3418
rect 2348 3368 4212 3432
rect 4148 2820 4212 3368
rect 3305 2623 3371 2624
rect 2816 2559 3306 2623
rect 3370 2559 3371 2623
rect 3305 2558 3371 2559
rect 4263 1642 4329 1643
rect 3083 1578 4264 1642
rect 4328 1578 4329 1642
rect 1378 749 1954 813
rect 3083 812 3147 1578
rect 4263 1577 4329 1578
rect 3943 1372 4007 1375
rect 3942 1371 4008 1372
rect 3942 1307 3943 1371
rect 4007 1307 4008 1371
rect 3942 1306 4008 1307
rect 3943 1007 4007 1306
rect 4876 844 4940 3915
rect 2812 748 3147 812
rect 4609 780 4940 844
rect 5041 616 5105 5247
rect 5706 4929 5770 5552
rect 5705 4928 5771 4929
rect 5705 4864 5706 4928
rect 5770 4864 5771 4928
rect 5705 4863 5771 4864
rect 5205 3980 5271 3981
rect 5205 3916 5206 3980
rect 5270 3916 5546 3980
rect 5205 3915 5271 3916
rect 5736 1643 5800 1953
rect 5735 1642 5801 1643
rect 5735 1578 5736 1642
rect 5800 1578 5801 1642
rect 5735 1577 5801 1578
rect 5041 552 5566 616
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/transmission_gate
timestamp 1652661863
transform -1 0 10282 0 1 7290
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1652661863
transform -1 0 10221 0 1 5421
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1652661863
transform -1 0 10323 0 1 -1685
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1652661863
transform -1 0 10241 0 1 3655
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1652661863
transform -1 0 10262 0 1 1868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1652661863
transform -1 0 10262 0 1 61
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1652661863
transform 1 0 -3806 0 1 7249
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1652661863
transform 1 0 -3745 0 1 5380
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1652661863
transform 1 0 -3765 0 1 3614
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1652661863
transform 1 0 -3786 0 1 1827
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1652661863
transform 1 0 -3786 0 1 20
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1652661863
transform 1 0 -3847 0 1 -1726
box -216 -51 1283 1063
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_0
timestamp 1653389200
transform 1 0 630 0 1 580
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_1
timestamp 1653389200
transform 1 0 2430 0 1 580
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_2
timestamp 1653389200
transform 1 0 4230 0 1 580
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_3
timestamp 1653389200
transform 1 0 6030 0 1 580
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_4
timestamp 1653389200
transform 1 0 6030 0 1 2380
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_5
timestamp 1653389200
transform 1 0 4230 0 1 2380
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_6
timestamp 1653389200
transform 1 0 2430 0 1 2380
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_7
timestamp 1653389200
transform 1 0 630 0 1 2380
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_8
timestamp 1653389200
transform 1 0 6030 0 1 4180
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_9
timestamp 1653389200
transform 1 0 4230 0 1 4180
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_10
timestamp 1653389200
transform 1 0 2430 0 1 4180
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_11
timestamp 1653389200
transform 1 0 630 0 1 4180
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_12
timestamp 1653389200
transform 1 0 6030 0 1 5980
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_13
timestamp 1653389200
transform 1 0 4230 0 1 5980
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_14
timestamp 1653389200
transform 1 0 2430 0 1 5980
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_15
timestamp 1653389200
transform 1 0 630 0 1 5980
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_16
timestamp 1653389200
transform 1 0 7830 0 1 5980
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_17
timestamp 1653389200
transform 1 0 7830 0 1 4180
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_18
timestamp 1653389200
transform 1 0 7830 0 1 2380
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_19
timestamp 1653389200
transform 1 0 7830 0 1 580
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_20
timestamp 1653389200
transform 1 0 -1170 0 1 5980
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_21
timestamp 1653389200
transform 1 0 -1170 0 1 4180
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_22
timestamp 1653389200
transform 1 0 -1170 0 1 2380
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_23
timestamp 1653389200
transform 1 0 -1170 0 1 580
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_24
timestamp 1653389200
transform 1 0 7830 0 1 7780
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_25
timestamp 1653389200
transform 1 0 6030 0 1 7780
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_26
timestamp 1653389200
transform 1 0 4230 0 1 7780
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_27
timestamp 1653389200
transform 1 0 2430 0 1 7780
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_28
timestamp 1653389200
transform 1 0 630 0 1 7780
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_29
timestamp 1653389200
transform 1 0 -1170 0 1 7780
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_30
timestamp 1653389200
transform 1 0 -1170 0 1 -1220
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_31
timestamp 1653389200
transform 1 0 630 0 1 -1220
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_32
timestamp 1653389200
transform 1 0 2430 0 1 -1220
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_33
timestamp 1653389200
transform 1 0 4230 0 1 -1220
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_34
timestamp 1653389200
transform 1 0 6030 0 1 -1220
box -630 -580 529 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_35
timestamp 1653389200
transform 1 0 7830 0 1 -1220
box -630 -580 529 580
<< end >>
