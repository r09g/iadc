magic
tech sky130A
magscale 1 2
timestamp 1655456512
<< metal3 >>
rect -12624 -25192 12470 25192
<< mimcap >>
rect -12524 25002 -6526 25042
rect -12524 19084 -12484 25002
rect -6566 19084 -6526 25002
rect -12524 19044 -6526 19084
rect -6207 25002 -209 25042
rect -6207 19084 -6167 25002
rect -249 19084 -209 25002
rect -6207 19044 -209 19084
rect 110 25002 6108 25042
rect 110 19084 150 25002
rect 6068 19084 6108 25002
rect 110 19044 6108 19084
rect 6427 25002 12425 25042
rect 6427 19084 6467 25002
rect 12385 19084 12425 25002
rect 6427 19044 12425 19084
rect -12524 18704 -6526 18744
rect -12524 12786 -12484 18704
rect -6566 12786 -6526 18704
rect -12524 12746 -6526 12786
rect -6207 18704 -209 18744
rect -6207 12786 -6167 18704
rect -249 12786 -209 18704
rect -6207 12746 -209 12786
rect 110 18704 6108 18744
rect 110 12786 150 18704
rect 6068 12786 6108 18704
rect 110 12746 6108 12786
rect 6427 18704 12425 18744
rect 6427 12786 6467 18704
rect 12385 12786 12425 18704
rect 6427 12746 12425 12786
rect -12524 12406 -6526 12446
rect -12524 6488 -12484 12406
rect -6566 6488 -6526 12406
rect -12524 6448 -6526 6488
rect -6207 12406 -209 12446
rect -6207 6488 -6167 12406
rect -249 6488 -209 12406
rect -6207 6448 -209 6488
rect 110 12406 6108 12446
rect 110 6488 150 12406
rect 6068 6488 6108 12406
rect 110 6448 6108 6488
rect 6427 12406 12425 12446
rect 6427 6488 6467 12406
rect 12385 6488 12425 12406
rect 6427 6448 12425 6488
rect -12524 6108 -6526 6148
rect -12524 190 -12484 6108
rect -6566 190 -6526 6108
rect -12524 150 -6526 190
rect -6207 6108 -209 6148
rect -6207 190 -6167 6108
rect -249 190 -209 6108
rect -6207 150 -209 190
rect 110 6108 6108 6148
rect 110 190 150 6108
rect 6068 190 6108 6108
rect 110 150 6108 190
rect 6427 6108 12425 6148
rect 6427 190 6467 6108
rect 12385 190 12425 6108
rect 6427 150 12425 190
rect -12524 -190 -6526 -150
rect -12524 -6108 -12484 -190
rect -6566 -6108 -6526 -190
rect -12524 -6148 -6526 -6108
rect -6207 -190 -209 -150
rect -6207 -6108 -6167 -190
rect -249 -6108 -209 -190
rect -6207 -6148 -209 -6108
rect 110 -190 6108 -150
rect 110 -6108 150 -190
rect 6068 -6108 6108 -190
rect 110 -6148 6108 -6108
rect 6427 -190 12425 -150
rect 6427 -6108 6467 -190
rect 12385 -6108 12425 -190
rect 6427 -6148 12425 -6108
rect -12524 -6488 -6526 -6448
rect -12524 -12406 -12484 -6488
rect -6566 -12406 -6526 -6488
rect -12524 -12446 -6526 -12406
rect -6207 -6488 -209 -6448
rect -6207 -12406 -6167 -6488
rect -249 -12406 -209 -6488
rect -6207 -12446 -209 -12406
rect 110 -6488 6108 -6448
rect 110 -12406 150 -6488
rect 6068 -12406 6108 -6488
rect 110 -12446 6108 -12406
rect 6427 -6488 12425 -6448
rect 6427 -12406 6467 -6488
rect 12385 -12406 12425 -6488
rect 6427 -12446 12425 -12406
rect -12524 -12786 -6526 -12746
rect -12524 -18704 -12484 -12786
rect -6566 -18704 -6526 -12786
rect -12524 -18744 -6526 -18704
rect -6207 -12786 -209 -12746
rect -6207 -18704 -6167 -12786
rect -249 -18704 -209 -12786
rect -6207 -18744 -209 -18704
rect 110 -12786 6108 -12746
rect 110 -18704 150 -12786
rect 6068 -18704 6108 -12786
rect 110 -18744 6108 -18704
rect 6427 -12786 12425 -12746
rect 6427 -18704 6467 -12786
rect 12385 -18704 12425 -12786
rect 6427 -18744 12425 -18704
rect -12524 -19084 -6526 -19044
rect -12524 -25002 -12484 -19084
rect -6566 -25002 -6526 -19084
rect -12524 -25042 -6526 -25002
rect -6207 -19084 -209 -19044
rect -6207 -25002 -6167 -19084
rect -249 -25002 -209 -19084
rect -6207 -25042 -209 -25002
rect 110 -19084 6108 -19044
rect 110 -25002 150 -19084
rect 6068 -25002 6108 -19084
rect 110 -25042 6108 -25002
rect 6427 -19084 12425 -19044
rect 6427 -25002 6467 -19084
rect 12385 -25002 12425 -19084
rect 6427 -25042 12425 -25002
<< mimcapcontact >>
rect -12484 19084 -6566 25002
rect -6167 19084 -249 25002
rect 150 19084 6068 25002
rect 6467 19084 12385 25002
rect -12484 12786 -6566 18704
rect -6167 12786 -249 18704
rect 150 12786 6068 18704
rect 6467 12786 12385 18704
rect -12484 6488 -6566 12406
rect -6167 6488 -249 12406
rect 150 6488 6068 12406
rect 6467 6488 12385 12406
rect -12484 190 -6566 6108
rect -6167 190 -249 6108
rect 150 190 6068 6108
rect 6467 190 12385 6108
rect -12484 -6108 -6566 -190
rect -6167 -6108 -249 -190
rect 150 -6108 6068 -190
rect 6467 -6108 12385 -190
rect -12484 -12406 -6566 -6488
rect -6167 -12406 -249 -6488
rect 150 -12406 6068 -6488
rect 6467 -12406 12385 -6488
rect -12484 -18704 -6566 -12786
rect -6167 -18704 -249 -12786
rect 150 -18704 6068 -12786
rect 6467 -18704 12385 -12786
rect -12484 -25002 -6566 -19084
rect -6167 -25002 -249 -19084
rect 150 -25002 6068 -19084
rect 6467 -25002 12385 -19084
<< metal4 >>
rect -12624 25002 12470 25192
rect -12624 19084 -12484 25002
rect -6566 19084 -6167 25002
rect -249 19084 150 25002
rect 6068 19084 6467 25002
rect 12385 19084 12470 25002
rect -12624 18704 12470 19084
rect -12624 12786 -12484 18704
rect -6566 12786 -6167 18704
rect -249 12786 150 18704
rect 6068 12786 6467 18704
rect 12385 12786 12470 18704
rect -12624 12406 12470 12786
rect -12624 6488 -12484 12406
rect -6566 6488 -6167 12406
rect -249 6488 150 12406
rect 6068 6488 6467 12406
rect 12385 6488 12470 12406
rect -12624 6108 12470 6488
rect -12624 190 -12484 6108
rect -6566 190 -6167 6108
rect -249 190 150 6108
rect 6068 190 6467 6108
rect 12385 190 12470 6108
rect -12624 -190 12470 190
rect -12624 -6108 -12484 -190
rect -6566 -6108 -6167 -190
rect -249 -6108 150 -190
rect 6068 -6108 6467 -190
rect 12385 -6108 12470 -190
rect -12624 -6488 12470 -6108
rect -12624 -12406 -12484 -6488
rect -6566 -12406 -6167 -6488
rect -249 -12406 150 -6488
rect 6068 -12406 6467 -6488
rect 12385 -12406 12470 -6488
rect -12624 -12786 12470 -12406
rect -12624 -18704 -12484 -12786
rect -6566 -18704 -6167 -12786
rect -249 -18704 150 -12786
rect 6068 -18704 6467 -12786
rect 12385 -18704 12470 -12786
rect -12624 -19084 12470 -18704
rect -12624 -25002 -12484 -19084
rect -6566 -25002 -6167 -19084
rect -249 -25002 150 -19084
rect 6068 -25002 6467 -19084
rect 12385 -25002 12470 -19084
rect -12624 -25192 12470 -25002
<< properties >>
string FIXED_BBOX 6327 18944 12525 25142
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 29.993 l 29.993 val 1.821k carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
