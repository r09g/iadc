magic
tech sky130A
magscale 1 2
timestamp 1653906530
<< nwell >>
rect -65 1501 3553 3095
<< pwell >>
rect -35 -65 3523 1451
<< mvnmos >>
rect 193 193 293 1193
rect 351 193 451 1193
rect 509 193 609 1193
rect 667 193 767 1193
rect 825 193 925 1193
rect 983 193 1083 1193
rect 1141 193 1241 1193
rect 1299 193 1399 1193
rect 1457 193 1557 1193
rect 1615 193 1715 1193
rect 1773 193 1873 1193
rect 1931 193 2031 1193
rect 2089 193 2189 1193
rect 2247 193 2347 1193
rect 2405 193 2505 1193
rect 2563 193 2663 1193
rect 2721 193 2821 1193
rect 2879 193 2979 1193
rect 3037 193 3137 1193
rect 3195 193 3295 1193
<< mvpmos >>
rect 193 1798 293 2798
rect 351 1798 451 2798
rect 509 1798 609 2798
rect 667 1798 767 2798
rect 825 1798 925 2798
rect 983 1798 1083 2798
rect 1141 1798 1241 2798
rect 1299 1798 1399 2798
rect 1457 1798 1557 2798
rect 1615 1798 1715 2798
rect 1773 1798 1873 2798
rect 1931 1798 2031 2798
rect 2089 1798 2189 2798
rect 2247 1798 2347 2798
rect 2405 1798 2505 2798
rect 2563 1798 2663 2798
rect 2721 1798 2821 2798
rect 2879 1798 2979 2798
rect 3037 1798 3137 2798
rect 3195 1798 3295 2798
<< mvndiff >>
rect 135 1181 193 1193
rect 135 205 147 1181
rect 181 205 193 1181
rect 135 193 193 205
rect 293 1181 351 1193
rect 293 205 305 1181
rect 339 205 351 1181
rect 293 193 351 205
rect 451 1181 509 1193
rect 451 205 463 1181
rect 497 205 509 1181
rect 451 193 509 205
rect 609 1181 667 1193
rect 609 205 621 1181
rect 655 205 667 1181
rect 609 193 667 205
rect 767 1181 825 1193
rect 767 205 779 1181
rect 813 205 825 1181
rect 767 193 825 205
rect 925 1181 983 1193
rect 925 205 937 1181
rect 971 205 983 1181
rect 925 193 983 205
rect 1083 1181 1141 1193
rect 1083 205 1095 1181
rect 1129 205 1141 1181
rect 1083 193 1141 205
rect 1241 1181 1299 1193
rect 1241 205 1253 1181
rect 1287 205 1299 1181
rect 1241 193 1299 205
rect 1399 1181 1457 1193
rect 1399 205 1411 1181
rect 1445 205 1457 1181
rect 1399 193 1457 205
rect 1557 1181 1615 1193
rect 1557 205 1569 1181
rect 1603 205 1615 1181
rect 1557 193 1615 205
rect 1715 1181 1773 1193
rect 1715 205 1727 1181
rect 1761 205 1773 1181
rect 1715 193 1773 205
rect 1873 1181 1931 1193
rect 1873 205 1885 1181
rect 1919 205 1931 1181
rect 1873 193 1931 205
rect 2031 1181 2089 1193
rect 2031 205 2043 1181
rect 2077 205 2089 1181
rect 2031 193 2089 205
rect 2189 1181 2247 1193
rect 2189 205 2201 1181
rect 2235 205 2247 1181
rect 2189 193 2247 205
rect 2347 1181 2405 1193
rect 2347 205 2359 1181
rect 2393 205 2405 1181
rect 2347 193 2405 205
rect 2505 1181 2563 1193
rect 2505 205 2517 1181
rect 2551 205 2563 1181
rect 2505 193 2563 205
rect 2663 1181 2721 1193
rect 2663 205 2675 1181
rect 2709 205 2721 1181
rect 2663 193 2721 205
rect 2821 1181 2879 1193
rect 2821 205 2833 1181
rect 2867 205 2879 1181
rect 2821 193 2879 205
rect 2979 1181 3037 1193
rect 2979 205 2991 1181
rect 3025 205 3037 1181
rect 2979 193 3037 205
rect 3137 1181 3195 1193
rect 3137 205 3149 1181
rect 3183 205 3195 1181
rect 3137 193 3195 205
rect 3295 1181 3353 1193
rect 3295 205 3307 1181
rect 3341 205 3353 1181
rect 3295 193 3353 205
<< mvpdiff >>
rect 135 2786 193 2798
rect 135 1810 147 2786
rect 181 1810 193 2786
rect 135 1798 193 1810
rect 293 2786 351 2798
rect 293 1810 305 2786
rect 339 1810 351 2786
rect 293 1798 351 1810
rect 451 2786 509 2798
rect 451 1810 463 2786
rect 497 1810 509 2786
rect 451 1798 509 1810
rect 609 2786 667 2798
rect 609 1810 621 2786
rect 655 1810 667 2786
rect 609 1798 667 1810
rect 767 2786 825 2798
rect 767 1810 779 2786
rect 813 1810 825 2786
rect 767 1798 825 1810
rect 925 2786 983 2798
rect 925 1810 937 2786
rect 971 1810 983 2786
rect 925 1798 983 1810
rect 1083 2786 1141 2798
rect 1083 1810 1095 2786
rect 1129 1810 1141 2786
rect 1083 1798 1141 1810
rect 1241 2786 1299 2798
rect 1241 1810 1253 2786
rect 1287 1810 1299 2786
rect 1241 1798 1299 1810
rect 1399 2786 1457 2798
rect 1399 1810 1411 2786
rect 1445 1810 1457 2786
rect 1399 1798 1457 1810
rect 1557 2786 1615 2798
rect 1557 1810 1569 2786
rect 1603 1810 1615 2786
rect 1557 1798 1615 1810
rect 1715 2786 1773 2798
rect 1715 1810 1727 2786
rect 1761 1810 1773 2786
rect 1715 1798 1773 1810
rect 1873 2786 1931 2798
rect 1873 1810 1885 2786
rect 1919 1810 1931 2786
rect 1873 1798 1931 1810
rect 2031 2786 2089 2798
rect 2031 1810 2043 2786
rect 2077 1810 2089 2786
rect 2031 1798 2089 1810
rect 2189 2786 2247 2798
rect 2189 1810 2201 2786
rect 2235 1810 2247 2786
rect 2189 1798 2247 1810
rect 2347 2786 2405 2798
rect 2347 1810 2359 2786
rect 2393 1810 2405 2786
rect 2347 1798 2405 1810
rect 2505 2786 2563 2798
rect 2505 1810 2517 2786
rect 2551 1810 2563 2786
rect 2505 1798 2563 1810
rect 2663 2786 2721 2798
rect 2663 1810 2675 2786
rect 2709 1810 2721 2786
rect 2663 1798 2721 1810
rect 2821 2786 2879 2798
rect 2821 1810 2833 2786
rect 2867 1810 2879 2786
rect 2821 1798 2879 1810
rect 2979 2786 3037 2798
rect 2979 1810 2991 2786
rect 3025 1810 3037 2786
rect 2979 1798 3037 1810
rect 3137 2786 3195 2798
rect 3137 1810 3149 2786
rect 3183 1810 3195 2786
rect 3137 1798 3195 1810
rect 3295 2786 3353 2798
rect 3295 1810 3307 2786
rect 3341 1810 3353 2786
rect 3295 1798 3353 1810
<< mvndiffc >>
rect 147 205 181 1181
rect 305 205 339 1181
rect 463 205 497 1181
rect 621 205 655 1181
rect 779 205 813 1181
rect 937 205 971 1181
rect 1095 205 1129 1181
rect 1253 205 1287 1181
rect 1411 205 1445 1181
rect 1569 205 1603 1181
rect 1727 205 1761 1181
rect 1885 205 1919 1181
rect 2043 205 2077 1181
rect 2201 205 2235 1181
rect 2359 205 2393 1181
rect 2517 205 2551 1181
rect 2675 205 2709 1181
rect 2833 205 2867 1181
rect 2991 205 3025 1181
rect 3149 205 3183 1181
rect 3307 205 3341 1181
<< mvpdiffc >>
rect 147 1810 181 2786
rect 305 1810 339 2786
rect 463 1810 497 2786
rect 621 1810 655 2786
rect 779 1810 813 2786
rect 937 1810 971 2786
rect 1095 1810 1129 2786
rect 1253 1810 1287 2786
rect 1411 1810 1445 2786
rect 1569 1810 1603 2786
rect 1727 1810 1761 2786
rect 1885 1810 1919 2786
rect 2043 1810 2077 2786
rect 2201 1810 2235 2786
rect 2359 1810 2393 2786
rect 2517 1810 2551 2786
rect 2675 1810 2709 2786
rect 2833 1810 2867 2786
rect 2991 1810 3025 2786
rect 3149 1810 3183 2786
rect 3307 1810 3341 2786
<< mvpsubdiff >>
rect 1 1403 3487 1415
rect 1 1369 109 1403
rect 3379 1369 3487 1403
rect 1 1357 3487 1369
rect 1 1307 59 1357
rect 1 79 13 1307
rect 47 79 59 1307
rect 3429 1307 3487 1357
rect 1 29 59 79
rect 3429 79 3441 1307
rect 3475 79 3487 1307
rect 3429 29 3487 79
rect 1 17 3487 29
rect 1 -17 109 17
rect 3379 -17 3487 17
rect 1 -29 3487 -17
<< mvnsubdiff >>
rect 1 3017 3487 3029
rect 1 2983 109 3017
rect 3379 2983 3487 3017
rect 1 2971 3487 2983
rect 1 2921 59 2971
rect 1 1675 13 2921
rect 47 1675 59 2921
rect 3429 2921 3487 2971
rect 1 1625 59 1675
rect 3429 1675 3441 2921
rect 3475 1675 3487 2921
rect 3429 1625 3487 1675
rect 1 1613 3487 1625
rect 1 1579 109 1613
rect 3379 1579 3487 1613
rect 1 1567 3487 1579
<< mvpsubdiffcont >>
rect 109 1369 3379 1403
rect 13 79 47 1307
rect 3441 79 3475 1307
rect 109 -17 3379 17
<< mvnsubdiffcont >>
rect 109 2983 3379 3017
rect 13 1675 47 2921
rect 3441 1675 3475 2921
rect 109 1579 3379 1613
<< poly >>
rect 193 2879 293 2895
rect 193 2845 209 2879
rect 277 2845 293 2879
rect 193 2798 293 2845
rect 351 2879 451 2895
rect 351 2845 367 2879
rect 435 2845 451 2879
rect 351 2798 451 2845
rect 509 2879 609 2895
rect 509 2845 525 2879
rect 593 2845 609 2879
rect 509 2798 609 2845
rect 667 2879 767 2895
rect 667 2845 683 2879
rect 751 2845 767 2879
rect 667 2798 767 2845
rect 825 2879 925 2895
rect 825 2845 841 2879
rect 909 2845 925 2879
rect 825 2798 925 2845
rect 983 2879 1083 2895
rect 983 2845 999 2879
rect 1067 2845 1083 2879
rect 983 2798 1083 2845
rect 1141 2879 1241 2895
rect 1141 2845 1157 2879
rect 1225 2845 1241 2879
rect 1141 2798 1241 2845
rect 1299 2879 1399 2895
rect 1299 2845 1315 2879
rect 1383 2845 1399 2879
rect 1299 2798 1399 2845
rect 1457 2879 1557 2895
rect 1457 2845 1473 2879
rect 1541 2845 1557 2879
rect 1457 2798 1557 2845
rect 1615 2879 1715 2895
rect 1615 2845 1631 2879
rect 1699 2845 1715 2879
rect 1615 2798 1715 2845
rect 1773 2879 1873 2895
rect 1773 2845 1789 2879
rect 1857 2845 1873 2879
rect 1773 2798 1873 2845
rect 1931 2879 2031 2895
rect 1931 2845 1947 2879
rect 2015 2845 2031 2879
rect 1931 2798 2031 2845
rect 2089 2879 2189 2895
rect 2089 2845 2105 2879
rect 2173 2845 2189 2879
rect 2089 2798 2189 2845
rect 2247 2879 2347 2895
rect 2247 2845 2263 2879
rect 2331 2845 2347 2879
rect 2247 2798 2347 2845
rect 2405 2879 2505 2895
rect 2405 2845 2421 2879
rect 2489 2845 2505 2879
rect 2405 2798 2505 2845
rect 2563 2879 2663 2895
rect 2563 2845 2579 2879
rect 2647 2845 2663 2879
rect 2563 2798 2663 2845
rect 2721 2879 2821 2895
rect 2721 2845 2737 2879
rect 2805 2845 2821 2879
rect 2721 2798 2821 2845
rect 2879 2879 2979 2895
rect 2879 2845 2895 2879
rect 2963 2845 2979 2879
rect 2879 2798 2979 2845
rect 3037 2879 3137 2895
rect 3037 2845 3053 2879
rect 3121 2845 3137 2879
rect 3037 2798 3137 2845
rect 3195 2879 3295 2895
rect 3195 2845 3211 2879
rect 3279 2845 3295 2879
rect 3195 2798 3295 2845
rect 193 1751 293 1798
rect 193 1717 209 1751
rect 277 1717 293 1751
rect 193 1701 293 1717
rect 351 1751 451 1798
rect 351 1717 367 1751
rect 435 1717 451 1751
rect 351 1701 451 1717
rect 509 1751 609 1798
rect 509 1717 525 1751
rect 593 1717 609 1751
rect 509 1701 609 1717
rect 667 1751 767 1798
rect 667 1717 683 1751
rect 751 1717 767 1751
rect 667 1701 767 1717
rect 825 1751 925 1798
rect 825 1717 841 1751
rect 909 1717 925 1751
rect 825 1701 925 1717
rect 983 1751 1083 1798
rect 983 1717 999 1751
rect 1067 1717 1083 1751
rect 983 1701 1083 1717
rect 1141 1751 1241 1798
rect 1141 1717 1157 1751
rect 1225 1717 1241 1751
rect 1141 1701 1241 1717
rect 1299 1751 1399 1798
rect 1299 1717 1315 1751
rect 1383 1717 1399 1751
rect 1299 1701 1399 1717
rect 1457 1751 1557 1798
rect 1457 1717 1473 1751
rect 1541 1717 1557 1751
rect 1457 1701 1557 1717
rect 1615 1751 1715 1798
rect 1615 1717 1631 1751
rect 1699 1717 1715 1751
rect 1615 1701 1715 1717
rect 1773 1751 1873 1798
rect 1773 1717 1789 1751
rect 1857 1717 1873 1751
rect 1773 1701 1873 1717
rect 1931 1751 2031 1798
rect 1931 1717 1947 1751
rect 2015 1717 2031 1751
rect 1931 1701 2031 1717
rect 2089 1751 2189 1798
rect 2089 1717 2105 1751
rect 2173 1717 2189 1751
rect 2089 1701 2189 1717
rect 2247 1751 2347 1798
rect 2247 1717 2263 1751
rect 2331 1717 2347 1751
rect 2247 1701 2347 1717
rect 2405 1751 2505 1798
rect 2405 1717 2421 1751
rect 2489 1717 2505 1751
rect 2405 1701 2505 1717
rect 2563 1751 2663 1798
rect 2563 1717 2579 1751
rect 2647 1717 2663 1751
rect 2563 1701 2663 1717
rect 2721 1751 2821 1798
rect 2721 1717 2737 1751
rect 2805 1717 2821 1751
rect 2721 1701 2821 1717
rect 2879 1751 2979 1798
rect 2879 1717 2895 1751
rect 2963 1717 2979 1751
rect 2879 1701 2979 1717
rect 3037 1751 3137 1798
rect 3037 1717 3053 1751
rect 3121 1717 3137 1751
rect 3037 1701 3137 1717
rect 3195 1751 3295 1798
rect 3195 1717 3211 1751
rect 3279 1717 3295 1751
rect 3195 1701 3295 1717
rect 193 1265 293 1281
rect 193 1231 209 1265
rect 277 1231 293 1265
rect 193 1193 293 1231
rect 351 1265 451 1281
rect 351 1231 367 1265
rect 435 1231 451 1265
rect 351 1193 451 1231
rect 509 1265 609 1281
rect 509 1231 525 1265
rect 593 1231 609 1265
rect 509 1193 609 1231
rect 667 1265 767 1281
rect 667 1231 683 1265
rect 751 1231 767 1265
rect 667 1193 767 1231
rect 825 1265 925 1281
rect 825 1231 841 1265
rect 909 1231 925 1265
rect 825 1193 925 1231
rect 983 1265 1083 1281
rect 983 1231 999 1265
rect 1067 1231 1083 1265
rect 983 1193 1083 1231
rect 1141 1265 1241 1281
rect 1141 1231 1157 1265
rect 1225 1231 1241 1265
rect 1141 1193 1241 1231
rect 1299 1265 1399 1281
rect 1299 1231 1315 1265
rect 1383 1231 1399 1265
rect 1299 1193 1399 1231
rect 1457 1265 1557 1281
rect 1457 1231 1473 1265
rect 1541 1231 1557 1265
rect 1457 1193 1557 1231
rect 1615 1265 1715 1281
rect 1615 1231 1631 1265
rect 1699 1231 1715 1265
rect 1615 1193 1715 1231
rect 1773 1265 1873 1281
rect 1773 1231 1789 1265
rect 1857 1231 1873 1265
rect 1773 1193 1873 1231
rect 1931 1265 2031 1281
rect 1931 1231 1947 1265
rect 2015 1231 2031 1265
rect 1931 1193 2031 1231
rect 2089 1265 2189 1281
rect 2089 1231 2105 1265
rect 2173 1231 2189 1265
rect 2089 1193 2189 1231
rect 2247 1265 2347 1281
rect 2247 1231 2263 1265
rect 2331 1231 2347 1265
rect 2247 1193 2347 1231
rect 2405 1265 2505 1281
rect 2405 1231 2421 1265
rect 2489 1231 2505 1265
rect 2405 1193 2505 1231
rect 2563 1265 2663 1281
rect 2563 1231 2579 1265
rect 2647 1231 2663 1265
rect 2563 1193 2663 1231
rect 2721 1265 2821 1281
rect 2721 1231 2737 1265
rect 2805 1231 2821 1265
rect 2721 1193 2821 1231
rect 2879 1265 2979 1281
rect 2879 1231 2895 1265
rect 2963 1231 2979 1265
rect 2879 1193 2979 1231
rect 3037 1265 3137 1281
rect 3037 1231 3053 1265
rect 3121 1231 3137 1265
rect 3037 1193 3137 1231
rect 3195 1265 3295 1281
rect 3195 1231 3211 1265
rect 3279 1231 3295 1265
rect 3195 1193 3295 1231
rect 193 155 293 193
rect 193 121 209 155
rect 277 121 293 155
rect 193 105 293 121
rect 351 155 451 193
rect 351 121 367 155
rect 435 121 451 155
rect 351 105 451 121
rect 509 155 609 193
rect 509 121 525 155
rect 593 121 609 155
rect 509 105 609 121
rect 667 155 767 193
rect 667 121 683 155
rect 751 121 767 155
rect 667 105 767 121
rect 825 155 925 193
rect 825 121 841 155
rect 909 121 925 155
rect 825 105 925 121
rect 983 155 1083 193
rect 983 121 999 155
rect 1067 121 1083 155
rect 983 105 1083 121
rect 1141 155 1241 193
rect 1141 121 1157 155
rect 1225 121 1241 155
rect 1141 105 1241 121
rect 1299 155 1399 193
rect 1299 121 1315 155
rect 1383 121 1399 155
rect 1299 105 1399 121
rect 1457 155 1557 193
rect 1457 121 1473 155
rect 1541 121 1557 155
rect 1457 105 1557 121
rect 1615 155 1715 193
rect 1615 121 1631 155
rect 1699 121 1715 155
rect 1615 105 1715 121
rect 1773 155 1873 193
rect 1773 121 1789 155
rect 1857 121 1873 155
rect 1773 105 1873 121
rect 1931 155 2031 193
rect 1931 121 1947 155
rect 2015 121 2031 155
rect 1931 105 2031 121
rect 2089 155 2189 193
rect 2089 121 2105 155
rect 2173 121 2189 155
rect 2089 105 2189 121
rect 2247 155 2347 193
rect 2247 121 2263 155
rect 2331 121 2347 155
rect 2247 105 2347 121
rect 2405 155 2505 193
rect 2405 121 2421 155
rect 2489 121 2505 155
rect 2405 105 2505 121
rect 2563 155 2663 193
rect 2563 121 2579 155
rect 2647 121 2663 155
rect 2563 105 2663 121
rect 2721 155 2821 193
rect 2721 121 2737 155
rect 2805 121 2821 155
rect 2721 105 2821 121
rect 2879 155 2979 193
rect 2879 121 2895 155
rect 2963 121 2979 155
rect 2879 105 2979 121
rect 3037 155 3137 193
rect 3037 121 3053 155
rect 3121 121 3137 155
rect 3037 105 3137 121
rect 3195 155 3295 193
rect 3195 121 3211 155
rect 3279 121 3295 155
rect 3195 105 3295 121
<< polycont >>
rect 209 2845 277 2879
rect 367 2845 435 2879
rect 525 2845 593 2879
rect 683 2845 751 2879
rect 841 2845 909 2879
rect 999 2845 1067 2879
rect 1157 2845 1225 2879
rect 1315 2845 1383 2879
rect 1473 2845 1541 2879
rect 1631 2845 1699 2879
rect 1789 2845 1857 2879
rect 1947 2845 2015 2879
rect 2105 2845 2173 2879
rect 2263 2845 2331 2879
rect 2421 2845 2489 2879
rect 2579 2845 2647 2879
rect 2737 2845 2805 2879
rect 2895 2845 2963 2879
rect 3053 2845 3121 2879
rect 3211 2845 3279 2879
rect 209 1717 277 1751
rect 367 1717 435 1751
rect 525 1717 593 1751
rect 683 1717 751 1751
rect 841 1717 909 1751
rect 999 1717 1067 1751
rect 1157 1717 1225 1751
rect 1315 1717 1383 1751
rect 1473 1717 1541 1751
rect 1631 1717 1699 1751
rect 1789 1717 1857 1751
rect 1947 1717 2015 1751
rect 2105 1717 2173 1751
rect 2263 1717 2331 1751
rect 2421 1717 2489 1751
rect 2579 1717 2647 1751
rect 2737 1717 2805 1751
rect 2895 1717 2963 1751
rect 3053 1717 3121 1751
rect 3211 1717 3279 1751
rect 209 1231 277 1265
rect 367 1231 435 1265
rect 525 1231 593 1265
rect 683 1231 751 1265
rect 841 1231 909 1265
rect 999 1231 1067 1265
rect 1157 1231 1225 1265
rect 1315 1231 1383 1265
rect 1473 1231 1541 1265
rect 1631 1231 1699 1265
rect 1789 1231 1857 1265
rect 1947 1231 2015 1265
rect 2105 1231 2173 1265
rect 2263 1231 2331 1265
rect 2421 1231 2489 1265
rect 2579 1231 2647 1265
rect 2737 1231 2805 1265
rect 2895 1231 2963 1265
rect 3053 1231 3121 1265
rect 3211 1231 3279 1265
rect 209 121 277 155
rect 367 121 435 155
rect 525 121 593 155
rect 683 121 751 155
rect 841 121 909 155
rect 999 121 1067 155
rect 1157 121 1225 155
rect 1315 121 1383 155
rect 1473 121 1541 155
rect 1631 121 1699 155
rect 1789 121 1857 155
rect 1947 121 2015 155
rect 2105 121 2173 155
rect 2263 121 2331 155
rect 2421 121 2489 155
rect 2579 121 2647 155
rect 2737 121 2805 155
rect 2895 121 2963 155
rect 3053 121 3121 155
rect 3211 121 3279 155
<< locali >>
rect 13 2983 109 3017
rect 3379 2983 3475 3017
rect 13 2921 47 2983
rect 3441 2921 3475 2983
rect 193 2845 209 2879
rect 277 2845 293 2879
rect 351 2845 367 2879
rect 435 2845 451 2879
rect 509 2845 525 2879
rect 593 2845 609 2879
rect 667 2845 683 2879
rect 751 2845 767 2879
rect 825 2845 841 2879
rect 909 2845 925 2879
rect 983 2845 999 2879
rect 1067 2845 1083 2879
rect 1141 2845 1157 2879
rect 1225 2845 1241 2879
rect 1299 2845 1315 2879
rect 1383 2845 1399 2879
rect 1457 2845 1473 2879
rect 1541 2845 1557 2879
rect 1615 2845 1631 2879
rect 1699 2845 1715 2879
rect 1773 2845 1789 2879
rect 1857 2845 1873 2879
rect 1931 2845 1947 2879
rect 2015 2845 2031 2879
rect 2089 2845 2105 2879
rect 2173 2845 2189 2879
rect 2247 2845 2263 2879
rect 2331 2845 2347 2879
rect 2405 2845 2421 2879
rect 2489 2845 2505 2879
rect 2563 2845 2579 2879
rect 2647 2845 2663 2879
rect 2721 2845 2737 2879
rect 2805 2845 2821 2879
rect 2879 2845 2895 2879
rect 2963 2845 2979 2879
rect 3037 2845 3053 2879
rect 3121 2845 3137 2879
rect 3195 2845 3211 2879
rect 3279 2845 3295 2879
rect 147 2786 181 2802
rect 147 1794 181 1810
rect 305 2786 339 2802
rect 305 1794 339 1810
rect 463 2786 497 2802
rect 463 1794 497 1810
rect 621 2786 655 2802
rect 621 1794 655 1810
rect 779 2786 813 2802
rect 779 1794 813 1810
rect 937 2786 971 2802
rect 937 1794 971 1810
rect 1095 2786 1129 2802
rect 1095 1794 1129 1810
rect 1253 2786 1287 2802
rect 1253 1794 1287 1810
rect 1411 2786 1445 2802
rect 1411 1794 1445 1810
rect 1569 2786 1603 2802
rect 1569 1794 1603 1810
rect 1727 2786 1761 2802
rect 1727 1794 1761 1810
rect 1885 2786 1919 2802
rect 1885 1794 1919 1810
rect 2043 2786 2077 2802
rect 2043 1794 2077 1810
rect 2201 2786 2235 2802
rect 2201 1794 2235 1810
rect 2359 2786 2393 2802
rect 2359 1794 2393 1810
rect 2517 2786 2551 2802
rect 2517 1794 2551 1810
rect 2675 2786 2709 2802
rect 2675 1794 2709 1810
rect 2833 2786 2867 2802
rect 2833 1794 2867 1810
rect 2991 2786 3025 2802
rect 2991 1794 3025 1810
rect 3149 2786 3183 2802
rect 3149 1794 3183 1810
rect 3307 2786 3341 2802
rect 3307 1794 3341 1810
rect 193 1717 209 1751
rect 277 1717 293 1751
rect 351 1717 367 1751
rect 435 1717 451 1751
rect 509 1717 525 1751
rect 593 1717 609 1751
rect 667 1717 683 1751
rect 751 1717 767 1751
rect 825 1717 841 1751
rect 909 1717 925 1751
rect 983 1717 999 1751
rect 1067 1717 1083 1751
rect 1141 1717 1157 1751
rect 1225 1717 1241 1751
rect 1299 1717 1315 1751
rect 1383 1717 1399 1751
rect 1457 1717 1473 1751
rect 1541 1717 1557 1751
rect 1615 1717 1631 1751
rect 1699 1717 1715 1751
rect 1773 1717 1789 1751
rect 1857 1717 1873 1751
rect 1931 1717 1947 1751
rect 2015 1717 2031 1751
rect 2089 1717 2105 1751
rect 2173 1717 2189 1751
rect 2247 1717 2263 1751
rect 2331 1717 2347 1751
rect 2405 1717 2421 1751
rect 2489 1717 2505 1751
rect 2563 1717 2579 1751
rect 2647 1717 2663 1751
rect 2721 1717 2737 1751
rect 2805 1717 2821 1751
rect 2879 1717 2895 1751
rect 2963 1717 2979 1751
rect 3037 1717 3053 1751
rect 3121 1717 3137 1751
rect 3195 1717 3211 1751
rect 3279 1717 3295 1751
rect 13 1613 47 1675
rect 3441 1613 3475 1675
rect 13 1579 109 1613
rect 3379 1579 3475 1613
rect 13 1369 109 1403
rect 3379 1369 3475 1403
rect 13 1307 47 1369
rect 3441 1307 3475 1369
rect 193 1231 209 1265
rect 277 1231 293 1265
rect 351 1231 367 1265
rect 435 1231 451 1265
rect 509 1231 525 1265
rect 593 1231 609 1265
rect 667 1231 683 1265
rect 751 1231 767 1265
rect 825 1231 841 1265
rect 909 1231 925 1265
rect 983 1231 999 1265
rect 1067 1231 1083 1265
rect 1141 1231 1157 1265
rect 1225 1231 1241 1265
rect 1299 1231 1315 1265
rect 1383 1231 1399 1265
rect 1457 1231 1473 1265
rect 1541 1231 1557 1265
rect 1615 1231 1631 1265
rect 1699 1231 1715 1265
rect 1773 1231 1789 1265
rect 1857 1231 1873 1265
rect 1931 1231 1947 1265
rect 2015 1231 2031 1265
rect 2089 1231 2105 1265
rect 2173 1231 2189 1265
rect 2247 1231 2263 1265
rect 2331 1231 2347 1265
rect 2405 1231 2421 1265
rect 2489 1231 2505 1265
rect 2563 1231 2579 1265
rect 2647 1231 2663 1265
rect 2721 1231 2737 1265
rect 2805 1231 2821 1265
rect 2879 1231 2895 1265
rect 2963 1231 2979 1265
rect 3037 1231 3053 1265
rect 3121 1231 3137 1265
rect 3195 1231 3211 1265
rect 3279 1231 3295 1265
rect 147 1181 181 1197
rect 147 189 181 205
rect 305 1181 339 1197
rect 305 189 339 205
rect 463 1181 497 1197
rect 463 189 497 205
rect 621 1181 655 1197
rect 621 189 655 205
rect 779 1181 813 1197
rect 779 189 813 205
rect 937 1181 971 1197
rect 937 189 971 205
rect 1095 1181 1129 1197
rect 1095 189 1129 205
rect 1253 1181 1287 1197
rect 1253 189 1287 205
rect 1411 1181 1445 1197
rect 1411 189 1445 205
rect 1569 1181 1603 1197
rect 1569 189 1603 205
rect 1727 1181 1761 1197
rect 1727 189 1761 205
rect 1885 1181 1919 1197
rect 1885 189 1919 205
rect 2043 1181 2077 1197
rect 2043 189 2077 205
rect 2201 1181 2235 1197
rect 2201 189 2235 205
rect 2359 1181 2393 1197
rect 2359 189 2393 205
rect 2517 1181 2551 1197
rect 2517 189 2551 205
rect 2675 1181 2709 1197
rect 2675 189 2709 205
rect 2833 1181 2867 1197
rect 2833 189 2867 205
rect 2991 1181 3025 1197
rect 2991 189 3025 205
rect 3149 1181 3183 1197
rect 3149 189 3183 205
rect 3307 1181 3341 1197
rect 3307 189 3341 205
rect 193 121 209 155
rect 277 121 293 155
rect 351 121 367 155
rect 435 121 451 155
rect 509 121 525 155
rect 593 121 609 155
rect 667 121 683 155
rect 751 121 767 155
rect 825 121 841 155
rect 909 121 925 155
rect 983 121 999 155
rect 1067 121 1083 155
rect 1141 121 1157 155
rect 1225 121 1241 155
rect 1299 121 1315 155
rect 1383 121 1399 155
rect 1457 121 1473 155
rect 1541 121 1557 155
rect 1615 121 1631 155
rect 1699 121 1715 155
rect 1773 121 1789 155
rect 1857 121 1873 155
rect 1931 121 1947 155
rect 2015 121 2031 155
rect 2089 121 2105 155
rect 2173 121 2189 155
rect 2247 121 2263 155
rect 2331 121 2347 155
rect 2405 121 2421 155
rect 2489 121 2505 155
rect 2563 121 2579 155
rect 2647 121 2663 155
rect 2721 121 2737 155
rect 2805 121 2821 155
rect 2879 121 2895 155
rect 2963 121 2979 155
rect 3037 121 3053 155
rect 3121 121 3137 155
rect 3195 121 3211 155
rect 3279 121 3295 155
rect 13 17 47 79
rect 3441 17 3475 79
rect 13 -17 109 17
rect 3379 -17 3475 17
<< viali >>
rect 13 1675 47 2921
rect 226 2845 260 2879
rect 384 2845 418 2879
rect 542 2845 576 2879
rect 700 2845 734 2879
rect 858 2845 892 2879
rect 1016 2845 1050 2879
rect 1174 2845 1208 2879
rect 1332 2845 1366 2879
rect 1490 2845 1524 2879
rect 1648 2845 1682 2879
rect 1806 2845 1840 2879
rect 1964 2845 1998 2879
rect 2122 2845 2156 2879
rect 2280 2845 2314 2879
rect 2438 2845 2472 2879
rect 2596 2845 2630 2879
rect 2754 2845 2788 2879
rect 2912 2845 2946 2879
rect 3070 2845 3104 2879
rect 3228 2845 3262 2879
rect 147 1810 181 2786
rect 305 1810 339 2786
rect 463 1810 497 2786
rect 621 1810 655 2786
rect 779 1810 813 2786
rect 937 1810 971 2786
rect 1095 1810 1129 2786
rect 1253 1810 1287 2786
rect 1411 1810 1445 2786
rect 1569 1810 1603 2786
rect 1727 1810 1761 2786
rect 1885 1810 1919 2786
rect 2043 1810 2077 2786
rect 2201 1810 2235 2786
rect 2359 1810 2393 2786
rect 2517 1810 2551 2786
rect 2675 1810 2709 2786
rect 2833 1810 2867 2786
rect 2991 1810 3025 2786
rect 3149 1810 3183 2786
rect 3307 1810 3341 2786
rect 226 1717 260 1751
rect 384 1717 418 1751
rect 542 1717 576 1751
rect 700 1717 734 1751
rect 858 1717 892 1751
rect 1016 1717 1050 1751
rect 1174 1717 1208 1751
rect 1332 1717 1366 1751
rect 1490 1717 1524 1751
rect 1648 1717 1682 1751
rect 1806 1717 1840 1751
rect 1964 1717 1998 1751
rect 2122 1717 2156 1751
rect 2280 1717 2314 1751
rect 2438 1717 2472 1751
rect 2596 1717 2630 1751
rect 2754 1717 2788 1751
rect 2912 1717 2946 1751
rect 3070 1717 3104 1751
rect 3228 1717 3262 1751
rect 3441 1675 3475 2921
rect 13 79 47 1307
rect 226 1231 260 1265
rect 384 1231 418 1265
rect 542 1231 576 1265
rect 700 1231 734 1265
rect 858 1231 892 1265
rect 1016 1231 1050 1265
rect 1174 1231 1208 1265
rect 1332 1231 1366 1265
rect 1490 1231 1524 1265
rect 1648 1231 1682 1265
rect 1806 1231 1840 1265
rect 1964 1231 1998 1265
rect 2122 1231 2156 1265
rect 2280 1231 2314 1265
rect 2438 1231 2472 1265
rect 2596 1231 2630 1265
rect 2754 1231 2788 1265
rect 2912 1231 2946 1265
rect 3070 1231 3104 1265
rect 3228 1231 3262 1265
rect 147 205 181 1181
rect 305 205 339 1181
rect 463 205 497 1181
rect 621 205 655 1181
rect 779 205 813 1181
rect 937 205 971 1181
rect 1095 205 1129 1181
rect 1253 205 1287 1181
rect 1411 205 1445 1181
rect 1569 205 1603 1181
rect 1727 205 1761 1181
rect 1885 205 1919 1181
rect 2043 205 2077 1181
rect 2201 205 2235 1181
rect 2359 205 2393 1181
rect 2517 205 2551 1181
rect 2675 205 2709 1181
rect 2833 205 2867 1181
rect 2991 205 3025 1181
rect 3149 205 3183 1181
rect 3307 205 3341 1181
rect 226 121 260 155
rect 384 121 418 155
rect 542 121 576 155
rect 700 121 734 155
rect 858 121 892 155
rect 1016 121 1050 155
rect 1174 121 1208 155
rect 1332 121 1366 155
rect 1490 121 1524 155
rect 1648 121 1682 155
rect 1806 121 1840 155
rect 1964 121 1998 155
rect 2122 121 2156 155
rect 2280 121 2314 155
rect 2438 121 2472 155
rect 2596 121 2630 155
rect 2754 121 2788 155
rect 2912 121 2946 155
rect 3070 121 3104 155
rect 3228 121 3262 155
rect 3441 79 3475 1307
<< metal1 >>
rect 7 2921 53 2933
rect 7 1675 13 2921
rect 47 2885 53 2921
rect 3435 2921 3481 2933
rect 3435 2885 3441 2921
rect 47 2879 3441 2885
rect 47 2845 226 2879
rect 260 2845 384 2879
rect 418 2845 542 2879
rect 576 2845 700 2879
rect 734 2845 858 2879
rect 892 2845 1016 2879
rect 1050 2845 1174 2879
rect 1208 2845 1332 2879
rect 1366 2845 1490 2879
rect 1524 2845 1648 2879
rect 1682 2845 1806 2879
rect 1840 2845 1964 2879
rect 1998 2845 2122 2879
rect 2156 2845 2280 2879
rect 2314 2845 2438 2879
rect 2472 2845 2596 2879
rect 2630 2845 2754 2879
rect 2788 2845 2912 2879
rect 2946 2845 3070 2879
rect 3104 2845 3228 2879
rect 3262 2845 3441 2879
rect 47 2839 3441 2845
rect 47 1757 59 2839
rect 141 2786 187 2839
rect 141 1810 147 2786
rect 181 1810 187 2786
rect 299 2786 345 2798
rect 299 1914 305 2786
rect 339 1914 345 2786
rect 457 2786 503 2839
rect 286 1810 296 1914
rect 348 1810 358 1914
rect 457 1810 463 2786
rect 497 1810 503 2786
rect 615 2786 661 2798
rect 615 1914 621 2786
rect 655 1914 661 2786
rect 773 2786 819 2839
rect 602 1810 612 1914
rect 664 1810 674 1914
rect 773 1810 779 2786
rect 813 1810 819 2786
rect 931 2786 977 2798
rect 931 1914 937 2786
rect 971 1914 977 2786
rect 1089 2786 1135 2839
rect 918 1810 928 1914
rect 980 1810 990 1914
rect 1089 1810 1095 2786
rect 1129 1810 1135 2786
rect 1247 2786 1293 2798
rect 1247 1914 1253 2786
rect 1287 1914 1293 2786
rect 1405 2786 1451 2839
rect 1234 1810 1244 1914
rect 1296 1810 1306 1914
rect 1405 1810 1411 2786
rect 1445 1810 1451 2786
rect 1563 2786 1609 2798
rect 1563 1914 1569 2786
rect 1603 1914 1609 2786
rect 1721 2786 1767 2839
rect 1550 1810 1560 1914
rect 1612 1810 1622 1914
rect 1721 1810 1727 2786
rect 1761 1810 1767 2786
rect 1879 2786 1925 2798
rect 1879 1914 1885 2786
rect 1919 1914 1925 2786
rect 2037 2786 2083 2839
rect 1866 1810 1876 1914
rect 1928 1810 1938 1914
rect 2037 1810 2043 2786
rect 2077 1810 2083 2786
rect 2195 2786 2241 2798
rect 2195 1914 2201 2786
rect 2235 1914 2241 2786
rect 2353 2786 2399 2839
rect 2182 1810 2192 1914
rect 2244 1810 2254 1914
rect 2353 1810 2359 2786
rect 2393 1810 2399 2786
rect 2511 2786 2557 2798
rect 2511 1914 2517 2786
rect 2551 1914 2557 2786
rect 2669 2786 2715 2839
rect 2498 1810 2508 1914
rect 2560 1810 2570 1914
rect 2669 1810 2675 2786
rect 2709 1810 2715 2786
rect 2827 2786 2873 2798
rect 2827 1914 2833 2786
rect 2867 1914 2873 2786
rect 2985 2786 3031 2839
rect 2814 1810 2824 1914
rect 2876 1810 2886 1914
rect 2985 1810 2991 2786
rect 3025 1810 3031 2786
rect 3143 2786 3189 2798
rect 3143 1914 3149 2786
rect 3183 1914 3189 2786
rect 3301 2786 3347 2839
rect 3130 1810 3140 1914
rect 3192 1810 3202 1914
rect 3301 1810 3307 2786
rect 3341 1810 3347 2786
rect 141 1757 187 1810
rect 299 1798 345 1810
rect 457 1798 503 1810
rect 615 1798 661 1810
rect 773 1798 819 1810
rect 931 1798 977 1810
rect 1089 1798 1135 1810
rect 1247 1798 1293 1810
rect 1405 1798 1451 1810
rect 1563 1798 1609 1810
rect 1721 1798 1767 1810
rect 1879 1798 1925 1810
rect 2037 1798 2083 1810
rect 2195 1798 2241 1810
rect 2353 1798 2399 1810
rect 2511 1798 2557 1810
rect 2669 1798 2715 1810
rect 2827 1798 2873 1810
rect 2985 1798 3031 1810
rect 3143 1798 3189 1810
rect 3301 1757 3347 1810
rect 3429 1757 3441 2839
rect 47 1751 3441 1757
rect 47 1717 226 1751
rect 260 1717 384 1751
rect 418 1717 542 1751
rect 576 1717 700 1751
rect 734 1717 858 1751
rect 892 1717 1016 1751
rect 1050 1717 1174 1751
rect 1208 1717 1332 1751
rect 1366 1717 1490 1751
rect 1524 1717 1648 1751
rect 1682 1717 1806 1751
rect 1840 1717 1964 1751
rect 1998 1717 2122 1751
rect 2156 1717 2280 1751
rect 2314 1717 2438 1751
rect 2472 1717 2596 1751
rect 2630 1717 2754 1751
rect 2788 1717 2912 1751
rect 2946 1717 3070 1751
rect 3104 1717 3228 1751
rect 3262 1717 3441 1751
rect 47 1711 3441 1717
rect 47 1675 53 1711
rect 7 1663 53 1675
rect 3435 1675 3441 1711
rect 3475 1675 3481 2921
rect 3435 1663 3481 1675
rect -65 1544 3553 1555
rect -65 1440 296 1544
rect 348 1440 612 1544
rect 664 1440 928 1544
rect 980 1440 1244 1544
rect 1296 1440 1560 1544
rect 1612 1440 1876 1544
rect 1928 1440 2192 1544
rect 2244 1440 2508 1544
rect 2560 1440 2824 1544
rect 2876 1440 3140 1544
rect 3192 1440 3553 1544
rect -65 1427 3553 1440
rect 7 1307 53 1319
rect 7 79 13 1307
rect 47 1271 53 1307
rect 3435 1307 3481 1319
rect 3435 1271 3441 1307
rect 47 1265 3441 1271
rect 47 1231 226 1265
rect 260 1231 384 1265
rect 418 1231 542 1265
rect 576 1231 700 1265
rect 734 1231 858 1265
rect 892 1231 1016 1265
rect 1050 1231 1174 1265
rect 1208 1231 1332 1265
rect 1366 1231 1490 1265
rect 1524 1231 1648 1265
rect 1682 1231 1806 1265
rect 1840 1231 1964 1265
rect 1998 1231 2122 1265
rect 2156 1231 2280 1265
rect 2314 1231 2438 1265
rect 2472 1231 2596 1265
rect 2630 1231 2754 1265
rect 2788 1231 2912 1265
rect 2946 1231 3070 1265
rect 3104 1231 3228 1265
rect 3262 1231 3441 1265
rect 47 1225 3441 1231
rect 47 161 53 1225
rect 141 1181 187 1193
rect 299 1181 345 1193
rect 457 1181 503 1193
rect 615 1181 661 1193
rect 773 1181 819 1193
rect 931 1181 977 1193
rect 1089 1181 1135 1193
rect 1247 1181 1293 1193
rect 1405 1181 1451 1193
rect 1563 1181 1609 1193
rect 1721 1181 1767 1193
rect 1879 1181 1925 1193
rect 2037 1181 2083 1193
rect 2195 1181 2241 1193
rect 2353 1181 2399 1193
rect 2511 1181 2557 1193
rect 2669 1181 2715 1193
rect 2827 1181 2873 1193
rect 2985 1181 3031 1193
rect 3143 1181 3189 1193
rect 3301 1181 3347 1225
rect 141 205 147 1181
rect 181 205 187 1181
rect 286 1077 296 1181
rect 348 1077 358 1181
rect 141 161 187 205
rect 299 205 305 1077
rect 339 205 345 1077
rect 299 193 345 205
rect 457 205 463 1181
rect 497 205 503 1181
rect 602 1077 612 1181
rect 664 1077 674 1181
rect 457 161 503 205
rect 615 205 621 1077
rect 655 205 661 1077
rect 615 193 661 205
rect 773 205 779 1181
rect 813 205 819 1181
rect 918 1077 928 1181
rect 980 1077 990 1181
rect 773 161 819 205
rect 931 205 937 1077
rect 971 205 977 1077
rect 931 193 977 205
rect 1089 205 1095 1181
rect 1129 205 1135 1181
rect 1234 1077 1244 1181
rect 1296 1077 1306 1181
rect 1089 161 1135 205
rect 1247 205 1253 1077
rect 1287 205 1293 1077
rect 1247 193 1293 205
rect 1405 205 1411 1181
rect 1445 205 1451 1181
rect 1550 1077 1560 1181
rect 1612 1077 1622 1181
rect 1405 161 1451 205
rect 1563 205 1569 1077
rect 1603 205 1609 1077
rect 1563 193 1609 205
rect 1721 205 1727 1181
rect 1761 205 1767 1181
rect 1866 1077 1876 1181
rect 1928 1077 1938 1181
rect 1721 161 1767 205
rect 1879 205 1885 1077
rect 1919 205 1925 1077
rect 1879 193 1925 205
rect 2037 205 2043 1181
rect 2077 205 2083 1181
rect 2182 1077 2192 1181
rect 2244 1077 2254 1181
rect 2037 161 2083 205
rect 2195 205 2201 1077
rect 2235 205 2241 1077
rect 2195 193 2241 205
rect 2353 205 2359 1181
rect 2393 205 2399 1181
rect 2498 1077 2508 1181
rect 2560 1077 2570 1181
rect 2353 161 2399 205
rect 2511 205 2517 1077
rect 2551 205 2557 1077
rect 2511 193 2557 205
rect 2669 205 2675 1181
rect 2709 205 2715 1181
rect 2814 1077 2824 1181
rect 2876 1077 2886 1181
rect 2669 161 2715 205
rect 2827 205 2833 1077
rect 2867 205 2873 1077
rect 2827 193 2873 205
rect 2985 205 2991 1181
rect 3025 205 3031 1181
rect 3130 1077 3140 1181
rect 3192 1077 3202 1181
rect 2985 161 3031 205
rect 3143 205 3149 1077
rect 3183 205 3189 1077
rect 3143 193 3189 205
rect 3301 205 3307 1181
rect 3341 205 3347 1181
rect 3301 161 3347 205
rect 3435 161 3441 1225
rect 47 155 3441 161
rect 47 121 226 155
rect 260 121 384 155
rect 418 121 542 155
rect 576 121 700 155
rect 734 121 858 155
rect 892 121 1016 155
rect 1050 121 1174 155
rect 1208 121 1332 155
rect 1366 121 1490 155
rect 1524 121 1648 155
rect 1682 121 1806 155
rect 1840 121 1964 155
rect 1998 121 2122 155
rect 2156 121 2280 155
rect 2314 121 2438 155
rect 2472 121 2596 155
rect 2630 121 2754 155
rect 2788 121 2912 155
rect 2946 121 3070 155
rect 3104 121 3228 155
rect 3262 121 3441 155
rect 47 115 3441 121
rect 47 79 53 115
rect 7 67 53 79
rect 3435 79 3441 115
rect 3475 79 3481 1307
rect 3435 67 3481 79
<< via1 >>
rect 296 1810 305 1914
rect 305 1810 339 1914
rect 339 1810 348 1914
rect 612 1810 621 1914
rect 621 1810 655 1914
rect 655 1810 664 1914
rect 928 1810 937 1914
rect 937 1810 971 1914
rect 971 1810 980 1914
rect 1244 1810 1253 1914
rect 1253 1810 1287 1914
rect 1287 1810 1296 1914
rect 1560 1810 1569 1914
rect 1569 1810 1603 1914
rect 1603 1810 1612 1914
rect 1876 1810 1885 1914
rect 1885 1810 1919 1914
rect 1919 1810 1928 1914
rect 2192 1810 2201 1914
rect 2201 1810 2235 1914
rect 2235 1810 2244 1914
rect 2508 1810 2517 1914
rect 2517 1810 2551 1914
rect 2551 1810 2560 1914
rect 2824 1810 2833 1914
rect 2833 1810 2867 1914
rect 2867 1810 2876 1914
rect 3140 1810 3149 1914
rect 3149 1810 3183 1914
rect 3183 1810 3192 1914
rect 296 1440 348 1544
rect 612 1440 664 1544
rect 928 1440 980 1544
rect 1244 1440 1296 1544
rect 1560 1440 1612 1544
rect 1876 1440 1928 1544
rect 2192 1440 2244 1544
rect 2508 1440 2560 1544
rect 2824 1440 2876 1544
rect 3140 1440 3192 1544
rect 296 1077 305 1181
rect 305 1077 339 1181
rect 339 1077 348 1181
rect 612 1077 621 1181
rect 621 1077 655 1181
rect 655 1077 664 1181
rect 928 1077 937 1181
rect 937 1077 971 1181
rect 971 1077 980 1181
rect 1244 1077 1253 1181
rect 1253 1077 1287 1181
rect 1287 1077 1296 1181
rect 1560 1077 1569 1181
rect 1569 1077 1603 1181
rect 1603 1077 1612 1181
rect 1876 1077 1885 1181
rect 1885 1077 1919 1181
rect 1919 1077 1928 1181
rect 2192 1077 2201 1181
rect 2201 1077 2235 1181
rect 2235 1077 2244 1181
rect 2508 1077 2517 1181
rect 2517 1077 2551 1181
rect 2551 1077 2560 1181
rect 2824 1077 2833 1181
rect 2833 1077 2867 1181
rect 2867 1077 2876 1181
rect 3140 1077 3149 1181
rect 3149 1077 3183 1181
rect 3183 1077 3192 1181
<< metal2 >>
rect 296 1914 348 1924
rect 296 1544 348 1810
rect 296 1181 348 1440
rect 296 1067 348 1077
rect 612 1914 664 1924
rect 612 1544 664 1810
rect 612 1181 664 1440
rect 612 1067 664 1077
rect 928 1914 980 1924
rect 928 1544 980 1810
rect 928 1181 980 1440
rect 928 1067 980 1077
rect 1244 1914 1296 1924
rect 1244 1544 1296 1810
rect 1244 1181 1296 1440
rect 1244 1067 1296 1077
rect 1560 1914 1612 1924
rect 1560 1544 1612 1810
rect 1560 1181 1612 1440
rect 1560 1067 1612 1077
rect 1876 1914 1928 1924
rect 1876 1544 1928 1810
rect 1876 1181 1928 1440
rect 1876 1067 1928 1077
rect 2192 1914 2244 1924
rect 2192 1544 2244 1810
rect 2192 1181 2244 1440
rect 2192 1067 2244 1077
rect 2508 1914 2560 1924
rect 2508 1544 2560 1810
rect 2508 1181 2560 1440
rect 2508 1067 2560 1077
rect 2824 1914 2876 1924
rect 2824 1544 2876 1810
rect 2824 1181 2876 1440
rect 2824 1067 2876 1077
rect 3140 1914 3192 1924
rect 3140 1544 3192 1810
rect 3140 1181 3192 1440
rect 3140 1067 3192 1077
<< labels >>
flabel metal1 -54 1487 -54 1487 1 FreeSans 400 0 0 0 esd
port 1 n
flabel metal1 30 2927 30 2927 1 FreeSans 400 0 0 0 VDD
port 2 n power bidirectional
flabel metal1 30 71 30 71 1 FreeSans 400 0 0 0 VSS
port 3 n power bidirectional
<< end >>
