magic
tech sky130A
magscale 1 2
timestamp 1654549423
<< nmos >>
rect -2997 -140 -2877 140
rect -2819 -140 -2699 140
rect -2641 -140 -2521 140
rect -2463 -140 -2343 140
rect -2285 -140 -2165 140
rect -2107 -140 -1987 140
rect -1929 -140 -1809 140
rect -1751 -140 -1631 140
rect -1573 -140 -1453 140
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
rect 1453 -140 1573 140
rect 1631 -140 1751 140
rect 1809 -140 1929 140
rect 1987 -140 2107 140
rect 2165 -140 2285 140
rect 2343 -140 2463 140
rect 2521 -140 2641 140
rect 2699 -140 2819 140
rect 2877 -140 2997 140
<< ndiff >>
rect -3055 128 -2997 140
rect -3055 -128 -3043 128
rect -3009 -128 -2997 128
rect -3055 -140 -2997 -128
rect -2877 128 -2819 140
rect -2877 -128 -2865 128
rect -2831 -128 -2819 128
rect -2877 -140 -2819 -128
rect -2699 128 -2641 140
rect -2699 -128 -2687 128
rect -2653 -128 -2641 128
rect -2699 -140 -2641 -128
rect -2521 128 -2463 140
rect -2521 -128 -2509 128
rect -2475 -128 -2463 128
rect -2521 -140 -2463 -128
rect -2343 128 -2285 140
rect -2343 -128 -2331 128
rect -2297 -128 -2285 128
rect -2343 -140 -2285 -128
rect -2165 128 -2107 140
rect -2165 -128 -2153 128
rect -2119 -128 -2107 128
rect -2165 -140 -2107 -128
rect -1987 128 -1929 140
rect -1987 -128 -1975 128
rect -1941 -128 -1929 128
rect -1987 -140 -1929 -128
rect -1809 128 -1751 140
rect -1809 -128 -1797 128
rect -1763 -128 -1751 128
rect -1809 -140 -1751 -128
rect -1631 128 -1573 140
rect -1631 -128 -1619 128
rect -1585 -128 -1573 128
rect -1631 -140 -1573 -128
rect -1453 128 -1395 140
rect -1453 -128 -1441 128
rect -1407 -128 -1395 128
rect -1453 -140 -1395 -128
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
rect 1395 128 1453 140
rect 1395 -128 1407 128
rect 1441 -128 1453 128
rect 1395 -140 1453 -128
rect 1573 128 1631 140
rect 1573 -128 1585 128
rect 1619 -128 1631 128
rect 1573 -140 1631 -128
rect 1751 128 1809 140
rect 1751 -128 1763 128
rect 1797 -128 1809 128
rect 1751 -140 1809 -128
rect 1929 128 1987 140
rect 1929 -128 1941 128
rect 1975 -128 1987 128
rect 1929 -140 1987 -128
rect 2107 128 2165 140
rect 2107 -128 2119 128
rect 2153 -128 2165 128
rect 2107 -140 2165 -128
rect 2285 128 2343 140
rect 2285 -128 2297 128
rect 2331 -128 2343 128
rect 2285 -140 2343 -128
rect 2463 128 2521 140
rect 2463 -128 2475 128
rect 2509 -128 2521 128
rect 2463 -140 2521 -128
rect 2641 128 2699 140
rect 2641 -128 2653 128
rect 2687 -128 2699 128
rect 2641 -140 2699 -128
rect 2819 128 2877 140
rect 2819 -128 2831 128
rect 2865 -128 2877 128
rect 2819 -140 2877 -128
rect 2997 128 3055 140
rect 2997 -128 3009 128
rect 3043 -128 3055 128
rect 2997 -140 3055 -128
<< ndiffc >>
rect -3043 -128 -3009 128
rect -2865 -128 -2831 128
rect -2687 -128 -2653 128
rect -2509 -128 -2475 128
rect -2331 -128 -2297 128
rect -2153 -128 -2119 128
rect -1975 -128 -1941 128
rect -1797 -128 -1763 128
rect -1619 -128 -1585 128
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
rect 1585 -128 1619 128
rect 1763 -128 1797 128
rect 1941 -128 1975 128
rect 2119 -128 2153 128
rect 2297 -128 2331 128
rect 2475 -128 2509 128
rect 2653 -128 2687 128
rect 2831 -128 2865 128
rect 3009 -128 3043 128
<< poly >>
rect -2979 212 -2895 228
rect -2979 195 -2963 212
rect -2997 178 -2963 195
rect -2911 195 -2895 212
rect -2801 212 -2717 228
rect -2801 195 -2785 212
rect -2911 178 -2877 195
rect -2997 140 -2877 178
rect -2819 178 -2785 195
rect -2733 195 -2717 212
rect -2623 212 -2539 228
rect -2623 195 -2607 212
rect -2733 178 -2699 195
rect -2819 140 -2699 178
rect -2641 178 -2607 195
rect -2555 195 -2539 212
rect -2445 212 -2361 228
rect -2445 195 -2429 212
rect -2555 178 -2521 195
rect -2641 140 -2521 178
rect -2463 178 -2429 195
rect -2377 195 -2361 212
rect -2267 212 -2183 228
rect -2267 195 -2251 212
rect -2377 178 -2343 195
rect -2463 140 -2343 178
rect -2285 178 -2251 195
rect -2199 195 -2183 212
rect -2089 212 -2005 228
rect -2089 195 -2073 212
rect -2199 178 -2165 195
rect -2285 140 -2165 178
rect -2107 178 -2073 195
rect -2021 195 -2005 212
rect -1911 212 -1827 228
rect -1911 195 -1895 212
rect -2021 178 -1987 195
rect -2107 140 -1987 178
rect -1929 178 -1895 195
rect -1843 195 -1827 212
rect -1733 212 -1649 228
rect -1733 195 -1717 212
rect -1843 178 -1809 195
rect -1929 140 -1809 178
rect -1751 178 -1717 195
rect -1665 195 -1649 212
rect -1555 212 -1471 228
rect -1555 195 -1539 212
rect -1665 178 -1631 195
rect -1751 140 -1631 178
rect -1573 178 -1539 195
rect -1487 195 -1471 212
rect -1377 212 -1293 228
rect -1377 195 -1361 212
rect -1487 178 -1453 195
rect -1573 140 -1453 178
rect -1395 178 -1361 195
rect -1309 195 -1293 212
rect -1199 212 -1115 228
rect -1199 195 -1183 212
rect -1309 178 -1275 195
rect -1395 140 -1275 178
rect -1217 178 -1183 195
rect -1131 195 -1115 212
rect -1021 212 -937 228
rect -1021 195 -1005 212
rect -1131 178 -1097 195
rect -1217 140 -1097 178
rect -1039 178 -1005 195
rect -953 195 -937 212
rect -843 212 -759 228
rect -843 195 -827 212
rect -953 178 -919 195
rect -1039 140 -919 178
rect -861 178 -827 195
rect -775 195 -759 212
rect -665 212 -581 228
rect -665 195 -649 212
rect -775 178 -741 195
rect -861 140 -741 178
rect -683 178 -649 195
rect -597 195 -581 212
rect -487 212 -403 228
rect -487 195 -471 212
rect -597 178 -563 195
rect -683 140 -563 178
rect -505 178 -471 195
rect -419 195 -403 212
rect -309 212 -225 228
rect -309 195 -293 212
rect -419 178 -385 195
rect -505 140 -385 178
rect -327 178 -293 195
rect -241 195 -225 212
rect -131 212 -47 228
rect -131 195 -115 212
rect -241 178 -207 195
rect -327 140 -207 178
rect -149 178 -115 195
rect -63 195 -47 212
rect 47 212 131 228
rect 47 195 63 212
rect -63 178 -29 195
rect -149 140 -29 178
rect 29 178 63 195
rect 115 195 131 212
rect 225 212 309 228
rect 225 195 241 212
rect 115 178 149 195
rect 29 140 149 178
rect 207 178 241 195
rect 293 195 309 212
rect 403 212 487 228
rect 403 195 419 212
rect 293 178 327 195
rect 207 140 327 178
rect 385 178 419 195
rect 471 195 487 212
rect 581 212 665 228
rect 581 195 597 212
rect 471 178 505 195
rect 385 140 505 178
rect 563 178 597 195
rect 649 195 665 212
rect 759 212 843 228
rect 759 195 775 212
rect 649 178 683 195
rect 563 140 683 178
rect 741 178 775 195
rect 827 195 843 212
rect 937 212 1021 228
rect 937 195 953 212
rect 827 178 861 195
rect 741 140 861 178
rect 919 178 953 195
rect 1005 195 1021 212
rect 1115 212 1199 228
rect 1115 195 1131 212
rect 1005 178 1039 195
rect 919 140 1039 178
rect 1097 178 1131 195
rect 1183 195 1199 212
rect 1293 212 1377 228
rect 1293 195 1309 212
rect 1183 178 1217 195
rect 1097 140 1217 178
rect 1275 178 1309 195
rect 1361 195 1377 212
rect 1471 212 1555 228
rect 1471 195 1487 212
rect 1361 178 1395 195
rect 1275 140 1395 178
rect 1453 178 1487 195
rect 1539 195 1555 212
rect 1649 212 1733 228
rect 1649 195 1665 212
rect 1539 178 1573 195
rect 1453 140 1573 178
rect 1631 178 1665 195
rect 1717 195 1733 212
rect 1827 212 1911 228
rect 1827 195 1843 212
rect 1717 178 1751 195
rect 1631 140 1751 178
rect 1809 178 1843 195
rect 1895 195 1911 212
rect 2005 212 2089 228
rect 2005 195 2021 212
rect 1895 178 1929 195
rect 1809 140 1929 178
rect 1987 178 2021 195
rect 2073 195 2089 212
rect 2183 212 2267 228
rect 2183 195 2199 212
rect 2073 178 2107 195
rect 1987 140 2107 178
rect 2165 178 2199 195
rect 2251 195 2267 212
rect 2361 212 2445 228
rect 2361 195 2377 212
rect 2251 178 2285 195
rect 2165 140 2285 178
rect 2343 178 2377 195
rect 2429 195 2445 212
rect 2539 212 2623 228
rect 2539 195 2555 212
rect 2429 178 2463 195
rect 2343 140 2463 178
rect 2521 178 2555 195
rect 2607 195 2623 212
rect 2717 212 2801 228
rect 2717 195 2733 212
rect 2607 178 2641 195
rect 2521 140 2641 178
rect 2699 178 2733 195
rect 2785 195 2801 212
rect 2895 212 2979 228
rect 2895 195 2911 212
rect 2785 178 2819 195
rect 2699 140 2819 178
rect 2877 178 2911 195
rect 2963 195 2979 212
rect 2963 178 2997 195
rect 2877 140 2997 178
rect -2997 -178 -2877 -140
rect -2997 -195 -2963 -178
rect -2979 -212 -2963 -195
rect -2911 -195 -2877 -178
rect -2819 -178 -2699 -140
rect -2819 -195 -2785 -178
rect -2911 -212 -2895 -195
rect -2979 -228 -2895 -212
rect -2801 -212 -2785 -195
rect -2733 -195 -2699 -178
rect -2641 -178 -2521 -140
rect -2641 -195 -2607 -178
rect -2733 -212 -2717 -195
rect -2801 -228 -2717 -212
rect -2623 -212 -2607 -195
rect -2555 -195 -2521 -178
rect -2463 -178 -2343 -140
rect -2463 -195 -2429 -178
rect -2555 -212 -2539 -195
rect -2623 -228 -2539 -212
rect -2445 -212 -2429 -195
rect -2377 -195 -2343 -178
rect -2285 -178 -2165 -140
rect -2285 -195 -2251 -178
rect -2377 -212 -2361 -195
rect -2445 -228 -2361 -212
rect -2267 -212 -2251 -195
rect -2199 -195 -2165 -178
rect -2107 -178 -1987 -140
rect -2107 -195 -2073 -178
rect -2199 -212 -2183 -195
rect -2267 -228 -2183 -212
rect -2089 -212 -2073 -195
rect -2021 -195 -1987 -178
rect -1929 -178 -1809 -140
rect -1929 -195 -1895 -178
rect -2021 -212 -2005 -195
rect -2089 -228 -2005 -212
rect -1911 -212 -1895 -195
rect -1843 -195 -1809 -178
rect -1751 -178 -1631 -140
rect -1751 -195 -1717 -178
rect -1843 -212 -1827 -195
rect -1911 -228 -1827 -212
rect -1733 -212 -1717 -195
rect -1665 -195 -1631 -178
rect -1573 -178 -1453 -140
rect -1573 -195 -1539 -178
rect -1665 -212 -1649 -195
rect -1733 -228 -1649 -212
rect -1555 -212 -1539 -195
rect -1487 -195 -1453 -178
rect -1395 -178 -1275 -140
rect -1395 -195 -1361 -178
rect -1487 -212 -1471 -195
rect -1555 -228 -1471 -212
rect -1377 -212 -1361 -195
rect -1309 -195 -1275 -178
rect -1217 -178 -1097 -140
rect -1217 -195 -1183 -178
rect -1309 -212 -1293 -195
rect -1377 -228 -1293 -212
rect -1199 -212 -1183 -195
rect -1131 -195 -1097 -178
rect -1039 -178 -919 -140
rect -1039 -195 -1005 -178
rect -1131 -212 -1115 -195
rect -1199 -228 -1115 -212
rect -1021 -212 -1005 -195
rect -953 -195 -919 -178
rect -861 -178 -741 -140
rect -861 -195 -827 -178
rect -953 -212 -937 -195
rect -1021 -228 -937 -212
rect -843 -212 -827 -195
rect -775 -195 -741 -178
rect -683 -178 -563 -140
rect -683 -195 -649 -178
rect -775 -212 -759 -195
rect -843 -228 -759 -212
rect -665 -212 -649 -195
rect -597 -195 -563 -178
rect -505 -178 -385 -140
rect -505 -195 -471 -178
rect -597 -212 -581 -195
rect -665 -228 -581 -212
rect -487 -212 -471 -195
rect -419 -195 -385 -178
rect -327 -178 -207 -140
rect -327 -195 -293 -178
rect -419 -212 -403 -195
rect -487 -228 -403 -212
rect -309 -212 -293 -195
rect -241 -195 -207 -178
rect -149 -178 -29 -140
rect -149 -195 -115 -178
rect -241 -212 -225 -195
rect -309 -228 -225 -212
rect -131 -212 -115 -195
rect -63 -195 -29 -178
rect 29 -178 149 -140
rect 29 -195 63 -178
rect -63 -212 -47 -195
rect -131 -228 -47 -212
rect 47 -212 63 -195
rect 115 -195 149 -178
rect 207 -178 327 -140
rect 207 -195 241 -178
rect 115 -212 131 -195
rect 47 -228 131 -212
rect 225 -212 241 -195
rect 293 -195 327 -178
rect 385 -178 505 -140
rect 385 -195 419 -178
rect 293 -212 309 -195
rect 225 -228 309 -212
rect 403 -212 419 -195
rect 471 -195 505 -178
rect 563 -178 683 -140
rect 563 -195 597 -178
rect 471 -212 487 -195
rect 403 -228 487 -212
rect 581 -212 597 -195
rect 649 -195 683 -178
rect 741 -178 861 -140
rect 741 -195 775 -178
rect 649 -212 665 -195
rect 581 -228 665 -212
rect 759 -212 775 -195
rect 827 -195 861 -178
rect 919 -178 1039 -140
rect 919 -195 953 -178
rect 827 -212 843 -195
rect 759 -228 843 -212
rect 937 -212 953 -195
rect 1005 -195 1039 -178
rect 1097 -178 1217 -140
rect 1097 -195 1131 -178
rect 1005 -212 1021 -195
rect 937 -228 1021 -212
rect 1115 -212 1131 -195
rect 1183 -195 1217 -178
rect 1275 -178 1395 -140
rect 1275 -195 1309 -178
rect 1183 -212 1199 -195
rect 1115 -228 1199 -212
rect 1293 -212 1309 -195
rect 1361 -195 1395 -178
rect 1453 -178 1573 -140
rect 1453 -195 1487 -178
rect 1361 -212 1377 -195
rect 1293 -228 1377 -212
rect 1471 -212 1487 -195
rect 1539 -195 1573 -178
rect 1631 -178 1751 -140
rect 1631 -195 1665 -178
rect 1539 -212 1555 -195
rect 1471 -228 1555 -212
rect 1649 -212 1665 -195
rect 1717 -195 1751 -178
rect 1809 -178 1929 -140
rect 1809 -195 1843 -178
rect 1717 -212 1733 -195
rect 1649 -228 1733 -212
rect 1827 -212 1843 -195
rect 1895 -195 1929 -178
rect 1987 -178 2107 -140
rect 1987 -195 2021 -178
rect 1895 -212 1911 -195
rect 1827 -228 1911 -212
rect 2005 -212 2021 -195
rect 2073 -195 2107 -178
rect 2165 -178 2285 -140
rect 2165 -195 2199 -178
rect 2073 -212 2089 -195
rect 2005 -228 2089 -212
rect 2183 -212 2199 -195
rect 2251 -195 2285 -178
rect 2343 -178 2463 -140
rect 2343 -195 2377 -178
rect 2251 -212 2267 -195
rect 2183 -228 2267 -212
rect 2361 -212 2377 -195
rect 2429 -195 2463 -178
rect 2521 -178 2641 -140
rect 2521 -195 2555 -178
rect 2429 -212 2445 -195
rect 2361 -228 2445 -212
rect 2539 -212 2555 -195
rect 2607 -195 2641 -178
rect 2699 -178 2819 -140
rect 2699 -195 2733 -178
rect 2607 -212 2623 -195
rect 2539 -228 2623 -212
rect 2717 -212 2733 -195
rect 2785 -195 2819 -178
rect 2877 -178 2997 -140
rect 2877 -195 2911 -178
rect 2785 -212 2801 -195
rect 2717 -228 2801 -212
rect 2895 -212 2911 -195
rect 2963 -195 2997 -178
rect 2963 -212 2979 -195
rect 2895 -228 2979 -212
<< polycont >>
rect -2963 178 -2911 212
rect -2785 178 -2733 212
rect -2607 178 -2555 212
rect -2429 178 -2377 212
rect -2251 178 -2199 212
rect -2073 178 -2021 212
rect -1895 178 -1843 212
rect -1717 178 -1665 212
rect -1539 178 -1487 212
rect -1361 178 -1309 212
rect -1183 178 -1131 212
rect -1005 178 -953 212
rect -827 178 -775 212
rect -649 178 -597 212
rect -471 178 -419 212
rect -293 178 -241 212
rect -115 178 -63 212
rect 63 178 115 212
rect 241 178 293 212
rect 419 178 471 212
rect 597 178 649 212
rect 775 178 827 212
rect 953 178 1005 212
rect 1131 178 1183 212
rect 1309 178 1361 212
rect 1487 178 1539 212
rect 1665 178 1717 212
rect 1843 178 1895 212
rect 2021 178 2073 212
rect 2199 178 2251 212
rect 2377 178 2429 212
rect 2555 178 2607 212
rect 2733 178 2785 212
rect 2911 178 2963 212
rect -2963 -212 -2911 -178
rect -2785 -212 -2733 -178
rect -2607 -212 -2555 -178
rect -2429 -212 -2377 -178
rect -2251 -212 -2199 -178
rect -2073 -212 -2021 -178
rect -1895 -212 -1843 -178
rect -1717 -212 -1665 -178
rect -1539 -212 -1487 -178
rect -1361 -212 -1309 -178
rect -1183 -212 -1131 -178
rect -1005 -212 -953 -178
rect -827 -212 -775 -178
rect -649 -212 -597 -178
rect -471 -212 -419 -178
rect -293 -212 -241 -178
rect -115 -212 -63 -178
rect 63 -212 115 -178
rect 241 -212 293 -178
rect 419 -212 471 -178
rect 597 -212 649 -178
rect 775 -212 827 -178
rect 953 -212 1005 -178
rect 1131 -212 1183 -178
rect 1309 -212 1361 -178
rect 1487 -212 1539 -178
rect 1665 -212 1717 -178
rect 1843 -212 1895 -178
rect 2021 -212 2073 -178
rect 2199 -212 2251 -178
rect 2377 -212 2429 -178
rect 2555 -212 2607 -178
rect 2733 -212 2785 -178
rect 2911 -212 2963 -178
<< locali >>
rect -2979 178 -2963 212
rect -2911 178 -2895 212
rect -2801 178 -2785 212
rect -2733 178 -2717 212
rect -2623 178 -2607 212
rect -2555 178 -2539 212
rect -2445 178 -2429 212
rect -2377 178 -2361 212
rect -2267 178 -2251 212
rect -2199 178 -2183 212
rect -2089 178 -2073 212
rect -2021 178 -2005 212
rect -1911 178 -1895 212
rect -1843 178 -1827 212
rect -1733 178 -1717 212
rect -1665 178 -1649 212
rect -1555 178 -1539 212
rect -1487 178 -1471 212
rect -1377 178 -1361 212
rect -1309 178 -1293 212
rect -1199 178 -1183 212
rect -1131 178 -1115 212
rect -1021 178 -1005 212
rect -953 178 -937 212
rect -843 178 -827 212
rect -775 178 -759 212
rect -665 178 -649 212
rect -597 178 -581 212
rect -487 178 -471 212
rect -419 178 -403 212
rect -309 178 -293 212
rect -241 178 -225 212
rect -131 178 -115 212
rect -63 178 -47 212
rect 47 178 63 212
rect 115 178 131 212
rect 225 178 241 212
rect 293 178 309 212
rect 403 178 419 212
rect 471 178 487 212
rect 581 178 597 212
rect 649 178 665 212
rect 759 178 775 212
rect 827 178 843 212
rect 937 178 953 212
rect 1005 178 1021 212
rect 1115 178 1131 212
rect 1183 178 1199 212
rect 1293 178 1309 212
rect 1361 178 1377 212
rect 1471 178 1487 212
rect 1539 178 1555 212
rect 1649 178 1665 212
rect 1717 178 1733 212
rect 1827 178 1843 212
rect 1895 178 1911 212
rect 2005 178 2021 212
rect 2073 178 2089 212
rect 2183 178 2199 212
rect 2251 178 2267 212
rect 2361 178 2377 212
rect 2429 178 2445 212
rect 2539 178 2555 212
rect 2607 178 2623 212
rect 2717 178 2733 212
rect 2785 178 2801 212
rect 2895 178 2911 212
rect 2963 178 2979 212
rect -3043 128 -3009 144
rect -3043 -144 -3009 -128
rect -2865 128 -2831 144
rect -2865 -144 -2831 -128
rect -2687 128 -2653 144
rect -2687 -144 -2653 -128
rect -2509 128 -2475 144
rect -2509 -144 -2475 -128
rect -2331 128 -2297 144
rect -2331 -144 -2297 -128
rect -2153 128 -2119 144
rect -2153 -144 -2119 -128
rect -1975 128 -1941 144
rect -1975 -144 -1941 -128
rect -1797 128 -1763 144
rect -1797 -144 -1763 -128
rect -1619 128 -1585 144
rect -1619 -144 -1585 -128
rect -1441 128 -1407 144
rect -1441 -144 -1407 -128
rect -1263 128 -1229 144
rect -1263 -144 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 144
rect 1229 -144 1263 -128
rect 1407 128 1441 144
rect 1407 -144 1441 -128
rect 1585 128 1619 144
rect 1585 -144 1619 -128
rect 1763 128 1797 144
rect 1763 -144 1797 -128
rect 1941 128 1975 144
rect 1941 -144 1975 -128
rect 2119 128 2153 144
rect 2119 -144 2153 -128
rect 2297 128 2331 144
rect 2297 -144 2331 -128
rect 2475 128 2509 144
rect 2475 -144 2509 -128
rect 2653 128 2687 144
rect 2653 -144 2687 -128
rect 2831 128 2865 144
rect 2831 -144 2865 -128
rect 3009 128 3043 144
rect 3009 -144 3043 -128
rect -2979 -212 -2963 -178
rect -2911 -212 -2895 -178
rect -2801 -212 -2785 -178
rect -2733 -212 -2717 -178
rect -2623 -212 -2607 -178
rect -2555 -212 -2539 -178
rect -2445 -212 -2429 -178
rect -2377 -212 -2361 -178
rect -2267 -212 -2251 -178
rect -2199 -212 -2183 -178
rect -2089 -212 -2073 -178
rect -2021 -212 -2005 -178
rect -1911 -212 -1895 -178
rect -1843 -212 -1827 -178
rect -1733 -212 -1717 -178
rect -1665 -212 -1649 -178
rect -1555 -212 -1539 -178
rect -1487 -212 -1471 -178
rect -1377 -212 -1361 -178
rect -1309 -212 -1293 -178
rect -1199 -212 -1183 -178
rect -1131 -212 -1115 -178
rect -1021 -212 -1005 -178
rect -953 -212 -937 -178
rect -843 -212 -827 -178
rect -775 -212 -759 -178
rect -665 -212 -649 -178
rect -597 -212 -581 -178
rect -487 -212 -471 -178
rect -419 -212 -403 -178
rect -309 -212 -293 -178
rect -241 -212 -225 -178
rect -131 -212 -115 -178
rect -63 -212 -47 -178
rect 47 -212 63 -178
rect 115 -212 131 -178
rect 225 -212 241 -178
rect 293 -212 309 -178
rect 403 -212 419 -178
rect 471 -212 487 -178
rect 581 -212 597 -178
rect 649 -212 665 -178
rect 759 -212 775 -178
rect 827 -212 843 -178
rect 937 -212 953 -178
rect 1005 -212 1021 -178
rect 1115 -212 1131 -178
rect 1183 -212 1199 -178
rect 1293 -212 1309 -178
rect 1361 -212 1377 -178
rect 1471 -212 1487 -178
rect 1539 -212 1555 -178
rect 1649 -212 1665 -178
rect 1717 -212 1733 -178
rect 1827 -212 1843 -178
rect 1895 -212 1911 -178
rect 2005 -212 2021 -178
rect 2073 -212 2089 -178
rect 2183 -212 2199 -178
rect 2251 -212 2267 -178
rect 2361 -212 2377 -178
rect 2429 -212 2445 -178
rect 2539 -212 2555 -178
rect 2607 -212 2623 -178
rect 2717 -212 2733 -178
rect 2785 -212 2801 -178
rect 2895 -212 2911 -178
rect 2963 -212 2979 -178
<< viali >>
rect -2963 178 -2911 212
rect -2785 178 -2733 212
rect -2607 178 -2555 212
rect -2429 178 -2377 212
rect -2251 178 -2199 212
rect -2073 178 -2021 212
rect -1895 178 -1843 212
rect -1717 178 -1665 212
rect -1539 178 -1487 212
rect -1361 178 -1309 212
rect -1183 178 -1131 212
rect -1005 178 -953 212
rect -827 178 -775 212
rect -649 178 -597 212
rect -471 178 -419 212
rect -293 178 -241 212
rect -115 178 -63 212
rect 63 178 115 212
rect 241 178 293 212
rect 419 178 471 212
rect 597 178 649 212
rect 775 178 827 212
rect 953 178 1005 212
rect 1131 178 1183 212
rect 1309 178 1361 212
rect 1487 178 1539 212
rect 1665 178 1717 212
rect 1843 178 1895 212
rect 2021 178 2073 212
rect 2199 178 2251 212
rect 2377 178 2429 212
rect 2555 178 2607 212
rect 2733 178 2785 212
rect 2911 178 2963 212
rect -2963 -212 -2911 -178
rect -2785 -212 -2733 -178
rect -2607 -212 -2555 -178
rect -2429 -212 -2377 -178
rect -2251 -212 -2199 -178
rect -2073 -212 -2021 -178
rect -1895 -212 -1843 -178
rect -1717 -212 -1665 -178
rect -1539 -212 -1487 -178
rect -1361 -212 -1309 -178
rect -1183 -212 -1131 -178
rect -1005 -212 -953 -178
rect -827 -212 -775 -178
rect -649 -212 -597 -178
rect -471 -212 -419 -178
rect -293 -212 -241 -178
rect -115 -212 -63 -178
rect 63 -212 115 -178
rect 241 -212 293 -178
rect 419 -212 471 -178
rect 597 -212 649 -178
rect 775 -212 827 -178
rect 953 -212 1005 -178
rect 1131 -212 1183 -178
rect 1309 -212 1361 -178
rect 1487 -212 1539 -178
rect 1665 -212 1717 -178
rect 1843 -212 1895 -178
rect 2021 -212 2073 -178
rect 2199 -212 2251 -178
rect 2377 -212 2429 -178
rect 2555 -212 2607 -178
rect 2733 -212 2785 -178
rect 2911 -212 2963 -178
<< metal1 >>
rect -2975 212 -2899 218
rect -2975 178 -2963 212
rect -2911 178 -2899 212
rect -2975 172 -2899 178
rect -2797 212 -2721 218
rect -2797 178 -2785 212
rect -2733 178 -2721 212
rect -2797 172 -2721 178
rect -2619 212 -2543 218
rect -2619 178 -2607 212
rect -2555 178 -2543 212
rect -2619 172 -2543 178
rect -2441 212 -2365 218
rect -2441 178 -2429 212
rect -2377 178 -2365 212
rect -2441 172 -2365 178
rect -2263 212 -2187 218
rect -2263 178 -2251 212
rect -2199 178 -2187 212
rect -2263 172 -2187 178
rect -2085 212 -2009 218
rect -2085 178 -2073 212
rect -2021 178 -2009 212
rect -2085 172 -2009 178
rect -1907 212 -1831 218
rect -1907 178 -1895 212
rect -1843 178 -1831 212
rect -1907 172 -1831 178
rect -1729 212 -1653 218
rect -1729 178 -1717 212
rect -1665 178 -1653 212
rect -1729 172 -1653 178
rect -1551 212 -1475 218
rect -1551 178 -1539 212
rect -1487 178 -1475 212
rect -1551 172 -1475 178
rect -1373 212 -1297 218
rect -1373 178 -1361 212
rect -1309 178 -1297 212
rect -1373 172 -1297 178
rect -1195 212 -1119 218
rect -1195 178 -1183 212
rect -1131 178 -1119 212
rect -1195 172 -1119 178
rect -1017 212 -941 218
rect -1017 178 -1005 212
rect -953 178 -941 212
rect -1017 172 -941 178
rect -839 212 -763 218
rect -839 178 -827 212
rect -775 178 -763 212
rect -839 172 -763 178
rect -661 212 -585 218
rect -661 178 -649 212
rect -597 178 -585 212
rect -661 172 -585 178
rect -483 212 -407 218
rect -483 178 -471 212
rect -419 178 -407 212
rect -483 172 -407 178
rect -305 212 -229 218
rect -305 178 -293 212
rect -241 178 -229 212
rect -305 172 -229 178
rect -127 212 -51 218
rect -127 178 -115 212
rect -63 178 -51 212
rect -127 172 -51 178
rect 51 212 127 218
rect 51 178 63 212
rect 115 178 127 212
rect 51 172 127 178
rect 229 212 305 218
rect 229 178 241 212
rect 293 178 305 212
rect 229 172 305 178
rect 407 212 483 218
rect 407 178 419 212
rect 471 178 483 212
rect 407 172 483 178
rect 585 212 661 218
rect 585 178 597 212
rect 649 178 661 212
rect 585 172 661 178
rect 763 212 839 218
rect 763 178 775 212
rect 827 178 839 212
rect 763 172 839 178
rect 941 212 1017 218
rect 941 178 953 212
rect 1005 178 1017 212
rect 941 172 1017 178
rect 1119 212 1195 218
rect 1119 178 1131 212
rect 1183 178 1195 212
rect 1119 172 1195 178
rect 1297 212 1373 218
rect 1297 178 1309 212
rect 1361 178 1373 212
rect 1297 172 1373 178
rect 1475 212 1551 218
rect 1475 178 1487 212
rect 1539 178 1551 212
rect 1475 172 1551 178
rect 1653 212 1729 218
rect 1653 178 1665 212
rect 1717 178 1729 212
rect 1653 172 1729 178
rect 1831 212 1907 218
rect 1831 178 1843 212
rect 1895 178 1907 212
rect 1831 172 1907 178
rect 2009 212 2085 218
rect 2009 178 2021 212
rect 2073 178 2085 212
rect 2009 172 2085 178
rect 2187 212 2263 218
rect 2187 178 2199 212
rect 2251 178 2263 212
rect 2187 172 2263 178
rect 2365 212 2441 218
rect 2365 178 2377 212
rect 2429 178 2441 212
rect 2365 172 2441 178
rect 2543 212 2619 218
rect 2543 178 2555 212
rect 2607 178 2619 212
rect 2543 172 2619 178
rect 2721 212 2797 218
rect 2721 178 2733 212
rect 2785 178 2797 212
rect 2721 172 2797 178
rect 2899 212 2975 218
rect 2899 178 2911 212
rect 2963 178 2975 212
rect 2899 172 2975 178
rect -2975 -178 -2899 -172
rect -2975 -212 -2963 -178
rect -2911 -212 -2899 -178
rect -2975 -218 -2899 -212
rect -2797 -178 -2721 -172
rect -2797 -212 -2785 -178
rect -2733 -212 -2721 -178
rect -2797 -218 -2721 -212
rect -2619 -178 -2543 -172
rect -2619 -212 -2607 -178
rect -2555 -212 -2543 -178
rect -2619 -218 -2543 -212
rect -2441 -178 -2365 -172
rect -2441 -212 -2429 -178
rect -2377 -212 -2365 -178
rect -2441 -218 -2365 -212
rect -2263 -178 -2187 -172
rect -2263 -212 -2251 -178
rect -2199 -212 -2187 -178
rect -2263 -218 -2187 -212
rect -2085 -178 -2009 -172
rect -2085 -212 -2073 -178
rect -2021 -212 -2009 -178
rect -2085 -218 -2009 -212
rect -1907 -178 -1831 -172
rect -1907 -212 -1895 -178
rect -1843 -212 -1831 -178
rect -1907 -218 -1831 -212
rect -1729 -178 -1653 -172
rect -1729 -212 -1717 -178
rect -1665 -212 -1653 -178
rect -1729 -218 -1653 -212
rect -1551 -178 -1475 -172
rect -1551 -212 -1539 -178
rect -1487 -212 -1475 -178
rect -1551 -218 -1475 -212
rect -1373 -178 -1297 -172
rect -1373 -212 -1361 -178
rect -1309 -212 -1297 -178
rect -1373 -218 -1297 -212
rect -1195 -178 -1119 -172
rect -1195 -212 -1183 -178
rect -1131 -212 -1119 -178
rect -1195 -218 -1119 -212
rect -1017 -178 -941 -172
rect -1017 -212 -1005 -178
rect -953 -212 -941 -178
rect -1017 -218 -941 -212
rect -839 -178 -763 -172
rect -839 -212 -827 -178
rect -775 -212 -763 -178
rect -839 -218 -763 -212
rect -661 -178 -585 -172
rect -661 -212 -649 -178
rect -597 -212 -585 -178
rect -661 -218 -585 -212
rect -483 -178 -407 -172
rect -483 -212 -471 -178
rect -419 -212 -407 -178
rect -483 -218 -407 -212
rect -305 -178 -229 -172
rect -305 -212 -293 -178
rect -241 -212 -229 -178
rect -305 -218 -229 -212
rect -127 -178 -51 -172
rect -127 -212 -115 -178
rect -63 -212 -51 -178
rect -127 -218 -51 -212
rect 51 -178 127 -172
rect 51 -212 63 -178
rect 115 -212 127 -178
rect 51 -218 127 -212
rect 229 -178 305 -172
rect 229 -212 241 -178
rect 293 -212 305 -178
rect 229 -218 305 -212
rect 407 -178 483 -172
rect 407 -212 419 -178
rect 471 -212 483 -178
rect 407 -218 483 -212
rect 585 -178 661 -172
rect 585 -212 597 -178
rect 649 -212 661 -178
rect 585 -218 661 -212
rect 763 -178 839 -172
rect 763 -212 775 -178
rect 827 -212 839 -178
rect 763 -218 839 -212
rect 941 -178 1017 -172
rect 941 -212 953 -178
rect 1005 -212 1017 -178
rect 941 -218 1017 -212
rect 1119 -178 1195 -172
rect 1119 -212 1131 -178
rect 1183 -212 1195 -178
rect 1119 -218 1195 -212
rect 1297 -178 1373 -172
rect 1297 -212 1309 -178
rect 1361 -212 1373 -178
rect 1297 -218 1373 -212
rect 1475 -178 1551 -172
rect 1475 -212 1487 -178
rect 1539 -212 1551 -178
rect 1475 -218 1551 -212
rect 1653 -178 1729 -172
rect 1653 -212 1665 -178
rect 1717 -212 1729 -178
rect 1653 -218 1729 -212
rect 1831 -178 1907 -172
rect 1831 -212 1843 -178
rect 1895 -212 1907 -178
rect 1831 -218 1907 -212
rect 2009 -178 2085 -172
rect 2009 -212 2021 -178
rect 2073 -212 2085 -178
rect 2009 -218 2085 -212
rect 2187 -178 2263 -172
rect 2187 -212 2199 -178
rect 2251 -212 2263 -178
rect 2187 -218 2263 -212
rect 2365 -178 2441 -172
rect 2365 -212 2377 -178
rect 2429 -212 2441 -178
rect 2365 -218 2441 -212
rect 2543 -178 2619 -172
rect 2543 -212 2555 -178
rect 2607 -212 2619 -178
rect 2543 -218 2619 -212
rect 2721 -178 2797 -172
rect 2721 -212 2733 -178
rect 2785 -212 2797 -178
rect 2721 -218 2797 -212
rect 2899 -178 2975 -172
rect 2899 -212 2911 -178
rect 2963 -212 2975 -178
rect 2899 -218 2975 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 34 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
