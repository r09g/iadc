magic
tech sky130A
timestamp 1653386003
<< nmos >>
rect -1765 -70 -1705 70
rect -1676 -70 -1616 70
rect -1587 -70 -1527 70
rect -1498 -70 -1438 70
rect -1409 -70 -1349 70
rect -1320 -70 -1260 70
rect -1231 -70 -1171 70
rect -1142 -70 -1082 70
rect -1053 -70 -993 70
rect -964 -70 -904 70
rect -875 -70 -815 70
rect -786 -70 -726 70
rect -697 -70 -637 70
rect -608 -70 -548 70
rect -519 -70 -459 70
rect -430 -70 -370 70
rect -341 -70 -281 70
rect -252 -70 -192 70
rect -163 -70 -103 70
rect -74 -70 -14 70
rect 14 -70 74 70
rect 103 -70 163 70
rect 192 -70 252 70
rect 281 -70 341 70
rect 370 -70 430 70
rect 459 -70 519 70
rect 548 -70 608 70
rect 637 -70 697 70
rect 726 -70 786 70
rect 815 -70 875 70
rect 904 -70 964 70
rect 993 -70 1053 70
rect 1082 -70 1142 70
rect 1171 -70 1231 70
rect 1260 -70 1320 70
rect 1349 -70 1409 70
rect 1438 -70 1498 70
rect 1527 -70 1587 70
rect 1616 -70 1676 70
rect 1705 -70 1765 70
<< ndiff >>
rect -1794 64 -1765 70
rect -1794 -64 -1788 64
rect -1771 -64 -1765 64
rect -1794 -70 -1765 -64
rect -1705 64 -1676 70
rect -1705 -64 -1699 64
rect -1682 -64 -1676 64
rect -1705 -70 -1676 -64
rect -1616 64 -1587 70
rect -1616 -64 -1610 64
rect -1593 -64 -1587 64
rect -1616 -70 -1587 -64
rect -1527 64 -1498 70
rect -1527 -64 -1521 64
rect -1504 -64 -1498 64
rect -1527 -70 -1498 -64
rect -1438 64 -1409 70
rect -1438 -64 -1432 64
rect -1415 -64 -1409 64
rect -1438 -70 -1409 -64
rect -1349 64 -1320 70
rect -1349 -64 -1343 64
rect -1326 -64 -1320 64
rect -1349 -70 -1320 -64
rect -1260 64 -1231 70
rect -1260 -64 -1254 64
rect -1237 -64 -1231 64
rect -1260 -70 -1231 -64
rect -1171 64 -1142 70
rect -1171 -64 -1165 64
rect -1148 -64 -1142 64
rect -1171 -70 -1142 -64
rect -1082 64 -1053 70
rect -1082 -64 -1076 64
rect -1059 -64 -1053 64
rect -1082 -70 -1053 -64
rect -993 64 -964 70
rect -993 -64 -987 64
rect -970 -64 -964 64
rect -993 -70 -964 -64
rect -904 64 -875 70
rect -904 -64 -898 64
rect -881 -64 -875 64
rect -904 -70 -875 -64
rect -815 64 -786 70
rect -815 -64 -809 64
rect -792 -64 -786 64
rect -815 -70 -786 -64
rect -726 64 -697 70
rect -726 -64 -720 64
rect -703 -64 -697 64
rect -726 -70 -697 -64
rect -637 64 -608 70
rect -637 -64 -631 64
rect -614 -64 -608 64
rect -637 -70 -608 -64
rect -548 64 -519 70
rect -548 -64 -542 64
rect -525 -64 -519 64
rect -548 -70 -519 -64
rect -459 64 -430 70
rect -459 -64 -453 64
rect -436 -64 -430 64
rect -459 -70 -430 -64
rect -370 64 -341 70
rect -370 -64 -364 64
rect -347 -64 -341 64
rect -370 -70 -341 -64
rect -281 64 -252 70
rect -281 -64 -275 64
rect -258 -64 -252 64
rect -281 -70 -252 -64
rect -192 64 -163 70
rect -192 -64 -186 64
rect -169 -64 -163 64
rect -192 -70 -163 -64
rect -103 64 -74 70
rect -103 -64 -97 64
rect -80 -64 -74 64
rect -103 -70 -74 -64
rect -14 64 14 70
rect -14 -64 -8 64
rect 8 -64 14 64
rect -14 -70 14 -64
rect 74 64 103 70
rect 74 -64 80 64
rect 97 -64 103 64
rect 74 -70 103 -64
rect 163 64 192 70
rect 163 -64 169 64
rect 186 -64 192 64
rect 163 -70 192 -64
rect 252 64 281 70
rect 252 -64 258 64
rect 275 -64 281 64
rect 252 -70 281 -64
rect 341 64 370 70
rect 341 -64 347 64
rect 364 -64 370 64
rect 341 -70 370 -64
rect 430 64 459 70
rect 430 -64 436 64
rect 453 -64 459 64
rect 430 -70 459 -64
rect 519 64 548 70
rect 519 -64 525 64
rect 542 -64 548 64
rect 519 -70 548 -64
rect 608 64 637 70
rect 608 -64 614 64
rect 631 -64 637 64
rect 608 -70 637 -64
rect 697 64 726 70
rect 697 -64 703 64
rect 720 -64 726 64
rect 697 -70 726 -64
rect 786 64 815 70
rect 786 -64 792 64
rect 809 -64 815 64
rect 786 -70 815 -64
rect 875 64 904 70
rect 875 -64 881 64
rect 898 -64 904 64
rect 875 -70 904 -64
rect 964 64 993 70
rect 964 -64 970 64
rect 987 -64 993 64
rect 964 -70 993 -64
rect 1053 64 1082 70
rect 1053 -64 1059 64
rect 1076 -64 1082 64
rect 1053 -70 1082 -64
rect 1142 64 1171 70
rect 1142 -64 1148 64
rect 1165 -64 1171 64
rect 1142 -70 1171 -64
rect 1231 64 1260 70
rect 1231 -64 1237 64
rect 1254 -64 1260 64
rect 1231 -70 1260 -64
rect 1320 64 1349 70
rect 1320 -64 1326 64
rect 1343 -64 1349 64
rect 1320 -70 1349 -64
rect 1409 64 1438 70
rect 1409 -64 1415 64
rect 1432 -64 1438 64
rect 1409 -70 1438 -64
rect 1498 64 1527 70
rect 1498 -64 1504 64
rect 1521 -64 1527 64
rect 1498 -70 1527 -64
rect 1587 64 1616 70
rect 1587 -64 1593 64
rect 1610 -64 1616 64
rect 1587 -70 1616 -64
rect 1676 64 1705 70
rect 1676 -64 1682 64
rect 1699 -64 1705 64
rect 1676 -70 1705 -64
rect 1765 64 1794 70
rect 1765 -64 1771 64
rect 1788 -64 1794 64
rect 1765 -70 1794 -64
<< ndiffc >>
rect -1788 -64 -1771 64
rect -1699 -64 -1682 64
rect -1610 -64 -1593 64
rect -1521 -64 -1504 64
rect -1432 -64 -1415 64
rect -1343 -64 -1326 64
rect -1254 -64 -1237 64
rect -1165 -64 -1148 64
rect -1076 -64 -1059 64
rect -987 -64 -970 64
rect -898 -64 -881 64
rect -809 -64 -792 64
rect -720 -64 -703 64
rect -631 -64 -614 64
rect -542 -64 -525 64
rect -453 -64 -436 64
rect -364 -64 -347 64
rect -275 -64 -258 64
rect -186 -64 -169 64
rect -97 -64 -80 64
rect -8 -64 8 64
rect 80 -64 97 64
rect 169 -64 186 64
rect 258 -64 275 64
rect 347 -64 364 64
rect 436 -64 453 64
rect 525 -64 542 64
rect 614 -64 631 64
rect 703 -64 720 64
rect 792 -64 809 64
rect 881 -64 898 64
rect 970 -64 987 64
rect 1059 -64 1076 64
rect 1148 -64 1165 64
rect 1237 -64 1254 64
rect 1326 -64 1343 64
rect 1415 -64 1432 64
rect 1504 -64 1521 64
rect 1593 -64 1610 64
rect 1682 -64 1699 64
rect 1771 -64 1788 64
<< poly >>
rect -1754 106 -1716 114
rect -1754 97 -1746 106
rect -1765 89 -1746 97
rect -1724 97 -1716 106
rect -1665 106 -1627 114
rect -1665 97 -1657 106
rect -1724 89 -1705 97
rect -1765 70 -1705 89
rect -1676 89 -1657 97
rect -1635 97 -1627 106
rect -1576 106 -1538 114
rect -1576 97 -1568 106
rect -1635 89 -1616 97
rect -1676 70 -1616 89
rect -1587 89 -1568 97
rect -1546 97 -1538 106
rect -1487 106 -1449 114
rect -1487 97 -1479 106
rect -1546 89 -1527 97
rect -1587 70 -1527 89
rect -1498 89 -1479 97
rect -1457 97 -1449 106
rect -1398 106 -1360 114
rect -1398 97 -1390 106
rect -1457 89 -1438 97
rect -1498 70 -1438 89
rect -1409 89 -1390 97
rect -1368 97 -1360 106
rect -1309 106 -1271 114
rect -1309 97 -1301 106
rect -1368 89 -1349 97
rect -1409 70 -1349 89
rect -1320 89 -1301 97
rect -1279 97 -1271 106
rect -1220 106 -1182 114
rect -1220 97 -1212 106
rect -1279 89 -1260 97
rect -1320 70 -1260 89
rect -1231 89 -1212 97
rect -1190 97 -1182 106
rect -1131 106 -1093 114
rect -1131 97 -1123 106
rect -1190 89 -1171 97
rect -1231 70 -1171 89
rect -1142 89 -1123 97
rect -1101 97 -1093 106
rect -1042 106 -1004 114
rect -1042 97 -1034 106
rect -1101 89 -1082 97
rect -1142 70 -1082 89
rect -1053 89 -1034 97
rect -1012 97 -1004 106
rect -953 106 -915 114
rect -953 97 -945 106
rect -1012 89 -993 97
rect -1053 70 -993 89
rect -964 89 -945 97
rect -923 97 -915 106
rect -864 106 -826 114
rect -864 97 -856 106
rect -923 89 -904 97
rect -964 70 -904 89
rect -875 89 -856 97
rect -834 97 -826 106
rect -775 106 -737 114
rect -775 97 -767 106
rect -834 89 -815 97
rect -875 70 -815 89
rect -786 89 -767 97
rect -745 97 -737 106
rect -686 106 -648 114
rect -686 97 -678 106
rect -745 89 -726 97
rect -786 70 -726 89
rect -697 89 -678 97
rect -656 97 -648 106
rect -597 106 -559 114
rect -597 97 -589 106
rect -656 89 -637 97
rect -697 70 -637 89
rect -608 89 -589 97
rect -567 97 -559 106
rect -508 106 -470 114
rect -508 97 -500 106
rect -567 89 -548 97
rect -608 70 -548 89
rect -519 89 -500 97
rect -478 97 -470 106
rect -419 106 -381 114
rect -419 97 -411 106
rect -478 89 -459 97
rect -519 70 -459 89
rect -430 89 -411 97
rect -389 97 -381 106
rect -330 106 -292 114
rect -330 97 -322 106
rect -389 89 -370 97
rect -430 70 -370 89
rect -341 89 -322 97
rect -300 97 -292 106
rect -241 106 -203 114
rect -241 97 -233 106
rect -300 89 -281 97
rect -341 70 -281 89
rect -252 89 -233 97
rect -211 97 -203 106
rect -152 106 -114 114
rect -152 97 -144 106
rect -211 89 -192 97
rect -252 70 -192 89
rect -163 89 -144 97
rect -122 97 -114 106
rect -63 106 -25 114
rect -63 97 -55 106
rect -122 89 -103 97
rect -163 70 -103 89
rect -74 89 -55 97
rect -33 97 -25 106
rect 25 106 63 114
rect 25 97 33 106
rect -33 89 -14 97
rect -74 70 -14 89
rect 14 89 33 97
rect 55 97 63 106
rect 114 106 152 114
rect 114 97 122 106
rect 55 89 74 97
rect 14 70 74 89
rect 103 89 122 97
rect 144 97 152 106
rect 203 106 241 114
rect 203 97 211 106
rect 144 89 163 97
rect 103 70 163 89
rect 192 89 211 97
rect 233 97 241 106
rect 292 106 330 114
rect 292 97 300 106
rect 233 89 252 97
rect 192 70 252 89
rect 281 89 300 97
rect 322 97 330 106
rect 381 106 419 114
rect 381 97 389 106
rect 322 89 341 97
rect 281 70 341 89
rect 370 89 389 97
rect 411 97 419 106
rect 470 106 508 114
rect 470 97 478 106
rect 411 89 430 97
rect 370 70 430 89
rect 459 89 478 97
rect 500 97 508 106
rect 559 106 597 114
rect 559 97 567 106
rect 500 89 519 97
rect 459 70 519 89
rect 548 89 567 97
rect 589 97 597 106
rect 648 106 686 114
rect 648 97 656 106
rect 589 89 608 97
rect 548 70 608 89
rect 637 89 656 97
rect 678 97 686 106
rect 737 106 775 114
rect 737 97 745 106
rect 678 89 697 97
rect 637 70 697 89
rect 726 89 745 97
rect 767 97 775 106
rect 826 106 864 114
rect 826 97 834 106
rect 767 89 786 97
rect 726 70 786 89
rect 815 89 834 97
rect 856 97 864 106
rect 915 106 953 114
rect 915 97 923 106
rect 856 89 875 97
rect 815 70 875 89
rect 904 89 923 97
rect 945 97 953 106
rect 1004 106 1042 114
rect 1004 97 1012 106
rect 945 89 964 97
rect 904 70 964 89
rect 993 89 1012 97
rect 1034 97 1042 106
rect 1093 106 1131 114
rect 1093 97 1101 106
rect 1034 89 1053 97
rect 993 70 1053 89
rect 1082 89 1101 97
rect 1123 97 1131 106
rect 1182 106 1220 114
rect 1182 97 1190 106
rect 1123 89 1142 97
rect 1082 70 1142 89
rect 1171 89 1190 97
rect 1212 97 1220 106
rect 1271 106 1309 114
rect 1271 97 1279 106
rect 1212 89 1231 97
rect 1171 70 1231 89
rect 1260 89 1279 97
rect 1301 97 1309 106
rect 1360 106 1398 114
rect 1360 97 1368 106
rect 1301 89 1320 97
rect 1260 70 1320 89
rect 1349 89 1368 97
rect 1390 97 1398 106
rect 1449 106 1487 114
rect 1449 97 1457 106
rect 1390 89 1409 97
rect 1349 70 1409 89
rect 1438 89 1457 97
rect 1479 97 1487 106
rect 1538 106 1576 114
rect 1538 97 1546 106
rect 1479 89 1498 97
rect 1438 70 1498 89
rect 1527 89 1546 97
rect 1568 97 1576 106
rect 1627 106 1665 114
rect 1627 97 1635 106
rect 1568 89 1587 97
rect 1527 70 1587 89
rect 1616 89 1635 97
rect 1657 97 1665 106
rect 1716 106 1754 114
rect 1716 97 1724 106
rect 1657 89 1676 97
rect 1616 70 1676 89
rect 1705 89 1724 97
rect 1746 97 1754 106
rect 1746 89 1765 97
rect 1705 70 1765 89
rect -1765 -89 -1705 -70
rect -1765 -97 -1746 -89
rect -1754 -106 -1746 -97
rect -1724 -97 -1705 -89
rect -1676 -89 -1616 -70
rect -1676 -97 -1657 -89
rect -1724 -106 -1716 -97
rect -1754 -114 -1716 -106
rect -1665 -106 -1657 -97
rect -1635 -97 -1616 -89
rect -1587 -89 -1527 -70
rect -1587 -97 -1568 -89
rect -1635 -106 -1627 -97
rect -1665 -114 -1627 -106
rect -1576 -106 -1568 -97
rect -1546 -97 -1527 -89
rect -1498 -89 -1438 -70
rect -1498 -97 -1479 -89
rect -1546 -106 -1538 -97
rect -1576 -114 -1538 -106
rect -1487 -106 -1479 -97
rect -1457 -97 -1438 -89
rect -1409 -89 -1349 -70
rect -1409 -97 -1390 -89
rect -1457 -106 -1449 -97
rect -1487 -114 -1449 -106
rect -1398 -106 -1390 -97
rect -1368 -97 -1349 -89
rect -1320 -89 -1260 -70
rect -1320 -97 -1301 -89
rect -1368 -106 -1360 -97
rect -1398 -114 -1360 -106
rect -1309 -106 -1301 -97
rect -1279 -97 -1260 -89
rect -1231 -89 -1171 -70
rect -1231 -97 -1212 -89
rect -1279 -106 -1271 -97
rect -1309 -114 -1271 -106
rect -1220 -106 -1212 -97
rect -1190 -97 -1171 -89
rect -1142 -89 -1082 -70
rect -1142 -97 -1123 -89
rect -1190 -106 -1182 -97
rect -1220 -114 -1182 -106
rect -1131 -106 -1123 -97
rect -1101 -97 -1082 -89
rect -1053 -89 -993 -70
rect -1053 -97 -1034 -89
rect -1101 -106 -1093 -97
rect -1131 -114 -1093 -106
rect -1042 -106 -1034 -97
rect -1012 -97 -993 -89
rect -964 -89 -904 -70
rect -964 -97 -945 -89
rect -1012 -106 -1004 -97
rect -1042 -114 -1004 -106
rect -953 -106 -945 -97
rect -923 -97 -904 -89
rect -875 -89 -815 -70
rect -875 -97 -856 -89
rect -923 -106 -915 -97
rect -953 -114 -915 -106
rect -864 -106 -856 -97
rect -834 -97 -815 -89
rect -786 -89 -726 -70
rect -786 -97 -767 -89
rect -834 -106 -826 -97
rect -864 -114 -826 -106
rect -775 -106 -767 -97
rect -745 -97 -726 -89
rect -697 -89 -637 -70
rect -697 -97 -678 -89
rect -745 -106 -737 -97
rect -775 -114 -737 -106
rect -686 -106 -678 -97
rect -656 -97 -637 -89
rect -608 -89 -548 -70
rect -608 -97 -589 -89
rect -656 -106 -648 -97
rect -686 -114 -648 -106
rect -597 -106 -589 -97
rect -567 -97 -548 -89
rect -519 -89 -459 -70
rect -519 -97 -500 -89
rect -567 -106 -559 -97
rect -597 -114 -559 -106
rect -508 -106 -500 -97
rect -478 -97 -459 -89
rect -430 -89 -370 -70
rect -430 -97 -411 -89
rect -478 -106 -470 -97
rect -508 -114 -470 -106
rect -419 -106 -411 -97
rect -389 -97 -370 -89
rect -341 -89 -281 -70
rect -341 -97 -322 -89
rect -389 -106 -381 -97
rect -419 -114 -381 -106
rect -330 -106 -322 -97
rect -300 -97 -281 -89
rect -252 -89 -192 -70
rect -252 -97 -233 -89
rect -300 -106 -292 -97
rect -330 -114 -292 -106
rect -241 -106 -233 -97
rect -211 -97 -192 -89
rect -163 -89 -103 -70
rect -163 -97 -144 -89
rect -211 -106 -203 -97
rect -241 -114 -203 -106
rect -152 -106 -144 -97
rect -122 -97 -103 -89
rect -74 -89 -14 -70
rect -74 -97 -55 -89
rect -122 -106 -114 -97
rect -152 -114 -114 -106
rect -63 -106 -55 -97
rect -33 -97 -14 -89
rect 14 -89 74 -70
rect 14 -97 33 -89
rect -33 -106 -25 -97
rect -63 -114 -25 -106
rect 25 -106 33 -97
rect 55 -97 74 -89
rect 103 -89 163 -70
rect 103 -97 122 -89
rect 55 -106 63 -97
rect 25 -114 63 -106
rect 114 -106 122 -97
rect 144 -97 163 -89
rect 192 -89 252 -70
rect 192 -97 211 -89
rect 144 -106 152 -97
rect 114 -114 152 -106
rect 203 -106 211 -97
rect 233 -97 252 -89
rect 281 -89 341 -70
rect 281 -97 300 -89
rect 233 -106 241 -97
rect 203 -114 241 -106
rect 292 -106 300 -97
rect 322 -97 341 -89
rect 370 -89 430 -70
rect 370 -97 389 -89
rect 322 -106 330 -97
rect 292 -114 330 -106
rect 381 -106 389 -97
rect 411 -97 430 -89
rect 459 -89 519 -70
rect 459 -97 478 -89
rect 411 -106 419 -97
rect 381 -114 419 -106
rect 470 -106 478 -97
rect 500 -97 519 -89
rect 548 -89 608 -70
rect 548 -97 567 -89
rect 500 -106 508 -97
rect 470 -114 508 -106
rect 559 -106 567 -97
rect 589 -97 608 -89
rect 637 -89 697 -70
rect 637 -97 656 -89
rect 589 -106 597 -97
rect 559 -114 597 -106
rect 648 -106 656 -97
rect 678 -97 697 -89
rect 726 -89 786 -70
rect 726 -97 745 -89
rect 678 -106 686 -97
rect 648 -114 686 -106
rect 737 -106 745 -97
rect 767 -97 786 -89
rect 815 -89 875 -70
rect 815 -97 834 -89
rect 767 -106 775 -97
rect 737 -114 775 -106
rect 826 -106 834 -97
rect 856 -97 875 -89
rect 904 -89 964 -70
rect 904 -97 923 -89
rect 856 -106 864 -97
rect 826 -114 864 -106
rect 915 -106 923 -97
rect 945 -97 964 -89
rect 993 -89 1053 -70
rect 993 -97 1012 -89
rect 945 -106 953 -97
rect 915 -114 953 -106
rect 1004 -106 1012 -97
rect 1034 -97 1053 -89
rect 1082 -89 1142 -70
rect 1082 -97 1101 -89
rect 1034 -106 1042 -97
rect 1004 -114 1042 -106
rect 1093 -106 1101 -97
rect 1123 -97 1142 -89
rect 1171 -89 1231 -70
rect 1171 -97 1190 -89
rect 1123 -106 1131 -97
rect 1093 -114 1131 -106
rect 1182 -106 1190 -97
rect 1212 -97 1231 -89
rect 1260 -89 1320 -70
rect 1260 -97 1279 -89
rect 1212 -106 1220 -97
rect 1182 -114 1220 -106
rect 1271 -106 1279 -97
rect 1301 -97 1320 -89
rect 1349 -89 1409 -70
rect 1349 -97 1368 -89
rect 1301 -106 1309 -97
rect 1271 -114 1309 -106
rect 1360 -106 1368 -97
rect 1390 -97 1409 -89
rect 1438 -89 1498 -70
rect 1438 -97 1457 -89
rect 1390 -106 1398 -97
rect 1360 -114 1398 -106
rect 1449 -106 1457 -97
rect 1479 -97 1498 -89
rect 1527 -89 1587 -70
rect 1527 -97 1546 -89
rect 1479 -106 1487 -97
rect 1449 -114 1487 -106
rect 1538 -106 1546 -97
rect 1568 -97 1587 -89
rect 1616 -89 1676 -70
rect 1616 -97 1635 -89
rect 1568 -106 1576 -97
rect 1538 -114 1576 -106
rect 1627 -106 1635 -97
rect 1657 -97 1676 -89
rect 1705 -89 1765 -70
rect 1705 -97 1724 -89
rect 1657 -106 1665 -97
rect 1627 -114 1665 -106
rect 1716 -106 1724 -97
rect 1746 -97 1765 -89
rect 1746 -106 1754 -97
rect 1716 -114 1754 -106
<< polycont >>
rect -1746 89 -1724 106
rect -1657 89 -1635 106
rect -1568 89 -1546 106
rect -1479 89 -1457 106
rect -1390 89 -1368 106
rect -1301 89 -1279 106
rect -1212 89 -1190 106
rect -1123 89 -1101 106
rect -1034 89 -1012 106
rect -945 89 -923 106
rect -856 89 -834 106
rect -767 89 -745 106
rect -678 89 -656 106
rect -589 89 -567 106
rect -500 89 -478 106
rect -411 89 -389 106
rect -322 89 -300 106
rect -233 89 -211 106
rect -144 89 -122 106
rect -55 89 -33 106
rect 33 89 55 106
rect 122 89 144 106
rect 211 89 233 106
rect 300 89 322 106
rect 389 89 411 106
rect 478 89 500 106
rect 567 89 589 106
rect 656 89 678 106
rect 745 89 767 106
rect 834 89 856 106
rect 923 89 945 106
rect 1012 89 1034 106
rect 1101 89 1123 106
rect 1190 89 1212 106
rect 1279 89 1301 106
rect 1368 89 1390 106
rect 1457 89 1479 106
rect 1546 89 1568 106
rect 1635 89 1657 106
rect 1724 89 1746 106
rect -1746 -106 -1724 -89
rect -1657 -106 -1635 -89
rect -1568 -106 -1546 -89
rect -1479 -106 -1457 -89
rect -1390 -106 -1368 -89
rect -1301 -106 -1279 -89
rect -1212 -106 -1190 -89
rect -1123 -106 -1101 -89
rect -1034 -106 -1012 -89
rect -945 -106 -923 -89
rect -856 -106 -834 -89
rect -767 -106 -745 -89
rect -678 -106 -656 -89
rect -589 -106 -567 -89
rect -500 -106 -478 -89
rect -411 -106 -389 -89
rect -322 -106 -300 -89
rect -233 -106 -211 -89
rect -144 -106 -122 -89
rect -55 -106 -33 -89
rect 33 -106 55 -89
rect 122 -106 144 -89
rect 211 -106 233 -89
rect 300 -106 322 -89
rect 389 -106 411 -89
rect 478 -106 500 -89
rect 567 -106 589 -89
rect 656 -106 678 -89
rect 745 -106 767 -89
rect 834 -106 856 -89
rect 923 -106 945 -89
rect 1012 -106 1034 -89
rect 1101 -106 1123 -89
rect 1190 -106 1212 -89
rect 1279 -106 1301 -89
rect 1368 -106 1390 -89
rect 1457 -106 1479 -89
rect 1546 -106 1568 -89
rect 1635 -106 1657 -89
rect 1724 -106 1746 -89
<< locali >>
rect -1754 89 -1746 106
rect -1724 89 -1716 106
rect -1665 89 -1657 106
rect -1635 89 -1627 106
rect -1576 89 -1568 106
rect -1546 89 -1538 106
rect -1487 89 -1479 106
rect -1457 89 -1449 106
rect -1398 89 -1390 106
rect -1368 89 -1360 106
rect -1309 89 -1301 106
rect -1279 89 -1271 106
rect -1220 89 -1212 106
rect -1190 89 -1182 106
rect -1131 89 -1123 106
rect -1101 89 -1093 106
rect -1042 89 -1034 106
rect -1012 89 -1004 106
rect -953 89 -945 106
rect -923 89 -915 106
rect -864 89 -856 106
rect -834 89 -826 106
rect -775 89 -767 106
rect -745 89 -737 106
rect -686 89 -678 106
rect -656 89 -648 106
rect -597 89 -589 106
rect -567 89 -559 106
rect -508 89 -500 106
rect -478 89 -470 106
rect -419 89 -411 106
rect -389 89 -381 106
rect -330 89 -322 106
rect -300 89 -292 106
rect -241 89 -233 106
rect -211 89 -203 106
rect -152 89 -144 106
rect -122 89 -114 106
rect -63 89 -55 106
rect -33 89 -25 106
rect 25 89 33 106
rect 55 89 63 106
rect 114 89 122 106
rect 144 89 152 106
rect 203 89 211 106
rect 233 89 241 106
rect 292 89 300 106
rect 322 89 330 106
rect 381 89 389 106
rect 411 89 419 106
rect 470 89 478 106
rect 500 89 508 106
rect 559 89 567 106
rect 589 89 597 106
rect 648 89 656 106
rect 678 89 686 106
rect 737 89 745 106
rect 767 89 775 106
rect 826 89 834 106
rect 856 89 864 106
rect 915 89 923 106
rect 945 89 953 106
rect 1004 89 1012 106
rect 1034 89 1042 106
rect 1093 89 1101 106
rect 1123 89 1131 106
rect 1182 89 1190 106
rect 1212 89 1220 106
rect 1271 89 1279 106
rect 1301 89 1309 106
rect 1360 89 1368 106
rect 1390 89 1398 106
rect 1449 89 1457 106
rect 1479 89 1487 106
rect 1538 89 1546 106
rect 1568 89 1576 106
rect 1627 89 1635 106
rect 1657 89 1665 106
rect 1716 89 1724 106
rect 1746 89 1754 106
rect -1788 64 -1771 72
rect -1788 -72 -1771 -64
rect -1699 64 -1682 72
rect -1699 -72 -1682 -64
rect -1610 64 -1593 72
rect -1610 -72 -1593 -64
rect -1521 64 -1504 72
rect -1521 -72 -1504 -64
rect -1432 64 -1415 72
rect -1432 -72 -1415 -64
rect -1343 64 -1326 72
rect -1343 -72 -1326 -64
rect -1254 64 -1237 72
rect -1254 -72 -1237 -64
rect -1165 64 -1148 72
rect -1165 -72 -1148 -64
rect -1076 64 -1059 72
rect -1076 -72 -1059 -64
rect -987 64 -970 72
rect -987 -72 -970 -64
rect -898 64 -881 72
rect -898 -72 -881 -64
rect -809 64 -792 72
rect -809 -72 -792 -64
rect -720 64 -703 72
rect -720 -72 -703 -64
rect -631 64 -614 72
rect -631 -72 -614 -64
rect -542 64 -525 72
rect -542 -72 -525 -64
rect -453 64 -436 72
rect -453 -72 -436 -64
rect -364 64 -347 72
rect -364 -72 -347 -64
rect -275 64 -258 72
rect -275 -72 -258 -64
rect -186 64 -169 72
rect -186 -72 -169 -64
rect -97 64 -80 72
rect -97 -72 -80 -64
rect -8 64 8 72
rect -8 -72 8 -64
rect 80 64 97 72
rect 80 -72 97 -64
rect 169 64 186 72
rect 169 -72 186 -64
rect 258 64 275 72
rect 258 -72 275 -64
rect 347 64 364 72
rect 347 -72 364 -64
rect 436 64 453 72
rect 436 -72 453 -64
rect 525 64 542 72
rect 525 -72 542 -64
rect 614 64 631 72
rect 614 -72 631 -64
rect 703 64 720 72
rect 703 -72 720 -64
rect 792 64 809 72
rect 792 -72 809 -64
rect 881 64 898 72
rect 881 -72 898 -64
rect 970 64 987 72
rect 970 -72 987 -64
rect 1059 64 1076 72
rect 1059 -72 1076 -64
rect 1148 64 1165 72
rect 1148 -72 1165 -64
rect 1237 64 1254 72
rect 1237 -72 1254 -64
rect 1326 64 1343 72
rect 1326 -72 1343 -64
rect 1415 64 1432 72
rect 1415 -72 1432 -64
rect 1504 64 1521 72
rect 1504 -72 1521 -64
rect 1593 64 1610 72
rect 1593 -72 1610 -64
rect 1682 64 1699 72
rect 1682 -72 1699 -64
rect 1771 64 1788 72
rect 1771 -72 1788 -64
rect -1754 -106 -1746 -89
rect -1724 -106 -1716 -89
rect -1665 -106 -1657 -89
rect -1635 -106 -1627 -89
rect -1576 -106 -1568 -89
rect -1546 -106 -1538 -89
rect -1487 -106 -1479 -89
rect -1457 -106 -1449 -89
rect -1398 -106 -1390 -89
rect -1368 -106 -1360 -89
rect -1309 -106 -1301 -89
rect -1279 -106 -1271 -89
rect -1220 -106 -1212 -89
rect -1190 -106 -1182 -89
rect -1131 -106 -1123 -89
rect -1101 -106 -1093 -89
rect -1042 -106 -1034 -89
rect -1012 -106 -1004 -89
rect -953 -106 -945 -89
rect -923 -106 -915 -89
rect -864 -106 -856 -89
rect -834 -106 -826 -89
rect -775 -106 -767 -89
rect -745 -106 -737 -89
rect -686 -106 -678 -89
rect -656 -106 -648 -89
rect -597 -106 -589 -89
rect -567 -106 -559 -89
rect -508 -106 -500 -89
rect -478 -106 -470 -89
rect -419 -106 -411 -89
rect -389 -106 -381 -89
rect -330 -106 -322 -89
rect -300 -106 -292 -89
rect -241 -106 -233 -89
rect -211 -106 -203 -89
rect -152 -106 -144 -89
rect -122 -106 -114 -89
rect -63 -106 -55 -89
rect -33 -106 -25 -89
rect 25 -106 33 -89
rect 55 -106 63 -89
rect 114 -106 122 -89
rect 144 -106 152 -89
rect 203 -106 211 -89
rect 233 -106 241 -89
rect 292 -106 300 -89
rect 322 -106 330 -89
rect 381 -106 389 -89
rect 411 -106 419 -89
rect 470 -106 478 -89
rect 500 -106 508 -89
rect 559 -106 567 -89
rect 589 -106 597 -89
rect 648 -106 656 -89
rect 678 -106 686 -89
rect 737 -106 745 -89
rect 767 -106 775 -89
rect 826 -106 834 -89
rect 856 -106 864 -89
rect 915 -106 923 -89
rect 945 -106 953 -89
rect 1004 -106 1012 -89
rect 1034 -106 1042 -89
rect 1093 -106 1101 -89
rect 1123 -106 1131 -89
rect 1182 -106 1190 -89
rect 1212 -106 1220 -89
rect 1271 -106 1279 -89
rect 1301 -106 1309 -89
rect 1360 -106 1368 -89
rect 1390 -106 1398 -89
rect 1449 -106 1457 -89
rect 1479 -106 1487 -89
rect 1538 -106 1546 -89
rect 1568 -106 1576 -89
rect 1627 -106 1635 -89
rect 1657 -106 1665 -89
rect 1716 -106 1724 -89
rect 1746 -106 1754 -89
<< viali >>
rect -1746 89 -1724 106
rect -1657 89 -1635 106
rect -1568 89 -1546 106
rect -1479 89 -1457 106
rect -1390 89 -1368 106
rect -1301 89 -1279 106
rect -1212 89 -1190 106
rect -1123 89 -1101 106
rect -1034 89 -1012 106
rect -945 89 -923 106
rect -856 89 -834 106
rect -767 89 -745 106
rect -678 89 -656 106
rect -589 89 -567 106
rect -500 89 -478 106
rect -411 89 -389 106
rect -322 89 -300 106
rect -233 89 -211 106
rect -144 89 -122 106
rect -55 89 -33 106
rect 33 89 55 106
rect 122 89 144 106
rect 211 89 233 106
rect 300 89 322 106
rect 389 89 411 106
rect 478 89 500 106
rect 567 89 589 106
rect 656 89 678 106
rect 745 89 767 106
rect 834 89 856 106
rect 923 89 945 106
rect 1012 89 1034 106
rect 1101 89 1123 106
rect 1190 89 1212 106
rect 1279 89 1301 106
rect 1368 89 1390 106
rect 1457 89 1479 106
rect 1546 89 1568 106
rect 1635 89 1657 106
rect 1724 89 1746 106
rect -1788 -64 -1771 64
rect -1699 -64 -1682 64
rect -1610 -64 -1593 64
rect -1521 -64 -1504 64
rect -1432 -64 -1415 64
rect -1343 -64 -1326 64
rect -1254 -64 -1237 64
rect -1165 -64 -1148 64
rect -1076 -64 -1059 64
rect -987 -64 -970 64
rect -898 -64 -881 64
rect -809 -64 -792 64
rect -720 -64 -703 64
rect -631 -64 -614 64
rect -542 -64 -525 64
rect -453 -64 -436 64
rect -364 -64 -347 64
rect -275 -64 -258 64
rect -186 -64 -169 64
rect -97 -64 -80 64
rect -8 -64 8 64
rect 80 -64 97 64
rect 169 -64 186 64
rect 258 -64 275 64
rect 347 -64 364 64
rect 436 -64 453 64
rect 525 -64 542 64
rect 614 -64 631 64
rect 703 -64 720 64
rect 792 -64 809 64
rect 881 -64 898 64
rect 970 -64 987 64
rect 1059 -64 1076 64
rect 1148 -64 1165 64
rect 1237 -64 1254 64
rect 1326 -64 1343 64
rect 1415 -64 1432 64
rect 1504 -64 1521 64
rect 1593 -64 1610 64
rect 1682 -64 1699 64
rect 1771 -64 1788 64
rect -1746 -106 -1724 -89
rect -1657 -106 -1635 -89
rect -1568 -106 -1546 -89
rect -1479 -106 -1457 -89
rect -1390 -106 -1368 -89
rect -1301 -106 -1279 -89
rect -1212 -106 -1190 -89
rect -1123 -106 -1101 -89
rect -1034 -106 -1012 -89
rect -945 -106 -923 -89
rect -856 -106 -834 -89
rect -767 -106 -745 -89
rect -678 -106 -656 -89
rect -589 -106 -567 -89
rect -500 -106 -478 -89
rect -411 -106 -389 -89
rect -322 -106 -300 -89
rect -233 -106 -211 -89
rect -144 -106 -122 -89
rect -55 -106 -33 -89
rect 33 -106 55 -89
rect 122 -106 144 -89
rect 211 -106 233 -89
rect 300 -106 322 -89
rect 389 -106 411 -89
rect 478 -106 500 -89
rect 567 -106 589 -89
rect 656 -106 678 -89
rect 745 -106 767 -89
rect 834 -106 856 -89
rect 923 -106 945 -89
rect 1012 -106 1034 -89
rect 1101 -106 1123 -89
rect 1190 -106 1212 -89
rect 1279 -106 1301 -89
rect 1368 -106 1390 -89
rect 1457 -106 1479 -89
rect 1546 -106 1568 -89
rect 1635 -106 1657 -89
rect 1724 -106 1746 -89
<< metal1 >>
rect -1754 106 -1716 114
rect -1754 89 -1746 106
rect -1724 89 -1716 106
rect -1754 86 -1716 89
rect -1665 106 -1627 114
rect -1665 89 -1657 106
rect -1635 89 -1627 106
rect -1665 86 -1627 89
rect -1576 106 -1538 114
rect -1576 89 -1568 106
rect -1546 89 -1538 106
rect -1576 86 -1538 89
rect -1487 106 -1449 114
rect -1487 89 -1479 106
rect -1457 89 -1449 106
rect -1487 86 -1449 89
rect -1398 106 -1360 114
rect -1398 89 -1390 106
rect -1368 89 -1360 106
rect -1398 86 -1360 89
rect -1309 106 -1271 114
rect -1309 89 -1301 106
rect -1279 89 -1271 106
rect -1309 86 -1271 89
rect -1220 106 -1182 114
rect -1220 89 -1212 106
rect -1190 89 -1182 106
rect -1220 86 -1182 89
rect -1131 106 -1093 114
rect -1131 89 -1123 106
rect -1101 89 -1093 106
rect -1131 86 -1093 89
rect -1042 106 -1004 114
rect -1042 89 -1034 106
rect -1012 89 -1004 106
rect -1042 86 -1004 89
rect -953 106 -915 114
rect -953 89 -945 106
rect -923 89 -915 106
rect -953 86 -915 89
rect -864 106 -826 114
rect -864 89 -856 106
rect -834 89 -826 106
rect -864 86 -826 89
rect -775 106 -737 114
rect -775 89 -767 106
rect -745 89 -737 106
rect -775 86 -737 89
rect -686 106 -648 114
rect -686 89 -678 106
rect -656 89 -648 106
rect -686 86 -648 89
rect -597 106 -559 114
rect -597 89 -589 106
rect -567 89 -559 106
rect -597 86 -559 89
rect -508 106 -470 114
rect -508 89 -500 106
rect -478 89 -470 106
rect -508 86 -470 89
rect -419 106 -381 114
rect -419 89 -411 106
rect -389 89 -381 106
rect -419 86 -381 89
rect -330 106 -292 114
rect -330 89 -322 106
rect -300 89 -292 106
rect -330 86 -292 89
rect -241 106 -203 114
rect -241 89 -233 106
rect -211 89 -203 106
rect -241 86 -203 89
rect -152 106 -114 114
rect -152 89 -144 106
rect -122 89 -114 106
rect -152 86 -114 89
rect -63 106 -25 114
rect -63 89 -55 106
rect -33 89 -25 106
rect -63 86 -25 89
rect 25 106 63 114
rect 25 89 33 106
rect 55 89 63 106
rect 25 86 63 89
rect 114 106 152 114
rect 114 89 122 106
rect 144 89 152 106
rect 114 86 152 89
rect 203 106 241 114
rect 203 89 211 106
rect 233 89 241 106
rect 203 86 241 89
rect 292 106 330 114
rect 292 89 300 106
rect 322 89 330 106
rect 292 86 330 89
rect 381 106 419 114
rect 381 89 389 106
rect 411 89 419 106
rect 381 86 419 89
rect 470 106 508 114
rect 470 89 478 106
rect 500 89 508 106
rect 470 86 508 89
rect 559 106 597 114
rect 559 89 567 106
rect 589 89 597 106
rect 559 86 597 89
rect 648 106 686 114
rect 648 89 656 106
rect 678 89 686 106
rect 648 86 686 89
rect 737 106 775 114
rect 737 89 745 106
rect 767 89 775 106
rect 737 86 775 89
rect 826 106 864 114
rect 826 89 834 106
rect 856 89 864 106
rect 826 86 864 89
rect 915 106 953 114
rect 915 89 923 106
rect 945 89 953 106
rect 915 86 953 89
rect 1004 106 1042 114
rect 1004 89 1012 106
rect 1034 89 1042 106
rect 1004 86 1042 89
rect 1093 106 1131 114
rect 1093 89 1101 106
rect 1123 89 1131 106
rect 1093 86 1131 89
rect 1182 106 1220 114
rect 1182 89 1190 106
rect 1212 89 1220 106
rect 1182 86 1220 89
rect 1271 106 1309 114
rect 1271 89 1279 106
rect 1301 89 1309 106
rect 1271 86 1309 89
rect 1360 106 1398 114
rect 1360 89 1368 106
rect 1390 89 1398 106
rect 1360 86 1398 89
rect 1449 106 1487 114
rect 1449 89 1457 106
rect 1479 89 1487 106
rect 1449 86 1487 89
rect 1538 106 1576 114
rect 1538 89 1546 106
rect 1568 89 1576 106
rect 1538 86 1576 89
rect 1627 106 1665 114
rect 1627 89 1635 106
rect 1657 89 1665 106
rect 1627 86 1665 89
rect 1716 106 1754 114
rect 1716 89 1724 106
rect 1746 89 1754 106
rect 1716 86 1754 89
rect -1791 64 -1768 70
rect -1791 -64 -1788 64
rect -1771 -64 -1768 64
rect -1791 -70 -1768 -64
rect -1702 64 -1679 70
rect -1702 -64 -1699 64
rect -1682 -64 -1679 64
rect -1702 -70 -1679 -64
rect -1613 64 -1590 70
rect -1613 -64 -1610 64
rect -1593 -64 -1590 64
rect -1613 -70 -1590 -64
rect -1524 64 -1501 70
rect -1524 -64 -1521 64
rect -1504 -64 -1501 64
rect -1524 -70 -1501 -64
rect -1435 64 -1412 70
rect -1435 -64 -1432 64
rect -1415 -64 -1412 64
rect -1435 -70 -1412 -64
rect -1346 64 -1323 70
rect -1346 -64 -1343 64
rect -1326 -64 -1323 64
rect -1346 -70 -1323 -64
rect -1257 64 -1234 70
rect -1257 -64 -1254 64
rect -1237 -64 -1234 64
rect -1257 -70 -1234 -64
rect -1168 64 -1145 70
rect -1168 -64 -1165 64
rect -1148 -64 -1145 64
rect -1168 -70 -1145 -64
rect -1079 64 -1056 70
rect -1079 -64 -1076 64
rect -1059 -64 -1056 64
rect -1079 -70 -1056 -64
rect -990 64 -967 70
rect -990 -64 -987 64
rect -970 -64 -967 64
rect -990 -70 -967 -64
rect -901 64 -878 70
rect -901 -64 -898 64
rect -881 -64 -878 64
rect -901 -70 -878 -64
rect -812 64 -789 70
rect -812 -64 -809 64
rect -792 -64 -789 64
rect -812 -70 -789 -64
rect -723 64 -700 70
rect -723 -64 -720 64
rect -703 -64 -700 64
rect -723 -70 -700 -64
rect -634 64 -611 70
rect -634 -64 -631 64
rect -614 -64 -611 64
rect -634 -70 -611 -64
rect -545 64 -522 70
rect -545 -64 -542 64
rect -525 -64 -522 64
rect -545 -70 -522 -64
rect -456 64 -433 70
rect -456 -64 -453 64
rect -436 -64 -433 64
rect -456 -70 -433 -64
rect -367 64 -344 70
rect -367 -64 -364 64
rect -347 -64 -344 64
rect -367 -70 -344 -64
rect -278 64 -255 70
rect -278 -64 -275 64
rect -258 -64 -255 64
rect -278 -70 -255 -64
rect -189 64 -166 70
rect -189 -64 -186 64
rect -169 -64 -166 64
rect -189 -70 -166 -64
rect -100 64 -77 70
rect -100 -64 -97 64
rect -80 -64 -77 64
rect -100 -70 -77 -64
rect -11 64 11 70
rect -11 -64 -8 64
rect 8 -64 11 64
rect -11 -70 11 -64
rect 77 64 100 70
rect 77 -64 80 64
rect 97 -64 100 64
rect 77 -70 100 -64
rect 166 64 189 70
rect 166 -64 169 64
rect 186 -64 189 64
rect 166 -70 189 -64
rect 255 64 278 70
rect 255 -64 258 64
rect 275 -64 278 64
rect 255 -70 278 -64
rect 344 64 367 70
rect 344 -64 347 64
rect 364 -64 367 64
rect 344 -70 367 -64
rect 433 64 456 70
rect 433 -64 436 64
rect 453 -64 456 64
rect 433 -70 456 -64
rect 522 64 545 70
rect 522 -64 525 64
rect 542 -64 545 64
rect 522 -70 545 -64
rect 611 64 634 70
rect 611 -64 614 64
rect 631 -64 634 64
rect 611 -70 634 -64
rect 700 64 723 70
rect 700 -64 703 64
rect 720 -64 723 64
rect 700 -70 723 -64
rect 789 64 812 70
rect 789 -64 792 64
rect 809 -64 812 64
rect 789 -70 812 -64
rect 878 64 901 70
rect 878 -64 881 64
rect 898 -64 901 64
rect 878 -70 901 -64
rect 967 64 990 70
rect 967 -64 970 64
rect 987 -64 990 64
rect 967 -70 990 -64
rect 1056 64 1079 70
rect 1056 -64 1059 64
rect 1076 -64 1079 64
rect 1056 -70 1079 -64
rect 1145 64 1168 70
rect 1145 -64 1148 64
rect 1165 -64 1168 64
rect 1145 -70 1168 -64
rect 1234 64 1257 70
rect 1234 -64 1237 64
rect 1254 -64 1257 64
rect 1234 -70 1257 -64
rect 1323 64 1346 70
rect 1323 -64 1326 64
rect 1343 -64 1346 64
rect 1323 -70 1346 -64
rect 1412 64 1435 70
rect 1412 -64 1415 64
rect 1432 -64 1435 64
rect 1412 -70 1435 -64
rect 1501 64 1524 70
rect 1501 -64 1504 64
rect 1521 -64 1524 64
rect 1501 -70 1524 -64
rect 1590 64 1613 70
rect 1590 -64 1593 64
rect 1610 -64 1613 64
rect 1590 -70 1613 -64
rect 1679 64 1702 70
rect 1679 -64 1682 64
rect 1699 -64 1702 64
rect 1679 -70 1702 -64
rect 1768 64 1791 70
rect 1768 -64 1771 64
rect 1788 -64 1791 64
rect 1768 -70 1791 -64
rect -1754 -89 -1716 -86
rect -1754 -106 -1746 -89
rect -1724 -106 -1716 -89
rect -1754 -114 -1716 -106
rect -1665 -89 -1627 -86
rect -1665 -106 -1657 -89
rect -1635 -106 -1627 -89
rect -1665 -114 -1627 -106
rect -1576 -89 -1538 -86
rect -1576 -106 -1568 -89
rect -1546 -106 -1538 -89
rect -1576 -114 -1538 -106
rect -1487 -89 -1449 -86
rect -1487 -106 -1479 -89
rect -1457 -106 -1449 -89
rect -1487 -114 -1449 -106
rect -1398 -89 -1360 -86
rect -1398 -106 -1390 -89
rect -1368 -106 -1360 -89
rect -1398 -114 -1360 -106
rect -1309 -89 -1271 -86
rect -1309 -106 -1301 -89
rect -1279 -106 -1271 -89
rect -1309 -114 -1271 -106
rect -1220 -89 -1182 -86
rect -1220 -106 -1212 -89
rect -1190 -106 -1182 -89
rect -1220 -114 -1182 -106
rect -1131 -89 -1093 -86
rect -1131 -106 -1123 -89
rect -1101 -106 -1093 -89
rect -1131 -114 -1093 -106
rect -1042 -89 -1004 -86
rect -1042 -106 -1034 -89
rect -1012 -106 -1004 -89
rect -1042 -114 -1004 -106
rect -953 -89 -915 -86
rect -953 -106 -945 -89
rect -923 -106 -915 -89
rect -953 -114 -915 -106
rect -864 -89 -826 -86
rect -864 -106 -856 -89
rect -834 -106 -826 -89
rect -864 -114 -826 -106
rect -775 -89 -737 -86
rect -775 -106 -767 -89
rect -745 -106 -737 -89
rect -775 -114 -737 -106
rect -686 -89 -648 -86
rect -686 -106 -678 -89
rect -656 -106 -648 -89
rect -686 -114 -648 -106
rect -597 -89 -559 -86
rect -597 -106 -589 -89
rect -567 -106 -559 -89
rect -597 -114 -559 -106
rect -508 -89 -470 -86
rect -508 -106 -500 -89
rect -478 -106 -470 -89
rect -508 -114 -470 -106
rect -419 -89 -381 -86
rect -419 -106 -411 -89
rect -389 -106 -381 -89
rect -419 -114 -381 -106
rect -330 -89 -292 -86
rect -330 -106 -322 -89
rect -300 -106 -292 -89
rect -330 -114 -292 -106
rect -241 -89 -203 -86
rect -241 -106 -233 -89
rect -211 -106 -203 -89
rect -241 -114 -203 -106
rect -152 -89 -114 -86
rect -152 -106 -144 -89
rect -122 -106 -114 -89
rect -152 -114 -114 -106
rect -63 -89 -25 -86
rect -63 -106 -55 -89
rect -33 -106 -25 -89
rect -63 -114 -25 -106
rect 25 -89 63 -86
rect 25 -106 33 -89
rect 55 -106 63 -89
rect 25 -114 63 -106
rect 114 -89 152 -86
rect 114 -106 122 -89
rect 144 -106 152 -89
rect 114 -114 152 -106
rect 203 -89 241 -86
rect 203 -106 211 -89
rect 233 -106 241 -89
rect 203 -114 241 -106
rect 292 -89 330 -86
rect 292 -106 300 -89
rect 322 -106 330 -89
rect 292 -114 330 -106
rect 381 -89 419 -86
rect 381 -106 389 -89
rect 411 -106 419 -89
rect 381 -114 419 -106
rect 470 -89 508 -86
rect 470 -106 478 -89
rect 500 -106 508 -89
rect 470 -114 508 -106
rect 559 -89 597 -86
rect 559 -106 567 -89
rect 589 -106 597 -89
rect 559 -114 597 -106
rect 648 -89 686 -86
rect 648 -106 656 -89
rect 678 -106 686 -89
rect 648 -114 686 -106
rect 737 -89 775 -86
rect 737 -106 745 -89
rect 767 -106 775 -89
rect 737 -114 775 -106
rect 826 -89 864 -86
rect 826 -106 834 -89
rect 856 -106 864 -89
rect 826 -114 864 -106
rect 915 -89 953 -86
rect 915 -106 923 -89
rect 945 -106 953 -89
rect 915 -114 953 -106
rect 1004 -89 1042 -86
rect 1004 -106 1012 -89
rect 1034 -106 1042 -89
rect 1004 -114 1042 -106
rect 1093 -89 1131 -86
rect 1093 -106 1101 -89
rect 1123 -106 1131 -89
rect 1093 -114 1131 -106
rect 1182 -89 1220 -86
rect 1182 -106 1190 -89
rect 1212 -106 1220 -89
rect 1182 -114 1220 -106
rect 1271 -89 1309 -86
rect 1271 -106 1279 -89
rect 1301 -106 1309 -89
rect 1271 -114 1309 -106
rect 1360 -89 1398 -86
rect 1360 -106 1368 -89
rect 1390 -106 1398 -89
rect 1360 -114 1398 -106
rect 1449 -89 1487 -86
rect 1449 -106 1457 -89
rect 1479 -106 1487 -89
rect 1449 -114 1487 -106
rect 1538 -89 1576 -86
rect 1538 -106 1546 -89
rect 1568 -106 1576 -89
rect 1538 -114 1576 -106
rect 1627 -89 1665 -86
rect 1627 -106 1635 -89
rect 1657 -106 1665 -89
rect 1627 -114 1665 -106
rect 1716 -89 1754 -86
rect 1716 -106 1724 -89
rect 1746 -106 1754 -89
rect 1716 -114 1754 -106
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 40 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
