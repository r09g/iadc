magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -29 82 29 88
rect -29 48 -17 82
rect -29 42 29 48
<< pwell >>
rect -99 -116 99 36
<< nmos >>
rect -15 -90 15 10
<< ndiff >>
rect -73 -23 -15 10
rect -73 -57 -61 -23
rect -27 -57 -15 -23
rect -73 -90 -15 -57
rect 15 -23 73 10
rect 15 -57 27 -23
rect 61 -57 73 -23
rect 15 -90 73 -57
<< ndiffc >>
rect -61 -57 -27 -23
rect 27 -57 61 -23
<< poly >>
rect -33 82 33 98
rect -33 48 -17 82
rect 17 48 33 82
rect -33 32 33 48
rect -15 10 15 32
rect -15 -116 15 -90
<< polycont >>
rect -17 48 17 82
<< locali >>
rect -33 48 -17 82
rect 17 48 33 82
rect -61 -23 -27 14
rect -61 -94 -27 -57
rect 27 -23 61 14
rect 27 -94 61 -57
<< viali >>
rect -17 48 17 82
rect -61 -57 -27 -23
rect 27 -57 61 -23
<< metal1 >>
rect -29 82 29 88
rect -29 48 -17 82
rect 17 48 29 82
rect -29 42 29 48
rect -67 -23 -21 10
rect -67 -57 -61 -23
rect -27 -57 -21 -23
rect -67 -90 -21 -57
rect 21 -23 67 10
rect 21 -57 27 -23
rect 61 -57 67 -23
rect 21 -90 67 -57
<< end >>
