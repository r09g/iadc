magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -28 82 30 88
rect -28 48 -16 82
rect -28 42 30 48
<< pwell >>
rect -98 -116 100 36
<< nmos >>
rect -14 -90 16 10
<< ndiff >>
rect -72 -23 -14 10
rect -72 -57 -60 -23
rect -26 -57 -14 -23
rect -72 -90 -14 -57
rect 16 -23 74 10
rect 16 -57 28 -23
rect 62 -57 74 -23
rect 16 -90 74 -57
<< ndiffc >>
rect -60 -57 -26 -23
rect 28 -57 62 -23
<< poly >>
rect -32 82 34 98
rect -32 48 -16 82
rect 18 48 34 82
rect -32 32 34 48
rect -14 10 16 32
rect -14 -116 16 -90
<< polycont >>
rect -16 48 18 82
<< locali >>
rect -32 48 -16 82
rect 18 48 34 82
rect -60 -23 -26 14
rect -60 -94 -26 -57
rect 28 -23 62 14
rect 28 -94 62 -57
<< viali >>
rect -16 48 18 82
rect -60 -57 -26 -23
rect 28 -57 62 -23
<< metal1 >>
rect -28 82 30 88
rect -28 48 -16 82
rect 18 48 30 82
rect -28 42 30 48
rect -66 -23 -20 10
rect -66 -57 -60 -23
rect -26 -57 -20 -23
rect -66 -90 -20 -57
rect 22 -23 68 10
rect 22 -57 28 -23
rect 62 -57 68 -23
rect 22 -90 68 -57
<< end >>
