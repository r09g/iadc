magic
tech sky130A
magscale 1 2
timestamp 1652661863
<< viali >>
rect 1171 545 1205 931
rect 1171 81 1205 281
<< metal1 >>
rect -87 993 995 1027
rect -216 883 -189 935
rect -137 883 -127 935
rect -87 430 -53 993
rect 78 883 88 935
rect 140 883 150 935
rect 193 832 227 993
rect 271 883 281 935
rect 333 883 343 935
rect 385 832 419 993
rect 462 883 472 935
rect 524 883 534 935
rect 577 832 611 993
rect 654 883 664 935
rect 716 883 726 935
rect 769 832 803 993
rect 846 883 856 935
rect 908 883 918 935
rect 961 832 995 993
rect 1038 883 1048 935
rect 1100 883 1110 935
rect 1165 931 1211 1063
rect -216 396 -53 430
rect -216 76 -189 128
rect -137 76 -127 128
rect -87 19 -53 396
rect 97 430 131 608
rect 289 430 323 608
rect 481 430 515 608
rect 673 430 707 608
rect 865 430 899 608
rect 1057 430 1091 608
rect 1165 545 1171 931
rect 1205 545 1211 931
rect 1165 533 1211 545
rect 97 396 1283 430
rect 97 253 131 396
rect 289 253 323 396
rect 481 253 515 396
rect 673 253 707 396
rect 865 253 899 396
rect 1057 253 1091 396
rect 1165 281 1211 293
rect 78 76 88 128
rect 140 76 150 128
rect 193 19 227 180
rect 269 76 279 128
rect 331 76 341 128
rect 385 19 419 180
rect 461 76 471 128
rect 523 76 533 128
rect 577 19 611 180
rect 653 76 663 128
rect 715 76 725 128
rect 769 19 803 180
rect 846 75 856 127
rect 908 75 918 127
rect 961 19 995 180
rect 1038 75 1048 127
rect 1100 75 1110 127
rect 1165 81 1171 281
rect 1205 81 1211 281
rect -87 -15 995 19
rect 1165 -51 1211 81
<< via1 >>
rect -189 883 -137 935
rect 88 883 140 935
rect 281 883 333 935
rect 472 883 524 935
rect 664 883 716 935
rect 856 883 908 935
rect 1048 883 1100 935
rect -189 76 -137 128
rect 88 76 140 128
rect 279 76 331 128
rect 471 76 523 128
rect 663 76 715 128
rect 856 75 908 127
rect 1048 75 1100 127
<< metal2 >>
rect -189 935 -137 945
rect 88 935 140 945
rect 281 935 333 945
rect 472 935 524 945
rect 664 935 716 945
rect 856 935 908 945
rect 1048 935 1100 945
rect -137 883 88 935
rect 140 883 281 935
rect 333 883 472 935
rect 524 883 664 935
rect 716 883 856 935
rect 908 883 1048 935
rect 1100 883 1107 935
rect -189 873 -137 883
rect 88 873 140 883
rect 281 873 333 883
rect 472 873 524 883
rect 664 873 716 883
rect 856 873 908 883
rect 1048 873 1100 883
rect -189 128 -137 138
rect 88 128 140 138
rect 279 128 331 138
rect 471 128 523 138
rect 663 128 715 138
rect 856 128 908 137
rect 1048 128 1100 137
rect -137 76 88 128
rect 140 76 279 128
rect 331 76 471 128
rect 523 76 663 128
rect 715 127 1107 128
rect 715 76 856 127
rect -189 66 -137 76
rect 88 66 140 76
rect 279 66 331 76
rect 471 66 523 76
rect 663 66 715 76
rect 908 76 1048 127
rect 856 65 908 75
rect 1100 76 1107 127
rect 1048 65 1100 75
use sky130_fd_pr__nfet_01v8_6J4AMR  sky130_fd_pr__nfet_01v8_6J4AMR_0
timestamp 1652660033
transform 1 0 594 0 1 212
box -647 -263 647 201
use sky130_fd_pr__pfet_01v8_UNG2NQ  sky130_fd_pr__pfet_01v8_UNG2NQ_0
timestamp 1652659422
transform -1 0 594 0 -1 707
box -647 -356 647 294
<< labels >>
flabel metal1 1188 -48 1188 -48 1 FreeSans 400 0 0 0 VSS
flabel metal1 1188 1058 1188 1058 5 FreeSans 400 0 0 0 VDD
flabel metal1 -211 909 -211 909 3 FreeSans 400 0 0 0 en_b
flabel metal1 -212 413 -212 413 3 FreeSans 400 0 0 0 in
flabel metal1 -212 102 -212 102 3 FreeSans 400 0 0 0 en
flabel metal1 1279 412 1279 412 7 FreeSans 400 0 0 0 out
<< end >>