magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< metal3 >>
rect -1310 -1260 1210 1260
<< mimcap >>
rect -1210 1112 1110 1160
rect -1210 -1112 -1162 1112
rect 1062 -1112 1110 1112
rect -1210 -1160 1110 -1112
<< mimcapcontact >>
rect -1162 -1112 1062 1112
<< metal4 >>
rect -1171 1112 1071 1121
rect -1171 -1112 -1162 1112
rect 1062 -1112 1071 1112
rect -1171 -1121 1071 -1112
<< properties >>
string FIXED_BBOX -1310 -1260 1210 1260
<< end >>
