magic
tech sky130A
timestamp 1654517900
<< nwell >>
rect -1056 -120 1056 120
<< pmos >>
rect -1009 -70 -949 70
rect -920 -70 -860 70
rect -831 -70 -771 70
rect -742 -70 -682 70
rect -653 -70 -593 70
rect -564 -70 -504 70
rect -475 -70 -415 70
rect -386 -70 -326 70
rect -297 -70 -237 70
rect -208 -70 -148 70
rect -119 -70 -59 70
rect -30 -70 30 70
rect 59 -70 119 70
rect 148 -70 208 70
rect 237 -70 297 70
rect 326 -70 386 70
rect 415 -70 475 70
rect 504 -70 564 70
rect 593 -70 653 70
rect 682 -70 742 70
rect 771 -70 831 70
rect 860 -70 920 70
rect 949 -70 1009 70
<< pdiff >>
rect -1038 64 -1009 70
rect -1038 -64 -1032 64
rect -1015 -64 -1009 64
rect -1038 -70 -1009 -64
rect -949 64 -920 70
rect -949 -64 -943 64
rect -926 -64 -920 64
rect -949 -70 -920 -64
rect -860 64 -831 70
rect -860 -64 -854 64
rect -837 -64 -831 64
rect -860 -70 -831 -64
rect -771 64 -742 70
rect -771 -64 -765 64
rect -748 -64 -742 64
rect -771 -70 -742 -64
rect -682 64 -653 70
rect -682 -64 -676 64
rect -659 -64 -653 64
rect -682 -70 -653 -64
rect -593 64 -564 70
rect -593 -64 -587 64
rect -570 -64 -564 64
rect -593 -70 -564 -64
rect -504 64 -475 70
rect -504 -64 -498 64
rect -481 -64 -475 64
rect -504 -70 -475 -64
rect -415 64 -386 70
rect -415 -64 -409 64
rect -392 -64 -386 64
rect -415 -70 -386 -64
rect -326 64 -297 70
rect -326 -64 -320 64
rect -303 -64 -297 64
rect -326 -70 -297 -64
rect -237 64 -208 70
rect -237 -64 -231 64
rect -214 -64 -208 64
rect -237 -70 -208 -64
rect -148 64 -119 70
rect -148 -64 -142 64
rect -125 -64 -119 64
rect -148 -70 -119 -64
rect -59 64 -30 70
rect -59 -64 -53 64
rect -36 -64 -30 64
rect -59 -70 -30 -64
rect 30 64 59 70
rect 30 -64 36 64
rect 53 -64 59 64
rect 30 -70 59 -64
rect 119 64 148 70
rect 119 -64 125 64
rect 142 -64 148 64
rect 119 -70 148 -64
rect 208 64 237 70
rect 208 -64 214 64
rect 231 -64 237 64
rect 208 -70 237 -64
rect 297 64 326 70
rect 297 -64 303 64
rect 320 -64 326 64
rect 297 -70 326 -64
rect 386 64 415 70
rect 386 -64 392 64
rect 409 -64 415 64
rect 386 -70 415 -64
rect 475 64 504 70
rect 475 -64 481 64
rect 498 -64 504 64
rect 475 -70 504 -64
rect 564 64 593 70
rect 564 -64 570 64
rect 587 -64 593 64
rect 564 -70 593 -64
rect 653 64 682 70
rect 653 -64 659 64
rect 676 -64 682 64
rect 653 -70 682 -64
rect 742 64 771 70
rect 742 -64 748 64
rect 765 -64 771 64
rect 742 -70 771 -64
rect 831 64 860 70
rect 831 -64 837 64
rect 854 -64 860 64
rect 831 -70 860 -64
rect 920 64 949 70
rect 920 -64 926 64
rect 943 -64 949 64
rect 920 -70 949 -64
rect 1009 64 1038 70
rect 1009 -64 1015 64
rect 1032 -64 1038 64
rect 1009 -70 1038 -64
<< pdiffc >>
rect -1032 -64 -1015 64
rect -943 -64 -926 64
rect -854 -64 -837 64
rect -765 -64 -748 64
rect -676 -64 -659 64
rect -587 -64 -570 64
rect -498 -64 -481 64
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
rect 481 -64 498 64
rect 570 -64 587 64
rect 659 -64 676 64
rect 748 -64 765 64
rect 837 -64 854 64
rect 926 -64 943 64
rect 1015 -64 1032 64
<< poly >>
rect -998 110 -960 118
rect -998 102 -990 110
rect -1009 93 -990 102
rect -968 102 -960 110
rect -909 110 -871 118
rect -909 102 -901 110
rect -968 93 -949 102
rect -1009 70 -949 93
rect -920 93 -901 102
rect -879 102 -871 110
rect -820 110 -782 118
rect -820 102 -812 110
rect -879 93 -860 102
rect -920 70 -860 93
rect -831 93 -812 102
rect -790 102 -782 110
rect -731 110 -693 118
rect -731 102 -723 110
rect -790 93 -771 102
rect -831 70 -771 93
rect -742 93 -723 102
rect -701 102 -693 110
rect -642 110 -604 118
rect -642 102 -634 110
rect -701 93 -682 102
rect -742 70 -682 93
rect -653 93 -634 102
rect -612 102 -604 110
rect -553 110 -515 118
rect -553 102 -545 110
rect -612 93 -593 102
rect -653 70 -593 93
rect -564 93 -545 102
rect -523 102 -515 110
rect -464 110 -426 118
rect -464 102 -456 110
rect -523 93 -504 102
rect -564 70 -504 93
rect -475 93 -456 102
rect -434 102 -426 110
rect -375 110 -337 118
rect -375 102 -367 110
rect -434 93 -415 102
rect -475 70 -415 93
rect -386 93 -367 102
rect -345 102 -337 110
rect -286 110 -248 118
rect -286 102 -278 110
rect -345 93 -326 102
rect -386 70 -326 93
rect -297 93 -278 102
rect -256 102 -248 110
rect -197 110 -159 118
rect -197 102 -189 110
rect -256 93 -237 102
rect -297 70 -237 93
rect -208 93 -189 102
rect -167 102 -159 110
rect -108 110 -70 118
rect -108 102 -100 110
rect -167 93 -148 102
rect -208 70 -148 93
rect -119 93 -100 102
rect -78 102 -70 110
rect -19 110 19 118
rect -19 102 -11 110
rect -78 93 -59 102
rect -119 70 -59 93
rect -30 93 -11 102
rect 11 102 19 110
rect 70 110 108 118
rect 70 102 78 110
rect 11 93 30 102
rect -30 70 30 93
rect 59 93 78 102
rect 100 102 108 110
rect 159 110 197 118
rect 159 102 167 110
rect 100 93 119 102
rect 59 70 119 93
rect 148 93 167 102
rect 189 102 197 110
rect 248 110 286 118
rect 248 102 256 110
rect 189 93 208 102
rect 148 70 208 93
rect 237 93 256 102
rect 278 102 286 110
rect 337 110 375 118
rect 337 102 345 110
rect 278 93 297 102
rect 237 70 297 93
rect 326 93 345 102
rect 367 102 375 110
rect 426 110 464 118
rect 426 102 434 110
rect 367 93 386 102
rect 326 70 386 93
rect 415 93 434 102
rect 456 102 464 110
rect 515 110 553 118
rect 515 102 523 110
rect 456 93 475 102
rect 415 70 475 93
rect 504 93 523 102
rect 545 102 553 110
rect 604 110 642 118
rect 604 102 612 110
rect 545 93 564 102
rect 504 70 564 93
rect 593 93 612 102
rect 634 102 642 110
rect 693 110 731 118
rect 693 102 701 110
rect 634 93 653 102
rect 593 70 653 93
rect 682 93 701 102
rect 723 102 731 110
rect 782 110 820 118
rect 782 102 790 110
rect 723 93 742 102
rect 682 70 742 93
rect 771 93 790 102
rect 812 102 820 110
rect 871 110 909 118
rect 871 102 879 110
rect 812 93 831 102
rect 771 70 831 93
rect 860 93 879 102
rect 901 102 909 110
rect 960 110 998 118
rect 960 102 968 110
rect 901 93 920 102
rect 860 70 920 93
rect 949 93 968 102
rect 990 102 998 110
rect 990 93 1009 102
rect 949 70 1009 93
rect -1009 -93 -949 -70
rect -1009 -102 -990 -93
rect -998 -110 -990 -102
rect -968 -102 -949 -93
rect -920 -93 -860 -70
rect -920 -102 -901 -93
rect -968 -110 -960 -102
rect -998 -118 -960 -110
rect -909 -110 -901 -102
rect -879 -102 -860 -93
rect -831 -93 -771 -70
rect -831 -102 -812 -93
rect -879 -110 -871 -102
rect -909 -118 -871 -110
rect -820 -110 -812 -102
rect -790 -102 -771 -93
rect -742 -93 -682 -70
rect -742 -102 -723 -93
rect -790 -110 -782 -102
rect -820 -118 -782 -110
rect -731 -110 -723 -102
rect -701 -102 -682 -93
rect -653 -93 -593 -70
rect -653 -102 -634 -93
rect -701 -110 -693 -102
rect -731 -118 -693 -110
rect -642 -110 -634 -102
rect -612 -102 -593 -93
rect -564 -93 -504 -70
rect -564 -102 -545 -93
rect -612 -110 -604 -102
rect -642 -118 -604 -110
rect -553 -110 -545 -102
rect -523 -102 -504 -93
rect -475 -93 -415 -70
rect -475 -102 -456 -93
rect -523 -110 -515 -102
rect -553 -118 -515 -110
rect -464 -110 -456 -102
rect -434 -102 -415 -93
rect -386 -93 -326 -70
rect -386 -102 -367 -93
rect -434 -110 -426 -102
rect -464 -118 -426 -110
rect -375 -110 -367 -102
rect -345 -102 -326 -93
rect -297 -93 -237 -70
rect -297 -102 -278 -93
rect -345 -110 -337 -102
rect -375 -118 -337 -110
rect -286 -110 -278 -102
rect -256 -102 -237 -93
rect -208 -93 -148 -70
rect -208 -102 -189 -93
rect -256 -110 -248 -102
rect -286 -118 -248 -110
rect -197 -110 -189 -102
rect -167 -102 -148 -93
rect -119 -93 -59 -70
rect -119 -102 -100 -93
rect -167 -110 -159 -102
rect -197 -118 -159 -110
rect -108 -110 -100 -102
rect -78 -102 -59 -93
rect -30 -93 30 -70
rect -30 -102 -11 -93
rect -78 -110 -70 -102
rect -108 -118 -70 -110
rect -19 -110 -11 -102
rect 11 -102 30 -93
rect 59 -93 119 -70
rect 59 -102 78 -93
rect 11 -110 19 -102
rect -19 -118 19 -110
rect 70 -110 78 -102
rect 100 -102 119 -93
rect 148 -93 208 -70
rect 148 -102 167 -93
rect 100 -110 108 -102
rect 70 -118 108 -110
rect 159 -110 167 -102
rect 189 -102 208 -93
rect 237 -93 297 -70
rect 237 -102 256 -93
rect 189 -110 197 -102
rect 159 -118 197 -110
rect 248 -110 256 -102
rect 278 -102 297 -93
rect 326 -93 386 -70
rect 326 -102 345 -93
rect 278 -110 286 -102
rect 248 -118 286 -110
rect 337 -110 345 -102
rect 367 -102 386 -93
rect 415 -93 475 -70
rect 415 -102 434 -93
rect 367 -110 375 -102
rect 337 -118 375 -110
rect 426 -110 434 -102
rect 456 -102 475 -93
rect 504 -93 564 -70
rect 504 -102 523 -93
rect 456 -110 464 -102
rect 426 -118 464 -110
rect 515 -110 523 -102
rect 545 -102 564 -93
rect 593 -93 653 -70
rect 593 -102 612 -93
rect 545 -110 553 -102
rect 515 -118 553 -110
rect 604 -110 612 -102
rect 634 -102 653 -93
rect 682 -93 742 -70
rect 682 -102 701 -93
rect 634 -110 642 -102
rect 604 -118 642 -110
rect 693 -110 701 -102
rect 723 -102 742 -93
rect 771 -93 831 -70
rect 771 -102 790 -93
rect 723 -110 731 -102
rect 693 -118 731 -110
rect 782 -110 790 -102
rect 812 -102 831 -93
rect 860 -93 920 -70
rect 860 -102 879 -93
rect 812 -110 820 -102
rect 782 -118 820 -110
rect 871 -110 879 -102
rect 901 -102 920 -93
rect 949 -93 1009 -70
rect 949 -102 968 -93
rect 901 -110 909 -102
rect 871 -118 909 -110
rect 960 -110 968 -102
rect 990 -102 1009 -93
rect 990 -110 998 -102
rect 960 -118 998 -110
<< polycont >>
rect -990 93 -968 110
rect -901 93 -879 110
rect -812 93 -790 110
rect -723 93 -701 110
rect -634 93 -612 110
rect -545 93 -523 110
rect -456 93 -434 110
rect -367 93 -345 110
rect -278 93 -256 110
rect -189 93 -167 110
rect -100 93 -78 110
rect -11 93 11 110
rect 78 93 100 110
rect 167 93 189 110
rect 256 93 278 110
rect 345 93 367 110
rect 434 93 456 110
rect 523 93 545 110
rect 612 93 634 110
rect 701 93 723 110
rect 790 93 812 110
rect 879 93 901 110
rect 968 93 990 110
rect -990 -110 -968 -93
rect -901 -110 -879 -93
rect -812 -110 -790 -93
rect -723 -110 -701 -93
rect -634 -110 -612 -93
rect -545 -110 -523 -93
rect -456 -110 -434 -93
rect -367 -110 -345 -93
rect -278 -110 -256 -93
rect -189 -110 -167 -93
rect -100 -110 -78 -93
rect -11 -110 11 -93
rect 78 -110 100 -93
rect 167 -110 189 -93
rect 256 -110 278 -93
rect 345 -110 367 -93
rect 434 -110 456 -93
rect 523 -110 545 -93
rect 612 -110 634 -93
rect 701 -110 723 -93
rect 790 -110 812 -93
rect 879 -110 901 -93
rect 968 -110 990 -93
<< locali >>
rect -998 93 -990 110
rect -968 93 -960 110
rect -909 93 -901 110
rect -879 93 -871 110
rect -820 93 -812 110
rect -790 93 -782 110
rect -731 93 -723 110
rect -701 93 -693 110
rect -642 93 -634 110
rect -612 93 -604 110
rect -553 93 -545 110
rect -523 93 -515 110
rect -464 93 -456 110
rect -434 93 -426 110
rect -375 93 -367 110
rect -345 93 -337 110
rect -286 93 -278 110
rect -256 93 -248 110
rect -197 93 -189 110
rect -167 93 -159 110
rect -108 93 -100 110
rect -78 93 -70 110
rect -19 93 -11 110
rect 11 93 19 110
rect 70 93 78 110
rect 100 93 108 110
rect 159 93 167 110
rect 189 93 197 110
rect 248 93 256 110
rect 278 93 286 110
rect 337 93 345 110
rect 367 93 375 110
rect 426 93 434 110
rect 456 93 464 110
rect 515 93 523 110
rect 545 93 553 110
rect 604 93 612 110
rect 634 93 642 110
rect 693 93 701 110
rect 723 93 731 110
rect 782 93 790 110
rect 812 93 820 110
rect 871 93 879 110
rect 901 93 909 110
rect 960 93 968 110
rect 990 93 998 110
rect -1032 64 -1015 72
rect -1032 -72 -1015 -64
rect -943 64 -926 72
rect -943 -72 -926 -64
rect -854 64 -837 72
rect -854 -72 -837 -64
rect -765 64 -748 72
rect -765 -72 -748 -64
rect -676 64 -659 72
rect -676 -72 -659 -64
rect -587 64 -570 72
rect -587 -72 -570 -64
rect -498 64 -481 72
rect -498 -72 -481 -64
rect -409 64 -392 72
rect -409 -72 -392 -64
rect -320 64 -303 72
rect -320 -72 -303 -64
rect -231 64 -214 72
rect -231 -72 -214 -64
rect -142 64 -125 72
rect -142 -72 -125 -64
rect -53 64 -36 72
rect -53 -72 -36 -64
rect 36 64 53 72
rect 36 -72 53 -64
rect 125 64 142 72
rect 125 -72 142 -64
rect 214 64 231 72
rect 214 -72 231 -64
rect 303 64 320 72
rect 303 -72 320 -64
rect 392 64 409 72
rect 392 -72 409 -64
rect 481 64 498 72
rect 481 -72 498 -64
rect 570 64 587 72
rect 570 -72 587 -64
rect 659 64 676 72
rect 659 -72 676 -64
rect 748 64 765 72
rect 748 -72 765 -64
rect 837 64 854 72
rect 837 -72 854 -64
rect 926 64 943 72
rect 926 -72 943 -64
rect 1015 64 1032 72
rect 1015 -72 1032 -64
rect -998 -110 -990 -93
rect -968 -110 -960 -93
rect -909 -110 -901 -93
rect -879 -110 -871 -93
rect -820 -110 -812 -93
rect -790 -110 -782 -93
rect -731 -110 -723 -93
rect -701 -110 -693 -93
rect -642 -110 -634 -93
rect -612 -110 -604 -93
rect -553 -110 -545 -93
rect -523 -110 -515 -93
rect -464 -110 -456 -93
rect -434 -110 -426 -93
rect -375 -110 -367 -93
rect -345 -110 -337 -93
rect -286 -110 -278 -93
rect -256 -110 -248 -93
rect -197 -110 -189 -93
rect -167 -110 -159 -93
rect -108 -110 -100 -93
rect -78 -110 -70 -93
rect -19 -110 -11 -93
rect 11 -110 19 -93
rect 70 -110 78 -93
rect 100 -110 108 -93
rect 159 -110 167 -93
rect 189 -110 197 -93
rect 248 -110 256 -93
rect 278 -110 286 -93
rect 337 -110 345 -93
rect 367 -110 375 -93
rect 426 -110 434 -93
rect 456 -110 464 -93
rect 515 -110 523 -93
rect 545 -110 553 -93
rect 604 -110 612 -93
rect 634 -110 642 -93
rect 693 -110 701 -93
rect 723 -110 731 -93
rect 782 -110 790 -93
rect 812 -110 820 -93
rect 871 -110 879 -93
rect 901 -110 909 -93
rect 960 -110 968 -93
rect 990 -110 998 -93
<< viali >>
rect -990 93 -968 110
rect -901 93 -879 110
rect -812 93 -790 110
rect -723 93 -701 110
rect -634 93 -612 110
rect -545 93 -523 110
rect -456 93 -434 110
rect -367 93 -345 110
rect -278 93 -256 110
rect -189 93 -167 110
rect -100 93 -78 110
rect -11 93 11 110
rect 78 93 100 110
rect 167 93 189 110
rect 256 93 278 110
rect 345 93 367 110
rect 434 93 456 110
rect 523 93 545 110
rect 612 93 634 110
rect 701 93 723 110
rect 790 93 812 110
rect 879 93 901 110
rect 968 93 990 110
rect -1032 -64 -1015 64
rect -943 -64 -926 64
rect -854 -64 -837 64
rect -765 -64 -748 64
rect -676 -64 -659 64
rect -587 -64 -570 64
rect -498 -64 -481 64
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
rect 481 -64 498 64
rect 570 -64 587 64
rect 659 -64 676 64
rect 748 -64 765 64
rect 837 -64 854 64
rect 926 -64 943 64
rect 1015 -64 1032 64
rect -990 -110 -968 -93
rect -901 -110 -879 -93
rect -812 -110 -790 -93
rect -723 -110 -701 -93
rect -634 -110 -612 -93
rect -545 -110 -523 -93
rect -456 -110 -434 -93
rect -367 -110 -345 -93
rect -278 -110 -256 -93
rect -189 -110 -167 -93
rect -100 -110 -78 -93
rect -11 -110 11 -93
rect 78 -110 100 -93
rect 167 -110 189 -93
rect 256 -110 278 -93
rect 345 -110 367 -93
rect 434 -110 456 -93
rect 523 -110 545 -93
rect 612 -110 634 -93
rect 701 -110 723 -93
rect 790 -110 812 -93
rect 879 -110 901 -93
rect 968 -110 990 -93
<< metal1 >>
rect -998 110 -960 118
rect -998 93 -990 110
rect -968 93 -960 110
rect -998 90 -960 93
rect -909 110 -871 118
rect -909 93 -901 110
rect -879 93 -871 110
rect -909 90 -871 93
rect -820 110 -782 118
rect -820 93 -812 110
rect -790 93 -782 110
rect -820 90 -782 93
rect -731 110 -693 118
rect -731 93 -723 110
rect -701 93 -693 110
rect -731 90 -693 93
rect -642 110 -604 118
rect -642 93 -634 110
rect -612 93 -604 110
rect -642 90 -604 93
rect -553 110 -515 118
rect -553 93 -545 110
rect -523 93 -515 110
rect -553 90 -515 93
rect -464 110 -426 118
rect -464 93 -456 110
rect -434 93 -426 110
rect -464 90 -426 93
rect -375 110 -337 118
rect -375 93 -367 110
rect -345 93 -337 110
rect -375 90 -337 93
rect -286 110 -248 118
rect -286 93 -278 110
rect -256 93 -248 110
rect -286 90 -248 93
rect -197 110 -159 118
rect -197 93 -189 110
rect -167 93 -159 110
rect -197 90 -159 93
rect -108 110 -70 118
rect -108 93 -100 110
rect -78 93 -70 110
rect -108 90 -70 93
rect -19 110 19 118
rect -19 93 -11 110
rect 11 93 19 110
rect -19 90 19 93
rect 70 110 108 118
rect 70 93 78 110
rect 100 93 108 110
rect 70 90 108 93
rect 159 110 197 118
rect 159 93 167 110
rect 189 93 197 110
rect 159 90 197 93
rect 248 110 286 118
rect 248 93 256 110
rect 278 93 286 110
rect 248 90 286 93
rect 337 110 375 118
rect 337 93 345 110
rect 367 93 375 110
rect 337 90 375 93
rect 426 110 464 118
rect 426 93 434 110
rect 456 93 464 110
rect 426 90 464 93
rect 515 110 553 118
rect 515 93 523 110
rect 545 93 553 110
rect 515 90 553 93
rect 604 110 642 118
rect 604 93 612 110
rect 634 93 642 110
rect 604 90 642 93
rect 693 110 731 118
rect 693 93 701 110
rect 723 93 731 110
rect 693 90 731 93
rect 782 110 820 118
rect 782 93 790 110
rect 812 93 820 110
rect 782 90 820 93
rect 871 110 909 118
rect 871 93 879 110
rect 901 93 909 110
rect 871 90 909 93
rect 960 110 998 118
rect 960 93 968 110
rect 990 93 998 110
rect 960 90 998 93
rect -1035 64 -1012 70
rect -1035 -64 -1032 64
rect -1015 -64 -1012 64
rect -1035 -70 -1012 -64
rect -946 64 -923 70
rect -946 -64 -943 64
rect -926 -64 -923 64
rect -946 -70 -923 -64
rect -857 64 -834 70
rect -857 -64 -854 64
rect -837 -64 -834 64
rect -857 -70 -834 -64
rect -768 64 -745 70
rect -768 -64 -765 64
rect -748 -64 -745 64
rect -768 -70 -745 -64
rect -679 64 -656 70
rect -679 -64 -676 64
rect -659 -64 -656 64
rect -679 -70 -656 -64
rect -590 64 -567 70
rect -590 -64 -587 64
rect -570 -64 -567 64
rect -590 -70 -567 -64
rect -501 64 -478 70
rect -501 -64 -498 64
rect -481 -64 -478 64
rect -501 -70 -478 -64
rect -412 64 -389 70
rect -412 -64 -409 64
rect -392 -64 -389 64
rect -412 -70 -389 -64
rect -323 64 -300 70
rect -323 -64 -320 64
rect -303 -64 -300 64
rect -323 -70 -300 -64
rect -234 64 -211 70
rect -234 -64 -231 64
rect -214 -64 -211 64
rect -234 -70 -211 -64
rect -145 64 -122 70
rect -145 -64 -142 64
rect -125 -64 -122 64
rect -145 -70 -122 -64
rect -56 64 -33 70
rect -56 -64 -53 64
rect -36 -64 -33 64
rect -56 -70 -33 -64
rect 33 64 56 70
rect 33 -64 36 64
rect 53 -64 56 64
rect 33 -70 56 -64
rect 122 64 145 70
rect 122 -64 125 64
rect 142 -64 145 64
rect 122 -70 145 -64
rect 211 64 234 70
rect 211 -64 214 64
rect 231 -64 234 64
rect 211 -70 234 -64
rect 300 64 323 70
rect 300 -64 303 64
rect 320 -64 323 64
rect 300 -70 323 -64
rect 389 64 412 70
rect 389 -64 392 64
rect 409 -64 412 64
rect 389 -70 412 -64
rect 478 64 501 70
rect 478 -64 481 64
rect 498 -64 501 64
rect 478 -70 501 -64
rect 567 64 590 70
rect 567 -64 570 64
rect 587 -64 590 64
rect 567 -70 590 -64
rect 656 64 679 70
rect 656 -64 659 64
rect 676 -64 679 64
rect 656 -70 679 -64
rect 745 64 768 70
rect 745 -64 748 64
rect 765 -64 768 64
rect 745 -70 768 -64
rect 834 64 857 70
rect 834 -64 837 64
rect 854 -64 857 64
rect 834 -70 857 -64
rect 923 64 946 70
rect 923 -64 926 64
rect 943 -64 946 64
rect 923 -70 946 -64
rect 1012 64 1035 70
rect 1012 -64 1015 64
rect 1032 -64 1035 64
rect 1012 -70 1035 -64
rect -998 -93 -960 -90
rect -998 -110 -990 -93
rect -968 -110 -960 -93
rect -998 -118 -960 -110
rect -909 -93 -871 -90
rect -909 -110 -901 -93
rect -879 -110 -871 -93
rect -909 -118 -871 -110
rect -820 -93 -782 -90
rect -820 -110 -812 -93
rect -790 -110 -782 -93
rect -820 -118 -782 -110
rect -731 -93 -693 -90
rect -731 -110 -723 -93
rect -701 -110 -693 -93
rect -731 -118 -693 -110
rect -642 -93 -604 -90
rect -642 -110 -634 -93
rect -612 -110 -604 -93
rect -642 -118 -604 -110
rect -553 -93 -515 -90
rect -553 -110 -545 -93
rect -523 -110 -515 -93
rect -553 -118 -515 -110
rect -464 -93 -426 -90
rect -464 -110 -456 -93
rect -434 -110 -426 -93
rect -464 -118 -426 -110
rect -375 -93 -337 -90
rect -375 -110 -367 -93
rect -345 -110 -337 -93
rect -375 -118 -337 -110
rect -286 -93 -248 -90
rect -286 -110 -278 -93
rect -256 -110 -248 -93
rect -286 -118 -248 -110
rect -197 -93 -159 -90
rect -197 -110 -189 -93
rect -167 -110 -159 -93
rect -197 -118 -159 -110
rect -108 -93 -70 -90
rect -108 -110 -100 -93
rect -78 -110 -70 -93
rect -108 -118 -70 -110
rect -19 -93 19 -90
rect -19 -110 -11 -93
rect 11 -110 19 -93
rect -19 -118 19 -110
rect 70 -93 108 -90
rect 70 -110 78 -93
rect 100 -110 108 -93
rect 70 -118 108 -110
rect 159 -93 197 -90
rect 159 -110 167 -93
rect 189 -110 197 -93
rect 159 -118 197 -110
rect 248 -93 286 -90
rect 248 -110 256 -93
rect 278 -110 286 -93
rect 248 -118 286 -110
rect 337 -93 375 -90
rect 337 -110 345 -93
rect 367 -110 375 -93
rect 337 -118 375 -110
rect 426 -93 464 -90
rect 426 -110 434 -93
rect 456 -110 464 -93
rect 426 -118 464 -110
rect 515 -93 553 -90
rect 515 -110 523 -93
rect 545 -110 553 -93
rect 515 -118 553 -110
rect 604 -93 642 -90
rect 604 -110 612 -93
rect 634 -110 642 -93
rect 604 -118 642 -110
rect 693 -93 731 -90
rect 693 -110 701 -93
rect 723 -110 731 -93
rect 693 -118 731 -110
rect 782 -93 820 -90
rect 782 -110 790 -93
rect 812 -110 820 -93
rect 782 -118 820 -110
rect 871 -93 909 -90
rect 871 -110 879 -93
rect 901 -110 909 -93
rect 871 -118 909 -110
rect 960 -93 998 -90
rect 960 -110 968 -93
rect 990 -110 998 -93
rect 960 -118 998 -110
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 23 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
