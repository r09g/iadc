magic
tech sky130A
magscale 1 2
timestamp 1654644491
<< pwell >>
rect -1591 -1097 1591 1097
<< nmoslvt >>
rect -1395 607 -1275 887
rect -1217 607 -1097 887
rect -1039 607 -919 887
rect -861 607 -741 887
rect -683 607 -563 887
rect -505 607 -385 887
rect -327 607 -207 887
rect -149 607 -29 887
rect 29 607 149 887
rect 207 607 327 887
rect 385 607 505 887
rect 563 607 683 887
rect 741 607 861 887
rect 919 607 1039 887
rect 1097 607 1217 887
rect 1275 607 1395 887
rect -1395 109 -1275 389
rect -1217 109 -1097 389
rect -1039 109 -919 389
rect -861 109 -741 389
rect -683 109 -563 389
rect -505 109 -385 389
rect -327 109 -207 389
rect -149 109 -29 389
rect 29 109 149 389
rect 207 109 327 389
rect 385 109 505 389
rect 563 109 683 389
rect 741 109 861 389
rect 919 109 1039 389
rect 1097 109 1217 389
rect 1275 109 1395 389
rect -1395 -389 -1275 -109
rect -1217 -389 -1097 -109
rect -1039 -389 -919 -109
rect -861 -389 -741 -109
rect -683 -389 -563 -109
rect -505 -389 -385 -109
rect -327 -389 -207 -109
rect -149 -389 -29 -109
rect 29 -389 149 -109
rect 207 -389 327 -109
rect 385 -389 505 -109
rect 563 -389 683 -109
rect 741 -389 861 -109
rect 919 -389 1039 -109
rect 1097 -389 1217 -109
rect 1275 -389 1395 -109
rect -1395 -887 -1275 -607
rect -1217 -887 -1097 -607
rect -1039 -887 -919 -607
rect -861 -887 -741 -607
rect -683 -887 -563 -607
rect -505 -887 -385 -607
rect -327 -887 -207 -607
rect -149 -887 -29 -607
rect 29 -887 149 -607
rect 207 -887 327 -607
rect 385 -887 505 -607
rect 563 -887 683 -607
rect 741 -887 861 -607
rect 919 -887 1039 -607
rect 1097 -887 1217 -607
rect 1275 -887 1395 -607
<< ndiff >>
rect -1453 875 -1395 887
rect -1453 619 -1441 875
rect -1407 619 -1395 875
rect -1453 607 -1395 619
rect -1275 875 -1217 887
rect -1275 619 -1263 875
rect -1229 619 -1217 875
rect -1275 607 -1217 619
rect -1097 875 -1039 887
rect -1097 619 -1085 875
rect -1051 619 -1039 875
rect -1097 607 -1039 619
rect -919 875 -861 887
rect -919 619 -907 875
rect -873 619 -861 875
rect -919 607 -861 619
rect -741 875 -683 887
rect -741 619 -729 875
rect -695 619 -683 875
rect -741 607 -683 619
rect -563 875 -505 887
rect -563 619 -551 875
rect -517 619 -505 875
rect -563 607 -505 619
rect -385 875 -327 887
rect -385 619 -373 875
rect -339 619 -327 875
rect -385 607 -327 619
rect -207 875 -149 887
rect -207 619 -195 875
rect -161 619 -149 875
rect -207 607 -149 619
rect -29 875 29 887
rect -29 619 -17 875
rect 17 619 29 875
rect -29 607 29 619
rect 149 875 207 887
rect 149 619 161 875
rect 195 619 207 875
rect 149 607 207 619
rect 327 875 385 887
rect 327 619 339 875
rect 373 619 385 875
rect 327 607 385 619
rect 505 875 563 887
rect 505 619 517 875
rect 551 619 563 875
rect 505 607 563 619
rect 683 875 741 887
rect 683 619 695 875
rect 729 619 741 875
rect 683 607 741 619
rect 861 875 919 887
rect 861 619 873 875
rect 907 619 919 875
rect 861 607 919 619
rect 1039 875 1097 887
rect 1039 619 1051 875
rect 1085 619 1097 875
rect 1039 607 1097 619
rect 1217 875 1275 887
rect 1217 619 1229 875
rect 1263 619 1275 875
rect 1217 607 1275 619
rect 1395 875 1453 887
rect 1395 619 1407 875
rect 1441 619 1453 875
rect 1395 607 1453 619
rect -1453 377 -1395 389
rect -1453 121 -1441 377
rect -1407 121 -1395 377
rect -1453 109 -1395 121
rect -1275 377 -1217 389
rect -1275 121 -1263 377
rect -1229 121 -1217 377
rect -1275 109 -1217 121
rect -1097 377 -1039 389
rect -1097 121 -1085 377
rect -1051 121 -1039 377
rect -1097 109 -1039 121
rect -919 377 -861 389
rect -919 121 -907 377
rect -873 121 -861 377
rect -919 109 -861 121
rect -741 377 -683 389
rect -741 121 -729 377
rect -695 121 -683 377
rect -741 109 -683 121
rect -563 377 -505 389
rect -563 121 -551 377
rect -517 121 -505 377
rect -563 109 -505 121
rect -385 377 -327 389
rect -385 121 -373 377
rect -339 121 -327 377
rect -385 109 -327 121
rect -207 377 -149 389
rect -207 121 -195 377
rect -161 121 -149 377
rect -207 109 -149 121
rect -29 377 29 389
rect -29 121 -17 377
rect 17 121 29 377
rect -29 109 29 121
rect 149 377 207 389
rect 149 121 161 377
rect 195 121 207 377
rect 149 109 207 121
rect 327 377 385 389
rect 327 121 339 377
rect 373 121 385 377
rect 327 109 385 121
rect 505 377 563 389
rect 505 121 517 377
rect 551 121 563 377
rect 505 109 563 121
rect 683 377 741 389
rect 683 121 695 377
rect 729 121 741 377
rect 683 109 741 121
rect 861 377 919 389
rect 861 121 873 377
rect 907 121 919 377
rect 861 109 919 121
rect 1039 377 1097 389
rect 1039 121 1051 377
rect 1085 121 1097 377
rect 1039 109 1097 121
rect 1217 377 1275 389
rect 1217 121 1229 377
rect 1263 121 1275 377
rect 1217 109 1275 121
rect 1395 377 1453 389
rect 1395 121 1407 377
rect 1441 121 1453 377
rect 1395 109 1453 121
rect -1453 -121 -1395 -109
rect -1453 -377 -1441 -121
rect -1407 -377 -1395 -121
rect -1453 -389 -1395 -377
rect -1275 -121 -1217 -109
rect -1275 -377 -1263 -121
rect -1229 -377 -1217 -121
rect -1275 -389 -1217 -377
rect -1097 -121 -1039 -109
rect -1097 -377 -1085 -121
rect -1051 -377 -1039 -121
rect -1097 -389 -1039 -377
rect -919 -121 -861 -109
rect -919 -377 -907 -121
rect -873 -377 -861 -121
rect -919 -389 -861 -377
rect -741 -121 -683 -109
rect -741 -377 -729 -121
rect -695 -377 -683 -121
rect -741 -389 -683 -377
rect -563 -121 -505 -109
rect -563 -377 -551 -121
rect -517 -377 -505 -121
rect -563 -389 -505 -377
rect -385 -121 -327 -109
rect -385 -377 -373 -121
rect -339 -377 -327 -121
rect -385 -389 -327 -377
rect -207 -121 -149 -109
rect -207 -377 -195 -121
rect -161 -377 -149 -121
rect -207 -389 -149 -377
rect -29 -121 29 -109
rect -29 -377 -17 -121
rect 17 -377 29 -121
rect -29 -389 29 -377
rect 149 -121 207 -109
rect 149 -377 161 -121
rect 195 -377 207 -121
rect 149 -389 207 -377
rect 327 -121 385 -109
rect 327 -377 339 -121
rect 373 -377 385 -121
rect 327 -389 385 -377
rect 505 -121 563 -109
rect 505 -377 517 -121
rect 551 -377 563 -121
rect 505 -389 563 -377
rect 683 -121 741 -109
rect 683 -377 695 -121
rect 729 -377 741 -121
rect 683 -389 741 -377
rect 861 -121 919 -109
rect 861 -377 873 -121
rect 907 -377 919 -121
rect 861 -389 919 -377
rect 1039 -121 1097 -109
rect 1039 -377 1051 -121
rect 1085 -377 1097 -121
rect 1039 -389 1097 -377
rect 1217 -121 1275 -109
rect 1217 -377 1229 -121
rect 1263 -377 1275 -121
rect 1217 -389 1275 -377
rect 1395 -121 1453 -109
rect 1395 -377 1407 -121
rect 1441 -377 1453 -121
rect 1395 -389 1453 -377
rect -1453 -619 -1395 -607
rect -1453 -875 -1441 -619
rect -1407 -875 -1395 -619
rect -1453 -887 -1395 -875
rect -1275 -619 -1217 -607
rect -1275 -875 -1263 -619
rect -1229 -875 -1217 -619
rect -1275 -887 -1217 -875
rect -1097 -619 -1039 -607
rect -1097 -875 -1085 -619
rect -1051 -875 -1039 -619
rect -1097 -887 -1039 -875
rect -919 -619 -861 -607
rect -919 -875 -907 -619
rect -873 -875 -861 -619
rect -919 -887 -861 -875
rect -741 -619 -683 -607
rect -741 -875 -729 -619
rect -695 -875 -683 -619
rect -741 -887 -683 -875
rect -563 -619 -505 -607
rect -563 -875 -551 -619
rect -517 -875 -505 -619
rect -563 -887 -505 -875
rect -385 -619 -327 -607
rect -385 -875 -373 -619
rect -339 -875 -327 -619
rect -385 -887 -327 -875
rect -207 -619 -149 -607
rect -207 -875 -195 -619
rect -161 -875 -149 -619
rect -207 -887 -149 -875
rect -29 -619 29 -607
rect -29 -875 -17 -619
rect 17 -875 29 -619
rect -29 -887 29 -875
rect 149 -619 207 -607
rect 149 -875 161 -619
rect 195 -875 207 -619
rect 149 -887 207 -875
rect 327 -619 385 -607
rect 327 -875 339 -619
rect 373 -875 385 -619
rect 327 -887 385 -875
rect 505 -619 563 -607
rect 505 -875 517 -619
rect 551 -875 563 -619
rect 505 -887 563 -875
rect 683 -619 741 -607
rect 683 -875 695 -619
rect 729 -875 741 -619
rect 683 -887 741 -875
rect 861 -619 919 -607
rect 861 -875 873 -619
rect 907 -875 919 -619
rect 861 -887 919 -875
rect 1039 -619 1097 -607
rect 1039 -875 1051 -619
rect 1085 -875 1097 -619
rect 1039 -887 1097 -875
rect 1217 -619 1275 -607
rect 1217 -875 1229 -619
rect 1263 -875 1275 -619
rect 1217 -887 1275 -875
rect 1395 -619 1453 -607
rect 1395 -875 1407 -619
rect 1441 -875 1453 -619
rect 1395 -887 1453 -875
<< ndiffc >>
rect -1441 619 -1407 875
rect -1263 619 -1229 875
rect -1085 619 -1051 875
rect -907 619 -873 875
rect -729 619 -695 875
rect -551 619 -517 875
rect -373 619 -339 875
rect -195 619 -161 875
rect -17 619 17 875
rect 161 619 195 875
rect 339 619 373 875
rect 517 619 551 875
rect 695 619 729 875
rect 873 619 907 875
rect 1051 619 1085 875
rect 1229 619 1263 875
rect 1407 619 1441 875
rect -1441 121 -1407 377
rect -1263 121 -1229 377
rect -1085 121 -1051 377
rect -907 121 -873 377
rect -729 121 -695 377
rect -551 121 -517 377
rect -373 121 -339 377
rect -195 121 -161 377
rect -17 121 17 377
rect 161 121 195 377
rect 339 121 373 377
rect 517 121 551 377
rect 695 121 729 377
rect 873 121 907 377
rect 1051 121 1085 377
rect 1229 121 1263 377
rect 1407 121 1441 377
rect -1441 -377 -1407 -121
rect -1263 -377 -1229 -121
rect -1085 -377 -1051 -121
rect -907 -377 -873 -121
rect -729 -377 -695 -121
rect -551 -377 -517 -121
rect -373 -377 -339 -121
rect -195 -377 -161 -121
rect -17 -377 17 -121
rect 161 -377 195 -121
rect 339 -377 373 -121
rect 517 -377 551 -121
rect 695 -377 729 -121
rect 873 -377 907 -121
rect 1051 -377 1085 -121
rect 1229 -377 1263 -121
rect 1407 -377 1441 -121
rect -1441 -875 -1407 -619
rect -1263 -875 -1229 -619
rect -1085 -875 -1051 -619
rect -907 -875 -873 -619
rect -729 -875 -695 -619
rect -551 -875 -517 -619
rect -373 -875 -339 -619
rect -195 -875 -161 -619
rect -17 -875 17 -619
rect 161 -875 195 -619
rect 339 -875 373 -619
rect 517 -875 551 -619
rect 695 -875 729 -619
rect 873 -875 907 -619
rect 1051 -875 1085 -619
rect 1229 -875 1263 -619
rect 1407 -875 1441 -619
<< psubdiff >>
rect -1555 1027 -1459 1061
rect 1459 1027 1555 1061
rect -1555 965 -1521 1027
rect 1521 965 1555 1027
rect -1555 -1027 -1521 -965
rect 1521 -1027 1555 -965
rect -1555 -1061 -1459 -1027
rect 1459 -1061 1555 -1027
<< psubdiffcont >>
rect -1459 1027 1459 1061
rect -1555 -965 -1521 965
rect 1521 -965 1555 965
rect -1459 -1061 1459 -1027
<< poly >>
rect -1377 959 -1293 975
rect -1377 942 -1361 959
rect -1395 925 -1361 942
rect -1309 942 -1293 959
rect -1199 959 -1115 975
rect -1199 942 -1183 959
rect -1309 925 -1275 942
rect -1395 887 -1275 925
rect -1217 925 -1183 942
rect -1131 942 -1115 959
rect -1021 959 -937 975
rect -1021 942 -1005 959
rect -1131 925 -1097 942
rect -1217 887 -1097 925
rect -1039 925 -1005 942
rect -953 942 -937 959
rect -843 959 -759 975
rect -843 942 -827 959
rect -953 925 -919 942
rect -1039 887 -919 925
rect -861 925 -827 942
rect -775 942 -759 959
rect -665 959 -581 975
rect -665 942 -649 959
rect -775 925 -741 942
rect -861 887 -741 925
rect -683 925 -649 942
rect -597 942 -581 959
rect -487 959 -403 975
rect -487 942 -471 959
rect -597 925 -563 942
rect -683 887 -563 925
rect -505 925 -471 942
rect -419 942 -403 959
rect -309 959 -225 975
rect -309 942 -293 959
rect -419 925 -385 942
rect -505 887 -385 925
rect -327 925 -293 942
rect -241 942 -225 959
rect -131 959 -47 975
rect -131 942 -115 959
rect -241 925 -207 942
rect -327 887 -207 925
rect -149 925 -115 942
rect -63 942 -47 959
rect 47 959 131 975
rect 47 942 63 959
rect -63 925 -29 942
rect -149 887 -29 925
rect 29 925 63 942
rect 115 942 131 959
rect 225 959 309 975
rect 225 942 241 959
rect 115 925 149 942
rect 29 887 149 925
rect 207 925 241 942
rect 293 942 309 959
rect 403 959 487 975
rect 403 942 419 959
rect 293 925 327 942
rect 207 887 327 925
rect 385 925 419 942
rect 471 942 487 959
rect 581 959 665 975
rect 581 942 597 959
rect 471 925 505 942
rect 385 887 505 925
rect 563 925 597 942
rect 649 942 665 959
rect 759 959 843 975
rect 759 942 775 959
rect 649 925 683 942
rect 563 887 683 925
rect 741 925 775 942
rect 827 942 843 959
rect 937 959 1021 975
rect 937 942 953 959
rect 827 925 861 942
rect 741 887 861 925
rect 919 925 953 942
rect 1005 942 1021 959
rect 1115 959 1199 975
rect 1115 942 1131 959
rect 1005 925 1039 942
rect 919 887 1039 925
rect 1097 925 1131 942
rect 1183 942 1199 959
rect 1293 959 1377 975
rect 1293 942 1309 959
rect 1183 925 1217 942
rect 1097 887 1217 925
rect 1275 925 1309 942
rect 1361 942 1377 959
rect 1361 925 1395 942
rect 1275 887 1395 925
rect -1395 569 -1275 607
rect -1395 552 -1361 569
rect -1377 535 -1361 552
rect -1309 552 -1275 569
rect -1217 569 -1097 607
rect -1217 552 -1183 569
rect -1309 535 -1293 552
rect -1377 519 -1293 535
rect -1199 535 -1183 552
rect -1131 552 -1097 569
rect -1039 569 -919 607
rect -1039 552 -1005 569
rect -1131 535 -1115 552
rect -1199 519 -1115 535
rect -1021 535 -1005 552
rect -953 552 -919 569
rect -861 569 -741 607
rect -861 552 -827 569
rect -953 535 -937 552
rect -1021 519 -937 535
rect -843 535 -827 552
rect -775 552 -741 569
rect -683 569 -563 607
rect -683 552 -649 569
rect -775 535 -759 552
rect -843 519 -759 535
rect -665 535 -649 552
rect -597 552 -563 569
rect -505 569 -385 607
rect -505 552 -471 569
rect -597 535 -581 552
rect -665 519 -581 535
rect -487 535 -471 552
rect -419 552 -385 569
rect -327 569 -207 607
rect -327 552 -293 569
rect -419 535 -403 552
rect -487 519 -403 535
rect -309 535 -293 552
rect -241 552 -207 569
rect -149 569 -29 607
rect -149 552 -115 569
rect -241 535 -225 552
rect -309 519 -225 535
rect -131 535 -115 552
rect -63 552 -29 569
rect 29 569 149 607
rect 29 552 63 569
rect -63 535 -47 552
rect -131 519 -47 535
rect 47 535 63 552
rect 115 552 149 569
rect 207 569 327 607
rect 207 552 241 569
rect 115 535 131 552
rect 47 519 131 535
rect 225 535 241 552
rect 293 552 327 569
rect 385 569 505 607
rect 385 552 419 569
rect 293 535 309 552
rect 225 519 309 535
rect 403 535 419 552
rect 471 552 505 569
rect 563 569 683 607
rect 563 552 597 569
rect 471 535 487 552
rect 403 519 487 535
rect 581 535 597 552
rect 649 552 683 569
rect 741 569 861 607
rect 741 552 775 569
rect 649 535 665 552
rect 581 519 665 535
rect 759 535 775 552
rect 827 552 861 569
rect 919 569 1039 607
rect 919 552 953 569
rect 827 535 843 552
rect 759 519 843 535
rect 937 535 953 552
rect 1005 552 1039 569
rect 1097 569 1217 607
rect 1097 552 1131 569
rect 1005 535 1021 552
rect 937 519 1021 535
rect 1115 535 1131 552
rect 1183 552 1217 569
rect 1275 569 1395 607
rect 1275 552 1309 569
rect 1183 535 1199 552
rect 1115 519 1199 535
rect 1293 535 1309 552
rect 1361 552 1395 569
rect 1361 535 1377 552
rect 1293 519 1377 535
rect -1377 461 -1293 477
rect -1377 444 -1361 461
rect -1395 427 -1361 444
rect -1309 444 -1293 461
rect -1199 461 -1115 477
rect -1199 444 -1183 461
rect -1309 427 -1275 444
rect -1395 389 -1275 427
rect -1217 427 -1183 444
rect -1131 444 -1115 461
rect -1021 461 -937 477
rect -1021 444 -1005 461
rect -1131 427 -1097 444
rect -1217 389 -1097 427
rect -1039 427 -1005 444
rect -953 444 -937 461
rect -843 461 -759 477
rect -843 444 -827 461
rect -953 427 -919 444
rect -1039 389 -919 427
rect -861 427 -827 444
rect -775 444 -759 461
rect -665 461 -581 477
rect -665 444 -649 461
rect -775 427 -741 444
rect -861 389 -741 427
rect -683 427 -649 444
rect -597 444 -581 461
rect -487 461 -403 477
rect -487 444 -471 461
rect -597 427 -563 444
rect -683 389 -563 427
rect -505 427 -471 444
rect -419 444 -403 461
rect -309 461 -225 477
rect -309 444 -293 461
rect -419 427 -385 444
rect -505 389 -385 427
rect -327 427 -293 444
rect -241 444 -225 461
rect -131 461 -47 477
rect -131 444 -115 461
rect -241 427 -207 444
rect -327 389 -207 427
rect -149 427 -115 444
rect -63 444 -47 461
rect 47 461 131 477
rect 47 444 63 461
rect -63 427 -29 444
rect -149 389 -29 427
rect 29 427 63 444
rect 115 444 131 461
rect 225 461 309 477
rect 225 444 241 461
rect 115 427 149 444
rect 29 389 149 427
rect 207 427 241 444
rect 293 444 309 461
rect 403 461 487 477
rect 403 444 419 461
rect 293 427 327 444
rect 207 389 327 427
rect 385 427 419 444
rect 471 444 487 461
rect 581 461 665 477
rect 581 444 597 461
rect 471 427 505 444
rect 385 389 505 427
rect 563 427 597 444
rect 649 444 665 461
rect 759 461 843 477
rect 759 444 775 461
rect 649 427 683 444
rect 563 389 683 427
rect 741 427 775 444
rect 827 444 843 461
rect 937 461 1021 477
rect 937 444 953 461
rect 827 427 861 444
rect 741 389 861 427
rect 919 427 953 444
rect 1005 444 1021 461
rect 1115 461 1199 477
rect 1115 444 1131 461
rect 1005 427 1039 444
rect 919 389 1039 427
rect 1097 427 1131 444
rect 1183 444 1199 461
rect 1293 461 1377 477
rect 1293 444 1309 461
rect 1183 427 1217 444
rect 1097 389 1217 427
rect 1275 427 1309 444
rect 1361 444 1377 461
rect 1361 427 1395 444
rect 1275 389 1395 427
rect -1395 71 -1275 109
rect -1395 54 -1361 71
rect -1377 37 -1361 54
rect -1309 54 -1275 71
rect -1217 71 -1097 109
rect -1217 54 -1183 71
rect -1309 37 -1293 54
rect -1377 21 -1293 37
rect -1199 37 -1183 54
rect -1131 54 -1097 71
rect -1039 71 -919 109
rect -1039 54 -1005 71
rect -1131 37 -1115 54
rect -1199 21 -1115 37
rect -1021 37 -1005 54
rect -953 54 -919 71
rect -861 71 -741 109
rect -861 54 -827 71
rect -953 37 -937 54
rect -1021 21 -937 37
rect -843 37 -827 54
rect -775 54 -741 71
rect -683 71 -563 109
rect -683 54 -649 71
rect -775 37 -759 54
rect -843 21 -759 37
rect -665 37 -649 54
rect -597 54 -563 71
rect -505 71 -385 109
rect -505 54 -471 71
rect -597 37 -581 54
rect -665 21 -581 37
rect -487 37 -471 54
rect -419 54 -385 71
rect -327 71 -207 109
rect -327 54 -293 71
rect -419 37 -403 54
rect -487 21 -403 37
rect -309 37 -293 54
rect -241 54 -207 71
rect -149 71 -29 109
rect -149 54 -115 71
rect -241 37 -225 54
rect -309 21 -225 37
rect -131 37 -115 54
rect -63 54 -29 71
rect 29 71 149 109
rect 29 54 63 71
rect -63 37 -47 54
rect -131 21 -47 37
rect 47 37 63 54
rect 115 54 149 71
rect 207 71 327 109
rect 207 54 241 71
rect 115 37 131 54
rect 47 21 131 37
rect 225 37 241 54
rect 293 54 327 71
rect 385 71 505 109
rect 385 54 419 71
rect 293 37 309 54
rect 225 21 309 37
rect 403 37 419 54
rect 471 54 505 71
rect 563 71 683 109
rect 563 54 597 71
rect 471 37 487 54
rect 403 21 487 37
rect 581 37 597 54
rect 649 54 683 71
rect 741 71 861 109
rect 741 54 775 71
rect 649 37 665 54
rect 581 21 665 37
rect 759 37 775 54
rect 827 54 861 71
rect 919 71 1039 109
rect 919 54 953 71
rect 827 37 843 54
rect 759 21 843 37
rect 937 37 953 54
rect 1005 54 1039 71
rect 1097 71 1217 109
rect 1097 54 1131 71
rect 1005 37 1021 54
rect 937 21 1021 37
rect 1115 37 1131 54
rect 1183 54 1217 71
rect 1275 71 1395 109
rect 1275 54 1309 71
rect 1183 37 1199 54
rect 1115 21 1199 37
rect 1293 37 1309 54
rect 1361 54 1395 71
rect 1361 37 1377 54
rect 1293 21 1377 37
rect -1377 -37 -1293 -21
rect -1377 -54 -1361 -37
rect -1395 -71 -1361 -54
rect -1309 -54 -1293 -37
rect -1199 -37 -1115 -21
rect -1199 -54 -1183 -37
rect -1309 -71 -1275 -54
rect -1395 -109 -1275 -71
rect -1217 -71 -1183 -54
rect -1131 -54 -1115 -37
rect -1021 -37 -937 -21
rect -1021 -54 -1005 -37
rect -1131 -71 -1097 -54
rect -1217 -109 -1097 -71
rect -1039 -71 -1005 -54
rect -953 -54 -937 -37
rect -843 -37 -759 -21
rect -843 -54 -827 -37
rect -953 -71 -919 -54
rect -1039 -109 -919 -71
rect -861 -71 -827 -54
rect -775 -54 -759 -37
rect -665 -37 -581 -21
rect -665 -54 -649 -37
rect -775 -71 -741 -54
rect -861 -109 -741 -71
rect -683 -71 -649 -54
rect -597 -54 -581 -37
rect -487 -37 -403 -21
rect -487 -54 -471 -37
rect -597 -71 -563 -54
rect -683 -109 -563 -71
rect -505 -71 -471 -54
rect -419 -54 -403 -37
rect -309 -37 -225 -21
rect -309 -54 -293 -37
rect -419 -71 -385 -54
rect -505 -109 -385 -71
rect -327 -71 -293 -54
rect -241 -54 -225 -37
rect -131 -37 -47 -21
rect -131 -54 -115 -37
rect -241 -71 -207 -54
rect -327 -109 -207 -71
rect -149 -71 -115 -54
rect -63 -54 -47 -37
rect 47 -37 131 -21
rect 47 -54 63 -37
rect -63 -71 -29 -54
rect -149 -109 -29 -71
rect 29 -71 63 -54
rect 115 -54 131 -37
rect 225 -37 309 -21
rect 225 -54 241 -37
rect 115 -71 149 -54
rect 29 -109 149 -71
rect 207 -71 241 -54
rect 293 -54 309 -37
rect 403 -37 487 -21
rect 403 -54 419 -37
rect 293 -71 327 -54
rect 207 -109 327 -71
rect 385 -71 419 -54
rect 471 -54 487 -37
rect 581 -37 665 -21
rect 581 -54 597 -37
rect 471 -71 505 -54
rect 385 -109 505 -71
rect 563 -71 597 -54
rect 649 -54 665 -37
rect 759 -37 843 -21
rect 759 -54 775 -37
rect 649 -71 683 -54
rect 563 -109 683 -71
rect 741 -71 775 -54
rect 827 -54 843 -37
rect 937 -37 1021 -21
rect 937 -54 953 -37
rect 827 -71 861 -54
rect 741 -109 861 -71
rect 919 -71 953 -54
rect 1005 -54 1021 -37
rect 1115 -37 1199 -21
rect 1115 -54 1131 -37
rect 1005 -71 1039 -54
rect 919 -109 1039 -71
rect 1097 -71 1131 -54
rect 1183 -54 1199 -37
rect 1293 -37 1377 -21
rect 1293 -54 1309 -37
rect 1183 -71 1217 -54
rect 1097 -109 1217 -71
rect 1275 -71 1309 -54
rect 1361 -54 1377 -37
rect 1361 -71 1395 -54
rect 1275 -109 1395 -71
rect -1395 -427 -1275 -389
rect -1395 -444 -1361 -427
rect -1377 -461 -1361 -444
rect -1309 -444 -1275 -427
rect -1217 -427 -1097 -389
rect -1217 -444 -1183 -427
rect -1309 -461 -1293 -444
rect -1377 -477 -1293 -461
rect -1199 -461 -1183 -444
rect -1131 -444 -1097 -427
rect -1039 -427 -919 -389
rect -1039 -444 -1005 -427
rect -1131 -461 -1115 -444
rect -1199 -477 -1115 -461
rect -1021 -461 -1005 -444
rect -953 -444 -919 -427
rect -861 -427 -741 -389
rect -861 -444 -827 -427
rect -953 -461 -937 -444
rect -1021 -477 -937 -461
rect -843 -461 -827 -444
rect -775 -444 -741 -427
rect -683 -427 -563 -389
rect -683 -444 -649 -427
rect -775 -461 -759 -444
rect -843 -477 -759 -461
rect -665 -461 -649 -444
rect -597 -444 -563 -427
rect -505 -427 -385 -389
rect -505 -444 -471 -427
rect -597 -461 -581 -444
rect -665 -477 -581 -461
rect -487 -461 -471 -444
rect -419 -444 -385 -427
rect -327 -427 -207 -389
rect -327 -444 -293 -427
rect -419 -461 -403 -444
rect -487 -477 -403 -461
rect -309 -461 -293 -444
rect -241 -444 -207 -427
rect -149 -427 -29 -389
rect -149 -444 -115 -427
rect -241 -461 -225 -444
rect -309 -477 -225 -461
rect -131 -461 -115 -444
rect -63 -444 -29 -427
rect 29 -427 149 -389
rect 29 -444 63 -427
rect -63 -461 -47 -444
rect -131 -477 -47 -461
rect 47 -461 63 -444
rect 115 -444 149 -427
rect 207 -427 327 -389
rect 207 -444 241 -427
rect 115 -461 131 -444
rect 47 -477 131 -461
rect 225 -461 241 -444
rect 293 -444 327 -427
rect 385 -427 505 -389
rect 385 -444 419 -427
rect 293 -461 309 -444
rect 225 -477 309 -461
rect 403 -461 419 -444
rect 471 -444 505 -427
rect 563 -427 683 -389
rect 563 -444 597 -427
rect 471 -461 487 -444
rect 403 -477 487 -461
rect 581 -461 597 -444
rect 649 -444 683 -427
rect 741 -427 861 -389
rect 741 -444 775 -427
rect 649 -461 665 -444
rect 581 -477 665 -461
rect 759 -461 775 -444
rect 827 -444 861 -427
rect 919 -427 1039 -389
rect 919 -444 953 -427
rect 827 -461 843 -444
rect 759 -477 843 -461
rect 937 -461 953 -444
rect 1005 -444 1039 -427
rect 1097 -427 1217 -389
rect 1097 -444 1131 -427
rect 1005 -461 1021 -444
rect 937 -477 1021 -461
rect 1115 -461 1131 -444
rect 1183 -444 1217 -427
rect 1275 -427 1395 -389
rect 1275 -444 1309 -427
rect 1183 -461 1199 -444
rect 1115 -477 1199 -461
rect 1293 -461 1309 -444
rect 1361 -444 1395 -427
rect 1361 -461 1377 -444
rect 1293 -477 1377 -461
rect -1377 -535 -1293 -519
rect -1377 -552 -1361 -535
rect -1395 -569 -1361 -552
rect -1309 -552 -1293 -535
rect -1199 -535 -1115 -519
rect -1199 -552 -1183 -535
rect -1309 -569 -1275 -552
rect -1395 -607 -1275 -569
rect -1217 -569 -1183 -552
rect -1131 -552 -1115 -535
rect -1021 -535 -937 -519
rect -1021 -552 -1005 -535
rect -1131 -569 -1097 -552
rect -1217 -607 -1097 -569
rect -1039 -569 -1005 -552
rect -953 -552 -937 -535
rect -843 -535 -759 -519
rect -843 -552 -827 -535
rect -953 -569 -919 -552
rect -1039 -607 -919 -569
rect -861 -569 -827 -552
rect -775 -552 -759 -535
rect -665 -535 -581 -519
rect -665 -552 -649 -535
rect -775 -569 -741 -552
rect -861 -607 -741 -569
rect -683 -569 -649 -552
rect -597 -552 -581 -535
rect -487 -535 -403 -519
rect -487 -552 -471 -535
rect -597 -569 -563 -552
rect -683 -607 -563 -569
rect -505 -569 -471 -552
rect -419 -552 -403 -535
rect -309 -535 -225 -519
rect -309 -552 -293 -535
rect -419 -569 -385 -552
rect -505 -607 -385 -569
rect -327 -569 -293 -552
rect -241 -552 -225 -535
rect -131 -535 -47 -519
rect -131 -552 -115 -535
rect -241 -569 -207 -552
rect -327 -607 -207 -569
rect -149 -569 -115 -552
rect -63 -552 -47 -535
rect 47 -535 131 -519
rect 47 -552 63 -535
rect -63 -569 -29 -552
rect -149 -607 -29 -569
rect 29 -569 63 -552
rect 115 -552 131 -535
rect 225 -535 309 -519
rect 225 -552 241 -535
rect 115 -569 149 -552
rect 29 -607 149 -569
rect 207 -569 241 -552
rect 293 -552 309 -535
rect 403 -535 487 -519
rect 403 -552 419 -535
rect 293 -569 327 -552
rect 207 -607 327 -569
rect 385 -569 419 -552
rect 471 -552 487 -535
rect 581 -535 665 -519
rect 581 -552 597 -535
rect 471 -569 505 -552
rect 385 -607 505 -569
rect 563 -569 597 -552
rect 649 -552 665 -535
rect 759 -535 843 -519
rect 759 -552 775 -535
rect 649 -569 683 -552
rect 563 -607 683 -569
rect 741 -569 775 -552
rect 827 -552 843 -535
rect 937 -535 1021 -519
rect 937 -552 953 -535
rect 827 -569 861 -552
rect 741 -607 861 -569
rect 919 -569 953 -552
rect 1005 -552 1021 -535
rect 1115 -535 1199 -519
rect 1115 -552 1131 -535
rect 1005 -569 1039 -552
rect 919 -607 1039 -569
rect 1097 -569 1131 -552
rect 1183 -552 1199 -535
rect 1293 -535 1377 -519
rect 1293 -552 1309 -535
rect 1183 -569 1217 -552
rect 1097 -607 1217 -569
rect 1275 -569 1309 -552
rect 1361 -552 1377 -535
rect 1361 -569 1395 -552
rect 1275 -607 1395 -569
rect -1395 -925 -1275 -887
rect -1395 -942 -1361 -925
rect -1377 -959 -1361 -942
rect -1309 -942 -1275 -925
rect -1217 -925 -1097 -887
rect -1217 -942 -1183 -925
rect -1309 -959 -1293 -942
rect -1377 -975 -1293 -959
rect -1199 -959 -1183 -942
rect -1131 -942 -1097 -925
rect -1039 -925 -919 -887
rect -1039 -942 -1005 -925
rect -1131 -959 -1115 -942
rect -1199 -975 -1115 -959
rect -1021 -959 -1005 -942
rect -953 -942 -919 -925
rect -861 -925 -741 -887
rect -861 -942 -827 -925
rect -953 -959 -937 -942
rect -1021 -975 -937 -959
rect -843 -959 -827 -942
rect -775 -942 -741 -925
rect -683 -925 -563 -887
rect -683 -942 -649 -925
rect -775 -959 -759 -942
rect -843 -975 -759 -959
rect -665 -959 -649 -942
rect -597 -942 -563 -925
rect -505 -925 -385 -887
rect -505 -942 -471 -925
rect -597 -959 -581 -942
rect -665 -975 -581 -959
rect -487 -959 -471 -942
rect -419 -942 -385 -925
rect -327 -925 -207 -887
rect -327 -942 -293 -925
rect -419 -959 -403 -942
rect -487 -975 -403 -959
rect -309 -959 -293 -942
rect -241 -942 -207 -925
rect -149 -925 -29 -887
rect -149 -942 -115 -925
rect -241 -959 -225 -942
rect -309 -975 -225 -959
rect -131 -959 -115 -942
rect -63 -942 -29 -925
rect 29 -925 149 -887
rect 29 -942 63 -925
rect -63 -959 -47 -942
rect -131 -975 -47 -959
rect 47 -959 63 -942
rect 115 -942 149 -925
rect 207 -925 327 -887
rect 207 -942 241 -925
rect 115 -959 131 -942
rect 47 -975 131 -959
rect 225 -959 241 -942
rect 293 -942 327 -925
rect 385 -925 505 -887
rect 385 -942 419 -925
rect 293 -959 309 -942
rect 225 -975 309 -959
rect 403 -959 419 -942
rect 471 -942 505 -925
rect 563 -925 683 -887
rect 563 -942 597 -925
rect 471 -959 487 -942
rect 403 -975 487 -959
rect 581 -959 597 -942
rect 649 -942 683 -925
rect 741 -925 861 -887
rect 741 -942 775 -925
rect 649 -959 665 -942
rect 581 -975 665 -959
rect 759 -959 775 -942
rect 827 -942 861 -925
rect 919 -925 1039 -887
rect 919 -942 953 -925
rect 827 -959 843 -942
rect 759 -975 843 -959
rect 937 -959 953 -942
rect 1005 -942 1039 -925
rect 1097 -925 1217 -887
rect 1097 -942 1131 -925
rect 1005 -959 1021 -942
rect 937 -975 1021 -959
rect 1115 -959 1131 -942
rect 1183 -942 1217 -925
rect 1275 -925 1395 -887
rect 1275 -942 1309 -925
rect 1183 -959 1199 -942
rect 1115 -975 1199 -959
rect 1293 -959 1309 -942
rect 1361 -942 1395 -925
rect 1361 -959 1377 -942
rect 1293 -975 1377 -959
<< polycont >>
rect -1361 925 -1309 959
rect -1183 925 -1131 959
rect -1005 925 -953 959
rect -827 925 -775 959
rect -649 925 -597 959
rect -471 925 -419 959
rect -293 925 -241 959
rect -115 925 -63 959
rect 63 925 115 959
rect 241 925 293 959
rect 419 925 471 959
rect 597 925 649 959
rect 775 925 827 959
rect 953 925 1005 959
rect 1131 925 1183 959
rect 1309 925 1361 959
rect -1361 535 -1309 569
rect -1183 535 -1131 569
rect -1005 535 -953 569
rect -827 535 -775 569
rect -649 535 -597 569
rect -471 535 -419 569
rect -293 535 -241 569
rect -115 535 -63 569
rect 63 535 115 569
rect 241 535 293 569
rect 419 535 471 569
rect 597 535 649 569
rect 775 535 827 569
rect 953 535 1005 569
rect 1131 535 1183 569
rect 1309 535 1361 569
rect -1361 427 -1309 461
rect -1183 427 -1131 461
rect -1005 427 -953 461
rect -827 427 -775 461
rect -649 427 -597 461
rect -471 427 -419 461
rect -293 427 -241 461
rect -115 427 -63 461
rect 63 427 115 461
rect 241 427 293 461
rect 419 427 471 461
rect 597 427 649 461
rect 775 427 827 461
rect 953 427 1005 461
rect 1131 427 1183 461
rect 1309 427 1361 461
rect -1361 37 -1309 71
rect -1183 37 -1131 71
rect -1005 37 -953 71
rect -827 37 -775 71
rect -649 37 -597 71
rect -471 37 -419 71
rect -293 37 -241 71
rect -115 37 -63 71
rect 63 37 115 71
rect 241 37 293 71
rect 419 37 471 71
rect 597 37 649 71
rect 775 37 827 71
rect 953 37 1005 71
rect 1131 37 1183 71
rect 1309 37 1361 71
rect -1361 -71 -1309 -37
rect -1183 -71 -1131 -37
rect -1005 -71 -953 -37
rect -827 -71 -775 -37
rect -649 -71 -597 -37
rect -471 -71 -419 -37
rect -293 -71 -241 -37
rect -115 -71 -63 -37
rect 63 -71 115 -37
rect 241 -71 293 -37
rect 419 -71 471 -37
rect 597 -71 649 -37
rect 775 -71 827 -37
rect 953 -71 1005 -37
rect 1131 -71 1183 -37
rect 1309 -71 1361 -37
rect -1361 -461 -1309 -427
rect -1183 -461 -1131 -427
rect -1005 -461 -953 -427
rect -827 -461 -775 -427
rect -649 -461 -597 -427
rect -471 -461 -419 -427
rect -293 -461 -241 -427
rect -115 -461 -63 -427
rect 63 -461 115 -427
rect 241 -461 293 -427
rect 419 -461 471 -427
rect 597 -461 649 -427
rect 775 -461 827 -427
rect 953 -461 1005 -427
rect 1131 -461 1183 -427
rect 1309 -461 1361 -427
rect -1361 -569 -1309 -535
rect -1183 -569 -1131 -535
rect -1005 -569 -953 -535
rect -827 -569 -775 -535
rect -649 -569 -597 -535
rect -471 -569 -419 -535
rect -293 -569 -241 -535
rect -115 -569 -63 -535
rect 63 -569 115 -535
rect 241 -569 293 -535
rect 419 -569 471 -535
rect 597 -569 649 -535
rect 775 -569 827 -535
rect 953 -569 1005 -535
rect 1131 -569 1183 -535
rect 1309 -569 1361 -535
rect -1361 -959 -1309 -925
rect -1183 -959 -1131 -925
rect -1005 -959 -953 -925
rect -827 -959 -775 -925
rect -649 -959 -597 -925
rect -471 -959 -419 -925
rect -293 -959 -241 -925
rect -115 -959 -63 -925
rect 63 -959 115 -925
rect 241 -959 293 -925
rect 419 -959 471 -925
rect 597 -959 649 -925
rect 775 -959 827 -925
rect 953 -959 1005 -925
rect 1131 -959 1183 -925
rect 1309 -959 1361 -925
<< locali >>
rect -1555 1027 -1459 1061
rect 1459 1027 1555 1061
rect -1555 965 -1521 1027
rect 1521 965 1555 1027
rect -1521 925 -1361 959
rect -1309 925 -1293 959
rect -1199 925 -1183 959
rect -1131 925 -1115 959
rect -1021 925 -1005 959
rect -953 925 -937 959
rect -843 925 -827 959
rect -775 925 -759 959
rect -665 925 -649 959
rect -597 925 -581 959
rect -487 925 -471 959
rect -419 925 -403 959
rect -309 925 -293 959
rect -241 925 -225 959
rect -131 925 -115 959
rect -63 925 -47 959
rect 47 925 63 959
rect 115 925 131 959
rect 225 925 241 959
rect 293 925 309 959
rect 403 925 419 959
rect 471 925 487 959
rect 581 925 597 959
rect 649 925 665 959
rect 759 925 775 959
rect 827 925 843 959
rect 937 925 953 959
rect 1005 925 1021 959
rect 1115 925 1131 959
rect 1183 925 1199 959
rect 1293 925 1309 959
rect 1361 925 1521 959
rect -1441 875 -1407 925
rect -1441 569 -1407 619
rect -1263 875 -1229 891
rect -1263 603 -1229 619
rect -1085 875 -1051 891
rect -1085 603 -1051 619
rect -907 875 -873 891
rect -907 603 -873 619
rect -729 875 -695 891
rect -729 603 -695 619
rect -551 875 -517 891
rect -551 603 -517 619
rect -373 875 -339 891
rect -373 603 -339 619
rect -195 875 -161 891
rect -195 603 -161 619
rect -17 875 17 891
rect -17 603 17 619
rect 161 875 195 891
rect 161 603 195 619
rect 339 875 373 891
rect 339 603 373 619
rect 517 875 551 891
rect 517 603 551 619
rect 695 875 729 891
rect 695 603 729 619
rect 873 875 907 891
rect 873 603 907 619
rect 1051 875 1085 891
rect 1051 603 1085 619
rect 1229 875 1263 891
rect 1229 603 1263 619
rect 1407 875 1441 925
rect 1407 569 1441 619
rect -1521 535 -1361 569
rect -1309 535 -1293 569
rect -1199 535 -1183 569
rect -1131 535 -1115 569
rect -1021 535 -1005 569
rect -953 535 -937 569
rect -843 535 -827 569
rect -775 535 -759 569
rect -665 535 -649 569
rect -597 535 -581 569
rect -487 535 -471 569
rect -419 535 -403 569
rect -309 535 -293 569
rect -241 535 -225 569
rect -131 535 -115 569
rect -63 535 -47 569
rect 47 535 63 569
rect 115 535 131 569
rect 225 535 241 569
rect 293 535 309 569
rect 403 535 419 569
rect 471 535 487 569
rect 581 535 597 569
rect 649 535 665 569
rect 759 535 775 569
rect 827 535 843 569
rect 937 535 953 569
rect 1005 535 1021 569
rect 1115 535 1131 569
rect 1183 535 1199 569
rect 1293 535 1309 569
rect 1361 535 1521 569
rect -1521 427 -1361 461
rect -1309 427 -1293 461
rect -1199 427 -1183 461
rect -1131 427 -1115 461
rect -1021 427 -1005 461
rect -953 427 -937 461
rect -843 427 -827 461
rect -775 427 -759 461
rect -665 427 -649 461
rect -597 427 -581 461
rect -487 427 -471 461
rect -419 427 -403 461
rect -309 427 -293 461
rect -241 427 -225 461
rect -131 427 -115 461
rect -63 427 -47 461
rect 47 427 63 461
rect 115 427 131 461
rect 225 427 241 461
rect 293 427 309 461
rect 403 427 419 461
rect 471 427 487 461
rect 581 427 597 461
rect 649 427 665 461
rect 759 427 775 461
rect 827 427 843 461
rect 937 427 953 461
rect 1005 427 1021 461
rect 1115 427 1131 461
rect 1183 427 1199 461
rect 1293 427 1309 461
rect 1361 427 1521 461
rect -1441 377 -1407 427
rect -1441 71 -1407 121
rect -1263 377 -1229 393
rect -1263 105 -1229 121
rect -1085 377 -1051 393
rect -1085 105 -1051 121
rect -907 377 -873 393
rect -907 105 -873 121
rect -729 377 -695 393
rect -729 105 -695 121
rect -551 377 -517 393
rect -551 105 -517 121
rect -373 377 -339 393
rect -373 105 -339 121
rect -195 377 -161 393
rect -195 105 -161 121
rect -17 377 17 393
rect -17 105 17 121
rect 161 377 195 393
rect 161 105 195 121
rect 339 377 373 393
rect 339 105 373 121
rect 517 377 551 393
rect 517 105 551 121
rect 695 377 729 393
rect 695 105 729 121
rect 873 377 907 393
rect 873 105 907 121
rect 1051 377 1085 393
rect 1051 105 1085 121
rect 1229 377 1263 393
rect 1229 105 1263 121
rect 1407 377 1441 427
rect 1407 71 1441 121
rect -1521 37 -1361 71
rect -1309 37 -1293 71
rect -1199 37 -1183 71
rect -1131 37 -1115 71
rect -1021 37 -1005 71
rect -953 37 -937 71
rect -843 37 -827 71
rect -775 37 -759 71
rect -665 37 -649 71
rect -597 37 -581 71
rect -487 37 -471 71
rect -419 37 -403 71
rect -309 37 -293 71
rect -241 37 -225 71
rect -131 37 -115 71
rect -63 37 -47 71
rect 47 37 63 71
rect 115 37 131 71
rect 225 37 241 71
rect 293 37 309 71
rect 403 37 419 71
rect 471 37 487 71
rect 581 37 597 71
rect 649 37 665 71
rect 759 37 775 71
rect 827 37 843 71
rect 937 37 953 71
rect 1005 37 1021 71
rect 1115 37 1131 71
rect 1183 37 1199 71
rect 1293 37 1309 71
rect 1361 37 1521 71
rect -1521 -71 -1361 -37
rect -1309 -71 -1293 -37
rect -1199 -71 -1183 -37
rect -1131 -71 -1115 -37
rect -1021 -71 -1005 -37
rect -953 -71 -937 -37
rect -843 -71 -827 -37
rect -775 -71 -759 -37
rect -665 -71 -649 -37
rect -597 -71 -581 -37
rect -487 -71 -471 -37
rect -419 -71 -403 -37
rect -309 -71 -293 -37
rect -241 -71 -225 -37
rect -131 -71 -115 -37
rect -63 -71 -47 -37
rect 47 -71 63 -37
rect 115 -71 131 -37
rect 225 -71 241 -37
rect 293 -71 309 -37
rect 403 -71 419 -37
rect 471 -71 487 -37
rect 581 -71 597 -37
rect 649 -71 665 -37
rect 759 -71 775 -37
rect 827 -71 843 -37
rect 937 -71 953 -37
rect 1005 -71 1021 -37
rect 1115 -71 1131 -37
rect 1183 -71 1199 -37
rect 1293 -71 1309 -37
rect 1361 -71 1521 -37
rect -1441 -121 -1407 -71
rect -1441 -427 -1407 -377
rect -1263 -121 -1229 -105
rect -1263 -393 -1229 -377
rect -1085 -121 -1051 -105
rect -1085 -393 -1051 -377
rect -907 -121 -873 -105
rect -907 -393 -873 -377
rect -729 -121 -695 -105
rect -729 -393 -695 -377
rect -551 -121 -517 -105
rect -551 -393 -517 -377
rect -373 -121 -339 -105
rect -373 -393 -339 -377
rect -195 -121 -161 -105
rect -195 -393 -161 -377
rect -17 -121 17 -105
rect -17 -393 17 -377
rect 161 -121 195 -105
rect 161 -393 195 -377
rect 339 -121 373 -105
rect 339 -393 373 -377
rect 517 -121 551 -105
rect 517 -393 551 -377
rect 695 -121 729 -105
rect 695 -393 729 -377
rect 873 -121 907 -105
rect 873 -393 907 -377
rect 1051 -121 1085 -105
rect 1051 -393 1085 -377
rect 1229 -121 1263 -105
rect 1229 -393 1263 -377
rect 1407 -121 1441 -71
rect 1407 -427 1441 -377
rect -1521 -461 -1361 -427
rect -1309 -461 -1293 -427
rect -1199 -461 -1183 -427
rect -1131 -461 -1115 -427
rect -1021 -461 -1005 -427
rect -953 -461 -937 -427
rect -843 -461 -827 -427
rect -775 -461 -759 -427
rect -665 -461 -649 -427
rect -597 -461 -581 -427
rect -487 -461 -471 -427
rect -419 -461 -403 -427
rect -309 -461 -293 -427
rect -241 -461 -225 -427
rect -131 -461 -115 -427
rect -63 -461 -47 -427
rect 47 -461 63 -427
rect 115 -461 131 -427
rect 225 -461 241 -427
rect 293 -461 309 -427
rect 403 -461 419 -427
rect 471 -461 487 -427
rect 581 -461 597 -427
rect 649 -461 665 -427
rect 759 -461 775 -427
rect 827 -461 843 -427
rect 937 -461 953 -427
rect 1005 -461 1021 -427
rect 1115 -461 1131 -427
rect 1183 -461 1199 -427
rect 1293 -461 1309 -427
rect 1361 -461 1521 -427
rect -1521 -569 -1361 -535
rect -1309 -569 -1293 -535
rect -1199 -569 -1183 -535
rect -1131 -569 -1115 -535
rect -1021 -569 -1005 -535
rect -953 -569 -937 -535
rect -843 -569 -827 -535
rect -775 -569 -759 -535
rect -665 -569 -649 -535
rect -597 -569 -581 -535
rect -487 -569 -471 -535
rect -419 -569 -403 -535
rect -309 -569 -293 -535
rect -241 -569 -225 -535
rect -131 -569 -115 -535
rect -63 -569 -47 -535
rect 47 -569 63 -535
rect 115 -569 131 -535
rect 225 -569 241 -535
rect 293 -569 309 -535
rect 403 -569 419 -535
rect 471 -569 487 -535
rect 581 -569 597 -535
rect 649 -569 665 -535
rect 759 -569 775 -535
rect 827 -569 843 -535
rect 937 -569 953 -535
rect 1005 -569 1021 -535
rect 1115 -569 1131 -535
rect 1183 -569 1199 -535
rect 1293 -569 1309 -535
rect 1361 -569 1521 -535
rect -1441 -619 -1407 -569
rect -1441 -925 -1407 -875
rect -1263 -619 -1229 -603
rect -1263 -891 -1229 -875
rect -1085 -619 -1051 -603
rect -1085 -891 -1051 -875
rect -907 -619 -873 -603
rect -907 -891 -873 -875
rect -729 -619 -695 -603
rect -729 -891 -695 -875
rect -551 -619 -517 -603
rect -551 -891 -517 -875
rect -373 -619 -339 -603
rect -373 -891 -339 -875
rect -195 -619 -161 -603
rect -195 -891 -161 -875
rect -17 -619 17 -603
rect -17 -891 17 -875
rect 161 -619 195 -603
rect 161 -891 195 -875
rect 339 -619 373 -603
rect 339 -891 373 -875
rect 517 -619 551 -603
rect 517 -891 551 -875
rect 695 -619 729 -603
rect 695 -891 729 -875
rect 873 -619 907 -603
rect 873 -891 907 -875
rect 1051 -619 1085 -603
rect 1051 -891 1085 -875
rect 1229 -619 1263 -603
rect 1229 -891 1263 -875
rect 1407 -619 1441 -569
rect 1407 -925 1441 -875
rect -1521 -959 -1361 -925
rect -1309 -959 -1293 -925
rect -1199 -959 -1183 -925
rect -1131 -959 -1115 -925
rect -1021 -959 -1005 -925
rect -953 -959 -937 -925
rect -843 -959 -827 -925
rect -775 -959 -759 -925
rect -665 -959 -649 -925
rect -597 -959 -581 -925
rect -487 -959 -471 -925
rect -419 -959 -403 -925
rect -309 -959 -293 -925
rect -241 -959 -225 -925
rect -131 -959 -115 -925
rect -63 -959 -47 -925
rect 47 -959 63 -925
rect 115 -959 131 -925
rect 225 -959 241 -925
rect 293 -959 309 -925
rect 403 -959 419 -925
rect 471 -959 487 -925
rect 581 -959 597 -925
rect 649 -959 665 -925
rect 759 -959 775 -925
rect 827 -959 843 -925
rect 937 -959 953 -925
rect 1005 -959 1021 -925
rect 1115 -959 1131 -925
rect 1183 -959 1199 -925
rect 1293 -959 1309 -925
rect 1361 -959 1521 -925
rect -1555 -1027 -1521 -965
rect 1521 -1027 1555 -965
rect -1555 -1061 -1459 -1027
rect 1459 -1061 1555 -1027
<< viali >>
rect -1183 925 -1131 959
rect -1005 925 -953 959
rect -827 925 -775 959
rect -649 925 -597 959
rect -471 925 -419 959
rect -293 925 -241 959
rect -115 925 -63 959
rect 63 925 115 959
rect 241 925 293 959
rect 419 925 471 959
rect 597 925 649 959
rect 775 925 827 959
rect 953 925 1005 959
rect 1131 925 1183 959
rect -1183 535 -1131 569
rect -1005 535 -953 569
rect -827 535 -775 569
rect -649 535 -597 569
rect -471 535 -419 569
rect -293 535 -241 569
rect -115 535 -63 569
rect 63 535 115 569
rect 241 535 293 569
rect 419 535 471 569
rect 597 535 649 569
rect 775 535 827 569
rect 953 535 1005 569
rect 1131 535 1183 569
rect -1183 427 -1131 461
rect -1005 427 -953 461
rect -827 427 -775 461
rect -649 427 -597 461
rect -471 427 -419 461
rect -293 427 -241 461
rect -115 427 -63 461
rect 63 427 115 461
rect 241 427 293 461
rect 419 427 471 461
rect 597 427 649 461
rect 775 427 827 461
rect 953 427 1005 461
rect 1131 427 1183 461
rect -1183 37 -1131 71
rect -1005 37 -953 71
rect -827 37 -775 71
rect -649 37 -597 71
rect -471 37 -419 71
rect -293 37 -241 71
rect -115 37 -63 71
rect 63 37 115 71
rect 241 37 293 71
rect 419 37 471 71
rect 597 37 649 71
rect 775 37 827 71
rect 953 37 1005 71
rect 1131 37 1183 71
rect -1183 -71 -1131 -37
rect -1005 -71 -953 -37
rect -827 -71 -775 -37
rect -649 -71 -597 -37
rect -471 -71 -419 -37
rect -293 -71 -241 -37
rect -115 -71 -63 -37
rect 63 -71 115 -37
rect 241 -71 293 -37
rect 419 -71 471 -37
rect 597 -71 649 -37
rect 775 -71 827 -37
rect 953 -71 1005 -37
rect 1131 -71 1183 -37
rect -1183 -461 -1131 -427
rect -1005 -461 -953 -427
rect -827 -461 -775 -427
rect -649 -461 -597 -427
rect -471 -461 -419 -427
rect -293 -461 -241 -427
rect -115 -461 -63 -427
rect 63 -461 115 -427
rect 241 -461 293 -427
rect 419 -461 471 -427
rect 597 -461 649 -427
rect 775 -461 827 -427
rect 953 -461 1005 -427
rect 1131 -461 1183 -427
rect -1183 -569 -1131 -535
rect -1005 -569 -953 -535
rect -827 -569 -775 -535
rect -649 -569 -597 -535
rect -471 -569 -419 -535
rect -293 -569 -241 -535
rect -115 -569 -63 -535
rect 63 -569 115 -535
rect 241 -569 293 -535
rect 419 -569 471 -535
rect 597 -569 649 -535
rect 775 -569 827 -535
rect 953 -569 1005 -535
rect 1131 -569 1183 -535
rect -1183 -959 -1131 -925
rect -1005 -959 -953 -925
rect -827 -959 -775 -925
rect -649 -959 -597 -925
rect -471 -959 -419 -925
rect -293 -959 -241 -925
rect -115 -959 -63 -925
rect 63 -959 115 -925
rect 241 -959 293 -925
rect 419 -959 471 -925
rect 597 -959 649 -925
rect 775 -959 827 -925
rect 953 -959 1005 -925
rect 1131 -959 1183 -925
<< metal1 >>
rect -1195 959 -1119 965
rect -1195 925 -1183 959
rect -1131 925 -1119 959
rect -1195 919 -1119 925
rect -1017 959 -941 965
rect -1017 925 -1005 959
rect -953 925 -941 959
rect -1017 919 -941 925
rect -839 959 -763 965
rect -839 925 -827 959
rect -775 925 -763 959
rect -839 919 -763 925
rect -661 959 -585 965
rect -661 925 -649 959
rect -597 925 -585 959
rect -661 919 -585 925
rect -483 959 -407 965
rect -483 925 -471 959
rect -419 925 -407 959
rect -483 919 -407 925
rect -305 959 -229 965
rect -305 925 -293 959
rect -241 925 -229 959
rect -305 919 -229 925
rect -127 959 -51 965
rect -127 925 -115 959
rect -63 925 -51 959
rect -127 919 -51 925
rect 51 959 127 965
rect 51 925 63 959
rect 115 925 127 959
rect 51 919 127 925
rect 229 959 305 965
rect 229 925 241 959
rect 293 925 305 959
rect 229 919 305 925
rect 407 959 483 965
rect 407 925 419 959
rect 471 925 483 959
rect 407 919 483 925
rect 585 959 661 965
rect 585 925 597 959
rect 649 925 661 959
rect 585 919 661 925
rect 763 959 839 965
rect 763 925 775 959
rect 827 925 839 959
rect 763 919 839 925
rect 941 959 1017 965
rect 941 925 953 959
rect 1005 925 1017 959
rect 941 919 1017 925
rect 1119 959 1195 965
rect 1119 925 1131 959
rect 1183 925 1195 959
rect 1119 919 1195 925
rect -1195 569 -1119 575
rect -1195 535 -1183 569
rect -1131 535 -1119 569
rect -1195 529 -1119 535
rect -1017 569 -941 575
rect -1017 535 -1005 569
rect -953 535 -941 569
rect -1017 529 -941 535
rect -839 569 -763 575
rect -839 535 -827 569
rect -775 535 -763 569
rect -839 529 -763 535
rect -661 569 -585 575
rect -661 535 -649 569
rect -597 535 -585 569
rect -661 529 -585 535
rect -483 569 -407 575
rect -483 535 -471 569
rect -419 535 -407 569
rect -483 529 -407 535
rect -305 569 -229 575
rect -305 535 -293 569
rect -241 535 -229 569
rect -305 529 -229 535
rect -127 569 -51 575
rect -127 535 -115 569
rect -63 535 -51 569
rect -127 529 -51 535
rect 51 569 127 575
rect 51 535 63 569
rect 115 535 127 569
rect 51 529 127 535
rect 229 569 305 575
rect 229 535 241 569
rect 293 535 305 569
rect 229 529 305 535
rect 407 569 483 575
rect 407 535 419 569
rect 471 535 483 569
rect 407 529 483 535
rect 585 569 661 575
rect 585 535 597 569
rect 649 535 661 569
rect 585 529 661 535
rect 763 569 839 575
rect 763 535 775 569
rect 827 535 839 569
rect 763 529 839 535
rect 941 569 1017 575
rect 941 535 953 569
rect 1005 535 1017 569
rect 941 529 1017 535
rect 1119 569 1195 575
rect 1119 535 1131 569
rect 1183 535 1195 569
rect 1119 529 1195 535
rect -1195 461 -1119 467
rect -1195 427 -1183 461
rect -1131 427 -1119 461
rect -1195 421 -1119 427
rect -1017 461 -941 467
rect -1017 427 -1005 461
rect -953 427 -941 461
rect -1017 421 -941 427
rect -839 461 -763 467
rect -839 427 -827 461
rect -775 427 -763 461
rect -839 421 -763 427
rect -661 461 -585 467
rect -661 427 -649 461
rect -597 427 -585 461
rect -661 421 -585 427
rect -483 461 -407 467
rect -483 427 -471 461
rect -419 427 -407 461
rect -483 421 -407 427
rect -305 461 -229 467
rect -305 427 -293 461
rect -241 427 -229 461
rect -305 421 -229 427
rect -127 461 -51 467
rect -127 427 -115 461
rect -63 427 -51 461
rect -127 421 -51 427
rect 51 461 127 467
rect 51 427 63 461
rect 115 427 127 461
rect 51 421 127 427
rect 229 461 305 467
rect 229 427 241 461
rect 293 427 305 461
rect 229 421 305 427
rect 407 461 483 467
rect 407 427 419 461
rect 471 427 483 461
rect 407 421 483 427
rect 585 461 661 467
rect 585 427 597 461
rect 649 427 661 461
rect 585 421 661 427
rect 763 461 839 467
rect 763 427 775 461
rect 827 427 839 461
rect 763 421 839 427
rect 941 461 1017 467
rect 941 427 953 461
rect 1005 427 1017 461
rect 941 421 1017 427
rect 1119 461 1195 467
rect 1119 427 1131 461
rect 1183 427 1195 461
rect 1119 421 1195 427
rect -1195 71 -1119 77
rect -1195 37 -1183 71
rect -1131 37 -1119 71
rect -1195 31 -1119 37
rect -1017 71 -941 77
rect -1017 37 -1005 71
rect -953 37 -941 71
rect -1017 31 -941 37
rect -839 71 -763 77
rect -839 37 -827 71
rect -775 37 -763 71
rect -839 31 -763 37
rect -661 71 -585 77
rect -661 37 -649 71
rect -597 37 -585 71
rect -661 31 -585 37
rect -483 71 -407 77
rect -483 37 -471 71
rect -419 37 -407 71
rect -483 31 -407 37
rect -305 71 -229 77
rect -305 37 -293 71
rect -241 37 -229 71
rect -305 31 -229 37
rect -127 71 -51 77
rect -127 37 -115 71
rect -63 37 -51 71
rect -127 31 -51 37
rect 51 71 127 77
rect 51 37 63 71
rect 115 37 127 71
rect 51 31 127 37
rect 229 71 305 77
rect 229 37 241 71
rect 293 37 305 71
rect 229 31 305 37
rect 407 71 483 77
rect 407 37 419 71
rect 471 37 483 71
rect 407 31 483 37
rect 585 71 661 77
rect 585 37 597 71
rect 649 37 661 71
rect 585 31 661 37
rect 763 71 839 77
rect 763 37 775 71
rect 827 37 839 71
rect 763 31 839 37
rect 941 71 1017 77
rect 941 37 953 71
rect 1005 37 1017 71
rect 941 31 1017 37
rect 1119 71 1195 77
rect 1119 37 1131 71
rect 1183 37 1195 71
rect 1119 31 1195 37
rect -1195 -37 -1119 -31
rect -1195 -71 -1183 -37
rect -1131 -71 -1119 -37
rect -1195 -77 -1119 -71
rect -1017 -37 -941 -31
rect -1017 -71 -1005 -37
rect -953 -71 -941 -37
rect -1017 -77 -941 -71
rect -839 -37 -763 -31
rect -839 -71 -827 -37
rect -775 -71 -763 -37
rect -839 -77 -763 -71
rect -661 -37 -585 -31
rect -661 -71 -649 -37
rect -597 -71 -585 -37
rect -661 -77 -585 -71
rect -483 -37 -407 -31
rect -483 -71 -471 -37
rect -419 -71 -407 -37
rect -483 -77 -407 -71
rect -305 -37 -229 -31
rect -305 -71 -293 -37
rect -241 -71 -229 -37
rect -305 -77 -229 -71
rect -127 -37 -51 -31
rect -127 -71 -115 -37
rect -63 -71 -51 -37
rect -127 -77 -51 -71
rect 51 -37 127 -31
rect 51 -71 63 -37
rect 115 -71 127 -37
rect 51 -77 127 -71
rect 229 -37 305 -31
rect 229 -71 241 -37
rect 293 -71 305 -37
rect 229 -77 305 -71
rect 407 -37 483 -31
rect 407 -71 419 -37
rect 471 -71 483 -37
rect 407 -77 483 -71
rect 585 -37 661 -31
rect 585 -71 597 -37
rect 649 -71 661 -37
rect 585 -77 661 -71
rect 763 -37 839 -31
rect 763 -71 775 -37
rect 827 -71 839 -37
rect 763 -77 839 -71
rect 941 -37 1017 -31
rect 941 -71 953 -37
rect 1005 -71 1017 -37
rect 941 -77 1017 -71
rect 1119 -37 1195 -31
rect 1119 -71 1131 -37
rect 1183 -71 1195 -37
rect 1119 -77 1195 -71
rect -1195 -427 -1119 -421
rect -1195 -461 -1183 -427
rect -1131 -461 -1119 -427
rect -1195 -467 -1119 -461
rect -1017 -427 -941 -421
rect -1017 -461 -1005 -427
rect -953 -461 -941 -427
rect -1017 -467 -941 -461
rect -839 -427 -763 -421
rect -839 -461 -827 -427
rect -775 -461 -763 -427
rect -839 -467 -763 -461
rect -661 -427 -585 -421
rect -661 -461 -649 -427
rect -597 -461 -585 -427
rect -661 -467 -585 -461
rect -483 -427 -407 -421
rect -483 -461 -471 -427
rect -419 -461 -407 -427
rect -483 -467 -407 -461
rect -305 -427 -229 -421
rect -305 -461 -293 -427
rect -241 -461 -229 -427
rect -305 -467 -229 -461
rect -127 -427 -51 -421
rect -127 -461 -115 -427
rect -63 -461 -51 -427
rect -127 -467 -51 -461
rect 51 -427 127 -421
rect 51 -461 63 -427
rect 115 -461 127 -427
rect 51 -467 127 -461
rect 229 -427 305 -421
rect 229 -461 241 -427
rect 293 -461 305 -427
rect 229 -467 305 -461
rect 407 -427 483 -421
rect 407 -461 419 -427
rect 471 -461 483 -427
rect 407 -467 483 -461
rect 585 -427 661 -421
rect 585 -461 597 -427
rect 649 -461 661 -427
rect 585 -467 661 -461
rect 763 -427 839 -421
rect 763 -461 775 -427
rect 827 -461 839 -427
rect 763 -467 839 -461
rect 941 -427 1017 -421
rect 941 -461 953 -427
rect 1005 -461 1017 -427
rect 941 -467 1017 -461
rect 1119 -427 1195 -421
rect 1119 -461 1131 -427
rect 1183 -461 1195 -427
rect 1119 -467 1195 -461
rect -1195 -535 -1119 -529
rect -1195 -569 -1183 -535
rect -1131 -569 -1119 -535
rect -1195 -575 -1119 -569
rect -1017 -535 -941 -529
rect -1017 -569 -1005 -535
rect -953 -569 -941 -535
rect -1017 -575 -941 -569
rect -839 -535 -763 -529
rect -839 -569 -827 -535
rect -775 -569 -763 -535
rect -839 -575 -763 -569
rect -661 -535 -585 -529
rect -661 -569 -649 -535
rect -597 -569 -585 -535
rect -661 -575 -585 -569
rect -483 -535 -407 -529
rect -483 -569 -471 -535
rect -419 -569 -407 -535
rect -483 -575 -407 -569
rect -305 -535 -229 -529
rect -305 -569 -293 -535
rect -241 -569 -229 -535
rect -305 -575 -229 -569
rect -127 -535 -51 -529
rect -127 -569 -115 -535
rect -63 -569 -51 -535
rect -127 -575 -51 -569
rect 51 -535 127 -529
rect 51 -569 63 -535
rect 115 -569 127 -535
rect 51 -575 127 -569
rect 229 -535 305 -529
rect 229 -569 241 -535
rect 293 -569 305 -535
rect 229 -575 305 -569
rect 407 -535 483 -529
rect 407 -569 419 -535
rect 471 -569 483 -535
rect 407 -575 483 -569
rect 585 -535 661 -529
rect 585 -569 597 -535
rect 649 -569 661 -535
rect 585 -575 661 -569
rect 763 -535 839 -529
rect 763 -569 775 -535
rect 827 -569 839 -535
rect 763 -575 839 -569
rect 941 -535 1017 -529
rect 941 -569 953 -535
rect 1005 -569 1017 -535
rect 941 -575 1017 -569
rect 1119 -535 1195 -529
rect 1119 -569 1131 -535
rect 1183 -569 1195 -535
rect 1119 -575 1195 -569
rect -1195 -925 -1119 -919
rect -1195 -959 -1183 -925
rect -1131 -959 -1119 -925
rect -1195 -965 -1119 -959
rect -1017 -925 -941 -919
rect -1017 -959 -1005 -925
rect -953 -959 -941 -925
rect -1017 -965 -941 -959
rect -839 -925 -763 -919
rect -839 -959 -827 -925
rect -775 -959 -763 -925
rect -839 -965 -763 -959
rect -661 -925 -585 -919
rect -661 -959 -649 -925
rect -597 -959 -585 -925
rect -661 -965 -585 -959
rect -483 -925 -407 -919
rect -483 -959 -471 -925
rect -419 -959 -407 -925
rect -483 -965 -407 -959
rect -305 -925 -229 -919
rect -305 -959 -293 -925
rect -241 -959 -229 -925
rect -305 -965 -229 -959
rect -127 -925 -51 -919
rect -127 -959 -115 -925
rect -63 -959 -51 -925
rect -127 -965 -51 -959
rect 51 -925 127 -919
rect 51 -959 63 -925
rect 115 -959 127 -925
rect 51 -965 127 -959
rect 229 -925 305 -919
rect 229 -959 241 -925
rect 293 -959 305 -925
rect 229 -965 305 -959
rect 407 -925 483 -919
rect 407 -959 419 -925
rect 471 -959 483 -925
rect 407 -965 483 -959
rect 585 -925 661 -919
rect 585 -959 597 -925
rect 649 -959 661 -925
rect 585 -965 661 -959
rect 763 -925 839 -919
rect 763 -959 775 -925
rect 827 -959 839 -925
rect 763 -965 839 -959
rect 941 -925 1017 -919
rect 941 -959 953 -925
rect 1005 -959 1017 -925
rect 941 -965 1017 -959
rect 1119 -925 1195 -919
rect 1119 -959 1131 -925
rect 1183 -959 1195 -925
rect 1119 -965 1195 -959
<< properties >>
string FIXED_BBOX -1538 -1044 1538 1044
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.4 l 0.6 m 4 nf 16 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
