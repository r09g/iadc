magic
tech sky130A
timestamp 1654711401
<< metal3 >>
rect -655 -630 605 630
<< mimcap >>
rect -605 560 555 580
rect -605 -560 -585 560
rect 535 -560 555 560
rect -605 -580 555 -560
<< mimcapcontact >>
rect -585 -560 535 560
<< metal4 >>
rect -585 560 535 560
rect -585 -560 -585 560
rect 535 -560 535 560
rect -585 -560 535 -560
<< properties >>
string FIXED_BBOX -655 -630 605 630
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 11.6 l 11.6 val 277.936 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
