magic
tech sky130A
timestamp 1654517900
<< nmoslvt >>
rect -10 -60 10 60
<< ndiff >>
rect -39 54 -10 60
rect -39 -54 -33 54
rect -16 -54 -10 54
rect -39 -60 -10 -54
rect 10 54 39 60
rect 10 -54 16 54
rect 33 -54 39 54
rect 10 -60 39 -54
<< ndiffc >>
rect -33 -54 -16 54
rect 16 -54 33 54
<< poly >>
rect -16 96 16 104
rect -16 79 -8 96
rect 8 79 16 96
rect -16 71 16 79
rect -10 60 10 71
rect -10 -71 10 -60
rect -16 -79 16 -71
rect -16 -96 -8 -79
rect 8 -96 16 -79
rect -16 -104 16 -96
<< polycont >>
rect -8 79 8 96
rect -8 -96 8 -79
<< locali >>
rect -16 79 -8 96
rect 8 79 16 96
rect -33 54 -16 62
rect -33 -62 -16 -54
rect 16 54 33 62
rect 16 -62 33 -54
rect -16 -96 -8 -79
rect 8 -96 16 -79
<< viali >>
rect -8 79 8 96
rect -33 -54 -16 54
rect 16 -54 33 54
rect -8 -96 8 -79
<< metal1 >>
rect -16 96 16 104
rect -16 79 -8 96
rect 8 79 16 96
rect -16 76 16 79
rect -36 54 -13 60
rect -36 -54 -33 54
rect -16 -54 -13 54
rect -36 -60 -13 -54
rect 13 54 36 60
rect 13 -54 16 54
rect 33 -54 36 54
rect 13 -60 36 -54
rect -16 -79 16 -76
rect -16 -96 -8 -79
rect 8 -96 16 -79
rect -16 -104 16 -96
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.2 l 0.2 m 1 nf 1 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
