magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect 230 447 288 453
rect 422 447 480 453
rect 614 447 672 453
rect 806 447 864 453
rect 998 447 1056 453
rect 1190 447 1248 453
rect 1382 447 1440 453
rect 1574 447 1632 453
rect 230 413 242 447
rect 422 413 434 447
rect 614 413 626 447
rect 806 413 818 447
rect 998 413 1010 447
rect 1190 413 1202 447
rect 1382 413 1394 447
rect 1574 413 1586 447
rect 230 407 288 413
rect 422 407 480 413
rect 614 407 672 413
rect 806 407 864 413
rect 998 407 1056 413
rect 1190 407 1248 413
rect 1382 407 1440 413
rect 1574 407 1632 413
rect 326 119 384 125
rect 518 119 576 125
rect 710 119 768 125
rect 902 119 960 125
rect 1094 119 1152 125
rect 1286 119 1344 125
rect 1478 119 1536 125
rect 1670 119 1728 125
rect 326 85 338 119
rect 518 85 530 119
rect 710 85 722 119
rect 902 85 914 119
rect 1094 85 1106 119
rect 1286 85 1298 119
rect 1478 85 1490 119
rect 1670 85 1682 119
rect 326 79 384 85
rect 518 79 576 85
rect 710 79 768 85
rect 902 79 960 85
rect 1094 79 1152 85
rect 1286 79 1344 85
rect 1478 79 1536 85
rect 1670 79 1728 85
use sky130_fd_pr__pfet_01v8_VCG74W  sky130_fd_pr__pfet_01v8_VCG74W_0
timestamp 1654583101
transform 1 0 979 0 1 266
box -1031 -319 1031 319
<< end >>
