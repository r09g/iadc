* NGSPICE file created from ota.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_VU7MNH a_n652_n140# a_652_n194# a_772_n140# a_n60_n194#
+ a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140# a_296_n194#
+ a_60_n140# a_416_n140# a_n118_n140# a_118_n194# a_238_n140# a_n772_n194# a_n830_n140#
+ a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_118_n194# a_n60_n194# 0.10fF
C1 a_296_n194# a_n238_n194# 0.02fF
C2 a_296_n194# a_n594_n194# 0.01fF
C3 a_n296_n140# a_594_n140# 0.02fF
C4 a_n296_n140# a_416_n140# 0.03fF
C5 a_296_n194# a_n772_n194# 0.01fF
C6 a_n296_n140# a_n830_n140# 0.04fF
C7 a_n238_n194# a_n60_n194# 0.10fF
C8 a_594_n140# a_238_n140# 0.06fF
C9 a_238_n140# a_416_n140# 0.13fF
C10 a_n60_n194# a_n594_n194# 0.02fF
C11 a_n474_n140# a_n296_n140# 0.13fF
C12 a_n118_n140# a_594_n140# 0.03fF
C13 a_n118_n140# a_416_n140# 0.04fF
C14 a_n296_n140# a_772_n140# 0.02fF
C15 a_n830_n140# a_238_n140# 0.02fF
C16 a_60_n140# a_n652_n140# 0.03fF
C17 a_n60_n194# a_n772_n194# 0.01fF
C18 a_n416_n194# a_652_n194# 0.01fF
C19 a_n118_n140# a_n830_n140# 0.03fF
C20 a_118_n194# a_474_n194# 0.03fF
C21 a_n474_n140# a_238_n140# 0.03fF
C22 a_772_n140# a_238_n140# 0.04fF
C23 a_n118_n140# a_n474_n140# 0.06fF
C24 a_n118_n140# a_772_n140# 0.02fF
C25 a_296_n194# a_652_n194# 0.03fF
C26 a_474_n194# a_n238_n194# 0.01fF
C27 a_474_n194# a_n594_n194# 0.01fF
C28 a_118_n194# a_n238_n194# 0.03fF
C29 a_118_n194# a_n594_n194# 0.01fF
C30 a_474_n194# a_n772_n194# 0.01fF
C31 a_n60_n194# a_652_n194# 0.01fF
C32 a_118_n194# a_n772_n194# 0.01fF
C33 a_60_n140# a_n296_n140# 0.06fF
C34 a_n652_n140# a_n296_n140# 0.06fF
C35 a_594_n140# a_416_n140# 0.13fF
C36 a_296_n194# a_n416_n194# 0.01fF
C37 a_n830_n140# a_594_n140# 0.01fF
C38 a_n830_n140# a_416_n140# 0.02fF
C39 a_60_n140# a_238_n140# 0.13fF
C40 a_n652_n140# a_238_n140# 0.02fF
C41 a_n238_n194# a_n594_n194# 0.03fF
C42 a_n118_n140# a_60_n140# 0.13fF
C43 a_n118_n140# a_n652_n140# 0.04fF
C44 a_n238_n194# a_n772_n194# 0.02fF
C45 a_n474_n140# a_594_n140# 0.02fF
C46 a_n474_n140# a_416_n140# 0.02fF
C47 a_594_n140# a_772_n140# 0.13fF
C48 a_772_n140# a_416_n140# 0.06fF
C49 a_n416_n194# a_n60_n194# 0.03fF
C50 a_n594_n194# a_n772_n194# 0.10fF
C51 a_n474_n140# a_n830_n140# 0.06fF
C52 a_n830_n140# a_772_n140# 0.01fF
C53 a_474_n194# a_652_n194# 0.10fF
C54 a_n474_n140# a_772_n140# 0.02fF
C55 a_118_n194# a_652_n194# 0.02fF
C56 a_296_n194# a_n60_n194# 0.03fF
C57 a_n238_n194# a_652_n194# 0.01fF
C58 a_n296_n140# a_238_n140# 0.04fF
C59 a_474_n194# a_n416_n194# 0.01fF
C60 a_652_n194# a_n594_n194# 0.01fF
C61 a_n118_n140# a_n296_n140# 0.13fF
C62 a_118_n194# a_n416_n194# 0.02fF
C63 a_60_n140# a_594_n140# 0.04fF
C64 a_60_n140# a_416_n140# 0.06fF
C65 a_n652_n140# a_594_n140# 0.02fF
C66 a_n652_n140# a_416_n140# 0.02fF
C67 a_652_n194# a_n772_n194# 0.01fF
C68 a_60_n140# a_n830_n140# 0.02fF
C69 a_n652_n140# a_n830_n140# 0.13fF
C70 a_n118_n140# a_238_n140# 0.06fF
C71 a_296_n194# a_474_n194# 0.10fF
C72 a_60_n140# a_n474_n140# 0.04fF
C73 a_n652_n140# a_n474_n140# 0.13fF
C74 a_60_n140# a_772_n140# 0.03fF
C75 a_n652_n140# a_772_n140# 0.01fF
C76 a_n416_n194# a_n238_n194# 0.10fF
C77 a_118_n194# a_296_n194# 0.10fF
C78 a_n416_n194# a_n594_n194# 0.10fF
C79 a_n416_n194# a_n772_n194# 0.03fF
C80 a_474_n194# a_n60_n194# 0.02fF
C81 a_772_n140# VSUBS 0.02fF
C82 a_594_n140# VSUBS 0.02fF
C83 a_416_n140# VSUBS 0.02fF
C84 a_238_n140# VSUBS 0.02fF
C85 a_60_n140# VSUBS 0.02fF
C86 a_n118_n140# VSUBS 0.02fF
C87 a_n296_n140# VSUBS 0.02fF
C88 a_n474_n140# VSUBS 0.02fF
C89 a_n652_n140# VSUBS 0.02fF
C90 a_n830_n140# VSUBS 0.02fF
C91 a_652_n194# VSUBS 0.29fF
C92 a_474_n194# VSUBS 0.23fF
C93 a_296_n194# VSUBS 0.24fF
C94 a_118_n194# VSUBS 0.25fF
C95 a_n60_n194# VSUBS 0.26fF
C96 a_n238_n194# VSUBS 0.27fF
C97 a_n416_n194# VSUBS 0.28fF
C98 a_n594_n194# VSUBS 0.28fF
C99 a_n772_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_TRAZV8 a_21_n120# a_n79_n120# a_n33_n208# VSUBS
X0 a_21_n120# a_n33_n208# a_n79_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=210000u
C0 a_n33_n208# a_n79_n120# 0.01fF
C1 a_n33_n208# a_21_n120# 0.01fF
C2 a_21_n120# a_n79_n120# 0.27fF
C3 a_21_n120# VSUBS 0.02fF
C4 a_n79_n120# VSUBS 0.02fF
C5 a_n33_n208# VSUBS 0.29fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BASQVB a_n1008_n140# a_n652_n140# a_652_n194# a_772_n140#
+ a_n60_n194# a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140#
+ a_296_n194# a_60_n140# a_416_n140# a_n950_n194# a_n118_n140# a_118_n194# a_238_n140#
+ a_n772_n194# a_n830_n140# a_830_n194# a_950_n140# a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n416_n194# a_n238_n194# 0.10fF
C1 a_60_n140# a_594_n140# 0.04fF
C2 a_n594_n194# a_n60_n194# 0.02fF
C3 a_238_n140# a_416_n140# 0.13fF
C4 a_n1008_n140# a_60_n140# 0.02fF
C5 a_950_n140# a_416_n140# 0.04fF
C6 a_n594_n194# a_296_n194# 0.01fF
C7 a_474_n194# a_n238_n194# 0.01fF
C8 a_n594_n194# a_830_n194# 0.01fF
C9 a_652_n194# a_n950_n194# 0.01fF
C10 a_60_n140# a_n474_n140# 0.04fF
C11 a_n60_n194# a_n238_n194# 0.10fF
C12 a_n830_n140# a_594_n140# 0.01fF
C13 a_n238_n194# a_296_n194# 0.02fF
C14 a_n1008_n140# a_n830_n140# 0.13fF
C15 a_n118_n140# a_594_n140# 0.03fF
C16 a_238_n140# a_772_n140# 0.04fF
C17 a_118_n194# a_n950_n194# 0.01fF
C18 a_830_n194# a_n238_n194# 0.01fF
C19 a_772_n140# a_950_n140# 0.13fF
C20 a_n1008_n140# a_n118_n140# 0.02fF
C21 a_594_n140# a_n652_n140# 0.02fF
C22 a_n296_n140# a_594_n140# 0.02fF
C23 a_n416_n194# a_n772_n194# 0.03fF
C24 a_n1008_n140# a_n652_n140# 0.06fF
C25 a_n830_n140# a_n474_n140# 0.06fF
C26 a_n1008_n140# a_n296_n140# 0.03fF
C27 a_652_n194# a_118_n194# 0.02fF
C28 a_n118_n140# a_n474_n140# 0.06fF
C29 a_238_n140# a_950_n140# 0.03fF
C30 a_474_n194# a_n772_n194# 0.01fF
C31 a_474_n194# a_n416_n194# 0.01fF
C32 a_n594_n194# a_n950_n194# 0.03fF
C33 a_n474_n140# a_n652_n140# 0.13fF
C34 a_594_n140# a_416_n140# 0.13fF
C35 a_n474_n140# a_n296_n140# 0.13fF
C36 a_n830_n140# a_60_n140# 0.02fF
C37 a_n772_n194# a_n60_n194# 0.01fF
C38 a_n1008_n140# a_416_n140# 0.01fF
C39 a_n118_n140# a_60_n140# 0.13fF
C40 a_n772_n194# a_296_n194# 0.01fF
C41 a_n416_n194# a_n60_n194# 0.03fF
C42 a_n594_n194# a_652_n194# 0.01fF
C43 a_n416_n194# a_296_n194# 0.01fF
C44 a_n238_n194# a_n950_n194# 0.01fF
C45 a_60_n140# a_n652_n140# 0.03fF
C46 a_60_n140# a_n296_n140# 0.06fF
C47 a_n772_n194# a_830_n194# 0.01fF
C48 a_474_n194# a_n60_n194# 0.02fF
C49 a_n474_n140# a_416_n140# 0.02fF
C50 a_n416_n194# a_830_n194# 0.01fF
C51 a_474_n194# a_296_n194# 0.10fF
C52 a_n594_n194# a_118_n194# 0.01fF
C53 a_772_n140# a_594_n140# 0.13fF
C54 a_652_n194# a_n238_n194# 0.01fF
C55 a_n118_n140# a_n830_n140# 0.03fF
C56 a_474_n194# a_830_n194# 0.03fF
C57 a_n60_n194# a_296_n194# 0.03fF
C58 a_60_n140# a_416_n140# 0.06fF
C59 a_n830_n140# a_n652_n140# 0.13fF
C60 a_n830_n140# a_n296_n140# 0.04fF
C61 a_238_n140# a_594_n140# 0.06fF
C62 a_118_n194# a_n238_n194# 0.03fF
C63 a_830_n194# a_n60_n194# 0.01fF
C64 a_950_n140# a_594_n140# 0.06fF
C65 a_n118_n140# a_n652_n140# 0.04fF
C66 a_n118_n140# a_n296_n140# 0.13fF
C67 a_772_n140# a_n474_n140# 0.02fF
C68 a_n1008_n140# a_238_n140# 0.02fF
C69 a_830_n194# a_296_n194# 0.02fF
C70 a_n296_n140# a_n652_n140# 0.06fF
C71 a_n772_n194# a_n950_n194# 0.10fF
C72 a_n830_n140# a_416_n140# 0.02fF
C73 a_n416_n194# a_n950_n194# 0.02fF
C74 a_238_n140# a_n474_n140# 0.03fF
C75 a_772_n140# a_60_n140# 0.03fF
C76 a_950_n140# a_n474_n140# 0.01fF
C77 a_n118_n140# a_416_n140# 0.04fF
C78 a_n594_n194# a_n238_n194# 0.03fF
C79 a_652_n194# a_n772_n194# 0.01fF
C80 a_474_n194# a_n950_n194# 0.01fF
C81 a_n652_n140# a_416_n140# 0.02fF
C82 a_n296_n140# a_416_n140# 0.03fF
C83 a_n416_n194# a_652_n194# 0.01fF
C84 a_238_n140# a_60_n140# 0.13fF
C85 a_950_n140# a_60_n140# 0.02fF
C86 a_n60_n194# a_n950_n194# 0.01fF
C87 a_n772_n194# a_118_n194# 0.01fF
C88 a_474_n194# a_652_n194# 0.10fF
C89 a_772_n140# a_n830_n140# 0.01fF
C90 a_n950_n194# a_296_n194# 0.01fF
C91 a_n416_n194# a_118_n194# 0.02fF
C92 a_n118_n140# a_772_n140# 0.02fF
C93 a_652_n194# a_n60_n194# 0.01fF
C94 a_772_n140# a_n652_n140# 0.01fF
C95 a_474_n194# a_118_n194# 0.03fF
C96 a_652_n194# a_296_n194# 0.03fF
C97 a_n1008_n140# a_594_n140# 0.01fF
C98 a_772_n140# a_n296_n140# 0.02fF
C99 a_238_n140# a_n830_n140# 0.02fF
C100 a_n594_n194# a_n772_n194# 0.10fF
C101 a_n118_n140# a_238_n140# 0.06fF
C102 a_n118_n140# a_950_n140# 0.02fF
C103 a_652_n194# a_830_n194# 0.10fF
C104 a_118_n194# a_n60_n194# 0.10fF
C105 a_n416_n194# a_n594_n194# 0.10fF
C106 a_n474_n140# a_594_n140# 0.02fF
C107 a_238_n140# a_n652_n140# 0.02fF
C108 a_238_n140# a_n296_n140# 0.04fF
C109 a_118_n194# a_296_n194# 0.10fF
C110 a_950_n140# a_n652_n140# 0.01fF
C111 a_950_n140# a_n296_n140# 0.02fF
C112 a_772_n140# a_416_n140# 0.06fF
C113 a_n1008_n140# a_n474_n140# 0.04fF
C114 a_474_n194# a_n594_n194# 0.01fF
C115 a_n772_n194# a_n238_n194# 0.02fF
C116 a_830_n194# a_118_n194# 0.01fF
C117 a_950_n140# VSUBS 0.02fF
C118 a_772_n140# VSUBS 0.02fF
C119 a_594_n140# VSUBS 0.02fF
C120 a_416_n140# VSUBS 0.02fF
C121 a_238_n140# VSUBS 0.02fF
C122 a_60_n140# VSUBS 0.02fF
C123 a_n118_n140# VSUBS 0.02fF
C124 a_n296_n140# VSUBS 0.02fF
C125 a_n474_n140# VSUBS 0.02fF
C126 a_n652_n140# VSUBS 0.02fF
C127 a_n830_n140# VSUBS 0.02fF
C128 a_n1008_n140# VSUBS 0.02fF
C129 a_830_n194# VSUBS 0.29fF
C130 a_652_n194# VSUBS 0.23fF
C131 a_474_n194# VSUBS 0.24fF
C132 a_296_n194# VSUBS 0.25fF
C133 a_118_n194# VSUBS 0.26fF
C134 a_n60_n194# VSUBS 0.27fF
C135 a_n238_n194# VSUBS 0.28fF
C136 a_n416_n194# VSUBS 0.28fF
C137 a_n594_n194# VSUBS 0.29fF
C138 a_n772_n194# VSUBS 0.29fF
C139 a_n950_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_UFQYRB a_1751_n140# a_n149_n194# a_1987_n194# a_n2819_n194#
+ a_n207_n140# a_n1809_n140# a_n2877_n140# a_207_n194# a_n2285_n194# a_1453_n194#
+ a_n1217_n194# a_n3353_n194# a_327_n140# a_n1275_n140# a_n2343_n140# a_2521_n194#
+ a_n861_n194# a_1573_n140# a_n3411_n140# a_2641_n140# a_n2699_n140# a_2877_n194#
+ a_1809_n194# a_2997_n140# a_n29_n140# a_n1039_n194# a_n3175_n194# a_1929_n140# a_149_n140#
+ a_n1097_n140# a_2343_n194# a_1275_n194# a_29_n194# a_n2107_n194# a_n2165_n140# a_n3233_n140#
+ a_3411_n194# a_n683_n194# a_1395_n140# a_3531_n140# a_2463_n140# a_n741_n140# a_2699_n194#
+ a_741_n194# a_n3589_n140# a_n1751_n194# a_861_n140# a_1097_n194# a_2819_n140# a_3233_n194#
+ a_2165_n194# a_n3055_n140# a_n505_n194# a_2285_n140# a_n563_n140# a_563_n194# a_3353_n140#
+ a_1217_n140# a_n1573_n194# a_n2641_n194# a_683_n140# a_n919_n140# a_n1631_n140#
+ a_919_n194# a_3055_n194# a_n2997_n194# a_n1987_n140# a_n327_n194# a_n1929_n194#
+ a_3175_n140# a_1039_n140# a_n385_n140# a_385_n194# a_2107_n140# a_n1395_n194# a_n2463_n194#
+ a_n3531_n194# a_505_n140# a_n1453_n140# a_1631_n194# a_n2521_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2165_n140# a_n2285_n194# a_n2343_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_3175_n140# a_3055_n194# a_2997_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n3233_n140# a_n3353_n194# a_n3411_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_2997_n140# a_2877_n194# a_2819_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1987_n140# a_n2107_n194# a_n2165_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1809_n140# a_n1929_n194# a_n1987_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n1453_n140# a_n1573_n194# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2463_n140# a_2343_n194# a_2285_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n2521_n140# a_n2641_n194# a_n2699_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_3531_n140# a_3411_n194# a_3353_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1751_n140# a_1631_n194# a_1573_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n3055_n140# a_n3175_n194# a_n3233_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_2819_n140# a_2699_n194# a_2641_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n2877_n140# a_n2997_n194# a_n3055_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_2285_n140# a_2165_n194# a_2107_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_n2699_n140# a_n2819_n194# a_n2877_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n2343_n140# a_n2463_n194# a_n2521_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_2107_n140# a_1987_n194# a_1929_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X31 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_3353_n140# a_3233_n194# a_3175_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_n3411_n140# a_n3531_n194# a_n3589_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X36 a_1573_n140# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_1929_n140# a_1809_n194# a_1751_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_n1631_n140# a_n1751_n194# a_n1809_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_2641_n140# a_2521_n194# a_2463_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_385_n194# a_1453_n194# 0.01fF
C1 a_919_n194# a_2521_n194# 0.01fF
C2 a_n919_n140# a_n1631_n140# 0.03fF
C3 a_n1217_n194# a_n1395_n194# 0.10fF
C4 a_n2343_n140# a_n3589_n140# 0.02fF
C5 a_3411_n194# a_2165_n194# 0.01fF
C6 a_2877_n194# a_1453_n194# 0.01fF
C7 a_2699_n194# a_1631_n194# 0.01fF
C8 a_1751_n140# a_683_n140# 0.02fF
C9 a_1453_n194# a_2521_n194# 0.01fF
C10 a_1809_n194# a_2165_n194# 0.03fF
C11 a_1631_n194# a_2343_n194# 0.01fF
C12 a_n3175_n194# a_n3531_n194# 0.03fF
C13 a_n1809_n140# a_n1097_n140# 0.03fF
C14 a_2641_n140# a_2997_n140# 0.06fF
C15 a_2641_n140# a_2107_n140# 0.04fF
C16 a_2819_n140# a_1929_n140# 0.02fF
C17 a_741_n194# a_207_n194# 0.02fF
C18 a_n1039_n194# a_n1573_n194# 0.02fF
C19 a_1395_n140# a_n29_n140# 0.01fF
C20 a_n3055_n140# a_n1631_n140# 0.01fF
C21 a_1395_n140# a_861_n140# 0.04fF
C22 a_n29_n140# a_n1275_n140# 0.02fF
C23 a_n207_n140# a_n1097_n140# 0.02fF
C24 a_149_n140# a_327_n140# 0.13fF
C25 a_n2877_n140# a_n2521_n140# 0.06fF
C26 a_n2641_n194# a_n3175_n194# 0.02fF
C27 a_1809_n194# a_563_n194# 0.01fF
C28 a_327_n140# a_1039_n140# 0.03fF
C29 a_n505_n194# a_207_n194# 0.01fF
C30 a_919_n194# a_1275_n194# 0.03fF
C31 a_n1039_n194# a_n505_n194# 0.02fF
C32 a_n563_n140# a_327_n140# 0.02fF
C33 a_n207_n140# a_505_n140# 0.03fF
C34 a_n1039_n194# a_n1929_n194# 0.01fF
C35 a_n2165_n140# a_n1987_n140# 0.13fF
C36 a_n2343_n140# a_n1809_n140# 0.04fF
C37 a_2285_n140# a_1039_n140# 0.02fF
C38 a_n2107_n194# a_n1395_n194# 0.01fF
C39 a_n2641_n194# a_n1217_n194# 0.01fF
C40 a_385_n194# a_1809_n194# 0.01fF
C41 a_1275_n194# a_1453_n194# 0.10fF
C42 a_n919_n140# a_n1275_n140# 0.06fF
C43 a_n563_n140# a_n1631_n140# 0.02fF
C44 a_n741_n140# a_n1453_n140# 0.03fF
C45 a_919_n194# a_n683_n194# 0.01fF
C46 a_3411_n194# a_2877_n194# 0.02fF
C47 a_1929_n140# a_327_n140# 0.01fF
C48 a_n2343_n140# a_n3233_n140# 0.02fF
C49 a_n1987_n140# a_n3589_n140# 0.01fF
C50 a_n2165_n140# a_n3411_n140# 0.02fF
C51 a_3411_n194# a_2521_n194# 0.01fF
C52 a_3055_n194# a_1631_n194# 0.01fF
C53 a_2877_n194# a_1809_n194# 0.01fF
C54 a_741_n194# a_1097_n194# 0.03fF
C55 a_1809_n194# a_2521_n194# 0.01fF
C56 a_1217_n140# a_2641_n140# 0.01fF
C57 a_2819_n140# a_3175_n140# 0.06fF
C58 a_207_n194# a_29_n194# 0.10fF
C59 a_2819_n140# a_2285_n140# 0.04fF
C60 a_3175_n140# a_1929_n140# 0.02fF
C61 a_2641_n140# a_2463_n140# 0.13fF
C62 a_1929_n140# a_2285_n140# 0.06fF
C63 a_2997_n140# a_2107_n140# 0.02fF
C64 a_n327_n194# a_207_n194# 0.02fF
C65 a_n1039_n194# a_29_n194# 0.01fF
C66 a_n2107_n194# a_n3531_n194# 0.01fF
C67 a_n1039_n194# a_n327_n194# 0.01fF
C68 a_n3589_n140# a_n3411_n140# 0.13fF
C69 a_n2699_n140# a_n1631_n140# 0.02fF
C70 a_1987_n194# a_2165_n194# 0.10fF
C71 a_n2877_n140# a_n1453_n140# 0.01fF
C72 a_1751_n140# a_861_n140# 0.02fF
C73 a_1097_n194# a_n505_n194# 0.01fF
C74 a_n1039_n194# a_n2463_n194# 0.01fF
C75 a_n2819_n194# a_n1395_n194# 0.01fF
C76 a_n2285_n194# a_n683_n194# 0.01fF
C77 a_n861_n194# a_n149_n194# 0.01fF
C78 a_n1573_n194# a_n1395_n194# 0.10fF
C79 a_n2107_n194# a_n2641_n194# 0.02fF
C80 a_919_n194# a_1453_n194# 0.02fF
C81 a_1395_n140# a_149_n140# 0.02fF
C82 a_1395_n140# a_1039_n140# 0.06fF
C83 a_149_n140# a_n1275_n140# 0.01fF
C84 a_n1987_n140# a_n1809_n140# 0.13fF
C85 a_1987_n194# a_563_n194# 0.01fF
C86 a_1217_n140# a_n385_n140# 0.01fF
C87 a_1275_n194# a_1809_n194# 0.02fF
C88 a_n741_n140# a_n1097_n140# 0.06fF
C89 a_n385_n140# a_n1453_n140# 0.02fF
C90 a_n2997_n194# a_n1395_n194# 0.01fF
C91 a_n563_n140# a_n1275_n140# 0.03fF
C92 a_n505_n194# a_n1395_n194# 0.01fF
C93 a_n1217_n194# a_n149_n194# 0.01fF
C94 a_n2819_n194# a_n3531_n194# 0.01fF
C95 a_741_n194# a_2343_n194# 0.01fF
C96 a_n1395_n194# a_n1929_n194# 0.02fF
C97 a_n207_n140# a_683_n140# 0.02fF
C98 a_3411_n194# a_3233_n194# 0.10fF
C99 a_1097_n194# a_29_n194# 0.01fF
C100 a_n1809_n140# a_n3411_n140# 0.01fF
C101 a_n1987_n140# a_n3233_n140# 0.02fF
C102 a_385_n194# a_1987_n194# 0.01fF
C103 a_3233_n194# a_1809_n194# 0.01fF
C104 a_1097_n194# a_n327_n194# 0.01fF
C105 a_n741_n140# a_505_n140# 0.02fF
C106 a_1395_n140# a_2819_n140# 0.01fF
C107 a_1573_n140# a_2641_n140# 0.02fF
C108 a_1395_n140# a_1929_n140# 0.04fF
C109 a_1217_n140# a_2107_n140# 0.02fF
C110 a_2997_n140# a_2463_n140# 0.04fF
C111 a_2107_n140# a_2463_n140# 0.06fF
C112 a_3175_n140# a_2285_n140# 0.02fF
C113 a_2877_n194# a_1987_n194# 0.01fF
C114 a_n2641_n194# a_n2819_n194# 0.10fF
C115 a_n2997_n194# a_n3531_n194# 0.02fF
C116 a_n3411_n140# a_n3233_n140# 0.13fF
C117 a_n2521_n140# a_n1453_n140# 0.02fF
C118 a_1987_n194# a_2521_n194# 0.02fF
C119 a_n2699_n140# a_n1275_n140# 0.01fF
C120 a_n2165_n140# a_n919_n140# 0.02fF
C121 a_n2343_n140# a_n741_n140# 0.01fF
C122 a_n1929_n194# a_n3531_n194# 0.01fF
C123 a_n2641_n194# a_n1573_n194# 0.01fF
C124 a_n1395_n194# a_29_n194# 0.01fF
C125 a_n1395_n194# a_n327_n194# 0.01fF
C126 a_919_n194# a_1809_n194# 0.01fF
C127 a_207_n194# a_563_n194# 0.03fF
C128 a_1751_n140# a_149_n140# 0.01fF
C129 a_n1751_n194# a_n683_n194# 0.01fF
C130 a_n2463_n194# a_n1395_n194# 0.01fF
C131 a_1751_n140# a_1039_n140# 0.03fF
C132 a_n1039_n194# a_563_n194# 0.01fF
C133 a_n2641_n194# a_n2997_n194# 0.03fF
C134 a_n2641_n194# a_n1929_n194# 0.01fF
C135 a_n385_n140# a_n1097_n140# 0.03fF
C136 a_1453_n194# a_1809_n194# 0.03fF
C137 a_n2343_n140# a_n2877_n140# 0.04fF
C138 a_n2165_n140# a_n3055_n140# 0.02fF
C139 a_385_n194# a_207_n194# 0.10fF
C140 a_1395_n140# a_327_n140# 0.02fF
C141 a_n1039_n194# a_385_n194# 0.01fF
C142 a_327_n140# a_n1275_n140# 0.01fF
C143 a_n1217_n194# a_n861_n194# 0.03fF
C144 a_n2285_n194# a_n3353_n194# 0.01fF
C145 a_1097_n194# a_2165_n194# 0.01fF
C146 a_1275_n194# a_1987_n194# 0.01fF
C147 a_n385_n140# a_505_n140# 0.02fF
C148 a_1751_n140# a_2819_n140# 0.02fF
C149 a_1573_n140# a_2997_n140# 0.01fF
C150 a_1217_n140# a_2463_n140# 0.02fF
C151 a_1751_n140# a_1929_n140# 0.13fF
C152 a_1395_n140# a_2285_n140# 0.02fF
C153 a_1573_n140# a_2107_n140# 0.04fF
C154 a_n2463_n194# a_n3531_n194# 0.01fF
C155 a_n207_n140# a_n29_n140# 0.13fF
C156 a_n1631_n140# a_n1275_n140# 0.06fF
C157 a_n3589_n140# a_n3055_n140# 0.04fF
C158 a_n207_n140# a_861_n140# 0.02fF
C159 a_3233_n194# a_1987_n194# 0.01fF
C160 a_n2521_n140# a_n1097_n140# 0.01fF
C161 a_n1809_n140# a_n919_n140# 0.02fF
C162 a_n1987_n140# a_n741_n140# 0.02fF
C163 a_n741_n140# a_683_n140# 0.01fF
C164 a_n2165_n140# a_n563_n140# 0.01fF
C165 a_741_n194# a_n149_n194# 0.01fF
C166 a_2107_n140# a_505_n140# 0.01fF
C167 a_1097_n194# a_563_n194# 0.02fF
C168 a_n2641_n194# a_n2463_n194# 0.10fF
C169 a_n1573_n194# a_n149_n194# 0.01fF
C170 a_n2285_n194# a_n1751_n194# 0.02fF
C171 a_n919_n140# a_n207_n140# 0.03fF
C172 a_3353_n140# a_3531_n140# 0.13fF
C173 a_1097_n194# a_385_n194# 0.01fF
C174 a_n505_n194# a_n149_n194# 0.03fF
C175 a_3411_n194# a_1809_n194# 0.01fF
C176 a_n2107_n194# a_n861_n194# 0.01fF
C177 a_919_n194# a_1987_n194# 0.01fF
C178 a_2699_n194# a_2165_n194# 0.02fF
C179 a_n2165_n140# a_n2699_n140# 0.04fF
C180 a_n1809_n140# a_n3055_n140# 0.02fF
C181 a_n2343_n140# a_n2521_n140# 0.13fF
C182 a_n1987_n140# a_n2877_n140# 0.02fF
C183 a_1275_n194# a_207_n194# 0.01fF
C184 a_n2107_n194# a_n3175_n194# 0.01fF
C185 a_1751_n140# a_327_n140# 0.01fF
C186 a_2165_n194# a_2343_n194# 0.10fF
C187 a_1097_n194# a_2521_n194# 0.01fF
C188 a_1217_n140# a_1573_n140# 0.06fF
C189 a_1751_n140# a_3175_n140# 0.01fF
C190 a_1453_n194# a_1987_n194# 0.02fF
C191 a_1751_n140# a_2285_n140# 0.04fF
C192 a_1573_n140# a_2463_n140# 0.02fF
C193 a_n1453_n140# a_n1097_n140# 0.06fF
C194 a_n2107_n194# a_n1217_n194# 0.01fF
C195 a_n3411_n140# a_n2877_n140# 0.04fF
C196 a_n3233_n140# a_n3055_n140# 0.13fF
C197 a_n3589_n140# a_n2699_n140# 0.02fF
C198 a_n3353_n194# a_n1751_n194# 0.01fF
C199 a_n683_n194# a_207_n194# 0.01fF
C200 a_n1039_n194# a_n683_n194# 0.03fF
C201 a_1217_n140# a_505_n140# 0.03fF
C202 a_n1809_n140# a_n563_n140# 0.02fF
C203 a_n1987_n140# a_n385_n140# 0.01fF
C204 a_n385_n140# a_683_n140# 0.02fF
C205 a_n149_n194# a_29_n194# 0.10fF
C206 a_n149_n194# a_n327_n194# 0.10fF
C207 a_n207_n140# a_149_n140# 0.06fF
C208 a_n207_n140# a_1039_n140# 0.02fF
C209 a_741_n194# a_n861_n194# 0.01fF
C210 a_n2819_n194# a_n3175_n194# 0.03fF
C211 a_n563_n140# a_n207_n140# 0.06fF
C212 a_n741_n140# a_n29_n140# 0.03fF
C213 a_n861_n194# a_n1573_n194# 0.01fF
C214 a_n741_n140# a_861_n140# 0.01fF
C215 a_919_n194# a_207_n194# 0.01fF
C216 a_741_n194# a_1631_n194# 0.01fF
C217 a_2107_n140# a_683_n140# 0.01fF
C218 a_n2343_n140# a_n1453_n140# 0.02fF
C219 a_n2165_n140# a_n1631_n140# 0.04fF
C220 a_n3175_n194# a_n1573_n194# 0.01fF
C221 a_1097_n194# a_1275_n194# 0.10fF
C222 a_2699_n194# a_2877_n194# 0.10fF
C223 a_2699_n194# a_2521_n194# 0.10fF
C224 a_3055_n194# a_2165_n194# 0.01fF
C225 a_2877_n194# a_2343_n194# 0.02fF
C226 a_n1809_n140# a_n2699_n140# 0.02fF
C227 a_n1987_n140# a_n2521_n140# 0.04fF
C228 a_n1217_n194# a_n2819_n194# 0.01fF
C229 a_2343_n194# a_2521_n194# 0.10fF
C230 a_n861_n194# a_n505_n194# 0.03fF
C231 a_1453_n194# a_207_n194# 0.01fF
C232 a_n2997_n194# a_n3175_n194# 0.10fF
C233 a_n861_n194# a_n1929_n194# 0.01fF
C234 a_3411_n194# a_1987_n194# 0.01fF
C235 a_n1217_n194# a_n1573_n194# 0.03fF
C236 a_1395_n140# a_1751_n140# 0.06fF
C237 a_n919_n140# a_n741_n140# 0.13fF
C238 a_1809_n194# a_1987_n194# 0.10fF
C239 a_n3175_n194# a_n1929_n194# 0.01fF
C240 a_n3233_n140# a_n2699_n140# 0.04fF
C241 a_n3411_n140# a_n2521_n140# 0.02fF
C242 a_3353_n140# a_2819_n140# 0.04fF
C243 a_3531_n140# a_2641_n140# 0.02fF
C244 a_3353_n140# a_1929_n140# 0.01fF
C245 a_n1217_n194# a_n505_n194# 0.01fF
C246 a_n1039_n194# a_n2285_n194# 0.01fF
C247 a_1573_n140# a_505_n140# 0.02fF
C248 a_n1217_n194# a_n1929_n194# 0.01fF
C249 a_n1097_n140# a_505_n140# 0.01fF
C250 a_919_n194# a_1097_n194# 0.10fF
C251 a_n861_n194# a_29_n194# 0.01fF
C252 a_n1395_n194# a_n683_n194# 0.01fF
C253 a_1275_n194# a_2699_n194# 0.01fF
C254 a_n861_n194# a_n327_n194# 0.02fF
C255 a_n385_n140# a_n29_n140# 0.06fF
C256 a_1275_n194# a_2343_n194# 0.01fF
C257 a_1631_n194# a_29_n194# 0.01fF
C258 a_1217_n140# a_683_n140# 0.04fF
C259 a_n385_n140# a_861_n140# 0.02fF
C260 a_n2107_n194# a_n2819_n194# 0.01fF
C261 a_n1987_n140# a_n1453_n140# 0.04fF
C262 a_n861_n194# a_n2463_n194# 0.01fF
C263 a_n2343_n140# a_n1097_n140# 0.02fF
C264 a_n2165_n140# a_n1275_n140# 0.02fF
C265 a_n1809_n140# a_n1631_n140# 0.13fF
C266 a_n207_n140# a_327_n140# 0.04fF
C267 a_2877_n194# a_3055_n194# 0.10fF
C268 a_2699_n194# a_3233_n194# 0.02fF
C269 a_n2463_n194# a_n3175_n194# 0.01fF
C270 a_1097_n194# a_1453_n194# 0.03fF
C271 a_n2107_n194# a_n1573_n194# 0.02fF
C272 a_n149_n194# a_563_n194# 0.01fF
C273 a_3055_n194# a_2521_n194# 0.02fF
C274 a_3233_n194# a_2343_n194# 0.01fF
C275 a_n1217_n194# a_29_n194# 0.01fF
C276 a_n741_n140# a_149_n140# 0.02fF
C277 a_n1217_n194# a_n327_n194# 0.01fF
C278 a_1809_n194# a_207_n194# 0.01fF
C279 a_n207_n140# a_n1631_n140# 0.01fF
C280 a_2107_n140# a_861_n140# 0.02fF
C281 a_n3233_n140# a_n1631_n140# 0.01fF
C282 a_n3055_n140# a_n2877_n140# 0.13fF
C283 a_n919_n140# a_n385_n140# 0.04fF
C284 a_n741_n140# a_n563_n140# 0.13fF
C285 a_n2107_n194# a_n505_n194# 0.01fF
C286 a_n2107_n194# a_n2997_n194# 0.01fF
C287 a_n1217_n194# a_n2463_n194# 0.01fF
C288 a_385_n194# a_n149_n194# 0.02fF
C289 a_n2107_n194# a_n1929_n194# 0.10fF
C290 a_3531_n140# a_2997_n140# 0.04fF
C291 a_3353_n140# a_3175_n140# 0.13fF
C292 a_3353_n140# a_2285_n140# 0.02fF
C293 a_3531_n140# a_2107_n140# 0.01fF
C294 a_2641_n140# a_1039_n140# 0.01fF
C295 a_919_n194# a_2343_n194# 0.01fF
C296 a_n1039_n194# a_n1751_n194# 0.01fF
C297 a_n2819_n194# a_n1573_n194# 0.01fF
C298 a_n2285_n194# a_n1395_n194# 0.01fF
C299 a_n2521_n140# a_n919_n140# 0.01fF
C300 a_2699_n194# a_1453_n194# 0.01fF
C301 a_1573_n140# a_683_n140# 0.02fF
C302 a_1453_n194# a_2343_n194# 0.01fF
C303 a_1631_n194# a_2165_n194# 0.02fF
C304 a_n1987_n140# a_n1097_n140# 0.02fF
C305 a_n1809_n140# a_n1275_n140# 0.04fF
C306 a_2641_n140# a_2819_n140# 0.13fF
C307 a_2641_n140# a_1929_n140# 0.03fF
C308 a_n2997_n194# a_n2819_n194# 0.10fF
C309 a_3055_n194# a_3233_n194# 0.10fF
C310 a_1097_n194# a_1809_n194# 0.01fF
C311 a_741_n194# a_n505_n194# 0.01fF
C312 a_n2819_n194# a_n1929_n194# 0.01fF
C313 a_n2107_n194# a_n2463_n194# 0.03fF
C314 a_1217_n140# a_n29_n140# 0.02fF
C315 a_1395_n140# a_n207_n140# 0.01fF
C316 a_n385_n140# a_149_n140# 0.04fF
C317 a_n2997_n194# a_n1573_n194# 0.01fF
C318 a_n505_n194# a_n1573_n194# 0.01fF
C319 a_505_n140# a_683_n140# 0.13fF
C320 a_1217_n140# a_861_n140# 0.06fF
C321 a_n385_n140# a_1039_n140# 0.01fF
C322 a_n207_n140# a_n1275_n140# 0.02fF
C323 a_n29_n140# a_n1453_n140# 0.01fF
C324 a_n861_n194# a_563_n194# 0.01fF
C325 a_2463_n140# a_861_n140# 0.01fF
C326 a_n1573_n194# a_n1929_n194# 0.03fF
C327 a_n2285_n194# a_n3531_n194# 0.01fF
C328 a_n563_n140# a_n385_n140# 0.13fF
C329 a_n3055_n140# a_n2521_n140# 0.04fF
C330 a_n2877_n140# a_n2699_n140# 0.13fF
C331 a_1631_n194# a_563_n194# 0.01fF
C332 a_1275_n194# a_n149_n194# 0.01fF
C333 a_3531_n140# a_2463_n140# 0.02fF
C334 a_n741_n140# a_327_n140# 0.02fF
C335 a_n861_n194# a_385_n194# 0.01fF
C336 a_n2343_n140# a_n1987_n140# 0.06fF
C337 a_n2997_n194# a_n1929_n194# 0.01fF
C338 a_n505_n194# a_n1929_n194# 0.01fF
C339 a_2107_n140# a_1039_n140# 0.02fF
C340 a_385_n194# a_1631_n194# 0.01fF
C341 a_n2641_n194# a_n2285_n194# 0.03fF
C342 a_n919_n140# a_n1453_n140# 0.04fF
C343 a_n741_n140# a_n1631_n140# 0.02fF
C344 a_741_n194# a_29_n194# 0.01fF
C345 a_n683_n194# a_n149_n194# 0.02fF
C346 a_741_n194# a_n327_n194# 0.01fF
C347 a_n1573_n194# a_29_n194# 0.01fF
C348 a_3411_n194# a_2699_n194# 0.01fF
C349 a_n2165_n140# a_n3589_n140# 0.01fF
C350 a_n2343_n140# a_n3411_n140# 0.02fF
C351 a_n2463_n194# a_n2819_n194# 0.03fF
C352 a_n1573_n194# a_n327_n194# 0.01fF
C353 a_3411_n194# a_2343_n194# 0.01fF
C354 a_n3353_n194# a_n3531_n194# 0.10fF
C355 a_3055_n194# a_1453_n194# 0.01fF
C356 a_2699_n194# a_1809_n194# 0.01fF
C357 a_2877_n194# a_1631_n194# 0.01fF
C358 a_n1217_n194# a_385_n194# 0.01fF
C359 a_1631_n194# a_2521_n194# 0.01fF
C360 a_1809_n194# a_2343_n194# 0.02fF
C361 a_n1751_n194# a_n1395_n194# 0.03fF
C362 a_n2463_n194# a_n1573_n194# 0.01fF
C363 a_2641_n140# a_3175_n140# 0.04fF
C364 a_2819_n140# a_2997_n140# 0.13fF
C365 a_2819_n140# a_2107_n140# 0.03fF
C366 a_1929_n140# a_2107_n140# 0.13fF
C367 a_2641_n140# a_2285_n140# 0.06fF
C368 a_2997_n140# a_1929_n140# 0.02fF
C369 a_n505_n194# a_29_n194# 0.02fF
C370 a_n505_n194# a_n327_n194# 0.10fF
C371 a_1573_n140# a_n29_n140# 0.01fF
C372 a_n2877_n140# a_n1631_n140# 0.02fF
C373 a_919_n194# a_n149_n194# 0.01fF
C374 a_n3055_n140# a_n1453_n140# 0.01fF
C375 a_1573_n140# a_861_n140# 0.03fF
C376 a_n1929_n194# a_n327_n194# 0.01fF
C377 a_n29_n140# a_n1097_n140# 0.02fF
C378 a_n2997_n194# a_n2463_n194# 0.02fF
C379 a_n2641_n194# a_n3353_n194# 0.01fF
C380 a_1097_n194# a_1987_n194# 0.01fF
C381 a_n2699_n140# a_n2521_n140# 0.13fF
C382 a_n2463_n194# a_n1929_n194# 0.02fF
C383 a_n1039_n194# a_207_n194# 0.01fF
C384 a_1751_n140# a_3353_n140# 0.01fF
C385 a_n149_n194# a_1453_n194# 0.01fF
C386 a_1217_n140# a_149_n140# 0.02fF
C387 a_n385_n140# a_327_n140# 0.03fF
C388 a_n29_n140# a_505_n140# 0.04fF
C389 a_149_n140# a_n1453_n140# 0.01fF
C390 a_505_n140# a_861_n140# 0.06fF
C391 a_1217_n140# a_1039_n140# 0.13fF
C392 a_n2165_n140# a_n1809_n140# 0.06fF
C393 a_2463_n140# a_1039_n140# 0.01fF
C394 a_1275_n194# a_1631_n194# 0.03fF
C395 a_n563_n140# a_n1453_n140# 0.02fF
C396 a_n741_n140# a_n1275_n140# 0.04fF
C397 a_n385_n140# a_n1631_n140# 0.02fF
C398 a_n919_n140# a_n1097_n140# 0.13fF
C399 a_n327_n194# a_29_n194# 0.03fF
C400 a_741_n194# a_2165_n194# 0.01fF
C401 a_3411_n194# a_3055_n194# 0.03fF
C402 a_n1987_n140# a_n3411_n140# 0.01fF
C403 a_n2165_n140# a_n3233_n140# 0.02fF
C404 a_n2641_n194# a_n1751_n194# 0.01fF
C405 a_3233_n194# a_1631_n194# 0.01fF
C406 a_3055_n194# a_1809_n194# 0.01fF
C407 a_n861_n194# a_n683_n194# 0.10fF
C408 a_n919_n140# a_505_n140# 0.01fF
C409 a_1217_n140# a_2819_n140# 0.01fF
C410 a_1395_n140# a_2641_n140# 0.02fF
C411 a_1217_n140# a_1929_n140# 0.03fF
C412 a_2997_n140# a_3175_n140# 0.13fF
C413 a_2997_n140# a_2285_n140# 0.03fF
C414 a_2819_n140# a_2463_n140# 0.06fF
C415 a_1929_n140# a_2463_n140# 0.04fF
C416 a_3175_n140# a_2107_n140# 0.02fF
C417 a_2107_n140# a_2285_n140# 0.13fF
C418 a_2699_n194# a_1987_n194# 0.01fF
C419 a_1097_n194# a_207_n194# 0.01fF
C420 a_n3589_n140# a_n3233_n140# 0.06fF
C421 a_1987_n194# a_2343_n194# 0.03fF
C422 a_n2521_n140# a_n1631_n140# 0.02fF
C423 a_n2877_n140# a_n1275_n140# 0.01fF
C424 a_n2699_n140# a_n1453_n140# 0.02fF
C425 a_741_n194# a_563_n194# 0.10fF
C426 a_n2343_n140# a_n919_n140# 0.01fF
C427 a_n1217_n194# a_n683_n194# 0.02fF
C428 a_919_n194# a_1631_n194# 0.01fF
C429 a_1573_n140# a_149_n140# 0.01fF
C430 a_741_n194# a_385_n194# 0.03fF
C431 a_1573_n140# a_1039_n140# 0.04fF
C432 a_149_n140# a_n1097_n140# 0.02fF
C433 a_n505_n194# a_563_n194# 0.01fF
C434 a_n1395_n194# a_207_n194# 0.01fF
C435 a_n1039_n194# a_n1395_n194# 0.03fF
C436 a_n385_n140# a_n1275_n140# 0.02fF
C437 a_n563_n140# a_n1097_n140# 0.04fF
C438 a_1453_n194# a_1631_n194# 0.10fF
C439 a_n2343_n140# a_n3055_n140# 0.03fF
C440 a_n29_n140# a_683_n140# 0.03fF
C441 a_1217_n140# a_327_n140# 0.02fF
C442 a_149_n140# a_505_n140# 0.06fF
C443 a_n1809_n140# a_n207_n140# 0.01fF
C444 a_505_n140# a_1039_n140# 0.04fF
C445 a_683_n140# a_861_n140# 0.13fF
C446 a_385_n194# a_n505_n194# 0.01fF
C447 a_n1809_n140# a_n3233_n140# 0.01fF
C448 a_n2285_n194# a_n861_n194# 0.01fF
C449 a_n563_n140# a_505_n140# 0.02fF
C450 a_n1751_n194# a_n149_n194# 0.01fF
C451 a_1395_n140# a_2997_n140# 0.01fF
C452 a_1573_n140# a_2819_n140# 0.02fF
C453 a_1751_n140# a_2641_n140# 0.02fF
C454 a_1217_n140# a_2285_n140# 0.02fF
C455 a_n2285_n194# a_n3175_n194# 0.01fF
C456 a_1573_n140# a_1929_n140# 0.06fF
C457 a_1395_n140# a_2107_n140# 0.03fF
C458 a_3175_n140# a_2463_n140# 0.03fF
C459 a_2285_n140# a_2463_n140# 0.13fF
C460 a_n1631_n140# a_n1453_n140# 0.13fF
C461 a_n2107_n194# a_n683_n194# 0.01fF
C462 a_3055_n194# a_1987_n194# 0.01fF
C463 a_29_n194# a_563_n194# 0.02fF
C464 a_n2699_n140# a_n1097_n140# 0.01fF
C465 a_n2521_n140# a_n1275_n140# 0.02fF
C466 a_n327_n194# a_563_n194# 0.01fF
C467 a_n2165_n140# a_n741_n140# 0.01fF
C468 a_n1987_n140# a_n919_n140# 0.02fF
C469 a_n919_n140# a_683_n140# 0.01fF
C470 a_n1217_n194# a_n2285_n194# 0.01fF
C471 a_1929_n140# a_505_n140# 0.01fF
C472 a_385_n194# a_29_n194# 0.03fF
C473 a_741_n194# a_1275_n194# 0.02fF
C474 a_385_n194# a_n327_n194# 0.01fF
C475 a_n2641_n194# a_n1039_n194# 0.01fF
C476 a_n3353_n194# a_n3175_n194# 0.10fF
C477 a_1631_n194# a_1809_n194# 0.10fF
C478 a_n2343_n140# a_n2699_n140# 0.06fF
C479 a_n1987_n140# a_n3055_n140# 0.02fF
C480 a_n2165_n140# a_n2877_n140# 0.03fF
C481 a_1573_n140# a_327_n140# 0.02fF
C482 a_327_n140# a_n1097_n140# 0.01fF
C483 a_1097_n194# a_2699_n194# 0.01fF
C484 a_741_n194# a_n683_n194# 0.01fF
C485 a_1097_n194# a_2343_n194# 0.01fF
C486 a_1217_n140# a_1395_n140# 0.13fF
C487 a_n1573_n194# a_n683_n194# 0.01fF
C488 a_1751_n140# a_2997_n140# 0.02fF
C489 a_1573_n140# a_3175_n140# 0.01fF
C490 a_1395_n140# a_2463_n140# 0.02fF
C491 a_1751_n140# a_2107_n140# 0.06fF
C492 a_1573_n140# a_2285_n140# 0.03fF
C493 a_n1453_n140# a_n1275_n140# 0.13fF
C494 a_n1631_n140# a_n1097_n140# 0.04fF
C495 a_n3411_n140# a_n3055_n140# 0.06fF
C496 a_n3589_n140# a_n2877_n140# 0.03fF
C497 a_n861_n194# a_n1751_n194# 0.01fF
C498 a_n2107_n194# a_n2285_n194# 0.10fF
C499 a_327_n140# a_505_n140# 0.13fF
C500 a_n29_n140# a_861_n140# 0.02fF
C501 a_149_n140# a_683_n140# 0.04fF
C502 a_683_n140# a_1039_n140# 0.06fF
C503 a_n1751_n194# a_n3175_n194# 0.01fF
C504 a_n505_n194# a_n683_n194# 0.10fF
C505 a_2165_n194# a_563_n194# 0.01fF
C506 a_n1809_n140# a_n741_n140# 0.02fF
C507 a_n1987_n140# a_n563_n140# 0.01fF
C508 a_n563_n140# a_683_n140# 0.02fF
C509 a_741_n194# a_919_n194# 0.10fF
C510 a_n683_n194# a_n1929_n194# 0.01fF
C511 a_n1217_n194# a_n1751_n194# 0.02fF
C512 a_1275_n194# a_29_n194# 0.01fF
C513 a_n741_n140# a_n207_n140# 0.04fF
C514 a_n919_n140# a_n29_n140# 0.02fF
C515 a_1275_n194# a_n327_n194# 0.01fF
C516 a_741_n194# a_1453_n194# 0.01fF
C517 a_n149_n194# a_207_n194# 0.03fF
C518 a_1929_n140# a_683_n140# 0.02fF
C519 a_n2343_n140# a_n1631_n140# 0.03fF
C520 a_919_n194# a_n505_n194# 0.01fF
C521 a_n1039_n194# a_n149_n194# 0.01fF
C522 a_n2107_n194# a_n3353_n194# 0.01fF
C523 a_2699_n194# a_2343_n194# 0.03fF
C524 a_2877_n194# a_2165_n194# 0.01fF
C525 a_n2165_n140# a_n2521_n140# 0.06fF
C526 a_n1987_n140# a_n2699_n140# 0.03fF
C527 a_n1809_n140# a_n2877_n140# 0.02fF
C528 a_n2285_n194# a_n2819_n194# 0.02fF
C529 a_2165_n194# a_2521_n194# 0.03fF
C530 a_n2641_n194# a_n1395_n194# 0.01fF
C531 a_n683_n194# a_29_n194# 0.01fF
C532 a_n683_n194# a_n327_n194# 0.03fF
C533 a_385_n194# a_563_n194# 0.10fF
C534 a_1217_n140# a_1751_n140# 0.04fF
C535 a_n2285_n194# a_n1573_n194# 0.01fF
C536 a_1395_n140# a_1573_n140# 0.13fF
C537 a_1631_n194# a_1987_n194# 0.03fF
C538 a_1751_n140# a_2463_n140# 0.03fF
C539 a_n1275_n140# a_n1097_n140# 0.13fF
C540 a_n3589_n140# a_n2521_n140# 0.02fF
C541 a_n3411_n140# a_n2699_n140# 0.03fF
C542 a_n3233_n140# a_n2877_n140# 0.06fF
C543 a_3353_n140# a_2641_n140# 0.03fF
C544 a_n2997_n194# a_n2285_n194# 0.01fF
C545 a_919_n194# a_29_n194# 0.01fF
C546 a_n1809_n140# a_n385_n140# 0.01fF
C547 a_1395_n140# a_505_n140# 0.02fF
C548 a_n2107_n194# a_n1751_n194# 0.03fF
C549 a_n2285_n194# a_n1929_n194# 0.03fF
C550 a_919_n194# a_n327_n194# 0.01fF
C551 a_n2641_n194# a_n3531_n194# 0.01fF
C552 a_n29_n140# a_149_n140# 0.13fF
C553 a_n3353_n194# a_n2819_n194# 0.02fF
C554 a_149_n140# a_861_n140# 0.03fF
C555 a_327_n140# a_683_n140# 0.06fF
C556 a_n29_n140# a_1039_n140# 0.02fF
C557 a_1097_n194# a_n149_n194# 0.01fF
C558 a_861_n140# a_1039_n140# 0.13fF
C559 a_n385_n140# a_n207_n140# 0.13fF
C560 a_n563_n140# a_n29_n140# 0.04fF
C561 a_1275_n194# a_2165_n194# 0.01fF
C562 a_1453_n194# a_29_n194# 0.01fF
C563 a_n563_n140# a_861_n140# 0.01fF
C564 a_741_n194# a_1809_n194# 0.01fF
C565 a_2285_n140# a_683_n140# 0.01fF
C566 a_n2165_n140# a_n1453_n140# 0.03fF
C567 a_n1987_n140# a_n1631_n140# 0.06fF
C568 a_n2343_n140# a_n1275_n140# 0.02fF
C569 a_2699_n194# a_3055_n194# 0.03fF
C570 a_n861_n194# a_207_n194# 0.01fF
C571 a_2877_n194# a_2521_n194# 0.03fF
C572 a_3055_n194# a_2343_n194# 0.01fF
C573 a_3233_n194# a_2165_n194# 0.01fF
C574 a_n1809_n140# a_n2521_n140# 0.03fF
C575 a_n2997_n194# a_n3353_n194# 0.03fF
C576 a_n1039_n194# a_n861_n194# 0.10fF
C577 a_n919_n140# a_149_n140# 0.02fF
C578 a_1631_n194# a_207_n194# 0.01fF
C579 a_n1395_n194# a_n149_n194# 0.01fF
C580 a_1929_n140# a_861_n140# 0.02fF
C581 a_n3353_n194# a_n1929_n194# 0.01fF
C582 a_1275_n194# a_563_n194# 0.01fF
C583 a_1573_n140# a_1751_n140# 0.13fF
C584 a_n919_n140# a_n563_n140# 0.06fF
C585 a_n1751_n194# a_n2819_n194# 0.01fF
C586 a_n2285_n194# a_n2463_n194# 0.10fF
C587 a_n3233_n140# a_n2521_n140# 0.03fF
C588 a_3353_n140# a_2997_n140# 0.06fF
C589 a_n1217_n194# a_207_n194# 0.01fF
C590 a_3531_n140# a_2819_n140# 0.03fF
C591 a_3531_n140# a_1929_n140# 0.01fF
C592 a_3353_n140# a_2107_n140# 0.02fF
C593 a_n1751_n194# a_n1573_n194# 0.10fF
C594 a_n1217_n194# a_n1039_n194# 0.10fF
C595 a_1275_n194# a_385_n194# 0.01fF
C596 a_1751_n140# a_505_n140# 0.02fF
C597 a_n683_n194# a_563_n194# 0.01fF
C598 a_919_n194# a_2165_n194# 0.01fF
C599 a_n2997_n194# a_n1751_n194# 0.01fF
C600 a_n505_n194# a_n1751_n194# 0.01fF
C601 a_1275_n194# a_2877_n194# 0.01fF
C602 a_n1751_n194# a_n1929_n194# 0.10fF
C603 a_1275_n194# a_2521_n194# 0.01fF
C604 a_1395_n140# a_683_n140# 0.03fF
C605 a_1453_n194# a_2165_n194# 0.01fF
C606 a_385_n194# a_n683_n194# 0.01fF
C607 a_n2463_n194# a_n3353_n194# 0.01fF
C608 a_n1987_n140# a_n1275_n140# 0.03fF
C609 a_n1809_n140# a_n1453_n140# 0.06fF
C610 a_n2165_n140# a_n1097_n140# 0.02fF
C611 a_n29_n140# a_327_n140# 0.06fF
C612 a_2877_n194# a_3233_n194# 0.03fF
C613 a_149_n140# a_1039_n140# 0.02fF
C614 a_1097_n194# a_1631_n194# 0.02fF
C615 a_327_n140# a_861_n140# 0.04fF
C616 a_919_n194# a_563_n194# 0.03fF
C617 a_3233_n194# a_2521_n194# 0.01fF
C618 a_741_n194# a_1987_n194# 0.01fF
C619 a_n563_n140# a_149_n140# 0.03fF
C620 a_1217_n140# a_n207_n140# 0.01fF
C621 a_n563_n140# a_1039_n140# 0.01fF
C622 a_n207_n140# a_n1453_n140# 0.02fF
C623 a_n29_n140# a_n1631_n140# 0.01fF
C624 a_2285_n140# a_861_n140# 0.01fF
C625 a_n741_n140# a_n385_n140# 0.06fF
C626 a_n2107_n194# a_n1039_n194# 0.01fF
C627 a_n3055_n140# a_n2699_n140# 0.06fF
C628 a_1453_n194# a_563_n194# 0.01fF
C629 a_919_n194# a_385_n194# 0.02fF
C630 a_n861_n194# a_n1395_n194# 0.02fF
C631 a_n1751_n194# a_n327_n194# 0.01fF
C632 a_3531_n140# a_3175_n140# 0.06fF
C633 a_3531_n140# a_2285_n140# 0.02fF
C634 a_3353_n140# a_2463_n140# 0.02fF
C635 a_n919_n140# a_327_n140# 0.02fF
C636 a_n2343_n140# a_n2165_n140# 0.13fF
C637 a_1929_n140# a_1039_n140# 0.02fF
C638 a_n2463_n194# a_n1751_n194# 0.01fF
C639 a_3531_n140# VSUBS 0.02fF
C640 a_3353_n140# VSUBS 0.02fF
C641 a_3175_n140# VSUBS 0.02fF
C642 a_2997_n140# VSUBS 0.02fF
C643 a_2819_n140# VSUBS 0.02fF
C644 a_2641_n140# VSUBS 0.02fF
C645 a_2463_n140# VSUBS 0.02fF
C646 a_2285_n140# VSUBS 0.02fF
C647 a_2107_n140# VSUBS 0.02fF
C648 a_1929_n140# VSUBS 0.02fF
C649 a_1751_n140# VSUBS 0.02fF
C650 a_1573_n140# VSUBS 0.02fF
C651 a_1395_n140# VSUBS 0.02fF
C652 a_1217_n140# VSUBS 0.02fF
C653 a_1039_n140# VSUBS 0.02fF
C654 a_861_n140# VSUBS 0.02fF
C655 a_683_n140# VSUBS 0.02fF
C656 a_505_n140# VSUBS 0.02fF
C657 a_327_n140# VSUBS 0.02fF
C658 a_149_n140# VSUBS 0.02fF
C659 a_n29_n140# VSUBS 0.02fF
C660 a_n207_n140# VSUBS 0.02fF
C661 a_n385_n140# VSUBS 0.02fF
C662 a_n563_n140# VSUBS 0.02fF
C663 a_n741_n140# VSUBS 0.02fF
C664 a_n919_n140# VSUBS 0.02fF
C665 a_n1097_n140# VSUBS 0.02fF
C666 a_n1275_n140# VSUBS 0.02fF
C667 a_n1453_n140# VSUBS 0.02fF
C668 a_n1631_n140# VSUBS 0.02fF
C669 a_n1809_n140# VSUBS 0.02fF
C670 a_n1987_n140# VSUBS 0.02fF
C671 a_n2165_n140# VSUBS 0.02fF
C672 a_n2343_n140# VSUBS 0.02fF
C673 a_n2521_n140# VSUBS 0.02fF
C674 a_n2699_n140# VSUBS 0.02fF
C675 a_n2877_n140# VSUBS 0.02fF
C676 a_n3055_n140# VSUBS 0.02fF
C677 a_n3233_n140# VSUBS 0.02fF
C678 a_n3411_n140# VSUBS 0.02fF
C679 a_n3589_n140# VSUBS 0.02fF
C680 a_3411_n194# VSUBS 0.29fF
C681 a_3233_n194# VSUBS 0.23fF
C682 a_3055_n194# VSUBS 0.24fF
C683 a_2877_n194# VSUBS 0.25fF
C684 a_2699_n194# VSUBS 0.26fF
C685 a_2521_n194# VSUBS 0.27fF
C686 a_2343_n194# VSUBS 0.28fF
C687 a_2165_n194# VSUBS 0.28fF
C688 a_1987_n194# VSUBS 0.29fF
C689 a_1809_n194# VSUBS 0.29fF
C690 a_1631_n194# VSUBS 0.29fF
C691 a_1453_n194# VSUBS 0.29fF
C692 a_1275_n194# VSUBS 0.29fF
C693 a_1097_n194# VSUBS 0.29fF
C694 a_919_n194# VSUBS 0.29fF
C695 a_741_n194# VSUBS 0.29fF
C696 a_563_n194# VSUBS 0.29fF
C697 a_385_n194# VSUBS 0.29fF
C698 a_207_n194# VSUBS 0.29fF
C699 a_29_n194# VSUBS 0.29fF
C700 a_n149_n194# VSUBS 0.29fF
C701 a_n327_n194# VSUBS 0.29fF
C702 a_n505_n194# VSUBS 0.29fF
C703 a_n683_n194# VSUBS 0.29fF
C704 a_n861_n194# VSUBS 0.29fF
C705 a_n1039_n194# VSUBS 0.29fF
C706 a_n1217_n194# VSUBS 0.29fF
C707 a_n1395_n194# VSUBS 0.29fF
C708 a_n1573_n194# VSUBS 0.29fF
C709 a_n1751_n194# VSUBS 0.29fF
C710 a_n1929_n194# VSUBS 0.29fF
C711 a_n2107_n194# VSUBS 0.29fF
C712 a_n2285_n194# VSUBS 0.29fF
C713 a_n2463_n194# VSUBS 0.29fF
C714 a_n2641_n194# VSUBS 0.29fF
C715 a_n2819_n194# VSUBS 0.29fF
C716 a_n2997_n194# VSUBS 0.29fF
C717 a_n3175_n194# VSUBS 0.29fF
C718 a_n3353_n194# VSUBS 0.29fF
C719 a_n3531_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_7P4E2J a_n149_n194# a_n207_n140# a_207_n194# a_n1217_n194#
+ a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140# a_n1097_n140#
+ a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194# a_861_n140#
+ a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140# a_n919_n140#
+ a_919_n194# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194# a_n1395_n194# a_505_n140#
+ a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n741_n140# a_n563_n140# 0.13fF
C1 a_n385_n140# a_149_n140# 0.04fF
C2 a_149_n140# a_1039_n140# 0.02fF
C3 a_n149_n194# a_741_n194# 0.01fF
C4 a_1217_n140# a_861_n140# 0.06fF
C5 a_n861_n194# a_n1217_n194# 0.03fF
C6 a_n861_n194# a_n505_n194# 0.03fF
C7 a_n1039_n194# a_n327_n194# 0.01fF
C8 a_n207_n140# a_n563_n140# 0.06fF
C9 a_29_n194# a_563_n194# 0.02fF
C10 a_1275_n194# a_1097_n194# 0.10fF
C11 a_1097_n194# a_385_n194# 0.01fF
C12 a_n1097_n140# a_n563_n140# 0.04fF
C13 a_n385_n140# a_n1275_n140# 0.02fF
C14 a_n327_n194# a_1097_n194# 0.01fF
C15 a_n385_n140# a_n29_n140# 0.06fF
C16 a_n29_n140# a_1039_n140# 0.02fF
C17 a_327_n140# a_861_n140# 0.04fF
C18 a_505_n140# a_1217_n140# 0.03fF
C19 a_327_n140# a_n919_n140# 0.02fF
C20 a_207_n194# a_n861_n194# 0.01fF
C21 a_n1217_n194# a_n505_n194# 0.01fF
C22 a_n861_n194# a_n683_n194# 0.10fF
C23 a_n149_n194# a_563_n194# 0.01fF
C24 a_29_n194# a_1275_n194# 0.01fF
C25 a_29_n194# a_385_n194# 0.03fF
C26 a_149_n140# a_1395_n140# 0.02fF
C27 a_327_n140# a_505_n140# 0.13fF
C28 a_207_n194# a_n1217_n194# 0.01fF
C29 a_29_n194# a_n1039_n194# 0.01fF
C30 a_207_n194# a_n505_n194# 0.01fF
C31 a_29_n194# a_n327_n194# 0.03fF
C32 a_n505_n194# a_n683_n194# 0.10fF
C33 a_n1217_n194# a_n683_n194# 0.02fF
C34 a_149_n140# a_n1453_n140# 0.01fF
C35 a_n385_n140# a_861_n140# 0.02fF
C36 a_1039_n140# a_861_n140# 0.13fF
C37 a_n385_n140# a_n919_n140# 0.04fF
C38 a_149_n140# a_683_n140# 0.04fF
C39 a_n149_n194# a_1275_n194# 0.01fF
C40 a_n149_n194# a_385_n194# 0.02fF
C41 a_149_n140# a_n741_n140# 0.02fF
C42 a_n29_n140# a_1395_n140# 0.01fF
C43 a_327_n140# a_1217_n140# 0.02fF
C44 a_29_n194# a_1097_n194# 0.01fF
C45 a_n149_n194# a_n1039_n194# 0.01fF
C46 a_n149_n194# a_n327_n194# 0.10fF
C47 a_207_n194# a_n683_n194# 0.01fF
C48 a_n1275_n140# a_n1453_n140# 0.13fF
C49 a_149_n140# a_n207_n140# 0.06fF
C50 a_n385_n140# a_505_n140# 0.02fF
C51 a_n29_n140# a_n1453_n140# 0.01fF
C52 a_505_n140# a_1039_n140# 0.04fF
C53 a_n505_n194# a_919_n194# 0.01fF
C54 a_n29_n140# a_683_n140# 0.03fF
C55 a_n741_n140# a_n1275_n140# 0.04fF
C56 a_149_n140# a_n1097_n140# 0.02fF
C57 a_n29_n140# a_n741_n140# 0.03fF
C58 a_n861_n194# a_741_n194# 0.01fF
C59 a_n149_n194# a_1097_n194# 0.01fF
C60 a_1395_n140# a_861_n140# 0.04fF
C61 a_n385_n140# a_1217_n140# 0.01fF
C62 a_1217_n140# a_1039_n140# 0.13fF
C63 a_n207_n140# a_n1275_n140# 0.02fF
C64 a_n29_n140# a_n207_n140# 0.13fF
C65 a_207_n194# a_919_n194# 0.01fF
C66 a_n683_n194# a_919_n194# 0.01fF
C67 a_n919_n140# a_n1453_n140# 0.04fF
C68 a_n1097_n140# a_n1275_n140# 0.13fF
C69 a_n29_n140# a_n1097_n140# 0.02fF
C70 a_n505_n194# a_741_n194# 0.01fF
C71 a_683_n140# a_861_n140# 0.13fF
C72 a_683_n140# a_n919_n140# 0.01fF
C73 a_1395_n140# a_505_n140# 0.02fF
C74 a_n385_n140# a_327_n140# 0.03fF
C75 a_n741_n140# a_861_n140# 0.01fF
C76 a_327_n140# a_1039_n140# 0.03fF
C77 a_n861_n194# a_563_n194# 0.01fF
C78 a_149_n140# a_n563_n140# 0.03fF
C79 a_29_n194# a_n149_n194# 0.10fF
C80 a_n741_n140# a_n919_n140# 0.13fF
C81 a_n1395_n194# a_n327_n194# 0.01fF
C82 a_n1395_n194# a_n1039_n194# 0.03fF
C83 a_n207_n140# a_861_n140# 0.02fF
C84 a_n207_n140# a_n919_n140# 0.03fF
C85 a_207_n194# a_741_n194# 0.02fF
C86 a_n683_n194# a_741_n194# 0.01fF
C87 a_683_n140# a_505_n140# 0.13fF
C88 a_1395_n140# a_1217_n140# 0.13fF
C89 a_505_n140# a_n741_n140# 0.02fF
C90 a_n1275_n140# a_n563_n140# 0.03fF
C91 a_n505_n194# a_563_n194# 0.01fF
C92 a_n29_n140# a_n563_n140# 0.04fF
C93 a_n919_n140# a_n1097_n140# 0.13fF
C94 a_n861_n194# a_385_n194# 0.01fF
C95 a_n385_n140# a_1039_n140# 0.01fF
C96 a_n207_n140# a_505_n140# 0.03fF
C97 a_683_n140# a_1217_n140# 0.04fF
C98 a_327_n140# a_1395_n140# 0.02fF
C99 a_n861_n194# a_n1039_n194# 0.10fF
C100 a_n861_n194# a_n327_n194# 0.02fF
C101 a_505_n140# a_n1097_n140# 0.01fF
C102 a_919_n194# a_741_n194# 0.10fF
C103 a_207_n194# a_563_n194# 0.03fF
C104 a_n683_n194# a_563_n194# 0.01fF
C105 a_29_n194# a_n1395_n194# 0.01fF
C106 a_n207_n140# a_1217_n140# 0.01fF
C107 a_n1217_n194# a_385_n194# 0.01fF
C108 a_n505_n194# a_385_n194# 0.01fF
C109 a_n563_n140# a_861_n140# 0.01fF
C110 a_n919_n140# a_n563_n140# 0.06fF
C111 a_327_n140# a_683_n140# 0.06fF
C112 a_327_n140# a_n741_n140# 0.02fF
C113 a_n1039_n194# a_n1217_n194# 0.10fF
C114 a_n327_n194# a_n505_n194# 0.10fF
C115 a_n1217_n194# a_n327_n194# 0.01fF
C116 a_n1039_n194# a_n505_n194# 0.02fF
C117 a_1395_n140# a_1039_n140# 0.06fF
C118 a_n149_n194# a_n1395_n194# 0.01fF
C119 a_327_n140# a_n207_n140# 0.04fF
C120 a_207_n194# a_1275_n194# 0.01fF
C121 a_207_n194# a_385_n194# 0.10fF
C122 a_919_n194# a_563_n194# 0.03fF
C123 a_505_n140# a_n563_n140# 0.02fF
C124 a_n683_n194# a_385_n194# 0.01fF
C125 a_n385_n140# a_n1453_n140# 0.02fF
C126 a_n505_n194# a_1097_n194# 0.01fF
C127 a_327_n140# a_n1097_n140# 0.01fF
C128 a_29_n194# a_n861_n194# 0.01fF
C129 a_207_n194# a_n1039_n194# 0.01fF
C130 a_207_n194# a_n327_n194# 0.02fF
C131 a_n327_n194# a_n683_n194# 0.03fF
C132 a_n1039_n194# a_n683_n194# 0.03fF
C133 a_149_n140# a_n1275_n140# 0.01fF
C134 a_n385_n140# a_683_n140# 0.02fF
C135 a_683_n140# a_1039_n140# 0.06fF
C136 a_149_n140# a_n29_n140# 0.13fF
C137 a_n385_n140# a_n741_n140# 0.06fF
C138 a_n385_n140# a_n207_n140# 0.13fF
C139 a_n207_n140# a_1039_n140# 0.02fF
C140 a_207_n194# a_1097_n194# 0.01fF
C141 a_1275_n194# a_919_n194# 0.03fF
C142 a_741_n194# a_563_n194# 0.10fF
C143 a_919_n194# a_385_n194# 0.02fF
C144 a_29_n194# a_n1217_n194# 0.01fF
C145 a_n149_n194# a_n861_n194# 0.01fF
C146 a_29_n194# a_n505_n194# 0.02fF
C147 a_n29_n140# a_n1275_n140# 0.02fF
C148 a_n385_n140# a_n1097_n140# 0.03fF
C149 a_n327_n194# a_919_n194# 0.01fF
C150 a_327_n140# a_n563_n140# 0.02fF
C151 a_149_n140# a_861_n140# 0.03fF
C152 a_149_n140# a_n919_n140# 0.02fF
C153 a_1395_n140# a_683_n140# 0.03fF
C154 a_207_n194# a_29_n194# 0.10fF
C155 a_n149_n194# a_n1217_n194# 0.01fF
C156 a_n149_n194# a_n505_n194# 0.03fF
C157 a_29_n194# a_n683_n194# 0.01fF
C158 a_1097_n194# a_919_n194# 0.10fF
C159 a_1275_n194# a_741_n194# 0.02fF
C160 a_741_n194# a_385_n194# 0.03fF
C161 a_149_n140# a_505_n140# 0.06fF
C162 a_n29_n140# a_861_n140# 0.02fF
C163 a_1395_n140# a_n207_n140# 0.01fF
C164 a_n919_n140# a_n1275_n140# 0.06fF
C165 a_n741_n140# a_n1453_n140# 0.03fF
C166 a_n29_n140# a_n919_n140# 0.02fF
C167 a_n327_n194# a_741_n194# 0.01fF
C168 a_n385_n140# a_n563_n140# 0.13fF
C169 a_n563_n140# a_1039_n140# 0.01fF
C170 a_683_n140# a_n741_n140# 0.01fF
C171 a_207_n194# a_n149_n194# 0.03fF
C172 a_n149_n194# a_n683_n194# 0.02fF
C173 a_n207_n140# a_n1453_n140# 0.02fF
C174 a_n1395_n194# a_n861_n194# 0.02fF
C175 a_29_n194# a_919_n194# 0.01fF
C176 a_149_n140# a_1217_n140# 0.02fF
C177 a_n207_n140# a_683_n140# 0.02fF
C178 a_1097_n194# a_741_n194# 0.03fF
C179 a_1275_n194# a_563_n194# 0.01fF
C180 a_n29_n140# a_505_n140# 0.04fF
C181 a_563_n194# a_385_n194# 0.10fF
C182 a_n207_n140# a_n741_n140# 0.04fF
C183 a_n1097_n140# a_n1453_n140# 0.06fF
C184 a_n327_n194# a_563_n194# 0.01fF
C185 a_n1039_n194# a_563_n194# 0.01fF
C186 a_n741_n140# a_n1097_n140# 0.06fF
C187 a_n1395_n194# a_n505_n194# 0.01fF
C188 a_n1395_n194# a_n1217_n194# 0.10fF
C189 a_327_n140# a_149_n140# 0.13fF
C190 a_n149_n194# a_919_n194# 0.01fF
C191 a_n29_n140# a_1217_n140# 0.02fF
C192 a_n207_n140# a_n1097_n140# 0.02fF
C193 a_29_n194# a_741_n194# 0.01fF
C194 a_1275_n194# a_385_n194# 0.01fF
C195 a_1097_n194# a_563_n194# 0.02fF
C196 a_505_n140# a_861_n140# 0.06fF
C197 a_505_n140# a_n919_n140# 0.01fF
C198 a_n1453_n140# a_n563_n140# 0.02fF
C199 a_207_n194# a_n1395_n194# 0.01fF
C200 a_n1395_n194# a_n683_n194# 0.01fF
C201 a_327_n140# a_n1275_n140# 0.01fF
C202 a_n327_n194# a_1275_n194# 0.01fF
C203 a_683_n140# a_n563_n140# 0.02fF
C204 a_n1039_n194# a_385_n194# 0.01fF
C205 a_327_n140# a_n29_n140# 0.06fF
C206 a_n327_n194# a_385_n194# 0.01fF
C207 a_1395_n140# VSUBS 0.02fF
C208 a_1217_n140# VSUBS 0.02fF
C209 a_1039_n140# VSUBS 0.02fF
C210 a_861_n140# VSUBS 0.02fF
C211 a_683_n140# VSUBS 0.02fF
C212 a_505_n140# VSUBS 0.02fF
C213 a_327_n140# VSUBS 0.02fF
C214 a_149_n140# VSUBS 0.02fF
C215 a_n29_n140# VSUBS 0.02fF
C216 a_n207_n140# VSUBS 0.02fF
C217 a_n385_n140# VSUBS 0.02fF
C218 a_n563_n140# VSUBS 0.02fF
C219 a_n741_n140# VSUBS 0.02fF
C220 a_n919_n140# VSUBS 0.02fF
C221 a_n1097_n140# VSUBS 0.02fF
C222 a_n1275_n140# VSUBS 0.02fF
C223 a_n1453_n140# VSUBS 0.02fF
C224 a_1275_n194# VSUBS 0.29fF
C225 a_1097_n194# VSUBS 0.23fF
C226 a_919_n194# VSUBS 0.24fF
C227 a_741_n194# VSUBS 0.25fF
C228 a_563_n194# VSUBS 0.26fF
C229 a_385_n194# VSUBS 0.27fF
C230 a_207_n194# VSUBS 0.28fF
C231 a_29_n194# VSUBS 0.28fF
C232 a_n149_n194# VSUBS 0.29fF
C233 a_n327_n194# VSUBS 0.29fF
C234 a_n505_n194# VSUBS 0.29fF
C235 a_n683_n194# VSUBS 0.29fF
C236 a_n861_n194# VSUBS 0.29fF
C237 a_n1039_n194# VSUBS 0.29fF
C238 a_n1217_n194# VSUBS 0.29fF
C239 a_n1395_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_KEEN2X a_n1008_n140# a_2374_n140# a_1306_n140# a_n652_n140#
+ a_652_n194# a_n1662_n194# a_772_n140# a_n2730_n194# a_n1720_n140# a_n60_n194# a_2076_n194#
+ a_1008_n194# a_2196_n140# a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194#
+ a_n2552_n194# a_594_n140# a_n1542_n140# a_n2610_n140# a_1720_n194# a_1840_n140#
+ a_n238_n194# a_n2908_n194# a_3086_n140# a_n296_n140# a_n1898_n140# a_n2966_n140#
+ a_296_n194# a_2018_n140# a_60_n140# a_n1306_n194# a_n2374_n194# a_n1364_n140# a_1542_n194#
+ a_416_n140# a_n2432_n140# a_2610_n194# a_n950_n194# a_1662_n140# a_2730_n140# a_2966_n194#
+ a_1898_n194# a_n2788_n140# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194#
+ a_238_n140# a_n1186_n140# a_n2254_n140# a_2432_n194# a_1364_n194# a_n772_n194# a_2552_n140#
+ a_1484_n140# a_n830_n140# a_2788_n194# a_830_n194# a_n1840_n194# a_950_n140# a_n3086_n194#
+ a_2908_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_n3144_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2374_n140# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2788_n140# a_n2908_n194# a_n2966_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n2432_n140# a_n2552_n194# a_n2610_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2966_n140# a_n3086_n194# a_n3144_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_2730_n140# a_2610_n194# a_2552_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n2610_n140# a_n2730_n194# a_n2788_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n2254_n140# a_n2374_n194# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_3086_n140# a_2966_n194# a_2908_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_2552_n140# a_2432_n194# a_2374_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_2908_n140# a_2788_n194# a_2730_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_1662_n140# a_3086_n140# 0.01fF
C1 a_n1128_n194# a_n1306_n194# 0.10fF
C2 a_2730_n140# a_2374_n140# 0.06fF
C3 a_1662_n140# a_1306_n140# 0.06fF
C4 a_2196_n140# a_1840_n140# 0.06fF
C5 a_n1484_n194# a_n2018_n194# 0.02fF
C6 a_n2018_n194# a_n2908_n194# 0.01fF
C7 a_n2254_n140# a_n1898_n140# 0.06fF
C8 a_1186_n194# a_296_n194# 0.01fF
C9 a_n3086_n194# a_n2730_n194# 0.03fF
C10 a_n118_n140# a_n830_n140# 0.03fF
C11 a_n1008_n140# a_60_n140# 0.02fF
C12 a_n296_n140# a_n1898_n140# 0.01fF
C13 a_n1662_n194# a_n60_n194# 0.01fF
C14 a_1898_n194# a_2254_n194# 0.03fF
C15 a_2076_n194# a_1364_n194# 0.01fF
C16 a_1898_n194# a_1542_n194# 0.03fF
C17 a_n1542_n140# a_n1008_n140# 0.04fF
C18 a_2018_n140# a_950_n140# 0.02fF
C19 a_1008_n194# a_n416_n194# 0.01fF
C20 a_n1662_n194# a_n1306_n194# 0.03fF
C21 a_1008_n194# a_474_n194# 0.02fF
C22 a_n296_n140# a_1128_n140# 0.01fF
C23 a_n1720_n140# a_n2254_n140# 0.04fF
C24 a_n3144_n140# a_n1898_n140# 0.02fF
C25 a_n238_n194# a_n60_n194# 0.10fF
C26 a_n1720_n140# a_n296_n140# 0.01fF
C27 a_950_n140# a_n652_n140# 0.01fF
C28 a_n60_n194# a_652_n194# 0.01fF
C29 a_1662_n140# a_1128_n140# 0.04fF
C30 a_1008_n194# a_2610_n194# 0.01fF
C31 a_n2076_n140# a_n1542_n140# 0.04fF
C32 a_950_n140# a_1306_n140# 0.06fF
C33 a_n594_n194# a_118_n194# 0.01fF
C34 a_n772_n194# a_n60_n194# 0.01fF
C35 a_n238_n194# a_n1306_n194# 0.01fF
C36 a_n1542_n140# a_n2432_n140# 0.02fF
C37 a_594_n140# a_772_n140# 0.13fF
C38 a_n1364_n140# a_n652_n140# 0.03fF
C39 a_n1720_n140# a_n3144_n140# 0.01fF
C40 a_n772_n194# a_n1306_n194# 0.02fF
C41 a_n1484_n194# a_n594_n194# 0.01fF
C42 a_1364_n194# a_n60_n194# 0.01fF
C43 a_n1484_n194# a_n1840_n194# 0.03fF
C44 a_n2196_n194# a_n2730_n194# 0.02fF
C45 a_n1840_n194# a_n2908_n194# 0.01fF
C46 a_n2374_n194# a_n3086_n194# 0.01fF
C47 a_n2196_n194# a_n950_n194# 0.01fF
C48 a_830_n194# a_1898_n194# 0.01fF
C49 a_1484_n140# a_2374_n140# 0.02fF
C50 a_60_n140# a_238_n140# 0.13fF
C51 a_2254_n194# a_1542_n194# 0.01fF
C52 a_1898_n194# a_1720_n194# 0.10fF
C53 a_416_n140# a_60_n140# 0.06fF
C54 a_n1364_n140# a_n1898_n140# 0.04fF
C55 a_2908_n140# a_2018_n140# 0.02fF
C56 a_2374_n140# a_2552_n140# 0.13fF
C57 a_950_n140# a_1128_n140# 0.13fF
C58 a_1186_n194# a_n416_n194# 0.01fF
C59 a_n474_n140# a_60_n140# 0.04fF
C60 a_1186_n194# a_474_n194# 0.01fF
C61 a_n1542_n140# a_n474_n140# 0.02fF
C62 a_n1008_n140# a_n652_n140# 0.06fF
C63 a_n2788_n140# a_n2966_n140# 0.13fF
C64 a_1840_n140# a_2374_n140# 0.04fF
C65 a_2908_n140# a_3086_n140# 0.13fF
C66 a_n296_n140# a_594_n140# 0.02fF
C67 a_1186_n194# a_2610_n194# 0.01fF
C68 a_2908_n140# a_1306_n140# 0.01fF
C69 a_n1364_n140# a_n1720_n140# 0.06fF
C70 a_1008_n194# a_n238_n194# 0.01fF
C71 a_1008_n194# a_652_n194# 0.03fF
C72 a_1662_n140# a_594_n140# 0.02fF
C73 a_n2076_n140# a_n652_n140# 0.01fF
C74 a_n118_n140# a_n1186_n140# 0.02fF
C75 a_2610_n194# a_2966_n194# 0.03fF
C76 a_n1008_n140# a_n1898_n140# 0.02fF
C77 a_n594_n194# a_296_n194# 0.01fF
C78 a_n2196_n194# a_n2374_n194# 0.10fF
C79 a_n296_n140# a_772_n140# 0.02fF
C80 a_n60_n194# a_n1306_n194# 0.01fF
C81 a_n2610_n140# a_n2966_n140# 0.06fF
C82 a_n950_n194# a_118_n194# 0.01fF
C83 a_1008_n194# a_2076_n194# 0.01fF
C84 a_830_n194# a_2254_n194# 0.01fF
C85 a_1662_n140# a_772_n140# 0.02fF
C86 a_1008_n194# a_1364_n194# 0.03fF
C87 a_830_n194# a_1542_n194# 0.01fF
C88 a_2610_n194# a_2788_n194# 0.10fF
C89 a_2254_n194# a_1720_n194# 0.02fF
C90 a_1542_n194# a_1720_n194# 0.10fF
C91 a_2018_n140# a_416_n140# 0.01fF
C92 a_n2018_n194# a_n416_n194# 0.01fF
C93 a_2018_n140# a_2730_n140# 0.03fF
C94 a_n1720_n140# a_n1008_n140# 0.03fF
C95 a_n2076_n140# a_n1898_n140# 0.13fF
C96 a_n1484_n194# a_n2730_n194# 0.01fF
C97 a_n2908_n194# a_n2730_n194# 0.10fF
C98 a_n1484_n194# a_n950_n194# 0.02fF
C99 a_n2432_n140# a_n1898_n140# 0.04fF
C100 a_950_n140# a_594_n140# 0.06fF
C101 a_n652_n140# a_238_n140# 0.02fF
C102 a_n652_n140# a_416_n140# 0.02fF
C103 a_1484_n140# a_60_n140# 0.01fF
C104 a_3086_n140# a_2730_n140# 0.06fF
C105 a_n2018_n194# a_n2552_n194# 0.02fF
C106 a_1306_n140# a_238_n140# 0.02fF
C107 a_416_n140# a_1306_n140# 0.02fF
C108 a_2730_n140# a_1306_n140# 0.01fF
C109 a_1186_n194# a_n238_n194# 0.01fF
C110 a_n474_n140# a_n652_n140# 0.13fF
C111 a_1186_n194# a_652_n194# 0.02fF
C112 a_n2018_n194# a_n1128_n194# 0.01fF
C113 a_n1720_n140# a_n2076_n140# 0.06fF
C114 a_n1720_n140# a_n2432_n140# 0.03fF
C115 a_n2196_n194# a_n3086_n194# 0.01fF
C116 a_950_n140# a_772_n140# 0.13fF
C117 a_1008_n194# a_n60_n194# 0.01fF
C118 a_n3144_n140# a_n2254_n140# 0.02fF
C119 a_n2788_n140# a_n2610_n140# 0.13fF
C120 a_n830_n140# a_n1186_n140# 0.06fF
C121 a_1186_n194# a_2076_n194# 0.01fF
C122 a_1186_n194# a_1364_n194# 0.10fF
C123 a_830_n194# a_1720_n194# 0.01fF
C124 a_n474_n140# a_n1898_n140# 0.01fF
C125 a_n594_n194# a_n416_n194# 0.10fF
C126 a_n2018_n194# a_n1662_n194# 0.03fF
C127 a_1128_n140# a_238_n140# 0.02fF
C128 a_n594_n194# a_474_n194# 0.01fF
C129 a_n1840_n194# a_n416_n194# 0.01fF
C130 a_n1484_n194# a_n2374_n194# 0.01fF
C131 a_1128_n140# a_416_n140# 0.03fF
C132 a_2730_n140# a_1128_n140# 0.01fF
C133 a_n2374_n194# a_n2908_n194# 0.02fF
C134 a_n1008_n140# a_594_n140# 0.01fF
C135 a_n950_n194# a_296_n194# 0.01fF
C136 a_2076_n194# a_2966_n194# 0.01fF
C137 a_n474_n140# a_1128_n140# 0.01fF
C138 a_1542_n194# a_118_n194# 0.01fF
C139 a_1364_n194# a_2966_n194# 0.01fF
C140 a_n118_n140# a_60_n140# 0.13fF
C141 a_n1720_n140# a_n474_n140# 0.02fF
C142 a_n118_n140# a_n1542_n140# 0.01fF
C143 a_2018_n140# a_1484_n140# 0.04fF
C144 a_n1840_n194# a_n2552_n194# 0.01fF
C145 a_n2788_n140# a_n1186_n140# 0.01fF
C146 a_n1128_n194# a_n594_n194# 0.02fF
C147 a_2018_n140# a_2552_n140# 0.04fF
C148 a_950_n140# a_n296_n140# 0.02fF
C149 a_2432_n194# a_2610_n194# 0.10fF
C150 a_2076_n194# a_2788_n194# 0.01fF
C151 a_2788_n194# a_1364_n194# 0.01fF
C152 a_n1840_n194# a_n1128_n194# 0.01fF
C153 a_n2018_n194# a_n772_n194# 0.01fF
C154 a_2196_n140# a_2374_n140# 0.13fF
C155 a_1898_n194# a_296_n194# 0.01fF
C156 a_n1364_n140# a_n2254_n140# 0.02fF
C157 a_1662_n140# a_950_n140# 0.03fF
C158 a_3086_n140# a_1484_n140# 0.01fF
C159 a_n1364_n140# a_n296_n140# 0.02fF
C160 a_2018_n140# a_1840_n140# 0.13fF
C161 a_1484_n140# a_1306_n140# 0.13fF
C162 a_1186_n194# a_n60_n194# 0.01fF
C163 a_3086_n140# a_2552_n140# 0.04fF
C164 a_1306_n140# a_2552_n140# 0.02fF
C165 a_n1484_n194# a_n3086_n194# 0.01fF
C166 a_n3086_n194# a_n2908_n194# 0.10fF
C167 a_n1662_n194# a_n594_n194# 0.01fF
C168 a_3086_n140# a_1840_n140# 0.02fF
C169 a_n1840_n194# a_n1662_n194# 0.10fF
C170 a_n2610_n140# a_n1186_n140# 0.01fF
C171 a_1306_n140# a_1840_n140# 0.04fF
C172 a_n1542_n140# a_n2966_n140# 0.01fF
C173 a_830_n194# a_118_n194# 0.01fF
C174 a_594_n140# a_238_n140# 0.06fF
C175 a_1720_n194# a_118_n194# 0.01fF
C176 a_594_n140# a_416_n140# 0.13fF
C177 a_n594_n194# a_n238_n194# 0.03fF
C178 a_n2254_n140# a_n1008_n140# 0.02fF
C179 a_n594_n194# a_652_n194# 0.01fF
C180 a_n1840_n194# a_n238_n194# 0.01fF
C181 a_1484_n140# a_1128_n140# 0.06fF
C182 a_n474_n140# a_594_n140# 0.02fF
C183 a_n1008_n140# a_n296_n140# 0.03fF
C184 a_n772_n194# a_n594_n194# 0.10fF
C185 a_n950_n194# a_n416_n194# 0.02fF
C186 a_n950_n194# a_474_n194# 0.01fF
C187 a_1128_n140# a_2552_n140# 0.01fF
C188 a_n1840_n194# a_n772_n194# 0.01fF
C189 a_n830_n140# a_60_n140# 0.02fF
C190 a_1542_n194# a_296_n194# 0.01fF
C191 a_n1542_n140# a_n830_n140# 0.03fF
C192 a_n118_n140# a_n652_n140# 0.04fF
C193 a_772_n140# a_238_n140# 0.04fF
C194 a_1662_n140# a_2908_n140# 0.02fF
C195 a_416_n140# a_772_n140# 0.06fF
C196 a_n2552_n194# a_n2730_n194# 0.10fF
C197 a_n118_n140# a_1306_n140# 0.01fF
C198 a_n2076_n140# a_n2254_n140# 0.13fF
C199 a_1128_n140# a_1840_n140# 0.03fF
C200 a_n2552_n194# a_n950_n194# 0.01fF
C201 a_n474_n140# a_772_n140# 0.02fF
C202 a_n1484_n194# a_n2196_n194# 0.01fF
C203 a_n1128_n194# a_n2730_n194# 0.01fF
C204 a_n2254_n140# a_n2432_n140# 0.13fF
C205 a_n2196_n194# a_n2908_n194# 0.01fF
C206 a_1898_n194# a_474_n194# 0.01fF
C207 a_n2018_n194# a_n1306_n194# 0.01fF
C208 a_1008_n194# a_1186_n194# 0.10fF
C209 a_n1128_n194# a_n950_n194# 0.10fF
C210 a_2610_n194# a_1898_n194# 0.01fF
C211 a_2432_n194# a_2076_n194# 0.03fF
C212 a_2432_n194# a_1364_n194# 0.01fF
C213 a_n2076_n140# a_n3144_n140# 0.02fF
C214 a_n1542_n140# a_n2788_n140# 0.02fF
C215 a_n3144_n140# a_n2432_n140# 0.03fF
C216 a_n1662_n194# a_n2730_n194# 0.01fF
C217 a_n118_n140# a_1128_n140# 0.02fF
C218 a_n1662_n194# a_n950_n194# 0.01fF
C219 a_n296_n140# a_238_n140# 0.04fF
C220 a_n118_n140# a_n1720_n140# 0.01fF
C221 a_830_n194# a_296_n194# 0.02fF
C222 a_n296_n140# a_416_n140# 0.03fF
C223 a_n1364_n140# a_n1008_n140# 0.06fF
C224 a_1720_n194# a_296_n194# 0.01fF
C225 a_1662_n140# a_238_n140# 0.01fF
C226 a_1484_n140# a_594_n140# 0.02fF
C227 a_n594_n194# a_n60_n194# 0.02fF
C228 a_n474_n140# a_n296_n140# 0.13fF
C229 a_1662_n140# a_416_n140# 0.02fF
C230 a_n2552_n194# a_n2374_n194# 0.10fF
C231 a_1662_n140# a_2730_n140# 0.02fF
C232 a_n1542_n140# a_n2610_n140# 0.02fF
C233 a_n950_n194# a_n238_n194# 0.01fF
C234 a_n2374_n194# a_n1128_n194# 0.01fF
C235 a_n950_n194# a_652_n194# 0.01fF
C236 a_n594_n194# a_n1306_n194# 0.01fF
C237 a_n1484_n194# a_118_n194# 0.01fF
C238 a_n830_n140# a_n652_n140# 0.13fF
C239 a_1542_n194# a_474_n194# 0.01fF
C240 a_n1840_n194# a_n1306_n194# 0.02fF
C241 a_n2966_n140# a_n1898_n140# 0.02fF
C242 a_n950_n194# a_n772_n194# 0.10fF
C243 a_n1364_n140# a_n2076_n140# 0.03fF
C244 a_2196_n140# a_2018_n140# 0.13fF
C245 a_594_n140# a_1840_n140# 0.02fF
C246 a_1484_n140# a_772_n140# 0.03fF
C247 a_n1364_n140# a_n2432_n140# 0.02fF
C248 a_2610_n194# a_2254_n194# 0.03fF
C249 a_2610_n194# a_1542_n194# 0.01fF
C250 a_n1484_n194# a_n2908_n194# 0.01fF
C251 a_1898_n194# a_652_n194# 0.01fF
C252 a_2196_n140# a_3086_n140# 0.02fF
C253 a_n1186_n140# a_60_n140# 0.02fF
C254 a_n1720_n140# a_n2966_n140# 0.02fF
C255 a_n1662_n194# a_n2374_n194# 0.01fF
C256 a_2196_n140# a_1306_n140# 0.02fF
C257 a_n1542_n140# a_n1186_n140# 0.06fF
C258 a_1840_n140# a_772_n140# 0.02fF
C259 a_n830_n140# a_n1898_n140# 0.02fF
C260 a_950_n140# a_238_n140# 0.03fF
C261 a_950_n140# a_416_n140# 0.04fF
C262 a_1186_n194# a_2788_n194# 0.01fF
C263 a_n2552_n194# a_n3086_n194# 0.02fF
C264 a_n474_n140# a_950_n140# 0.01fF
C265 a_n118_n140# a_594_n140# 0.03fF
C266 a_n1364_n140# a_238_n140# 0.01fF
C267 a_1898_n194# a_2076_n194# 0.10fF
C268 a_1898_n194# a_1364_n194# 0.02fF
C269 a_n2076_n140# a_n1008_n140# 0.02fF
C270 a_n1720_n140# a_n830_n140# 0.02fF
C271 a_n1008_n140# a_n2432_n140# 0.01fF
C272 a_n1364_n140# a_n474_n140# 0.02fF
C273 a_830_n194# a_n416_n194# 0.01fF
C274 a_1008_n194# a_n594_n194# 0.01fF
C275 a_2788_n194# a_2966_n194# 0.10fF
C276 a_n2374_n194# a_n772_n194# 0.01fF
C277 a_118_n194# a_296_n194# 0.10fF
C278 a_830_n194# a_474_n194# 0.03fF
C279 a_1720_n194# a_474_n194# 0.01fF
C280 a_n2788_n140# a_n1898_n140# 0.02fF
C281 a_n118_n140# a_772_n140# 0.02fF
C282 a_1662_n140# a_1484_n140# 0.13fF
C283 a_2196_n140# a_1128_n140# 0.02fF
C284 a_1008_n194# a_2432_n194# 0.01fF
C285 a_2610_n194# a_1720_n194# 0.01fF
C286 a_1662_n140# a_2552_n140# 0.02fF
C287 a_n950_n194# a_n60_n194# 0.01fF
C288 a_n1662_n194# a_n3086_n194# 0.01fF
C289 a_2254_n194# a_652_n194# 0.01fF
C290 a_n2076_n140# a_n2432_n140# 0.06fF
C291 a_1542_n194# a_652_n194# 0.01fF
C292 a_n1306_n194# a_n2730_n194# 0.01fF
C293 a_n1720_n140# a_n2788_n140# 0.02fF
C294 a_n1008_n140# a_238_n140# 0.02fF
C295 a_n950_n194# a_n1306_n194# 0.03fF
C296 a_n1008_n140# a_416_n140# 0.01fF
C297 a_1662_n140# a_1840_n140# 0.13fF
C298 a_2908_n140# a_2730_n140# 0.13fF
C299 a_n2196_n194# a_n2552_n194# 0.03fF
C300 a_n474_n140# a_n1008_n140# 0.04fF
C301 a_n2610_n140# a_n1898_n140# 0.03fF
C302 a_n2196_n194# a_n1128_n194# 0.01fF
C303 a_2018_n140# a_2374_n140# 0.06fF
C304 a_n1186_n140# a_n652_n140# 0.04fF
C305 a_2076_n194# a_2254_n194# 0.10fF
C306 a_2254_n194# a_1364_n194# 0.01fF
C307 a_2076_n194# a_1542_n194# 0.02fF
C308 a_1364_n194# a_1542_n194# 0.10fF
C309 a_950_n140# a_1484_n140# 0.04fF
C310 a_n118_n140# a_n296_n140# 0.13fF
C311 a_n830_n140# a_594_n140# 0.01fF
C312 a_950_n140# a_2552_n140# 0.01fF
C313 a_n1720_n140# a_n2610_n140# 0.02fF
C314 a_n2076_n140# a_n474_n140# 0.01fF
C315 a_3086_n140# a_2374_n140# 0.03fF
C316 a_1306_n140# a_2374_n140# 0.02fF
C317 a_n1542_n140# a_60_n140# 0.01fF
C318 a_1186_n194# a_2432_n194# 0.01fF
C319 a_950_n140# a_1840_n140# 0.02fF
C320 a_n2196_n194# a_n1662_n194# 0.02fF
C321 a_n1186_n140# a_n1898_n140# 0.03fF
C322 a_830_n194# a_n238_n194# 0.01fF
C323 a_n416_n194# a_118_n194# 0.02fF
C324 a_118_n194# a_474_n194# 0.03fF
C325 a_830_n194# a_652_n194# 0.10fF
C326 a_n2374_n194# a_n1306_n194# 0.01fF
C327 a_2196_n140# a_594_n140# 0.01fF
C328 a_1720_n194# a_652_n194# 0.01fF
C329 a_n830_n140# a_772_n140# 0.01fF
C330 a_830_n194# a_n772_n194# 0.01fF
C331 a_2432_n194# a_2966_n194# 0.02fF
C332 a_416_n140# a_238_n140# 0.13fF
C333 a_n1484_n194# a_n416_n194# 0.01fF
C334 a_1542_n194# a_n60_n194# 0.01fF
C335 a_n1720_n140# a_n1186_n140# 0.04fF
C336 a_n474_n140# a_238_n140# 0.03fF
C337 a_n2254_n140# a_n2966_n140# 0.03fF
C338 a_n474_n140# a_416_n140# 0.02fF
C339 a_n1128_n194# a_118_n194# 0.01fF
C340 a_n2196_n194# a_n772_n194# 0.01fF
C341 a_830_n194# a_2076_n194# 0.01fF
C342 a_2196_n140# a_772_n140# 0.01fF
C343 a_1008_n194# a_1898_n194# 0.01fF
C344 a_830_n194# a_1364_n194# 0.02fF
C345 a_1128_n140# a_2374_n140# 0.02fF
C346 a_2432_n194# a_2788_n194# 0.03fF
C347 a_2076_n194# a_1720_n194# 0.03fF
C348 a_1364_n194# a_1720_n194# 0.03fF
C349 a_n118_n140# a_950_n140# 0.02fF
C350 a_n2018_n194# a_n594_n194# 0.01fF
C351 a_2908_n140# a_1484_n140# 0.01fF
C352 a_n1484_n194# a_n2552_n194# 0.01fF
C353 a_n2552_n194# a_n2908_n194# 0.03fF
C354 a_n2018_n194# a_n1840_n194# 0.10fF
C355 a_2908_n140# a_2552_n140# 0.06fF
C356 a_n1484_n194# a_n1128_n194# 0.03fF
C357 a_n118_n140# a_n1364_n140# 0.02fF
C358 a_n3144_n140# a_n2966_n140# 0.13fF
C359 a_n2254_n140# a_n830_n140# 0.01fF
C360 a_n830_n140# a_n296_n140# 0.04fF
C361 a_2908_n140# a_1840_n140# 0.02fF
C362 a_n652_n140# a_60_n140# 0.03fF
C363 a_n1542_n140# a_n652_n140# 0.02fF
C364 a_1306_n140# a_60_n140# 0.02fF
C365 a_n1484_n194# a_n1662_n194# 0.10fF
C366 a_n1662_n194# a_n2908_n194# 0.01fF
C367 a_830_n194# a_n60_n194# 0.01fF
C368 a_n238_n194# a_118_n194# 0.03fF
C369 a_n416_n194# a_296_n194# 0.01fF
C370 a_118_n194# a_652_n194# 0.02fF
C371 a_296_n194# a_474_n194# 0.10fF
C372 a_n2788_n140# a_n2254_n140# 0.04fF
C373 a_n772_n194# a_118_n194# 0.01fF
C374 a_2196_n140# a_1662_n140# 0.04fF
C375 a_1186_n194# a_1898_n194# 0.01fF
C376 a_1008_n194# a_2254_n194# 0.01fF
C377 a_1008_n194# a_1542_n194# 0.02fF
C378 a_n118_n140# a_n1008_n140# 0.02fF
C379 a_1484_n140# a_238_n140# 0.02fF
C380 a_n1364_n140# a_n2966_n140# 0.01fF
C381 a_n1484_n194# a_n238_n194# 0.01fF
C382 a_n1840_n194# a_n594_n194# 0.01fF
C383 a_1484_n140# a_416_n140# 0.02fF
C384 a_2730_n140# a_1484_n140# 0.02fF
C385 a_n1542_n140# a_n1898_n140# 0.06fF
C386 a_2730_n140# a_2552_n140# 0.13fF
C387 a_n1128_n194# a_296_n194# 0.01fF
C388 a_n1484_n194# a_n772_n194# 0.01fF
C389 a_n3144_n140# a_n2788_n140# 0.06fF
C390 a_1898_n194# a_2966_n194# 0.01fF
C391 a_1364_n194# a_118_n194# 0.01fF
C392 a_n2196_n194# a_n1306_n194# 0.01fF
C393 a_1128_n140# a_60_n140# 0.02fF
C394 a_1840_n140# a_238_n140# 0.01fF
C395 a_416_n140# a_1840_n140# 0.01fF
C396 a_2730_n140# a_1840_n140# 0.02fF
C397 a_n2018_n194# a_n2730_n194# 0.01fF
C398 a_n2254_n140# a_n2610_n140# 0.06fF
C399 a_n1364_n140# a_n830_n140# 0.04fF
C400 a_1898_n194# a_2788_n194# 0.01fF
C401 a_n1720_n140# a_n1542_n140# 0.13fF
C402 a_n2018_n194# a_n950_n194# 0.01fF
C403 a_772_n140# a_2374_n140# 0.01fF
C404 a_2196_n140# a_950_n140# 0.02fF
C405 a_3086_n140# a_2018_n140# 0.02fF
C406 a_2018_n140# a_1306_n140# 0.03fF
C407 a_n3144_n140# a_n2610_n140# 0.04fF
C408 a_830_n194# a_1008_n194# 0.10fF
C409 a_1186_n194# a_2254_n194# 0.01fF
C410 a_1186_n194# a_1542_n194# 0.03fF
C411 a_1008_n194# a_1720_n194# 0.01fF
C412 a_n118_n140# a_238_n140# 0.06fF
C413 a_n118_n140# a_416_n140# 0.04fF
C414 a_n1364_n140# a_n2788_n140# 0.01fF
C415 a_n2254_n140# a_n1186_n140# 0.02fF
C416 a_n60_n194# a_118_n194# 0.10fF
C417 a_n416_n194# a_474_n194# 0.01fF
C418 a_n238_n194# a_296_n194# 0.02fF
C419 a_296_n194# a_652_n194# 0.03fF
C420 a_n1186_n140# a_n296_n140# 0.02fF
C421 a_n2076_n140# a_n2966_n140# 0.02fF
C422 a_n118_n140# a_n474_n140# 0.06fF
C423 a_n830_n140# a_n1008_n140# 0.13fF
C424 a_n772_n194# a_296_n194# 0.01fF
C425 a_2254_n194# a_2966_n194# 0.01fF
C426 a_1542_n194# a_2966_n194# 0.01fF
C427 a_n2966_n140# a_n2432_n140# 0.04fF
C428 a_n1306_n194# a_118_n194# 0.01fF
C429 a_n1484_n194# a_n60_n194# 0.01fF
C430 a_2018_n140# a_1128_n140# 0.02fF
C431 a_n652_n140# a_n1898_n140# 0.02fF
C432 a_n2018_n194# a_n2374_n194# 0.03fF
C433 a_n1840_n194# a_n2730_n194# 0.01fF
C434 a_n950_n194# a_n594_n194# 0.03fF
C435 a_n1128_n194# a_n416_n194# 0.01fF
C436 a_n1128_n194# a_474_n194# 0.01fF
C437 a_1484_n140# a_2552_n140# 0.02fF
C438 a_2788_n194# a_1542_n194# 0.01fF
C439 a_2254_n194# a_2788_n194# 0.02fF
C440 a_594_n140# a_60_n140# 0.04fF
C441 a_n1840_n194# a_n950_n194# 0.01fF
C442 a_1662_n140# a_2374_n140# 0.03fF
C443 a_1364_n194# a_296_n194# 0.01fF
C444 a_n1484_n194# a_n1306_n194# 0.10fF
C445 a_n1306_n194# a_n2908_n194# 0.01fF
C446 a_n2076_n140# a_n830_n140# 0.02fF
C447 a_2196_n140# a_2908_n140# 0.03fF
C448 a_n1364_n140# a_n2610_n140# 0.02fF
C449 a_n830_n140# a_n2432_n140# 0.01fF
C450 a_1484_n140# a_1840_n140# 0.06fF
C451 a_1128_n140# a_1306_n140# 0.13fF
C452 a_n1720_n140# a_n652_n140# 0.02fF
C453 a_n2552_n194# a_n1128_n194# 0.01fF
C454 a_1840_n140# a_2552_n140# 0.03fF
C455 a_830_n194# a_1186_n194# 0.03fF
C456 a_772_n140# a_60_n140# 0.03fF
C457 a_1186_n194# a_1720_n194# 0.02fF
C458 a_n1662_n194# a_n416_n194# 0.01fF
C459 a_2432_n194# a_1898_n194# 0.02fF
C460 a_n2076_n140# a_n2788_n140# 0.03fF
C461 a_1008_n194# a_118_n194# 0.01fF
C462 a_n2018_n194# a_n3086_n194# 0.01fF
C463 a_n830_n140# a_238_n140# 0.02fF
C464 a_n1364_n140# a_n1186_n140# 0.13fF
C465 a_1720_n194# a_2966_n194# 0.01fF
C466 a_n1720_n140# a_n1898_n140# 0.13fF
C467 a_n2788_n140# a_n2432_n140# 0.06fF
C468 a_n830_n140# a_416_n140# 0.02fF
C469 a_950_n140# a_2374_n140# 0.01fF
C470 a_n1662_n194# a_n2552_n194# 0.01fF
C471 a_n416_n194# a_n238_n194# 0.10fF
C472 a_n2610_n140# a_n1008_n140# 0.01fF
C473 a_n118_n140# a_1484_n140# 0.01fF
C474 a_n416_n194# a_652_n194# 0.01fF
C475 a_n60_n194# a_296_n194# 0.03fF
C476 a_n238_n194# a_474_n194# 0.01fF
C477 a_n1840_n194# a_n2374_n194# 0.02fF
C478 a_474_n194# a_652_n194# 0.10fF
C479 a_n474_n140# a_n830_n140# 0.06fF
C480 a_n1662_n194# a_n1128_n194# 0.02fF
C481 a_n772_n194# a_n416_n194# 0.03fF
C482 a_n772_n194# a_474_n194# 0.01fF
C483 a_2788_n194# a_1720_n194# 0.01fF
C484 a_n1306_n194# a_296_n194# 0.01fF
C485 a_2018_n140# a_594_n140# 0.01fF
C486 a_2196_n140# a_2730_n140# 0.04fF
C487 a_n2076_n140# a_n2610_n140# 0.04fF
C488 a_n1542_n140# a_n2254_n140# 0.03fF
C489 a_n296_n140# a_60_n140# 0.06fF
C490 a_n1128_n194# a_n238_n194# 0.01fF
C491 a_n1542_n140# a_n296_n140# 0.02fF
C492 a_n652_n140# a_594_n140# 0.02fF
C493 a_2076_n194# a_474_n194# 0.01fF
C494 a_1364_n194# a_474_n194# 0.01fF
C495 a_n2610_n140# a_n2432_n140# 0.13fF
C496 a_1662_n140# a_60_n140# 0.01fF
C497 a_n1128_n194# a_n772_n194# 0.03fF
C498 a_n1186_n140# a_n1008_n140# 0.13fF
C499 a_594_n140# a_1306_n140# 0.03fF
C500 a_2018_n140# a_772_n140# 0.02fF
C501 a_2432_n194# a_2254_n194# 0.10fF
C502 a_2610_n194# a_2076_n194# 0.02fF
C503 a_2432_n194# a_1542_n194# 0.01fF
C504 a_2610_n194# a_1364_n194# 0.01fF
C505 a_n3144_n140# a_n1542_n140# 0.01fF
C506 a_n2196_n194# a_n2018_n194# 0.10fF
C507 a_1186_n194# a_118_n194# 0.01fF
C508 a_n1840_n194# a_n3086_n194# 0.01fF
C509 a_n652_n140# a_772_n140# 0.01fF
C510 a_2908_n140# a_2374_n140# 0.04fF
C511 a_n1662_n194# a_n238_n194# 0.01fF
C512 a_n2076_n140# a_n1186_n140# 0.02fF
C513 a_1306_n140# a_772_n140# 0.04fF
C514 a_n1662_n194# a_n772_n194# 0.01fF
C515 a_n1186_n140# a_n2432_n140# 0.02fF
C516 a_1008_n194# a_296_n194# 0.01fF
C517 a_1128_n140# a_594_n140# 0.04fF
C518 a_n416_n194# a_n60_n194# 0.03fF
C519 a_950_n140# a_60_n140# 0.02fF
C520 a_n238_n194# a_652_n194# 0.01fF
C521 a_n60_n194# a_474_n194# 0.02fF
C522 a_n2374_n194# a_n2730_n194# 0.03fF
C523 a_n772_n194# a_n238_n194# 0.02fF
C524 a_830_n194# a_n594_n194# 0.01fF
C525 a_n2374_n194# a_n950_n194# 0.01fF
C526 a_n772_n194# a_652_n194# 0.01fF
C527 a_n416_n194# a_n1306_n194# 0.01fF
C528 a_n1364_n140# a_60_n140# 0.01fF
C529 a_n1364_n140# a_n1542_n140# 0.13fF
C530 a_1662_n140# a_2018_n140# 0.06fF
C531 a_n1186_n140# a_238_n140# 0.01fF
C532 a_2196_n140# a_1484_n140# 0.03fF
C533 a_1128_n140# a_772_n140# 0.06fF
C534 a_n2254_n140# a_n652_n140# 0.01fF
C535 a_n1186_n140# a_416_n140# 0.01fF
C536 a_830_n194# a_2432_n194# 0.01fF
C537 a_2196_n140# a_2552_n140# 0.06fF
C538 a_2432_n194# a_1720_n194# 0.01fF
C539 a_n296_n140# a_n652_n140# 0.06fF
C540 a_n1128_n194# a_n60_n194# 0.01fF
C541 a_n2196_n194# a_n594_n194# 0.01fF
C542 a_1364_n194# a_n238_n194# 0.01fF
C543 a_n2552_n194# a_n1306_n194# 0.01fF
C544 a_2076_n194# a_652_n194# 0.01fF
C545 a_n2196_n194# a_n1840_n194# 0.03fF
C546 a_n474_n140# a_n1186_n140# 0.03fF
C547 a_1364_n194# a_652_n194# 0.01fF
C548 a_n296_n140# a_1306_n140# 0.01fF
C549 a_3086_n140# VSUBS 0.02fF
C550 a_2908_n140# VSUBS 0.02fF
C551 a_2730_n140# VSUBS 0.02fF
C552 a_2552_n140# VSUBS 0.02fF
C553 a_2374_n140# VSUBS 0.02fF
C554 a_2196_n140# VSUBS 0.02fF
C555 a_2018_n140# VSUBS 0.02fF
C556 a_1840_n140# VSUBS 0.02fF
C557 a_1662_n140# VSUBS 0.02fF
C558 a_1484_n140# VSUBS 0.02fF
C559 a_1306_n140# VSUBS 0.02fF
C560 a_1128_n140# VSUBS 0.02fF
C561 a_950_n140# VSUBS 0.02fF
C562 a_772_n140# VSUBS 0.02fF
C563 a_594_n140# VSUBS 0.02fF
C564 a_416_n140# VSUBS 0.02fF
C565 a_238_n140# VSUBS 0.02fF
C566 a_60_n140# VSUBS 0.02fF
C567 a_n118_n140# VSUBS 0.02fF
C568 a_n296_n140# VSUBS 0.02fF
C569 a_n474_n140# VSUBS 0.02fF
C570 a_n652_n140# VSUBS 0.02fF
C571 a_n830_n140# VSUBS 0.02fF
C572 a_n1008_n140# VSUBS 0.02fF
C573 a_n1186_n140# VSUBS 0.02fF
C574 a_n1364_n140# VSUBS 0.02fF
C575 a_n1542_n140# VSUBS 0.02fF
C576 a_n1720_n140# VSUBS 0.02fF
C577 a_n1898_n140# VSUBS 0.02fF
C578 a_n2076_n140# VSUBS 0.02fF
C579 a_n2254_n140# VSUBS 0.02fF
C580 a_n2432_n140# VSUBS 0.02fF
C581 a_n2610_n140# VSUBS 0.02fF
C582 a_n2788_n140# VSUBS 0.02fF
C583 a_n2966_n140# VSUBS 0.02fF
C584 a_n3144_n140# VSUBS 0.02fF
C585 a_2966_n194# VSUBS 0.29fF
C586 a_2788_n194# VSUBS 0.23fF
C587 a_2610_n194# VSUBS 0.24fF
C588 a_2432_n194# VSUBS 0.25fF
C589 a_2254_n194# VSUBS 0.26fF
C590 a_2076_n194# VSUBS 0.27fF
C591 a_1898_n194# VSUBS 0.28fF
C592 a_1720_n194# VSUBS 0.28fF
C593 a_1542_n194# VSUBS 0.29fF
C594 a_1364_n194# VSUBS 0.29fF
C595 a_1186_n194# VSUBS 0.29fF
C596 a_1008_n194# VSUBS 0.29fF
C597 a_830_n194# VSUBS 0.29fF
C598 a_652_n194# VSUBS 0.29fF
C599 a_474_n194# VSUBS 0.29fF
C600 a_296_n194# VSUBS 0.29fF
C601 a_118_n194# VSUBS 0.29fF
C602 a_n60_n194# VSUBS 0.29fF
C603 a_n238_n194# VSUBS 0.29fF
C604 a_n416_n194# VSUBS 0.29fF
C605 a_n594_n194# VSUBS 0.29fF
C606 a_n772_n194# VSUBS 0.29fF
C607 a_n950_n194# VSUBS 0.29fF
C608 a_n1128_n194# VSUBS 0.29fF
C609 a_n1306_n194# VSUBS 0.29fF
C610 a_n1484_n194# VSUBS 0.29fF
C611 a_n1662_n194# VSUBS 0.29fF
C612 a_n1840_n194# VSUBS 0.29fF
C613 a_n2018_n194# VSUBS 0.29fF
C614 a_n2196_n194# VSUBS 0.29fF
C615 a_n2374_n194# VSUBS 0.29fF
C616 a_n2552_n194# VSUBS 0.29fF
C617 a_n2730_n194# VSUBS 0.29fF
C618 a_n2908_n194# VSUBS 0.29fF
C619 a_n3086_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_VJ4JGY a_n352_n194# a_n60_n194# a_n644_n194# a_n936_n194#
+ a_n410_n140# a_n994_n140# a_n702_n140# a_n232_n140# a_n524_n140# a_524_n194# a_232_n194#
+ a_n816_n140# a_816_n194# a_644_n140# a_352_n140# a_936_n140# a_60_n140# a_174_n140#
+ a_466_n140# a_758_n140# a_n118_n140# VSUBS
X0 a_n232_n140# a_n352_n194# a_n410_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n524_n140# a_n644_n194# a_n702_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n816_n140# a_n936_n194# a_n994_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_352_n140# a_232_n194# a_174_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_644_n140# a_524_n194# a_466_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_936_n140# a_816_n194# a_758_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n936_n194# a_n644_n194# 0.04fF
C1 a_232_n194# a_816_n194# 0.02fF
C2 a_758_n140# a_466_n140# 0.07fF
C3 a_n816_n140# a_466_n140# 0.01fF
C4 a_174_n140# a_n232_n140# 0.05fF
C5 a_n816_n140# a_n994_n140# 0.13fF
C6 a_352_n140# a_758_n140# 0.05fF
C7 a_352_n140# a_n816_n140# 0.02fF
C8 a_644_n140# a_174_n140# 0.04fF
C9 a_174_n140# a_936_n140# 0.03fF
C10 a_60_n140# a_n524_n140# 0.03fF
C11 a_524_n194# a_n644_n194# 0.01fF
C12 a_60_n140# a_466_n140# 0.05fF
C13 a_174_n140# a_n702_n140# 0.02fF
C14 a_n232_n140# a_n524_n140# 0.07fF
C15 a_60_n140# a_n994_n140# 0.02fF
C16 a_60_n140# a_352_n140# 0.07fF
C17 a_644_n140# a_n524_n140# 0.02fF
C18 a_n232_n140# a_466_n140# 0.03fF
C19 a_n524_n140# a_936_n140# 0.01fF
C20 a_n232_n140# a_n994_n140# 0.03fF
C21 a_n60_n194# a_n936_n194# 0.01fF
C22 a_352_n140# a_n232_n140# 0.03fF
C23 a_644_n140# a_466_n140# 0.13fF
C24 a_936_n140# a_466_n140# 0.04fF
C25 a_644_n140# a_n994_n140# 0.01fF
C26 a_n702_n140# a_n524_n140# 0.13fF
C27 a_352_n140# a_644_n140# 0.07fF
C28 a_758_n140# a_n816_n140# 0.01fF
C29 a_352_n140# a_936_n140# 0.03fF
C30 a_n410_n140# a_n118_n140# 0.07fF
C31 a_n702_n140# a_466_n140# 0.02fF
C32 a_n702_n140# a_n994_n140# 0.07fF
C33 a_352_n140# a_n702_n140# 0.02fF
C34 a_n60_n194# a_524_n194# 0.02fF
C35 a_n352_n194# a_n644_n194# 0.04fF
C36 a_60_n140# a_758_n140# 0.03fF
C37 a_60_n140# a_n816_n140# 0.02fF
C38 a_524_n194# a_816_n194# 0.04fF
C39 a_758_n140# a_n232_n140# 0.02fF
C40 a_n232_n140# a_n816_n140# 0.03fF
C41 a_174_n140# a_n410_n140# 0.03fF
C42 a_644_n140# a_758_n140# 0.25fF
C43 a_644_n140# a_n816_n140# 0.01fF
C44 a_758_n140# a_936_n140# 0.13fF
C45 a_60_n140# a_n232_n140# 0.07fF
C46 a_758_n140# a_n702_n140# 0.01fF
C47 a_n702_n140# a_n816_n140# 0.25fF
C48 a_232_n194# a_n936_n194# 0.01fF
C49 a_n410_n140# a_n524_n140# 0.25fF
C50 a_60_n140# a_644_n140# 0.03fF
C51 a_n352_n194# a_n60_n194# 0.04fF
C52 a_60_n140# a_936_n140# 0.02fF
C53 a_n352_n194# a_816_n194# 0.01fF
C54 a_174_n140# a_n118_n140# 0.07fF
C55 a_n410_n140# a_466_n140# 0.02fF
C56 a_n410_n140# a_n994_n140# 0.03fF
C57 a_644_n140# a_n232_n140# 0.02fF
C58 a_352_n140# a_n410_n140# 0.03fF
C59 a_n232_n140# a_936_n140# 0.02fF
C60 a_60_n140# a_n702_n140# 0.03fF
C61 a_232_n194# a_524_n194# 0.04fF
C62 a_644_n140# a_936_n140# 0.07fF
C63 a_n702_n140# a_n232_n140# 0.04fF
C64 a_n118_n140# a_n524_n140# 0.05fF
C65 a_n60_n194# a_n644_n194# 0.02fF
C66 a_644_n140# a_n702_n140# 0.01fF
C67 a_816_n194# a_n644_n194# 0.01fF
C68 a_n702_n140# a_936_n140# 0.01fF
C69 a_n118_n140# a_466_n140# 0.03fF
C70 a_n118_n140# a_n994_n140# 0.02fF
C71 a_352_n140# a_n118_n140# 0.04fF
C72 a_758_n140# a_n410_n140# 0.02fF
C73 a_n410_n140# a_n816_n140# 0.05fF
C74 a_174_n140# a_n524_n140# 0.03fF
C75 a_n352_n194# a_232_n194# 0.02fF
C76 a_n936_n194# a_524_n194# 0.01fF
C77 a_174_n140# a_466_n140# 0.07fF
C78 a_174_n140# a_n994_n140# 0.02fF
C79 a_60_n140# a_n410_n140# 0.04fF
C80 a_352_n140# a_174_n140# 0.13fF
C81 a_n60_n194# a_816_n194# 0.01fF
C82 a_758_n140# a_n118_n140# 0.02fF
C83 a_n118_n140# a_n816_n140# 0.03fF
C84 a_n410_n140# a_n232_n140# 0.13fF
C85 a_n524_n140# a_466_n140# 0.02fF
C86 a_232_n194# a_n644_n194# 0.01fF
C87 a_644_n140# a_n410_n140# 0.02fF
C88 a_n524_n140# a_n994_n140# 0.04fF
C89 a_n410_n140# a_936_n140# 0.01fF
C90 a_352_n140# a_n524_n140# 0.02fF
C91 a_n994_n140# a_466_n140# 0.01fF
C92 a_60_n140# a_n118_n140# 0.13fF
C93 a_352_n140# a_466_n140# 0.25fF
C94 a_n702_n140# a_n410_n140# 0.07fF
C95 a_352_n140# a_n994_n140# 0.01fF
C96 a_n352_n194# a_n936_n194# 0.02fF
C97 a_174_n140# a_758_n140# 0.03fF
C98 a_174_n140# a_n816_n140# 0.02fF
C99 a_n118_n140# a_n232_n140# 0.25fF
C100 a_644_n140# a_n118_n140# 0.03fF
C101 a_n118_n140# a_936_n140# 0.02fF
C102 a_60_n140# a_174_n140# 0.25fF
C103 a_232_n194# a_n60_n194# 0.04fF
C104 a_n352_n194# a_524_n194# 0.01fF
C105 a_758_n140# a_n524_n140# 0.01fF
C106 a_n816_n140# a_n524_n140# 0.07fF
C107 a_n702_n140# a_n118_n140# 0.03fF
C108 a_936_n140# VSUBS 0.02fF
C109 a_758_n140# VSUBS 0.02fF
C110 a_644_n140# VSUBS 0.02fF
C111 a_466_n140# VSUBS 0.02fF
C112 a_352_n140# VSUBS 0.02fF
C113 a_174_n140# VSUBS 0.02fF
C114 a_60_n140# VSUBS 0.02fF
C115 a_n118_n140# VSUBS 0.02fF
C116 a_n232_n140# VSUBS 0.02fF
C117 a_n410_n140# VSUBS 0.02fF
C118 a_n524_n140# VSUBS 0.02fF
C119 a_n702_n140# VSUBS 0.02fF
C120 a_n816_n140# VSUBS 0.02fF
C121 a_n994_n140# VSUBS 0.02fF
C122 a_816_n194# VSUBS 0.29fF
C123 a_524_n194# VSUBS 0.24fF
C124 a_232_n194# VSUBS 0.26fF
C125 a_n60_n194# VSUBS 0.27fF
C126 a_n352_n194# VSUBS 0.29fF
C127 a_n644_n194# VSUBS 0.29fF
C128 a_n936_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_E4DCBA a_n1008_n140# a_n416_n205# a_1306_n140# a_n652_n140#
+ a_474_n205# a_n1484_n205# a_772_n140# a_n1720_n140# a_1720_n205# a_n238_n205# a_n474_n140#
+ a_296_n205# a_1128_n140# a_594_n140# a_1542_n205# a_n1306_n205# a_n1542_n140# a_n950_n205#
+ w_n2112_n241# a_1840_n140# a_1898_n205# a_n296_n140# a_n1898_n140# a_2018_n140#
+ a_60_n140# a_118_n205# a_n1128_n205# a_n1364_n140# a_1364_n205# a_416_n140# a_n772_n205#
+ a_1662_n140# a_830_n205# a_n1840_n205# a_n118_n140# a_1186_n205# a_n2018_n205# a_238_n140#
+ a_n1186_n140# a_n594_n205# a_1484_n140# a_n830_n140# a_652_n205# a_n1662_n205# a_950_n140#
+ a_n60_n205# a_n2076_n140# a_1008_n205# VSUBS
X0 a_1662_n140# a_1542_n205# a_1484_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n205# a_n296_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n205# a_n830_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_2018_n140# a_1898_n205# a_1840_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1008_n140# a_n1128_n205# a_n1186_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_594_n140# a_474_n205# a_416_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_60_n140# a_n60_n205# a_n118_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1484_n140# a_1364_n205# a_1306_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1542_n140# a_n1662_n205# a_n1720_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_950_n140# a_830_n205# a_772_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n830_n140# a_n950_n205# a_n1008_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n474_n140# a_n594_n205# a_n652_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_1840_n140# a_1720_n205# a_1662_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_416_n140# a_296_n205# a_238_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1898_n140# a_n2018_n205# a_n2076_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n296_n140# a_n416_n205# a_n474_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n1720_n140# a_n1840_n205# a_n1898_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1306_n140# a_1186_n205# a_1128_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1364_n140# a_n1484_n205# a_n1542_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_238_n140# a_118_n205# a_60_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_1128_n140# a_1008_n205# a_950_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_n1186_n140# a_n1306_n205# a_n1364_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_772_n140# a_652_n205# a_594_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_772_n140# a_60_n140# 0.03fF
C1 a_n594_n205# a_n2018_n205# 0.01fF
C2 a_n1720_n140# a_n1542_n140# 0.13fF
C3 a_950_n140# a_n296_n140# 0.02fF
C4 a_n1364_n140# a_n830_n140# 0.04fF
C5 a_n830_n140# a_60_n140# 0.02fF
C6 a_950_n140# a_1306_n140# 0.06fF
C7 a_118_n205# a_1008_n205# 0.01fF
C8 a_238_n140# a_n118_n140# 0.06fF
C9 a_n594_n205# a_n950_n205# 0.03fF
C10 a_n594_n205# a_n238_n205# 0.03fF
C11 a_n772_n205# a_n60_n205# 0.01fF
C12 a_n1306_n205# a_n1840_n205# 0.02fF
C13 a_1840_n140# a_416_n140# 0.01fF
C14 a_296_n205# a_1720_n205# 0.01fF
C15 a_n1186_n140# a_n1542_n140# 0.06fF
C16 a_296_n205# a_830_n205# 0.02fF
C17 w_n2112_n241# a_n118_n140# 0.02fF
C18 a_1484_n140# a_950_n140# 0.04fF
C19 w_n2112_n241# a_n1898_n140# 0.02fF
C20 a_1542_n205# a_1364_n205# 0.11fF
C21 a_1364_n205# a_652_n205# 0.01fF
C22 a_1128_n140# a_1662_n140# 0.04fF
C23 a_296_n205# a_n1306_n205# 0.01fF
C24 a_1898_n205# a_1186_n205# 0.01fF
C25 a_1662_n140# a_772_n140# 0.02fF
C26 w_n2112_n241# a_n594_n205# 0.24fF
C27 a_n950_n205# a_n2018_n205# 0.01fF
C28 a_n2076_n140# a_n1542_n140# 0.04fF
C29 a_594_n140# a_n118_n140# 0.03fF
C30 a_n60_n205# a_1364_n205# 0.01fF
C31 a_n1364_n140# a_n1008_n140# 0.06fF
C32 a_n652_n140# a_n118_n140# 0.04fF
C33 a_n1008_n140# a_60_n140# 0.02fF
C34 a_n474_n140# a_238_n140# 0.03fF
C35 a_n652_n140# a_n1898_n140# 0.02fF
C36 a_474_n205# a_n594_n205# 0.01fF
C37 a_n594_n205# a_n416_n205# 0.11fF
C38 a_n950_n205# a_n238_n205# 0.01fF
C39 a_1840_n140# a_1306_n140# 0.04fF
C40 w_n2112_n241# a_n474_n140# 0.02fF
C41 a_118_n205# a_1720_n205# 0.01fF
C42 a_118_n205# a_830_n205# 0.01fF
C43 a_1128_n140# a_416_n140# 0.03fF
C44 w_n2112_n241# a_n2018_n205# 0.31fF
C45 a_416_n140# a_772_n140# 0.06fF
C46 a_118_n205# a_n1306_n205# 0.01fF
C47 a_1840_n140# a_1484_n140# 0.06fF
C48 a_296_n205# a_1542_n205# 0.01fF
C49 a_296_n205# a_652_n205# 0.03fF
C50 a_n830_n140# a_416_n140# 0.02fF
C51 a_n1840_n205# a_n772_n205# 0.01fF
C52 a_n474_n140# a_594_n140# 0.02fF
C53 w_n2112_n241# a_n950_n205# 0.24fF
C54 w_n2112_n241# a_n238_n205# 0.24fF
C55 a_n416_n205# a_n2018_n205# 0.01fF
C56 a_n1306_n205# a_n1662_n205# 0.03fF
C57 a_1898_n205# a_1008_n205# 0.01fF
C58 a_n652_n140# a_n474_n140# 0.13fF
C59 a_474_n205# a_n950_n205# 0.01fF
C60 a_296_n205# a_n772_n205# 0.01fF
C61 a_296_n205# a_n60_n205# 0.03fF
C62 a_474_n205# a_n238_n205# 0.01fF
C63 a_n1306_n205# a_n1484_n205# 0.11fF
C64 a_n950_n205# a_n416_n205# 0.02fF
C65 a_n238_n205# a_n416_n205# 0.11fF
C66 w_n2112_n241# a_238_n140# 0.02fF
C67 a_1128_n140# a_n296_n140# 0.01fF
C68 a_1128_n140# a_1306_n140# 0.13fF
C69 a_n296_n140# a_772_n140# 0.02fF
C70 a_n1364_n140# a_n118_n140# 0.02fF
C71 a_60_n140# a_n118_n140# 0.13fF
C72 a_n1364_n140# a_n1898_n140# 0.04fF
C73 a_772_n140# a_1306_n140# 0.04fF
C74 a_n830_n140# a_n296_n140# 0.04fF
C75 a_118_n205# a_1542_n205# 0.01fF
C76 a_594_n140# a_238_n140# 0.06fF
C77 a_118_n205# a_652_n205# 0.02fF
C78 a_1484_n140# a_1128_n140# 0.06fF
C79 a_n830_n140# a_n1720_n140# 0.02fF
C80 a_n1008_n140# a_416_n140# 0.01fF
C81 a_474_n205# w_n2112_n241# 0.24fF
C82 a_1484_n140# a_772_n140# 0.03fF
C83 a_n652_n140# a_238_n140# 0.02fF
C84 w_n2112_n241# a_n416_n205# 0.24fF
C85 w_n2112_n241# a_594_n140# 0.02fF
C86 a_296_n205# a_1364_n205# 0.01fF
C87 a_n652_n140# w_n2112_n241# 0.02fF
C88 a_118_n205# a_n772_n205# 0.01fF
C89 a_474_n205# a_n416_n205# 0.01fF
C90 a_118_n205# a_n60_n205# 0.11fF
C91 a_1898_n205# a_1720_n205# 0.11fF
C92 a_n830_n140# a_n1186_n140# 0.06fF
C93 a_1898_n205# a_830_n205# 0.01fF
C94 a_n1364_n140# a_n474_n140# 0.02fF
C95 a_n474_n140# a_60_n140# 0.04fF
C96 a_n772_n205# a_n1662_n205# 0.01fF
C97 a_n60_n205# a_n1662_n205# 0.01fF
C98 a_n238_n205# a_1186_n205# 0.01fF
C99 a_n652_n140# a_594_n140# 0.02fF
C100 a_n1008_n140# a_n296_n140# 0.03fF
C101 w_n2112_n241# a_2018_n140# 0.02fF
C102 a_n1484_n205# a_n60_n205# 0.01fF
C103 a_n1128_n205# a_n1306_n205# 0.11fF
C104 a_n772_n205# a_n1484_n205# 0.01fF
C105 a_n830_n140# a_n2076_n140# 0.02fF
C106 a_n1008_n140# a_n1720_n140# 0.03fF
C107 a_n594_n205# a_1008_n205# 0.01fF
C108 a_1840_n140# a_950_n140# 0.02fF
C109 a_118_n205# a_1364_n205# 0.01fF
C110 a_416_n140# a_n118_n140# 0.04fF
C111 w_n2112_n241# a_1186_n205# 0.21fF
C112 a_2018_n140# a_594_n140# 0.01fF
C113 a_n1364_n140# a_238_n140# 0.01fF
C114 a_238_n140# a_60_n140# 0.13fF
C115 a_n1008_n140# a_n1186_n140# 0.13fF
C116 a_n1364_n140# w_n2112_n241# 0.02fF
C117 a_474_n205# a_1186_n205# 0.01fF
C118 w_n2112_n241# a_60_n140# 0.02fF
C119 a_n416_n205# a_1186_n205# 0.01fF
C120 a_1898_n205# a_1542_n205# 0.03fF
C121 a_1898_n205# a_652_n205# 0.01fF
C122 a_n1008_n140# a_n2076_n140# 0.02fF
C123 a_n238_n205# a_1008_n205# 0.01fF
C124 a_594_n140# a_60_n140# 0.04fF
C125 a_n296_n140# a_n118_n140# 0.13fF
C126 a_1128_n140# a_950_n140# 0.13fF
C127 a_n296_n140# a_n1898_n140# 0.01fF
C128 a_416_n140# a_n474_n140# 0.02fF
C129 a_n118_n140# a_1306_n140# 0.01fF
C130 a_n1364_n140# a_n652_n140# 0.03fF
C131 a_n1720_n140# a_n118_n140# 0.01fF
C132 a_950_n140# a_772_n140# 0.13fF
C133 a_n594_n205# a_830_n205# 0.01fF
C134 a_1662_n140# a_238_n140# 0.01fF
C135 a_n652_n140# a_60_n140# 0.03fF
C136 a_n1840_n205# a_n1662_n205# 0.11fF
C137 a_n830_n140# a_n1542_n140# 0.03fF
C138 a_296_n205# a_118_n205# 0.11fF
C139 a_n1720_n140# a_n1898_n140# 0.13fF
C140 a_n1128_n205# a_n60_n205# 0.01fF
C141 a_n1306_n205# a_n594_n205# 0.01fF
C142 a_n1128_n205# a_n772_n205# 0.03fF
C143 a_n1840_n205# a_n1484_n205# 0.03fF
C144 a_1662_n140# w_n2112_n241# 0.02fF
C145 w_n2112_n241# a_1008_n205# 0.22fF
C146 a_1484_n140# a_n118_n140# 0.01fF
C147 a_n1186_n140# a_n118_n140# 0.02fF
C148 a_n1186_n140# a_n1898_n140# 0.03fF
C149 a_474_n205# a_1008_n205# 0.02fF
C150 a_n416_n205# a_1008_n205# 0.01fF
C151 a_1662_n140# a_594_n140# 0.02fF
C152 a_1898_n205# a_1364_n205# 0.02fF
C153 a_n296_n140# a_n474_n140# 0.13fF
C154 a_416_n140# a_238_n140# 0.13fF
C155 a_n1306_n205# a_n2018_n205# 0.01fF
C156 a_n474_n140# a_n1720_n140# 0.02fF
C157 a_n238_n205# a_830_n205# 0.01fF
C158 a_n1008_n140# a_n1542_n140# 0.04fF
C159 a_n1898_n140# a_n2076_n140# 0.13fF
C160 a_1840_n140# a_1128_n140# 0.03fF
C161 w_n2112_n241# a_416_n140# 0.02fF
C162 a_1840_n140# a_772_n140# 0.02fF
C163 a_n1306_n205# a_n950_n205# 0.03fF
C164 a_n1306_n205# a_n238_n205# 0.01fF
C165 a_n594_n205# a_652_n205# 0.01fF
C166 a_n1364_n140# a_60_n140# 0.01fF
C167 a_n1186_n140# a_n474_n140# 0.03fF
C168 a_1662_n140# a_2018_n140# 0.06fF
C169 a_416_n140# a_594_n140# 0.13fF
C170 w_n2112_n241# a_1720_n205# 0.18fF
C171 a_118_n205# a_n1484_n205# 0.01fF
C172 a_n296_n140# a_238_n140# 0.04fF
C173 w_n2112_n241# a_830_n205# 0.23fF
C174 a_n652_n140# a_416_n140# 0.02fF
C175 a_n594_n205# a_n772_n205# 0.11fF
C176 a_238_n140# a_1306_n140# 0.02fF
C177 a_n594_n205# a_n60_n205# 0.02fF
C178 a_n1128_n205# a_n1840_n205# 0.01fF
C179 a_n1306_n205# w_n2112_n241# 0.24fF
C180 w_n2112_n241# a_n296_n140# 0.02fF
C181 a_474_n205# a_1720_n205# 0.01fF
C182 a_296_n205# a_1898_n205# 0.01fF
C183 a_n1484_n205# a_n1662_n205# 0.11fF
C184 a_n474_n140# a_n2076_n140# 0.01fF
C185 a_474_n205# a_830_n205# 0.03fF
C186 a_1186_n205# a_1008_n205# 0.11fF
C187 a_n416_n205# a_830_n205# 0.01fF
C188 w_n2112_n241# a_1306_n140# 0.02fF
C189 w_n2112_n241# a_n1720_n140# 0.02fF
C190 a_1484_n140# a_238_n140# 0.02fF
C191 a_296_n205# a_n1128_n205# 0.01fF
C192 a_n1306_n205# a_n416_n205# 0.01fF
C193 a_1662_n140# a_60_n140# 0.01fF
C194 a_416_n140# a_2018_n140# 0.01fF
C195 a_n1186_n140# a_238_n140# 0.01fF
C196 a_1128_n140# a_772_n140# 0.06fF
C197 a_n950_n205# a_652_n205# 0.01fF
C198 a_n238_n205# a_652_n205# 0.01fF
C199 a_n1542_n140# a_n118_n140# 0.01fF
C200 a_n296_n140# a_594_n140# 0.02fF
C201 a_n772_n205# a_n2018_n205# 0.01fF
C202 a_1484_n140# w_n2112_n241# 0.02fF
C203 a_n1898_n140# a_n1542_n140# 0.06fF
C204 a_594_n140# a_1306_n140# 0.03fF
C205 a_n652_n140# a_n296_n140# 0.06fF
C206 w_n2112_n241# a_n1186_n140# 0.02fF
C207 a_950_n140# a_n118_n140# 0.02fF
C208 a_n830_n140# a_772_n140# 0.01fF
C209 a_n652_n140# a_n1720_n140# 0.02fF
C210 a_n772_n205# a_n950_n205# 0.11fF
C211 a_n772_n205# a_n238_n205# 0.02fF
C212 a_n950_n205# a_n60_n205# 0.01fF
C213 a_n60_n205# a_n238_n205# 0.11fF
C214 a_1484_n140# a_594_n140# 0.02fF
C215 w_n2112_n241# a_1542_n205# 0.19fF
C216 w_n2112_n241# a_652_n205# 0.24fF
C217 a_416_n140# a_60_n140# 0.06fF
C218 w_n2112_n241# a_n2076_n140# 0.02fF
C219 a_118_n205# a_n1128_n205# 0.01fF
C220 a_n652_n140# a_n1186_n140# 0.04fF
C221 a_474_n205# a_1542_n205# 0.01fF
C222 a_2018_n140# a_1306_n140# 0.03fF
C223 a_1720_n205# a_1186_n205# 0.02fF
C224 a_1186_n205# a_830_n205# 0.03fF
C225 a_474_n205# a_652_n205# 0.11fF
C226 a_n474_n140# a_n1542_n140# 0.02fF
C227 a_n416_n205# a_652_n205# 0.01fF
C228 a_n1840_n205# a_n594_n205# 0.01fF
C229 w_n2112_n241# a_n60_n205# 0.24fF
C230 w_n2112_n241# a_n772_n205# 0.24fF
C231 a_n1128_n205# a_n1662_n205# 0.02fF
C232 a_950_n140# a_n474_n140# 0.01fF
C233 a_n238_n205# a_1364_n205# 0.01fF
C234 a_1484_n140# a_2018_n140# 0.04fF
C235 a_n652_n140# a_n2076_n140# 0.01fF
C236 a_474_n205# a_n772_n205# 0.01fF
C237 a_296_n205# a_n594_n205# 0.01fF
C238 a_474_n205# a_n60_n205# 0.02fF
C239 a_n1128_n205# a_n1484_n205# 0.03fF
C240 a_n772_n205# a_n416_n205# 0.03fF
C241 a_n60_n205# a_n416_n205# 0.03fF
C242 a_n1364_n140# a_n296_n140# 0.02fF
C243 a_n296_n140# a_60_n140# 0.06fF
C244 a_n830_n140# a_n1008_n140# 0.13fF
C245 a_1662_n140# a_416_n140# 0.02fF
C246 a_60_n140# a_1306_n140# 0.02fF
C247 a_n1364_n140# a_n1720_n140# 0.06fF
C248 a_n1840_n205# a_n2018_n205# 0.11fF
C249 w_n2112_n241# a_1364_n205# 0.20fF
C250 a_950_n140# a_238_n140# 0.03fF
C251 a_1484_n140# a_60_n140# 0.01fF
C252 a_n1840_n205# a_n238_n205# 0.01fF
C253 a_n1840_n205# a_n950_n205# 0.01fF
C254 w_n2112_n241# a_n1542_n140# 0.02fF
C255 a_n1364_n140# a_n1186_n140# 0.13fF
C256 a_n1186_n140# a_60_n140# 0.02fF
C257 a_1542_n205# a_1186_n205# 0.03fF
C258 a_474_n205# a_1364_n205# 0.01fF
C259 a_1720_n205# a_1008_n205# 0.01fF
C260 a_1186_n205# a_652_n205# 0.02fF
C261 a_1008_n205# a_830_n205# 0.11fF
C262 w_n2112_n241# a_950_n140# 0.02fF
C263 a_296_n205# a_n950_n205# 0.01fF
C264 a_118_n205# a_n594_n205# 0.01fF
C265 a_296_n205# a_n238_n205# 0.02fF
C266 a_1128_n140# a_n118_n140# 0.02fF
C267 a_1662_n140# a_1306_n140# 0.06fF
C268 a_772_n140# a_n118_n140# 0.02fF
C269 a_n1364_n140# a_n2076_n140# 0.03fF
C270 a_n1840_n205# w_n2112_n241# 0.24fF
C271 a_n594_n205# a_n1662_n205# 0.01fF
C272 a_n60_n205# a_1186_n205# 0.01fF
C273 a_n652_n140# a_n1542_n140# 0.02fF
C274 a_950_n140# a_594_n140# 0.06fF
C275 a_n830_n140# a_n118_n140# 0.03fF
C276 a_n652_n140# a_950_n140# 0.01fF
C277 a_1484_n140# a_1662_n140# 0.13fF
C278 a_n594_n205# a_n1484_n205# 0.01fF
C279 a_n830_n140# a_n1898_n140# 0.02fF
C280 a_296_n205# w_n2112_n241# 0.24fF
C281 a_n1840_n205# a_n416_n205# 0.01fF
C282 a_1840_n140# a_238_n140# 0.01fF
C283 a_416_n140# a_n296_n140# 0.03fF
C284 a_n1662_n205# a_n2018_n205# 0.03fF
C285 a_474_n205# a_296_n205# 0.11fF
C286 a_416_n140# a_1306_n140# 0.02fF
C287 a_118_n205# a_n950_n205# 0.01fF
C288 a_118_n205# a_n238_n205# 0.03fF
C289 a_296_n205# a_n416_n205# 0.01fF
C290 a_1128_n140# a_n474_n140# 0.01fF
C291 a_950_n140# a_2018_n140# 0.02fF
C292 a_1840_n140# w_n2112_n241# 0.02fF
C293 a_1720_n205# a_830_n205# 0.01fF
C294 a_1364_n205# a_1186_n205# 0.11fF
C295 a_1542_n205# a_1008_n205# 0.02fF
C296 a_1008_n205# a_652_n205# 0.03fF
C297 a_n474_n140# a_772_n140# 0.02fF
C298 a_n1484_n205# a_n2018_n205# 0.02fF
C299 a_n950_n205# a_n1662_n205# 0.01fF
C300 a_n238_n205# a_n1662_n205# 0.01fF
C301 a_1484_n140# a_416_n140# 0.02fF
C302 a_n830_n140# a_n474_n140# 0.06fF
C303 a_416_n140# a_n1186_n140# 0.01fF
C304 a_n1008_n140# a_n118_n140# 0.02fF
C305 a_1840_n140# a_594_n140# 0.02fF
C306 a_n950_n205# a_n1484_n205# 0.02fF
C307 a_n1484_n205# a_n238_n205# 0.01fF
C308 a_n1008_n140# a_n1898_n140# 0.02fF
C309 a_n60_n205# a_1008_n205# 0.01fF
C310 a_n1364_n140# a_n1542_n140# 0.13fF
C311 a_n1542_n140# a_60_n140# 0.01fF
C312 a_118_n205# w_n2112_n241# 0.24fF
C313 a_n296_n140# a_1306_n140# 0.01fF
C314 a_n296_n140# a_n1720_n140# 0.01fF
C315 a_950_n140# a_60_n140# 0.02fF
C316 a_1128_n140# a_238_n140# 0.02fF
C317 a_474_n205# a_118_n205# 0.03fF
C318 w_n2112_n241# a_n1662_n205# 0.24fF
C319 a_118_n205# a_n416_n205# 0.02fF
C320 a_772_n140# a_238_n140# 0.04fF
C321 a_n1128_n205# a_n594_n205# 0.02fF
C322 w_n2112_n241# a_n1484_n205# 0.24fF
C323 a_1128_n140# w_n2112_n241# 0.02fF
C324 a_296_n205# a_1186_n205# 0.01fF
C325 a_n830_n140# a_238_n140# 0.02fF
C326 a_1840_n140# a_2018_n140# 0.13fF
C327 w_n2112_n241# a_772_n140# 0.02fF
C328 a_n416_n205# a_n1662_n205# 0.01fF
C329 a_1484_n140# a_1306_n140# 0.13fF
C330 a_n1186_n140# a_n296_n140# 0.02fF
C331 a_1720_n205# a_1542_n205# 0.11fF
C332 a_1542_n205# a_830_n205# 0.01fF
C333 a_1720_n205# a_652_n205# 0.01fF
C334 a_1364_n205# a_1008_n205# 0.03fF
C335 a_n1008_n140# a_n474_n140# 0.04fF
C336 a_830_n205# a_652_n205# 0.11fF
C337 a_n1186_n140# a_n1720_n140# 0.04fF
C338 a_n830_n140# w_n2112_n241# 0.02fF
C339 a_n1484_n205# a_n416_n205# 0.01fF
C340 a_1128_n140# a_594_n140# 0.04fF
C341 a_594_n140# a_772_n140# 0.13fF
C342 a_n1128_n205# a_n2018_n205# 0.01fF
C343 a_1662_n140# a_950_n140# 0.03fF
C344 a_n772_n205# a_830_n205# 0.01fF
C345 a_n60_n205# a_830_n205# 0.01fF
C346 a_n652_n140# a_772_n140# 0.01fF
C347 a_n1720_n140# a_n2076_n140# 0.06fF
C348 a_n830_n140# a_594_n140# 0.01fF
C349 a_n1306_n205# a_n772_n205# 0.02fF
C350 a_n1306_n205# a_n60_n205# 0.01fF
C351 a_n1128_n205# a_n950_n205# 0.11fF
C352 a_n1128_n205# a_n238_n205# 0.01fF
C353 a_n652_n140# a_n830_n140# 0.13fF
C354 a_118_n205# a_1186_n205# 0.01fF
C355 a_n1008_n140# a_238_n140# 0.02fF
C356 a_1128_n140# a_2018_n140# 0.02fF
C357 a_n1186_n140# a_n2076_n140# 0.02fF
C358 a_2018_n140# a_772_n140# 0.02fF
C359 w_n2112_n241# a_1898_n205# 0.24fF
C360 a_296_n205# a_1008_n205# 0.01fF
C361 a_n1008_n140# w_n2112_n241# 0.02fF
C362 a_950_n140# a_416_n140# 0.04fF
C363 a_1720_n205# a_1364_n205# 0.03fF
C364 a_1364_n205# a_830_n205# 0.02fF
C365 a_1542_n205# a_652_n205# 0.01fF
C366 a_n1128_n205# w_n2112_n241# 0.24fF
C367 a_n474_n140# a_n118_n140# 0.06fF
C368 a_474_n205# a_1898_n205# 0.01fF
C369 a_n474_n140# a_n1898_n140# 0.01fF
C370 a_1840_n140# a_1662_n140# 0.13fF
C371 a_n1008_n140# a_594_n140# 0.01fF
C372 a_474_n205# a_n1128_n205# 0.01fF
C373 a_n1128_n205# a_n416_n205# 0.01fF
C374 a_1128_n140# a_60_n140# 0.02fF
C375 a_n60_n205# a_1542_n205# 0.01fF
C376 a_n296_n140# a_n1542_n140# 0.02fF
C377 a_n652_n140# a_n1008_n140# 0.06fF
C378 a_n772_n205# a_652_n205# 0.01fF
C379 a_n60_n205# a_652_n205# 0.01fF
C380 w_n2112_n241# VSUBS 6.11fF
.ends

.subckt sky130_fd_pr__pfet_01v8_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136# VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_n128_n136# a_256_n136# 0.05fF
C1 a_n224_n136# a_448_n136# 0.03fF
C2 a_n224_n136# a_n416_n136# 0.12fF
C3 a_160_n136# a_352_n136# 0.12fF
C4 w_n646_n356# a_64_n136# 0.05fF
C5 a_n508_n136# a_n224_n136# 0.07fF
C6 a_n320_n136# a_n512_n234# 0.06fF
C7 a_n512_n234# a_n128_n136# 0.06fF
C8 a_n32_n136# a_352_n136# 0.05fF
C9 w_n646_n356# a_448_n136# 0.13fF
C10 w_n646_n356# a_n416_n136# 0.08fF
C11 a_n320_n136# a_64_n136# 0.05fF
C12 a_64_n136# a_n128_n136# 0.12fF
C13 w_n646_n356# a_n508_n136# 0.13fF
C14 a_n320_n136# a_448_n136# 0.02fF
C15 a_n320_n136# a_n416_n136# 0.33fF
C16 a_448_n136# a_n128_n136# 0.03fF
C17 a_256_n136# a_352_n136# 0.33fF
C18 a_n128_n136# a_n416_n136# 0.07fF
C19 a_n32_n136# a_160_n136# 0.12fF
C20 a_n508_n136# a_n320_n136# 0.12fF
C21 a_n508_n136# a_n128_n136# 0.05fF
C22 w_n646_n356# a_n224_n136# 0.06fF
C23 a_64_n136# a_352_n136# 0.07fF
C24 a_160_n136# a_256_n136# 0.33fF
C25 a_n32_n136# a_256_n136# 0.07fF
C26 a_448_n136# a_352_n136# 0.33fF
C27 a_n320_n136# a_n224_n136# 0.33fF
C28 a_352_n136# a_n416_n136# 0.02fF
C29 a_n224_n136# a_n128_n136# 0.33fF
C30 a_n508_n136# a_352_n136# 0.02fF
C31 a_64_n136# a_160_n136# 0.33fF
C32 w_n646_n356# a_n320_n136# 0.06fF
C33 w_n646_n356# a_n128_n136# 0.05fF
C34 a_64_n136# a_n32_n136# 0.33fF
C35 a_448_n136# a_160_n136# 0.07fF
C36 a_160_n136# a_n416_n136# 0.03fF
C37 a_n508_n136# a_160_n136# 0.03fF
C38 a_n512_n234# a_256_n136# 0.06fF
C39 a_n320_n136# a_n128_n136# 0.12fF
C40 a_448_n136# a_n32_n136# 0.04fF
C41 a_n32_n136# a_n416_n136# 0.05fF
C42 a_n224_n136# a_352_n136# 0.03fF
C43 a_n508_n136# a_n32_n136# 0.04fF
C44 a_64_n136# a_256_n136# 0.12fF
C45 w_n646_n356# a_352_n136# 0.08fF
C46 a_448_n136# a_256_n136# 0.12fF
C47 a_n512_n234# a_64_n136# 0.06fF
C48 a_256_n136# a_n416_n136# 0.03fF
C49 a_n508_n136# a_256_n136# 0.02fF
C50 a_n224_n136# a_160_n136# 0.05fF
C51 a_n512_n234# a_448_n136# 0.06fF
C52 a_n320_n136# a_352_n136# 0.03fF
C53 a_n128_n136# a_352_n136# 0.04fF
C54 a_n224_n136# a_n32_n136# 0.12fF
C55 a_n508_n136# a_n512_n234# 0.06fF
C56 w_n646_n356# a_160_n136# 0.06fF
C57 a_64_n136# a_448_n136# 0.05fF
C58 a_64_n136# a_n416_n136# 0.04fF
C59 a_n508_n136# a_64_n136# 0.03fF
C60 w_n646_n356# a_n32_n136# 0.05fF
C61 a_448_n136# a_n416_n136# 0.02fF
C62 a_n224_n136# a_256_n136# 0.04fF
C63 a_n320_n136# a_160_n136# 0.04fF
C64 a_n128_n136# a_160_n136# 0.07fF
C65 a_n508_n136# a_448_n136# 0.02fF
C66 a_n508_n136# a_n416_n136# 0.33fF
C67 a_n320_n136# a_n32_n136# 0.07fF
C68 a_n32_n136# a_n128_n136# 0.33fF
C69 w_n646_n356# a_256_n136# 0.06fF
C70 a_n224_n136# a_64_n136# 0.07fF
C71 w_n646_n356# a_n512_n234# 1.13fF
C72 a_n320_n136# a_256_n136# 0.03fF
C73 w_n646_n356# VSUBS 2.52fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
X0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_n32_n52# a_n128_n52# 0.13fF
C1 a_n224_n52# a_n508_n52# 0.03fF
C2 a_n320_n52# a_n128_n52# 0.05fF
C3 a_448_n52# a_n128_n52# 0.01fF
C4 a_160_n52# a_n128_n52# 0.03fF
C5 a_n224_n52# a_256_n52# 0.02fF
C6 a_n224_n52# a_n416_n52# 0.05fF
C7 a_n512_n140# a_64_n52# 0.09fF
C8 a_n508_n52# a_352_n52# 0.01fF
C9 a_n224_n52# a_64_n52# 0.03fF
C10 a_n508_n52# a_n32_n52# 0.02fF
C11 a_256_n52# a_352_n52# 0.13fF
C12 a_n508_n52# a_n320_n52# 0.05fF
C13 a_n416_n52# a_352_n52# 0.01fF
C14 a_n508_n52# a_448_n52# 0.01fF
C15 a_n32_n52# a_256_n52# 0.03fF
C16 a_n508_n52# a_160_n52# 0.01fF
C17 a_n416_n52# a_n32_n52# 0.02fF
C18 a_n320_n52# a_256_n52# 0.01fF
C19 a_n416_n52# a_n320_n52# 0.13fF
C20 a_256_n52# a_448_n52# 0.05fF
C21 a_n416_n52# a_448_n52# 0.01fF
C22 a_64_n52# a_352_n52# 0.03fF
C23 a_160_n52# a_256_n52# 0.13fF
C24 a_n416_n52# a_160_n52# 0.01fF
C25 a_n508_n52# a_n128_n52# 0.02fF
C26 a_n32_n52# a_64_n52# 0.13fF
C27 a_n320_n52# a_64_n52# 0.02fF
C28 a_64_n52# a_448_n52# 0.02fF
C29 a_256_n52# a_n128_n52# 0.02fF
C30 a_n416_n52# a_n128_n52# 0.03fF
C31 a_64_n52# a_160_n52# 0.13fF
C32 a_64_n52# a_n128_n52# 0.05fF
C33 a_n512_n140# a_n320_n52# 0.09fF
C34 a_n224_n52# a_352_n52# 0.01fF
C35 a_n512_n140# a_448_n52# 0.09fF
C36 a_n508_n52# a_256_n52# 0.01fF
C37 a_n508_n52# a_n416_n52# 0.13fF
C38 a_n224_n52# a_n32_n52# 0.05fF
C39 a_n224_n52# a_n320_n52# 0.13fF
C40 a_n416_n52# a_256_n52# 0.01fF
C41 a_n224_n52# a_448_n52# 0.01fF
C42 a_n224_n52# a_160_n52# 0.02fF
C43 a_n512_n140# a_n128_n52# 0.09fF
C44 a_n508_n52# a_64_n52# 0.01fF
C45 a_64_n52# a_256_n52# 0.05fF
C46 a_n32_n52# a_352_n52# 0.02fF
C47 a_n416_n52# a_64_n52# 0.02fF
C48 a_n224_n52# a_n128_n52# 0.13fF
C49 a_n320_n52# a_352_n52# 0.01fF
C50 a_352_n52# a_448_n52# 0.13fF
C51 a_n320_n52# a_n32_n52# 0.03fF
C52 a_160_n52# a_352_n52# 0.05fF
C53 a_n32_n52# a_448_n52# 0.02fF
C54 a_n32_n52# a_160_n52# 0.05fF
C55 a_n512_n140# a_n508_n52# 0.09fF
C56 a_n320_n52# a_448_n52# 0.01fF
C57 a_n320_n52# a_160_n52# 0.02fF
C58 a_160_n52# a_448_n52# 0.03fF
C59 a_352_n52# a_n128_n52# 0.02fF
C60 a_n512_n140# a_256_n52# 0.09fF
C61 a_448_n52# a_n610_n226# 0.07fF
C62 a_352_n52# a_n610_n226# 0.05fF
C63 a_256_n52# a_n610_n226# 0.04fF
C64 a_160_n52# a_n610_n226# 0.04fF
C65 a_64_n52# a_n610_n226# 0.04fF
C66 a_n32_n52# a_n610_n226# 0.04fF
C67 a_n128_n52# a_n610_n226# 0.04fF
C68 a_n224_n52# a_n610_n226# 0.04fF
C69 a_n320_n52# a_n610_n226# 0.04fF
C70 a_n416_n52# a_n610_n226# 0.05fF
C71 a_n508_n52# a_n610_n226# 0.07fF
C72 a_n512_n140# a_n610_n226# 1.45fF
.ends

.subckt transmission_gate en VDD in out VSS en_b
Xsky130_fd_pr__pfet_01v8_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ VSS sky130_fd_pr__pfet_01v8_UNG2NQ
Xsky130_fd_pr__nfet_01v8_6J4AMR_0 out in in out in in VSS out en in out out out sky130_fd_pr__nfet_01v8_6J4AMR
C0 out VDD 0.40fF
C1 out en_b 0.03fF
C2 en out 0.05fF
C3 VDD en_b 0.10fF
C4 in out 0.71fF
C5 en VDD 0.05fF
C6 en en_b 0.14fF
C7 in VDD 0.92fF
C8 in en_b 1.18fF
C9 en in 1.30fF
C10 en VSS 1.66fF
C11 out VSS 1.04fF
C12 in VSS 1.15fF
C13 en_b VSS 0.24fF
C14 VDD VSS 3.18fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 c1_n530_n480# m3_n630_n580# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb cmc unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580#
+ on unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_8/in transmission_gate_4/out
+ bias_a p2_b p1 cm transmission_gate_9/in p2 VDD transmission_gate_3/out transmission_gate_7/in
+ op VSS p1_b
Xtransmission_gate_10 p1 VDD transmission_gate_3/out on VSS p1_b transmission_gate
Xtransmission_gate_11 p1 VDD transmission_gate_4/out op VSS p1_b transmission_gate
Xtransmission_gate_0 p1 VDD cm transmission_gate_7/in VSS p1_b transmission_gate
Xtransmission_gate_1 p1 VDD cm transmission_gate_6/in VSS p1_b transmission_gate
Xtransmission_gate_2 p1 VDD bias_a transmission_gate_8/in VSS p1_b transmission_gate
Xtransmission_gate_3 p2 VDD cm transmission_gate_3/out VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 VDD cm transmission_gate_4/out VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 VDD bias_a transmission_gate_9/in VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 VDD transmission_gate_6/in op VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 VDD transmission_gate_7/in on VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 VDD transmission_gate_8/in cmc VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 VDD transmission_gate_9/in cmc VSS p1_b transmission_gate
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_4/out 0.57fF
C1 transmission_gate_9/in p1_b 0.00fF
C2 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_34/c1_n530_n480# -0.19fF
C3 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_25/c1_n530_n480# -0.19fF
C4 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# 0.10fF
C5 transmission_gate_7/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.63fF
C6 VDD transmission_gate_3/out 0.27fF
C7 transmission_gate_8/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C8 transmission_gate_7/in p2 -0.01fF
C9 cmc unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C10 bias_a p1_b 0.04fF
C11 transmission_gate_4/out unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C12 VDD unit_cap_mim_m3m4_35/c1_n530_n480# -0.06fF
C13 transmission_gate_7/in unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C14 p2 transmission_gate_8/in -0.01fF
C15 cmc unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C16 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_24/c1_n530_n480# -0.24fF
C17 p1 unit_cap_mim_m3m4_23/m3_n630_n580# -0.71fF
C18 transmission_gate_6/in p1_b 0.04fF
C19 unit_cap_mim_m3m4_17/c1_n530_n480# p2_b -0.07fF
C20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C21 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C22 transmission_gate_9/in p2_b 0.03fF
C23 on unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C24 transmission_gate_7/in op 2.64fF
C25 cm unit_cap_mim_m3m4_19/c1_n530_n480# -0.22fF
C26 unit_cap_mim_m3m4_20/m3_n630_n580# p2_b -0.65fF
C27 transmission_gate_9/in on 0.79fF
C28 transmission_gate_8/in op 0.88fF
C29 VDD unit_cap_mim_m3m4_22/m3_n630_n580# 0.33fF
C30 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_23/c1_n530_n480# -0.20fF
C31 cmc p1_b 0.31fF
C32 bias_a p2_b 0.06fF
C33 unit_cap_mim_m3m4_20/m3_n630_n580# on 0.40fF
C34 VDD unit_cap_mim_m3m4_35/m3_n630_n580# -0.40fF
C35 transmission_gate_7/in transmission_gate_3/out 0.28fF
C36 transmission_gate_7/in VDD 0.25fF
C37 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580# -0.33fF
C38 transmission_gate_3/out transmission_gate_8/in 0.24fF
C39 VDD transmission_gate_8/in 0.21fF
C40 unit_cap_mim_m3m4_17/c1_n530_n480# p2 -0.25fF
C41 unit_cap_mim_m3m4_35/c1_n530_n480# transmission_gate_8/in -0.01fF
C42 transmission_gate_6/in p2_b 0.02fF
C43 p2 transmission_gate_9/in 0.02fF
C44 transmission_gate_6/in on 0.40fF
C45 unit_cap_mim_m3m4_30/m3_n630_n580# p1_b -0.72fF
C46 unit_cap_mim_m3m4_20/m3_n630_n580# p2 -0.71fF
C47 cm p1 0.12fF
C48 cmc p2_b 0.03fF
C49 p2 bias_a 0.05fF
C50 unit_cap_mim_m3m4_32/c1_n530_n480# on 0.06fF
C51 unit_cap_mim_m3m4_17/c1_n530_n480# op 0.06fF
C52 transmission_gate_4/out p1 0.01fF
C53 unit_cap_mim_m3m4_21/m3_n630_n580# p2_b -0.72fF
C54 cmc on 2.26fF
C55 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C56 transmission_gate_9/in op 0.68fF
C57 transmission_gate_6/in p2 0.00fF
C58 transmission_gate_6/in unit_cap_mim_m3m4_28/c1_n530_n480# -0.32fF
C59 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C60 unit_cap_mim_m3m4_31/m3_n630_n580# op 0.02fF
C61 VDD unit_cap_mim_m3m4_18/c1_n530_n480# -0.06fF
C62 transmission_gate_8/in unit_cap_mim_m3m4_35/m3_n630_n580# 0.58fF
C63 transmission_gate_7/in transmission_gate_8/in -0.06fF
C64 unit_cap_mim_m3m4_17/c1_n530_n480# transmission_gate_3/out -0.03fF
C65 unit_cap_mim_m3m4_17/c1_n530_n480# VDD -0.06fF
C66 transmission_gate_4/out unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C67 transmission_gate_3/out transmission_gate_9/in 2.49fF
C68 VDD transmission_gate_9/in 0.21fF
C69 p2 cmc 0.61fF
C70 VDD unit_cap_mim_m3m4_20/m3_n630_n580# 0.33fF
C71 unit_cap_mim_m3m4_31/c1_n530_n480# transmission_gate_4/out 0.06fF
C72 transmission_gate_6/in unit_cap_mim_m3m4_27/c1_n530_n480# -0.04fF
C73 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C74 unit_cap_mim_m3m4_21/m3_n630_n580# p2 -1.16fF
C75 transmission_gate_6/in op 0.68fF
C76 VDD bias_a -0.01fF
C77 transmission_gate_3/out bias_a 0.05fF
C78 unit_cap_mim_m3m4_35/c1_n530_n480# bias_a -0.22fF
C79 unit_cap_mim_m3m4_19/c1_n530_n480# p1_b 0.07fF
C80 p1 unit_cap_mim_m3m4_18/m3_n630_n580# -0.55fF
C81 unit_cap_mim_m3m4_24/c1_n530_n480# p2_b -0.07fF
C82 transmission_gate_6/in transmission_gate_3/out 0.76fF
C83 transmission_gate_6/in VDD 0.31fF
C84 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C85 cmc op 4.31fF
C86 transmission_gate_4/out cm 0.08fF
C87 unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_9/in 0.59fF
C88 unit_cap_mim_m3m4_17/m3_n630_n580# cm 0.41fF
C89 cm unit_cap_mim_m3m4_16/c1_n530_n480# -0.22fF
C90 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C91 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C92 transmission_gate_7/in transmission_gate_9/in 0.02fF
C93 transmission_gate_3/out cmc 0.79fF
C94 VDD cmc 0.66fF
C95 transmission_gate_9/in transmission_gate_8/in 3.34fF
C96 transmission_gate_7/in unit_cap_mim_m3m4_20/m3_n630_n580# 0.64fF
C97 transmission_gate_4/out unit_cap_mim_m3m4_16/c1_n530_n480# 0.03fF
C98 p1 p1_b 2.54fF
C99 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_8/in 0.17fF
C100 unit_cap_mim_m3m4_24/c1_n530_n480# p2 -0.30fF
C101 VDD unit_cap_mim_m3m4_21/m3_n630_n580# 0.33fF
C102 unit_cap_mim_m3m4_30/m3_n630_n580# op 0.31fF
C103 bias_a unit_cap_mim_m3m4_35/m3_n630_n580# 0.33fF
C104 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_28/c1_n530_n480# -0.17fF
C105 unit_cap_mim_m3m4_23/m3_n630_n580# p1_b -1.03fF
C106 unit_cap_mim_m3m4_16/m3_n630_n580# cm 0.36fF
C107 transmission_gate_7/in bias_a 0.09fF
C108 unit_cap_mim_m3m4_29/m3_n630_n580# p2_b -0.58fF
C109 bias_a transmission_gate_8/in 0.04fF
C110 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.17fF
C111 unit_cap_mim_m3m4_23/c1_n530_n480# p1_b 0.13fF
C112 unit_cap_mim_m3m4_16/m3_n630_n580# transmission_gate_4/out 0.62fF
C113 unit_cap_mim_m3m4_30/m3_n630_n580# VDD 0.28fF
C114 transmission_gate_6/in transmission_gate_7/in 0.44fF
C115 cm unit_cap_mim_m3m4_18/m3_n630_n580# 0.39fF
C116 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.12fF
C117 unit_cap_mim_m3m4_30/c1_n530_n480# op 0.05fF
C118 transmission_gate_6/in transmission_gate_8/in -0.10fF
C119 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.10fF
C120 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_16/c1_n530_n480# -0.35fF
C121 unit_cap_mim_m3m4_22/m3_n630_n580# cmc 0.60fF
C122 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C123 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_19/c1_n530_n480# -0.34fF
C124 unit_cap_mim_m3m4_28/m3_n630_n580# op 0.66fF
C125 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C126 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.17fF
C127 transmission_gate_7/in cmc 0.07fF
C128 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C129 p2 unit_cap_mim_m3m4_29/m3_n630_n580# -0.78fF
C130 cmc transmission_gate_8/in 8.00fF
C131 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C132 on p1 0.22fF
C133 VDD unit_cap_mim_m3m4_24/c1_n530_n480# -0.06fF
C134 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_27/c1_n530_n480# -0.13fF
C135 on unit_cap_mim_m3m4_23/m3_n630_n580# 0.02fF
C136 unit_cap_mim_m3m4_21/m3_n630_n580# transmission_gate_8/in 0.59fF
C137 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C138 unit_cap_mim_m3m4_27/m3_n630_n580# op 0.28fF
C139 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_32/c1_n530_n480# -0.15fF
C140 unit_cap_mim_m3m4_31/m3_n630_n580# transmission_gate_9/in 0.10fF
C141 unit_cap_mim_m3m4_32/m3_n630_n580# cmc 0.10fF
C142 unit_cap_mim_m3m4_33/c1_n530_n480# op 0.06fF
C143 cm p1_b 0.27fF
C144 transmission_gate_9/in bias_a 0.02fF
C145 cmc unit_cap_mim_m3m4_33/m3_n630_n580# 0.10fF
C146 p1 unit_cap_mim_m3m4_19/m3_n630_n580# -0.29fF
C147 transmission_gate_6/in unit_cap_mim_m3m4_18/c1_n530_n480# -0.03fF
C148 unit_cap_mim_m3m4_29/m3_n630_n580# op 0.42fF
C149 transmission_gate_4/out p1_b -0.01fF
C150 p2 p1 0.01fF
C151 transmission_gate_6/in transmission_gate_9/in 0.09fF
C152 VDD unit_cap_mim_m3m4_19/c1_n530_n480# -0.06fF
C153 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_29/c1_n530_n480# -0.13fF
C154 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C155 VDD unit_cap_mim_m3m4_29/m3_n630_n580# 0.35fF
C156 cm p2_b 0.16fF
C157 transmission_gate_6/in bias_a 0.05fF
C158 transmission_gate_9/in cmc 6.71fF
C159 transmission_gate_7/in unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C160 transmission_gate_7/in unit_cap_mim_m3m4_20/c1_n530_n480# 0.07fF
C161 transmission_gate_8/in unit_cap_mim_m3m4_28/m3_n630_n580# 0.12fF
C162 p1 op 0.10fF
C163 transmission_gate_4/out p2_b 0.03fF
C164 unit_cap_mim_m3m4_24/m3_n630_n580# p2_b -0.55fF
C165 unit_cap_mim_m3m4_17/m3_n630_n580# p2_b -0.46fF
C166 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.10fF
C167 unit_cap_mim_m3m4_16/c1_n530_n480# p2_b -0.07fF
C168 unit_cap_mim_m3m4_18/m3_n630_n580# p1_b -0.41fF
C169 transmission_gate_3/out p1 -0.00fF
C170 VDD p1 0.08fF
C171 transmission_gate_4/out on 3.14fF
C172 unit_cap_mim_m3m4_23/c1_n530_n480# op 0.13fF
C173 unit_cap_mim_m3m4_21/c1_n530_n480# on 0.06fF
C174 unit_cap_mim_m3m4_35/c1_n530_n480# p1 -0.30fF
C175 VDD unit_cap_mim_m3m4_23/m3_n630_n580# 0.33fF
C176 transmission_gate_3/out unit_cap_mim_m3m4_23/m3_n630_n580# 0.61fF
C177 cm unit_cap_mim_m3m4_19/m3_n630_n580# 0.38fF
C178 transmission_gate_6/in cmc 0.92fF
C179 p2 cm 0.21fF
C180 transmission_gate_7/in unit_cap_mim_m3m4_19/c1_n530_n480# 0.03fF
C181 unit_cap_mim_m3m4_31/c1_n530_n480# op 0.05fF
C182 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.17fF
C183 unit_cap_mim_m3m4_16/m3_n630_n580# p2_b -0.37fF
C184 p2 transmission_gate_4/out 0.02fF
C185 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_33/c1_n530_n480# -0.20fF
C186 unit_cap_mim_m3m4_24/m3_n630_n580# p2 -0.47fF
C187 unit_cap_mim_m3m4_21/c1_n530_n480# p2 0.03fF
C188 unit_cap_mim_m3m4_17/m3_n630_n580# p2 -0.56fF
C189 p2 unit_cap_mim_m3m4_16/c1_n530_n480# -0.30fF
C190 unit_cap_mim_m3m4_24/c1_n530_n480# transmission_gate_9/in -0.01fF
C191 unit_cap_mim_m3m4_22/m3_n630_n580# p1 -0.76fF
C192 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580# -0.20fF
C193 unit_cap_mim_m3m4_21/m3_n630_n580# cmc 0.58fF
C194 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.17fF
C195 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_20/c1_n530_n480# -0.20fF
C196 p1 unit_cap_mim_m3m4_35/m3_n630_n580# -0.25fF
C197 unit_cap_mim_m3m4_22/c1_n530_n480# op 0.07fF
C198 transmission_gate_7/in p1 0.02fF
C199 unit_cap_mim_m3m4_24/c1_n530_n480# bias_a -0.22fF
C200 transmission_gate_8/in p1 0.02fF
C201 transmission_gate_4/out op 1.08fF
C202 unit_cap_mim_m3m4_16/m3_n630_n580# p2 -0.29fF
C203 transmission_gate_3/out cm 0.19fF
C204 VDD cm 0.00fF
C205 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C206 transmission_gate_6/in unit_cap_mim_m3m4_28/m3_n630_n580# -1.01fF
C207 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C208 p2_b p1_b 0.01fF
C209 transmission_gate_3/out transmission_gate_4/out 0.37fF
C210 VDD transmission_gate_4/out 0.20fF
C211 unit_cap_mim_m3m4_24/m3_n630_n580# VDD -0.50fF
C212 unit_cap_mim_m3m4_17/m3_n630_n580# VDD -0.16fF
C213 unit_cap_mim_m3m4_17/m3_n630_n580# transmission_gate_3/out 0.62fF
C214 VDD unit_cap_mim_m3m4_16/c1_n530_n480# -0.06fF
C215 on p1_b 0.12fF
C216 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.12fF
C217 transmission_gate_6/in unit_cap_mim_m3m4_27/m3_n630_n580# 0.21fF
C218 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# 0.17fF
C219 p1 unit_cap_mim_m3m4_18/c1_n530_n480# -0.30fF
C220 VDD unit_cap_mim_m3m4_16/m3_n630_n580# -0.43fF
C221 unit_cap_mim_m3m4_34/m3_n630_n580# transmission_gate_8/in 0.56fF
C222 unit_cap_mim_m3m4_19/m3_n630_n580# p1_b -0.65fF
C223 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480# -0.20fF
C224 transmission_gate_7/in cm 0.11fF
C225 transmission_gate_9/in p1 0.01fF
C226 p2 p1_b 0.29fF
C227 transmission_gate_6/in unit_cap_mim_m3m4_29/m3_n630_n580# 0.63fF
C228 cm transmission_gate_8/in 0.03fF
C229 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_30/c1_n530_n480# -0.13fF
C230 unit_cap_mim_m3m4_27/m3_n630_n580# cmc 0.12fF
C231 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C232 transmission_gate_9/in unit_cap_mim_m3m4_23/m3_n630_n580# 0.17fF
C233 unit_cap_mim_m3m4_26/c1_n530_n480# on 0.06fF
C234 on p2_b 0.11fF
C235 VDD unit_cap_mim_m3m4_18/m3_n630_n580# -0.26fF
C236 transmission_gate_7/in transmission_gate_4/out 0.61fF
C237 bias_a p1 0.06fF
C238 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C239 transmission_gate_4/out transmission_gate_8/in 0.26fF
C240 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C241 p1_b op 0.10fF
C242 p2 p2_b 2.48fF
C243 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# -0.49fF
C244 transmission_gate_3/out p1_b 0.08fF
C245 VDD p1_b 0.07fF
C246 p2 on 0.28fF
C247 cm unit_cap_mim_m3m4_18/c1_n530_n480# -0.22fF
C248 unit_cap_mim_m3m4_35/c1_n530_n480# p1_b -0.07fF
C249 cmc p1 0.03fF
C250 unit_cap_mim_m3m4_17/c1_n530_n480# cm -0.22fF
C251 cm transmission_gate_9/in 0.04fF
C252 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C253 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.17fF
C254 unit_cap_mim_m3m4_25/m3_n630_n580# transmission_gate_9/in 0.43fF
C255 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C256 p2_b op 0.17fF
C257 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_17/c1_n530_n480# -0.15fF
C258 transmission_gate_4/out transmission_gate_9/in 3.03fF
C259 cm bias_a 0.91fF
C260 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C261 unit_cap_mim_m3m4_24/m3_n630_n580# transmission_gate_9/in 0.58fF
C262 on op 1.88fF
C263 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.17fF
C264 unit_cap_mim_m3m4_30/m3_n630_n580# p1 -0.67fF
C265 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C266 unit_cap_mim_m3m4_31/m3_n630_n580# transmission_gate_4/out 0.53fF
C267 unit_cap_mim_m3m4_22/m3_n630_n580# p1_b -0.63fF
C268 VDD p2_b 0.27fF
C269 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.10fF
C270 transmission_gate_6/in cm 0.19fF
C271 transmission_gate_4/out bias_a 0.09fF
C272 unit_cap_mim_m3m4_24/m3_n630_n580# bias_a 0.35fF
C273 unit_cap_mim_m3m4_35/m3_n630_n580# p1_b -0.40fF
C274 transmission_gate_3/out on 0.48fF
C275 VDD on 0.45fF
C276 transmission_gate_7/in p1_b 0.03fF
C277 transmission_gate_8/in p1_b 0.02fF
C278 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C279 unit_cap_mim_m3m4_16/m3_n630_n580# transmission_gate_9/in 0.17fF
C280 p2 op 0.04fF
C281 unit_cap_mim_m3m4_28/c1_n530_n480# op 0.17fF
C282 transmission_gate_6/in transmission_gate_4/out 0.46fF
C283 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580# -0.15fF
C284 VDD unit_cap_mim_m3m4_19/m3_n630_n580# -0.52fF
C285 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C286 transmission_gate_3/out p2 0.02fF
C287 VDD p2 0.15fF
C288 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C289 transmission_gate_4/out cmc 0.10fF
C290 unit_cap_mim_m3m4_17/m3_n630_n580# cmc 0.17fF
C291 unit_cap_mim_m3m4_27/c1_n530_n480# op -0.09fF
C292 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C293 transmission_gate_7/in p2_b 0.00fF
C294 transmission_gate_8/in p2_b -0.02fF
C295 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_21/c1_n530_n480# -0.20fF
C296 p1 unit_cap_mim_m3m4_19/c1_n530_n480# -0.30fF
C297 transmission_gate_7/in on 3.18fF
C298 unit_cap_mim_m3m4_18/c1_n530_n480# p1_b -0.07fF
C299 transmission_gate_8/in on 0.83fF
C300 VDD op 0.19fF
C301 transmission_gate_3/out op 0.42fF
C302 transmission_gate_6/in unit_cap_mim_m3m4_18/m3_n630_n580# 0.62fF
C303 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 0.98fF
C304 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.16fF
C305 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.56fF
C306 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.16fF
C307 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C308 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 0.98fF
C309 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C310 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C311 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C312 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.12fF
C313 cmc VSS -12.06fF
C314 transmission_gate_9/in VSS -27.53fF
C315 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.20fF
C316 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C317 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C318 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.55fF
C319 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.56fF
C320 p2 VSS 9.30fF
C321 p2_b VSS 1.84fF
C322 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C323 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.55fF
C324 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C325 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.55fF
C326 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.53fF
C327 transmission_gate_4/out VSS 1.26fF
C328 transmission_gate_3/out VSS -4.23fF
C329 transmission_gate_8/in VSS -0.18fF
C330 bias_a VSS 7.51fF
C331 transmission_gate_6/in VSS 2.86fF
C332 transmission_gate_7/in VSS 2.35fF
C333 cm VSS 0.43fF
C334 p1 VSS 10.10fF
C335 op VSS 11.93fF
C336 p1_b VSS 2.50fF
C337 VDD VSS 16.22fF
C338 on VSS -9.15fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6QKDBA a_n207_n140# a_n1039_n205# a_1275_n205#
+ a_29_n205# a_327_n140# a_n1275_n140# a_n683_n205# a_741_n205# a_n29_n140# a_149_n140#
+ a_n1097_n140# a_1097_n205# a_1395_n140# a_n505_n205# a_n741_n140# a_563_n205# a_861_n140#
+ a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_1217_n140# a_n1395_n205# a_683_n140#
+ a_n919_n140# a_n149_n205# w_n1489_n241# a_1039_n140# a_n385_n140# a_207_n205# a_n1217_n205#
+ a_505_n140# a_n1453_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1395_n140# a_1275_n205# a_1217_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_327_n140# a_207_n205# a_149_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_149_n140# a_29_n205# a_n29_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_861_n140# a_741_n205# a_683_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n207_n140# a_n327_n205# a_n385_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_1217_n140# a_1097_n205# a_1039_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n1275_n140# a_n1395_n205# a_n1453_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n205# a_n919_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1217_n205# a_n1275_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n205# a_505_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n205# a_861_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n29_n140# a_n149_n205# a_n207_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_n563_n140# a_n683_n205# a_n741_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_563_n205# a_n1039_n205# 0.01fF
C1 a_1217_n140# a_1039_n140# 0.13fF
C2 a_n741_n140# a_n1097_n140# 0.06fF
C3 a_n1097_n140# w_n1489_n241# 0.02fF
C4 a_n29_n140# a_683_n140# 0.03fF
C5 a_505_n140# a_n563_n140# 0.02fF
C6 a_n207_n140# a_n919_n140# 0.03fF
C7 a_n505_n205# a_n861_n205# 0.03fF
C8 a_861_n140# a_149_n140# 0.03fF
C9 a_n563_n140# a_n1453_n140# 0.02fF
C10 a_n1275_n140# a_327_n140# 0.01fF
C11 a_n29_n140# a_n741_n140# 0.03fF
C12 a_n385_n140# a_149_n140# 0.04fF
C13 a_n29_n140# w_n1489_n241# 0.02fF
C14 a_n683_n205# a_n861_n205# 0.11fF
C15 a_n327_n205# a_1275_n205# 0.01fF
C16 a_n861_n205# a_n1395_n205# 0.02fF
C17 a_1395_n140# a_1039_n140# 0.06fF
C18 a_n1217_n205# a_n505_n205# 0.01fF
C19 a_741_n205# a_1275_n205# 0.02fF
C20 a_1217_n140# a_149_n140# 0.02fF
C21 a_207_n205# a_1275_n205# 0.01fF
C22 a_29_n205# a_n327_n205# 0.03fF
C23 a_919_n205# w_n1489_n241# 0.19fF
C24 a_n683_n205# a_n1217_n205# 0.02fF
C25 a_861_n140# a_505_n140# 0.06fF
C26 a_n1217_n205# a_n1395_n205# 0.11fF
C27 a_1039_n140# a_683_n140# 0.06fF
C28 a_n505_n205# w_n1489_n241# 0.24fF
C29 a_505_n140# a_n385_n140# 0.02fF
C30 a_741_n205# a_29_n205# 0.01fF
C31 a_n385_n140# a_n1453_n140# 0.02fF
C32 a_29_n205# a_207_n205# 0.11fF
C33 a_n919_n140# a_n563_n140# 0.06fF
C34 a_1039_n140# w_n1489_n241# 0.02fF
C35 a_n683_n205# w_n1489_n241# 0.24fF
C36 a_n29_n140# a_n1097_n140# 0.02fF
C37 a_n861_n205# a_n1039_n205# 0.11fF
C38 a_n1395_n205# w_n1489_n241# 0.31fF
C39 a_1395_n140# a_149_n140# 0.02fF
C40 a_919_n205# a_1097_n205# 0.11fF
C41 a_1217_n140# a_505_n140# 0.03fF
C42 a_n207_n140# a_n1275_n140# 0.02fF
C43 a_n505_n205# a_1097_n205# 0.01fF
C44 a_149_n140# a_683_n140# 0.04fF
C45 a_741_n205# a_n327_n205# 0.01fF
C46 a_n207_n140# a_327_n140# 0.04fF
C47 a_n1217_n205# a_n1039_n205# 0.11fF
C48 a_n327_n205# a_207_n205# 0.02fF
C49 a_n741_n140# a_149_n140# 0.02fF
C50 a_n149_n205# a_1275_n205# 0.01fF
C51 w_n1489_n241# a_149_n140# 0.02fF
C52 a_n385_n140# a_n919_n140# 0.04fF
C53 a_741_n205# a_207_n205# 0.02fF
C54 a_n1039_n205# w_n1489_n241# 0.24fF
C55 a_505_n140# a_1395_n140# 0.02fF
C56 a_385_n205# a_1275_n205# 0.01fF
C57 a_n149_n205# a_29_n205# 0.11fF
C58 a_n29_n140# a_1039_n140# 0.02fF
C59 a_563_n205# a_1275_n205# 0.01fF
C60 a_505_n140# a_683_n140# 0.13fF
C61 a_29_n205# a_385_n205# 0.03fF
C62 a_n1275_n140# a_n563_n140# 0.03fF
C63 a_505_n140# a_n741_n140# 0.02fF
C64 a_n741_n140# a_n1453_n140# 0.03fF
C65 a_505_n140# w_n1489_n241# 0.02fF
C66 a_n505_n205# a_919_n205# 0.01fF
C67 w_n1489_n241# a_n1453_n140# 0.02fF
C68 a_327_n140# a_n563_n140# 0.02fF
C69 a_563_n205# a_29_n205# 0.02fF
C70 a_n1097_n140# a_149_n140# 0.02fF
C71 a_n683_n205# a_919_n205# 0.01fF
C72 a_n149_n205# a_n327_n205# 0.11fF
C73 a_n683_n205# a_n505_n205# 0.11fF
C74 a_n505_n205# a_n1395_n205# 0.01fF
C75 a_n29_n140# a_149_n140# 0.13fF
C76 a_n327_n205# a_385_n205# 0.01fF
C77 a_741_n205# a_n149_n205# 0.01fF
C78 a_n683_n205# a_n1395_n205# 0.01fF
C79 a_n149_n205# a_207_n205# 0.03fF
C80 a_n1275_n140# a_n385_n140# 0.02fF
C81 a_n919_n140# a_683_n140# 0.01fF
C82 a_741_n205# a_385_n205# 0.03fF
C83 a_861_n140# a_327_n140# 0.04fF
C84 a_385_n205# a_207_n205# 0.11fF
C85 a_563_n205# a_n327_n205# 0.01fF
C86 a_505_n140# a_n1097_n140# 0.01fF
C87 a_n1097_n140# a_n1453_n140# 0.06fF
C88 a_n385_n140# a_327_n140# 0.03fF
C89 a_n741_n140# a_n919_n140# 0.13fF
C90 a_n919_n140# w_n1489_n241# 0.02fF
C91 a_563_n205# a_741_n205# 0.11fF
C92 a_563_n205# a_207_n205# 0.03fF
C93 a_505_n140# a_n29_n140# 0.04fF
C94 a_n29_n140# a_n1453_n140# 0.01fF
C95 a_n505_n205# a_n1039_n205# 0.02fF
C96 a_1217_n140# a_327_n140# 0.02fF
C97 a_1039_n140# a_149_n140# 0.02fF
C98 a_n207_n140# a_n563_n140# 0.06fF
C99 a_n683_n205# a_n1039_n205# 0.03fF
C100 a_n1039_n205# a_n1395_n205# 0.03fF
C101 a_29_n205# a_n861_n205# 0.01fF
C102 a_n1097_n140# a_n919_n140# 0.13fF
C103 a_1395_n140# a_327_n140# 0.02fF
C104 a_505_n140# a_1039_n140# 0.04fF
C105 a_n149_n205# a_385_n205# 0.02fF
C106 a_n1217_n205# a_29_n205# 0.01fF
C107 w_n1489_n241# a_1275_n205# 0.24fF
C108 a_861_n140# a_n207_n140# 0.02fF
C109 a_n29_n140# a_n919_n140# 0.02fF
C110 a_n207_n140# a_n385_n140# 0.13fF
C111 a_n327_n205# a_n861_n205# 0.02fF
C112 a_n741_n140# a_n1275_n140# 0.04fF
C113 a_327_n140# a_683_n140# 0.06fF
C114 a_563_n205# a_n149_n205# 0.01fF
C115 a_n1275_n140# w_n1489_n241# 0.02fF
C116 a_29_n205# w_n1489_n241# 0.24fF
C117 a_563_n205# a_385_n205# 0.11fF
C118 a_n741_n140# a_327_n140# 0.02fF
C119 a_741_n205# a_n861_n205# 0.01fF
C120 w_n1489_n241# a_327_n140# 0.02fF
C121 a_n861_n205# a_207_n205# 0.01fF
C122 a_1097_n205# a_1275_n205# 0.11fF
C123 a_1217_n140# a_n207_n140# 0.01fF
C124 a_n1217_n205# a_n327_n205# 0.01fF
C125 a_505_n140# a_149_n140# 0.06fF
C126 a_n1453_n140# a_149_n140# 0.01fF
C127 a_29_n205# a_1097_n205# 0.01fF
C128 a_861_n140# a_n563_n140# 0.01fF
C129 a_n1217_n205# a_207_n205# 0.01fF
C130 a_n327_n205# w_n1489_n241# 0.24fF
C131 a_n385_n140# a_n563_n140# 0.13fF
C132 a_n1275_n140# a_n1097_n140# 0.13fF
C133 a_n207_n140# a_1395_n140# 0.01fF
C134 a_741_n205# w_n1489_n241# 0.20fF
C135 a_207_n205# w_n1489_n241# 0.23fF
C136 a_n1097_n140# a_327_n140# 0.01fF
C137 a_n29_n140# a_n1275_n140# 0.02fF
C138 a_n207_n140# a_683_n140# 0.02fF
C139 a_n327_n205# a_1097_n205# 0.01fF
C140 a_919_n205# a_1275_n205# 0.03fF
C141 a_n29_n140# a_327_n140# 0.06fF
C142 a_n149_n205# a_n861_n205# 0.01fF
C143 a_n919_n140# a_149_n140# 0.02fF
C144 a_n207_n140# a_n741_n140# 0.04fF
C145 a_n207_n140# w_n1489_n241# 0.02fF
C146 a_861_n140# a_n385_n140# 0.02fF
C147 a_741_n205# a_1097_n205# 0.03fF
C148 a_n861_n205# a_385_n205# 0.01fF
C149 a_207_n205# a_1097_n205# 0.01fF
C150 a_29_n205# a_919_n205# 0.01fF
C151 a_29_n205# a_n505_n205# 0.02fF
C152 a_563_n205# a_n861_n205# 0.01fF
C153 a_n149_n205# a_n1217_n205# 0.01fF
C154 a_861_n140# a_1217_n140# 0.06fF
C155 a_n683_n205# a_29_n205# 0.01fF
C156 a_n1217_n205# a_385_n205# 0.01fF
C157 a_1217_n140# a_n385_n140# 0.01fF
C158 a_505_n140# a_n919_n140# 0.01fF
C159 a_29_n205# a_n1395_n205# 0.01fF
C160 a_n919_n140# a_n1453_n140# 0.04fF
C161 a_1039_n140# a_327_n140# 0.03fF
C162 a_n563_n140# a_683_n140# 0.02fF
C163 a_n149_n205# w_n1489_n241# 0.24fF
C164 a_n207_n140# a_n1097_n140# 0.02fF
C165 a_385_n205# w_n1489_n241# 0.22fF
C166 a_n327_n205# a_919_n205# 0.01fF
C167 a_n741_n140# a_n563_n140# 0.13fF
C168 w_n1489_n241# a_n563_n140# 0.02fF
C169 a_n327_n205# a_n505_n205# 0.11fF
C170 a_861_n140# a_1395_n140# 0.04fF
C171 a_741_n205# a_919_n205# 0.11fF
C172 a_n207_n140# a_n29_n140# 0.13fF
C173 a_563_n205# w_n1489_n241# 0.21fF
C174 a_919_n205# a_207_n205# 0.01fF
C175 a_n683_n205# a_n327_n205# 0.03fF
C176 a_741_n205# a_n505_n205# 0.01fF
C177 a_n149_n205# a_1097_n205# 0.01fF
C178 a_n1275_n140# a_149_n140# 0.01fF
C179 a_n327_n205# a_n1395_n205# 0.01fF
C180 a_n505_n205# a_207_n205# 0.01fF
C181 a_29_n205# a_n1039_n205# 0.01fF
C182 a_861_n140# a_683_n140# 0.13fF
C183 a_385_n205# a_1097_n205# 0.01fF
C184 a_n683_n205# a_741_n205# 0.01fF
C185 a_327_n140# a_149_n140# 0.13fF
C186 a_n683_n205# a_207_n205# 0.01fF
C187 a_n385_n140# a_683_n140# 0.02fF
C188 a_861_n140# a_n741_n140# 0.01fF
C189 a_207_n205# a_n1395_n205# 0.01fF
C190 a_1217_n140# a_1395_n140# 0.13fF
C191 a_861_n140# w_n1489_n241# 0.02fF
C192 a_n741_n140# a_n385_n140# 0.06fF
C193 a_563_n205# a_1097_n205# 0.02fF
C194 a_n1097_n140# a_n563_n140# 0.04fF
C195 a_n385_n140# w_n1489_n241# 0.02fF
C196 a_1217_n140# a_683_n140# 0.04fF
C197 a_n207_n140# a_1039_n140# 0.02fF
C198 a_n1275_n140# a_n1453_n140# 0.13fF
C199 a_n29_n140# a_n563_n140# 0.04fF
C200 a_n327_n205# a_n1039_n205# 0.01fF
C201 a_505_n140# a_327_n140# 0.13fF
C202 a_1217_n140# w_n1489_n241# 0.02fF
C203 a_n1217_n205# a_n861_n205# 0.03fF
C204 a_n149_n205# a_919_n205# 0.01fF
C205 a_207_n205# a_n1039_n205# 0.01fF
C206 a_919_n205# a_385_n205# 0.02fF
C207 a_n149_n205# a_n505_n205# 0.03fF
C208 a_n861_n205# w_n1489_n241# 0.24fF
C209 a_1395_n140# a_683_n140# 0.03fF
C210 a_n1097_n140# a_n385_n140# 0.03fF
C211 a_n505_n205# a_385_n205# 0.01fF
C212 a_n683_n205# a_n149_n205# 0.02fF
C213 a_n207_n140# a_149_n140# 0.06fF
C214 a_n149_n205# a_n1395_n205# 0.01fF
C215 a_861_n140# a_n29_n140# 0.02fF
C216 a_563_n205# a_919_n205# 0.03fF
C217 a_1395_n140# w_n1489_n241# 0.02fF
C218 a_n683_n205# a_385_n205# 0.01fF
C219 a_1039_n140# a_n563_n140# 0.01fF
C220 a_n1275_n140# a_n919_n140# 0.06fF
C221 a_n29_n140# a_n385_n140# 0.06fF
C222 a_563_n205# a_n505_n205# 0.01fF
C223 a_n1217_n205# w_n1489_n241# 0.24fF
C224 a_n919_n140# a_327_n140# 0.02fF
C225 a_n741_n140# a_683_n140# 0.01fF
C226 w_n1489_n241# a_683_n140# 0.02fF
C227 a_n683_n205# a_563_n205# 0.01fF
C228 a_n741_n140# w_n1489_n241# 0.02fF
C229 a_1217_n140# a_n29_n140# 0.02fF
C230 a_n207_n140# a_505_n140# 0.03fF
C231 a_n207_n140# a_n1453_n140# 0.02fF
C232 a_n149_n205# a_n1039_n205# 0.01fF
C233 a_861_n140# a_1039_n140# 0.13fF
C234 a_n563_n140# a_149_n140# 0.03fF
C235 a_385_n205# a_n1039_n205# 0.01fF
C236 a_n385_n140# a_1039_n140# 0.01fF
C237 a_1097_n205# w_n1489_n241# 0.18fF
C238 a_29_n205# a_1275_n205# 0.01fF
C239 a_n29_n140# a_1395_n140# 0.01fF
C240 w_n1489_n241# VSUBS 4.31fF
.ends

.subckt ota ip in p1 p1_b p2 p2_b op on i_bias cm VDD VSS
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_0 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_1 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_2 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_3 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_4 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_0 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_1 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_5 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_2 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_BASQVB_0 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias
+ i_bias i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_6 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_3 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_0 m1_n1659_n11581# bias_d VSS bias_d bias_a m1_n947_n12836#
+ m1_n1659_n11581# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# on op bias_d
+ bias_d op op on op bias_d VSS on m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n947_n12836#
+ bias_d bias_d bias_d VSS m1_n1659_n11581# m1_n1659_n11581# on VSS m1_n1659_n11581#
+ on m1_n947_n12836# m1_n947_n12836# bias_d bias_d op bias_d op bias_d m1_n947_n12836#
+ bias_d bias_d op VSS on VSS VSS on op bias_d bias_d m1_n1659_n11581# on on bias_d
+ bias_d bias_d VSS bias_d VSS m1_n947_n12836# m1_n1659_n11581# m1_n2176_n12171# VSS
+ m1_n947_n12836# bias_d bias_d op VSS m1_n947_n12836# bias_d m1_n1659_n11581# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_1 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias
+ bias_c i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_7 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_4 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_1 m1_n947_n12836# bias_d bias_d bias_d op m1_n947_n12836#
+ m1_n2176_n12171# bias_d VSS bias_d VSS bias_d m1_n1659_n11581# on VSS bias_d bias_d
+ on bias_a bias_a bias_a bias_d bias_d bias_a m1_n1659_n11581# VSS bias_d on op VSS
+ VSS bias_d bias_d bias_d m1_n947_n12836# m1_n2176_n12171# bias_a bias_d m1_n947_n12836#
+ bias_a m1_n2176_n12171# m1_n1659_n11581# bias_d bias_d bias_a bias_d op VSS m1_n2176_n12171#
+ bias_d VSS bias_a bias_d VSS op bias_d bias_a on bias_d bias_d m1_n1659_n11581#
+ op on VSS bias_d bias_d on bias_d bias_d m1_n2176_n12171# VSS m1_n1659_n11581# bias_d
+ m1_n947_n12836# bias_d VSS bias_a op m1_n947_n12836# bias_d m1_n2176_n12171# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_2 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias
+ bias_c i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_5 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_2 m1_n947_n12836# bias_d VSS bias_d bias_a m1_n1659_n11581#
+ m1_n947_n12836# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# op on bias_d
+ bias_d on on op on bias_d VSS op m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n1659_n11581#
+ bias_d bias_d bias_d VSS m1_n947_n12836# m1_n947_n12836# op VSS m1_n947_n12836#
+ op m1_n1659_n11581# m1_n1659_n11581# bias_d bias_d on bias_d on bias_d m1_n1659_n11581#
+ bias_d bias_d on VSS op VSS VSS op on bias_d bias_d m1_n947_n12836# op op bias_d
+ bias_d bias_d VSS bias_d VSS m1_n1659_n11581# m1_n947_n12836# m1_n2176_n12171# VSS
+ m1_n1659_n11581# bias_d bias_d on VSS m1_n1659_n11581# bias_d m1_n947_n12836# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_3 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias
+ i_bias i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_10 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_11 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_6 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_12 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_7 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_7P4E2J_0 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_KEEN2X_10 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS cmc cmc bias_a VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS cmc bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_13 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_8 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_KEEN2X_11 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS bias_a bias_a cmc VSS m1_n5574_n13620# cmc VSS bias_a bias_a
+ cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS bias_a cmc VSS VSS
+ m1_n5574_n13620# m1_n5574_n13620# bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc
+ VSS VSS bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620#
+ bias_a bias_a cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# bias_a cmc
+ cmc VSS VSS m1_n5574_n13620# bias_a cmc bias_a m1_n5574_n13620# m1_n5574_n13620#
+ VSS cmc bias_a VSS m1_n5574_n13620# bias_a cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_7P4E2J_1 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d bias_a m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_a m1_6690_n8907# bias_a VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_9 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_14 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_7P4E2J_2 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_a
+ m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_7P4E2J_3 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d
+ m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_15 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_KEEN2X_12 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS bias_a bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# bias_a VSS bias_a bias_a VSS
+ VSS m1_n5574_n13620# m1_n5574_n13620# cmc m1_n5574_n13620# VSS cmc bias_a VSS bias_a
+ VSS VSS cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620#
+ bias_a bias_a cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc bias_a
+ bias_a VSS VSS m1_n5574_n13620# cmc cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS
+ cmc bias_a VSS m1_n5574_n13620# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_VJ4JGY_0 cm cm cm cm cm cm cm m1_11534_n9706# m1_11242_n9716#
+ cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# cm cm cm cm VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_1 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490#
+ m1_11534_n9706# m1_11242_n9716# cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711#
+ m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_2 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490#
+ m1_11534_n11258# m1_11244_n11260# cm cm cm cm m1_12410_n11263# m1_12118_n11263#
+ cm m1_11826_n11260# m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_3 cm cm cm cm VSS cm VSS m1_11534_n11258# m1_11244_n11260#
+ cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260# VSS VSS cm VSS
+ VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__pfet_01v8_E4DCBA_0 VDD bias_c m1_6690_n8907# op bias_c bias_c m1_1038_n2886#
+ bias_b bias_c VDD m1_n208_n2883# bias_c VDD on bias_c VDD m1_2463_n5585# VDD VDD
+ m1_2462_n3318# m1_2462_n3318# op m1_2463_n5585# m1_2462_n3318# VDD VDD VDD bias_b
+ bias_c m1_1038_n2886# bias_c m1_6690_n8907# VDD bias_c VDD VDD m1_2463_n5585# on
+ VDD bias_c m1_2462_n3318# m1_n208_n2883# bias_c bias_c VDD VDD m1_2463_n5585# VDD
+ VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_2 on VDD op on VDD bias_c m1_n208_n2883# on bias_c
+ bias_c VDD VDD m1_n208_n2883# op bias_c bias_c m1_1038_n2886# bias_c VDD m1_n208_n2883#
+ m1_n208_n2883# m1_n6302_n3889# m1_1038_n2886# m1_n208_n2883# m1_n6302_n3889# bias_c
+ bias_c on bias_c VDD bias_c op bias_c bias_c cm bias_c m1_1038_n2886# cm m1_1038_n2886#
+ VDD m1_n208_n2883# m1_1038_n2886# bias_c bias_c op bias_c m1_1038_n2886# bias_c
+ VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_1 op VDD on op VDD bias_c m1_1038_n2886# op bias_c
+ bias_c VDD VDD m1_1038_n2886# on bias_c bias_c m1_n208_n2883# bias_c VDD m1_1038_n2886#
+ m1_1038_n2886# m1_n6302_n3889# m1_n208_n2883# m1_1038_n2886# m1_n6302_n3889# bias_c
+ bias_c op bias_c VDD bias_c on bias_c bias_c cm bias_c m1_n208_n2883# cm m1_n208_n2883#
+ VDD m1_1038_n2886# m1_n208_n2883# bias_c bias_c on bias_c m1_n208_n2883# bias_c
+ VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_3 VDD bias_c bias_b on bias_c bias_c m1_n208_n2883#
+ m1_6690_n8907# bias_c VDD m1_1038_n2886# bias_c VDD op bias_c VDD m1_2462_n3318#
+ VDD VDD m1_2463_n5585# m1_2463_n5585# on m1_2462_n3318# m1_2463_n5585# VDD VDD VDD
+ m1_6690_n8907# bias_c m1_n208_n2883# bias_c bias_b VDD bias_c VDD VDD m1_2462_n3318#
+ op VDD bias_c m1_2463_n5585# m1_1038_n2886# bias_c bias_c VDD VDD m1_2462_n3318#
+ VDD VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsc_cmfb_0 cmc sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580#
+ on sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_8/in
+ sc_cmfb_0/transmission_gate_4/out bias_a p2_b p1 cm sc_cmfb_0/transmission_gate_9/in
+ p2 VDD sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_7/in op VSS
+ p1_b sc_cmfb
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_0 m1_n208_n2883# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_1038_n2886# VDD VDD VDD bias_b VDD bias_b m1_1038_n2886# bias_b bias_b
+ m1_1038_n2886# bias_b VDD VDD VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b VDD m1_n208_n2883#
+ VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_4 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS cmc cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS cmc cmc VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# bias_a m1_n5574_n13620# VSS bias_a cmc VSS cmc VSS VSS bias_a bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ bias_a bias_a m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_1 m1_2463_n5585# bias_b m1_2462_n3318# bias_b
+ VDD m1_2463_n5585# bias_b bias_b VDD m1_2462_n3318# VDD bias_b m1_2462_n3318# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2462_n3318# m1_2463_n5585#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2463_n5585#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_5 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS VSS bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS VSS bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS VSS VSS cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS m1_n5574_n13620# bias_a
+ bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_3 m1_2462_n3318# bias_b m1_2463_n5585# bias_b
+ VDD m1_2462_n3318# bias_b bias_b VDD m1_2463_n5585# VDD bias_b m1_2463_n5585# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2463_n5585# m1_2462_n3318#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2462_n3318#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_2 m1_n6302_n3889# bias_b m1_n6302_n3889# bias_b
+ VDD m1_n6302_n3889# bias_b bias_b VDD m1_n6302_n3889# VDD bias_b m1_n6302_n3889#
+ bias_b VDD bias_b m1_n208_n2883# bias_b bias_b m1_1038_n2886# bias_b m1_n6302_n3889#
+ m1_n6302_n3889# VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b bias_b m1_1038_n2886#
+ m1_n6302_n3889# bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_6 VSS VSS VSS VSS bias_a bias_a m1_n947_n12836# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n1659_n11581# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n947_n12836# bias_a m1_n1659_n11581# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n1659_n11581# m1_n947_n12836# bias_a bias_a bias_a
+ m1_n1659_n11581# m1_n2176_n12171# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_4 m1_1038_n2886# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_n208_n2883# VDD VDD VDD bias_b VDD bias_b m1_n208_n2883# bias_b bias_b
+ m1_n208_n2883# bias_b VDD VDD VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b VDD m1_1038_n2886#
+ VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_7 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n947_n12836# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n1659_n11581# m1_n2176_n12171# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n2176_n12171# m1_n1659_n11581# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_KEEN2X_9 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS VSS cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS VSS cmc VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ bias_a bias_a m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a VSS m1_n5574_n13620#
+ cmc cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_KEEN2X_8 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n947_n12836# m1_n947_n12836# bias_a m1_n1659_n11581# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n1659_n11581# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n1659_n11581# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n1659_n11581# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n947_n12836# m1_n2176_n12171# m1_n947_n12836# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
C0 bias_b m1_n208_n2883# 9.15fF
C1 m1_11534_n9706# m1_12410_n9718# 0.02fF
C2 m1_2462_n3318# m1_2463_n5585# 4.55fF
C3 m1_2462_n3318# bias_a 0.11fF
C4 cm m1_11534_n9706# 0.65fF
C5 cm m1_n208_n2883# 0.17fF
C6 bias_a cmc 12.13fF
C7 bias_a m1_n1659_n11581# 20.90fF
C8 bias_b m1_2463_n5585# 6.62fF
C9 m1_11940_n10482# m1_12232_n10488# 0.07fF
C10 p2_b cmc 0.01fF
C11 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# p1 -0.00fF
C12 m1_11242_n9716# m1_12410_n9718# 0.02fF
C13 m1_1038_n2886# i_bias 0.27fF
C14 m1_n6302_n3889# bias_c 3.58fF
C15 m1_2463_n5585# cm 0.52fF
C16 cm bias_a 0.62fF
C17 m1_11242_n9716# cm 0.68fF
C18 m1_11534_n11258# m1_11534_n9706# 0.01fF
C19 m1_11825_n9711# m1_12410_n9718# 0.03fF
C20 cm m1_11940_n10482# 0.59fF
C21 cm sc_cmfb_0/transmission_gate_8/in 0.04fF
C22 in i_bias 0.29fF
C23 m1_6690_n8907# sc_cmfb_0/transmission_gate_4/out 0.01fF
C24 m1_n2176_n12171# m1_6690_n8907# 0.00fF
C25 cm m1_11825_n9711# 0.65fF
C26 m1_12118_n9704# m1_12410_n9718# 0.07fF
C27 m1_n2176_n12171# m1_n947_n12836# 10.60fF
C28 m1_1038_n2886# on 3.37fF
C29 cm m1_12118_n9704# 0.64fF
C30 m1_n208_n2883# i_bias 0.24fF
C31 p1 op 0.00fF
C32 bias_a p1_b 0.01fF
C33 m1_2462_n3318# m1_6690_n8907# 2.72fF
C34 m1_6690_n8907# cmc 0.46fF
C35 m1_n947_n12836# cmc 0.37fF
C36 m1_n208_n2883# on 0.40fF
C37 m1_n1659_n11581# m1_n947_n12836# 9.35fF
C38 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# sc_cmfb_0/transmission_gate_7/in 0.02fF
C39 bias_b m1_6690_n8907# 0.39fF
C40 m1_1038_n2886# m1_n5574_n13620# 2.47fF
C41 bias_d bias_a 8.20fF
C42 m1_2463_n5585# on 0.09fF
C43 cm m1_6690_n8907# 4.14fF
C44 bias_a on 4.51fF
C45 m1_n2176_n12171# cmc 1.14fF
C46 m1_n2176_n12171# m1_n1659_n11581# 10.31fF
C47 m1_12410_n11263# m1_11244_n11260# 0.02fF
C48 m1_11826_n11260# m1_11825_n9711# 0.01fF
C49 sc_cmfb_0/transmission_gate_9/in on 0.00fF
C50 m1_1038_n2886# VDD 15.44fF
C51 m1_n5574_n13620# in 2.07fF
C52 cm m1_11244_n11260# 0.55fF
C53 m1_n208_n2883# m1_n5574_n13620# 2.51fF
C54 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# p1 0.00fF
C55 m1_12410_n11263# m1_12410_n9718# 0.01fF
C56 bias_b m1_2462_n3318# 3.43fF
C57 m1_n1659_n11581# cmc 0.44fF
C58 cm m1_12232_n10488# 0.57fF
C59 cm m1_12410_n11263# 0.58fF
C60 m1_n5574_n13620# bias_a 21.14fF
C61 ip m1_1038_n2886# 1.69fF
C62 m1_2462_n3318# cm 1.44fF
C63 m1_1038_n2886# op 0.78fF
C64 cm cmc 0.85fF
C65 m1_n208_n2883# VDD 15.21fF
C66 m1_11534_n11258# m1_11244_n11260# 0.07fF
C67 bias_b cm 0.36fF
C68 cm m1_12410_n9718# 0.64fF
C69 m1_2463_n5585# VDD 7.71fF
C70 m1_11534_n11258# m1_12410_n11263# 0.02fF
C71 bias_d m1_6690_n8907# 35.88fF
C72 bias_d m1_n947_n12836# 16.58fF
C73 bias_a VDD 0.11fF
C74 ip in 3.13fF
C75 m1_6690_n8907# on 1.68fF
C76 m1_n947_n12836# on 8.70fF
C77 m1_11063_n10490# m1_11356_n10481# 0.07fF
C78 p2_b VDD 0.00fF
C79 m1_1038_n2886# bias_c 7.06fF
C80 ip m1_n208_n2883# 1.08fF
C81 m1_1038_n2886# m1_n6302_n3889# 2.81fF
C82 m1_n208_n2883# op 3.85fF
C83 bias_d m1_n2176_n12171# 8.59fF
C84 p2 p2_b 0.00fF
C85 cm m1_11534_n11258# 0.58fF
C86 m1_n2176_n12171# on 8.63fF
C87 m1_11826_n11260# m1_11244_n11260# 0.03fF
C88 cmc p1_b 0.04fF
C89 m1_2463_n5585# op 0.25fF
C90 bias_a op 2.42fF
C91 in bias_c 0.44fF
C92 m1_11826_n11260# m1_12410_n11263# 0.03fF
C93 m1_11063_n10490# m1_11648_n10486# 0.03fF
C94 cm p1_b 0.09fF
C95 m1_n208_n2883# bias_c 8.21fF
C96 m1_6690_n8907# m1_n5574_n13620# 0.08fF
C97 m1_n5574_n13620# m1_n947_n12836# 0.12fF
C98 m1_n208_n2883# m1_n6302_n3889# 3.54fF
C99 bias_d cmc 0.03fF
C100 m1_2462_n3318# on 0.27fF
C101 bias_d m1_n1659_n11581# 12.63fF
C102 m1_12118_n11263# m1_12118_n9704# 0.01fF
C103 cmc on 0.96fF
C104 m1_n1659_n11581# on 1.52fF
C105 m1_2463_n5585# bias_c 2.57fF
C106 cm m1_11826_n11260# 0.58fF
C107 bias_b on 0.07fF
C108 m1_2463_n5585# m1_n6302_n3889# 0.56fF
C109 bias_a bias_c 0.00fF
C110 bias_d cm 0.08fF
C111 m1_n2176_n12171# m1_n5574_n13620# 0.57fF
C112 m1_6690_n8907# VDD 3.64fF
C113 cm on 1.01fF
C114 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_4/out 0.00fF
C115 m1_11356_n10481# m1_11648_n10486# 0.07fF
C116 m1_11534_n11258# m1_11826_n11260# 0.07fF
C117 sc_cmfb_0/transmission_gate_4/out VDD 0.01fF
C118 m1_n5574_n13620# cmc 54.64fF
C119 m1_n5574_n13620# m1_n1659_n11581# 0.14fF
C120 m1_6690_n8907# op 2.49fF
C121 m1_n947_n12836# op 1.19fF
C122 bias_b m1_n5574_n13620# 0.11fF
C123 cm m1_n5574_n13620# 0.02fF
C124 m1_2462_n3318# VDD 7.06fF
C125 m1_n2176_n12171# op 1.95fF
C126 cmc VDD 0.08fF
C127 m1_12118_n11263# m1_11244_n11260# 0.02fF
C128 bias_b VDD 41.27fF
C129 m1_11063_n10490# m1_11940_n10482# 0.02fF
C130 m1_6690_n8907# bias_c 1.61fF
C131 p2 cmc 0.00fF
C132 bias_a p1 0.04fF
C133 m1_12118_n11263# m1_12410_n11263# 0.07fF
C134 cm VDD 3.70fF
C135 bias_d on 13.96fF
C136 m1_2462_n3318# op 0.28fF
C137 m1_n2176_n12171# bias_c 0.02fF
C138 cmc op 1.20fF
C139 m1_n1659_n11581# op 8.09fF
C140 bias_b ip 0.07fF
C141 bias_b op 0.14fF
C142 cm m1_12118_n11263# 0.57fF
C143 m1_n5574_n13620# i_bias 0.12fF
C144 m1_11356_n10481# m1_11940_n10482# 0.03fF
C145 cm op 0.76fF
C146 m1_2462_n3318# bias_c 4.04fF
C147 VDD p1_b -0.01fF
C148 m1_2462_n3318# m1_n6302_n3889# 0.57fF
C149 m1_11534_n11258# m1_12118_n11263# 0.03fF
C150 bias_c cmc 0.07fF
C151 m1_n5574_n13620# on 0.06fF
C152 m1_1038_n2886# in 1.59fF
C153 bias_b bias_c 25.24fF
C154 bias_b m1_n6302_n3889# 2.49fF
C155 cm bias_c 3.39fF
C156 m1_1038_n2886# m1_n208_n2883# 17.20fF
C157 cm m1_n6302_n3889# 2.61fF
C158 m1_11648_n10486# m1_11940_n10482# 0.07fF
C159 on VDD 5.69fF
C160 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# p1 0.00fF
C161 ip i_bias 0.17fF
C162 m1_2463_n5585# m1_1038_n2886# 3.88fF
C163 m1_1038_n2886# bias_a 0.07fF
C164 m1_11826_n11260# m1_12118_n11263# 0.07fF
C165 p1 sc_cmfb_0/transmission_gate_4/out -0.00fF
C166 m1_n208_n2883# in 3.19fF
C167 cm sc_cmfb_0/transmission_gate_7/in 0.04fF
C168 m1_11063_n10490# m1_12232_n10488# 0.02fF
C169 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# cm 0.01fF
C170 bias_d op 12.45fF
C171 sc_cmfb_0/transmission_gate_3/out op 0.00fF
C172 op on 7.65fF
C173 i_bias bias_c 12.15fF
C174 m1_2463_n5585# m1_n208_n2883# 3.39fF
C175 m1_n208_n2883# bias_a 0.04fF
C176 m1_n5574_n13620# VDD 0.03fF
C177 m1_11242_n9716# m1_11534_n9706# 0.07fF
C178 cm m1_11063_n10490# 0.61fF
C179 cmc p1 0.00fF
C180 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VDD 0.02fF
C181 m1_11356_n10481# m1_12232_n10488# 0.02fF
C182 bias_c on 4.92fF
C183 m1_11534_n9706# m1_11825_n9711# 0.07fF
C184 cm p1 0.17fF
C185 m1_n6302_n3889# on 0.08fF
C186 m1_11534_n9706# m1_12118_n9704# 0.03fF
C187 bias_a sc_cmfb_0/transmission_gate_8/in 0.02fF
C188 ip m1_n5574_n13620# 1.03fF
C189 m1_n5574_n13620# op 0.17fF
C190 m1_1038_n2886# m1_6690_n8907# 0.28fF
C191 m1_11242_n9716# m1_11825_n9711# 0.03fF
C192 cm m1_11356_n10481# 0.58fF
C193 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# op 0.00fF
C194 m1_11242_n9716# m1_12118_n9704# 0.02fF
C195 m1_n2176_n12171# m1_1038_n2886# 0.11fF
C196 m1_11648_n10486# m1_12232_n10488# 0.03fF
C197 op VDD 5.61fF
C198 m1_n5574_n13620# bias_c 0.50fF
C199 p1 p1_b -0.00fF
C200 m1_11825_n9711# m1_12118_n9704# 0.07fF
C201 m1_n208_n2883# m1_6690_n8907# 0.10fF
C202 cm m1_11648_n10486# 0.59fF
C203 m1_2462_n3318# m1_1038_n2886# 4.36fF
C204 m1_2463_n5585# m1_6690_n8907# 0.36fF
C205 bias_c VDD 10.56fF
C206 m1_6690_n8907# bias_a 2.54fF
C207 bias_a m1_n947_n12836# 21.86fF
C208 m1_1038_n2886# cmc 0.17fF
C209 m1_n6302_n3889# VDD 3.85fF
C210 m1_n2176_n12171# m1_n208_n2883# 0.09fF
C211 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# bias_a 0.05fF
C212 bias_b m1_1038_n2886# 10.79fF
C213 p1 on 0.01fF
C214 m1_1038_n2886# cm 1.34fF
C215 m1_n2176_n12171# bias_a 23.78fF
C216 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/transmission_gate_8/in 0.08fF
C217 in cmc 0.04fF
C218 bias_b in 0.09fF
C219 ip bias_c 0.11fF
C220 m1_2462_n3318# m1_n208_n2883# 3.03fF
C221 m1_11242_n9716# m1_11244_n11260# 0.01fF
C222 bias_c op 5.30fF
C223 m1_n6302_n3889# op 0.17fF
C224 m1_n208_n2883# cmc 0.14fF
C225 m1_1038_n2886# VSS -48.90fF
C226 m1_n208_n2883# VSS -43.69fF
C227 m1_n6302_n3889# VSS 10.46fF
C228 m1_2463_n5585# VSS 0.31fF
C229 cmc VSS 34.44fF
C230 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C231 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C232 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C233 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C234 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C235 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C236 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C237 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C238 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C239 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.37fF
C240 sc_cmfb_0/transmission_gate_9/in VSS -27.59fF
C241 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C242 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C243 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C244 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C245 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C246 p2 VSS 9.74fF
C247 p2_b VSS 3.15fF
C248 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C249 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C250 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C251 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C252 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.35fF
C253 sc_cmfb_0/transmission_gate_4/out VSS 1.19fF
C254 sc_cmfb_0/transmission_gate_3/out VSS -4.31fF
C255 sc_cmfb_0/transmission_gate_8/in VSS -0.19fF
C256 sc_cmfb_0/transmission_gate_6/in VSS 2.79fF
C257 sc_cmfb_0/transmission_gate_7/in VSS 2.28fF
C258 cm VSS -12.35fF
C259 p1 VSS 10.06fF
C260 op VSS -11.29fF
C261 p1_b VSS 1.49fF
C262 VDD VSS 364.32fF
C263 on VSS -76.04fF
C264 m1_2462_n3318# VSS -13.18fF
C265 m1_12410_n11263# VSS 0.18fF
C266 m1_12118_n11263# VSS 0.31fF
C267 m1_11826_n11260# VSS 0.32fF
C268 m1_11534_n11258# VSS 0.24fF
C269 m1_11244_n11260# VSS 0.25fF
C270 m1_12232_n10488# VSS 0.24fF
C271 m1_11940_n10482# VSS 0.35fF
C272 m1_11648_n10486# VSS 0.25fF
C273 m1_11356_n10481# VSS 0.27fF
C274 m1_11063_n10490# VSS 0.27fF
C275 m1_12410_n9718# VSS 0.17fF
C276 m1_12118_n9704# VSS 0.28fF
C277 m1_11825_n9711# VSS 0.29fF
C278 m1_11534_n9706# VSS 0.23fF
C279 m1_11242_n9716# VSS 0.24fF
C280 bias_a VSS -228.03fF
C281 m1_n5574_n13620# VSS 239.91fF
C282 m1_6690_n8907# VSS -73.13fF
C283 bias_c VSS 46.85fF
C284 i_bias VSS 34.76fF
C285 m1_n1659_n11581# VSS 8.91fF
C286 m1_n947_n12836# VSS 15.61fF
C287 in VSS 2.41fF
C288 m1_n2176_n12171# VSS 17.30fF
C289 bias_d VSS 120.62fF
C290 ip VSS 2.33fF
C291 bias_b VSS 13.05fF
.ends

