magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< pwell >>
rect 5643 23633 5707 23697
rect 5284 9365 5337 9418
<< viali >>
rect -20380 33278 -20346 33564
rect -20380 32634 -20346 33008
<< metal1 >>
rect -13123 71958 -12995 78096
rect -13893 52998 -13765 66326
rect -12552 53600 -12424 66338
rect -12563 53536 -12553 53600
rect -12425 53536 -12415 53600
rect -7560 53536 -7550 53600
rect -7486 53536 -7476 53600
rect -6999 53536 -6989 53600
rect -6861 53536 -6851 53600
rect -12552 53520 -12424 53536
rect -13893 52992 -9120 52998
rect -13893 52928 -9398 52992
rect -9270 52928 -9120 52992
rect -13893 52923 -9120 52928
rect -9408 49923 -9398 49987
rect -9270 49923 -8690 49987
rect -7544 49921 -6989 49985
rect -6861 49921 -6851 49985
rect 93 45365 157 45366
rect -569 45313 157 45365
rect -6989 39805 -6861 39806
rect -9408 39741 -9398 39805
rect -9270 39741 -9260 39805
rect -6999 39741 -6989 39805
rect -6861 39741 -6851 39805
rect -14182 33901 -14172 33965
rect -14108 33901 -14098 33965
rect -20386 33564 -20340 33576
rect -20386 33439 -20380 33564
rect -20416 33405 -20380 33439
rect -20386 33278 -20380 33405
rect -20346 33439 -20340 33564
rect -19731 33558 -19667 33573
rect -20134 33524 -19667 33558
rect -20346 33405 -20295 33439
rect -20346 33278 -20340 33405
rect -19731 33318 -19667 33524
rect -14172 33373 -14108 33901
rect -20138 33284 -19667 33318
rect -20386 33266 -20340 33278
rect -20386 33008 -20340 33020
rect -20386 32839 -20380 33008
rect -20416 32805 -20380 32839
rect -20386 32634 -20380 32805
rect -20346 32839 -20340 33008
rect -19731 33002 -19667 33284
rect -14157 33020 -14123 33373
rect -20138 32968 -19667 33002
rect -20346 32805 -20288 32839
rect -20346 32634 -20340 32805
rect -19731 32688 -19667 32968
rect -19744 32674 -19353 32688
rect -20138 32640 -19353 32674
rect -20386 32622 -20340 32634
rect -19744 32624 -19353 32640
rect -19289 32674 -17888 32688
rect -19289 32640 -17603 32674
rect -19289 32624 -17888 32640
rect -18532 31791 -18522 31855
rect -18458 31840 -17895 31855
rect -18458 31806 -17529 31840
rect -18458 31791 -17895 31806
rect -14225 31099 -14191 31504
rect -14240 30534 -14176 31099
rect -14250 30470 -14240 30534
rect -14176 30470 -14166 30534
rect -9398 29481 -9270 39741
rect -6989 34999 -6861 39741
rect 93 37446 157 45313
rect 5361 37448 5425 40438
rect 83 37382 93 37446
rect 157 37382 167 37446
rect 1220 37382 1230 37446
rect 1294 37382 1304 37446
rect 2439 37384 2626 37448
rect 2690 37384 2700 37448
rect 5351 37384 5361 37448
rect 5425 37384 5435 37448
rect 93 36531 157 37382
rect 5361 37035 5425 37384
rect 5351 36971 5361 37035
rect 5425 36971 5435 37035
rect 83 36467 93 36531
rect 157 36467 167 36531
rect 3417 36467 3427 36531
rect 3491 36467 3501 36531
rect 93 35696 157 36467
rect 2324 36023 2334 36087
rect 2398 36023 2408 36087
rect 2334 35696 2398 36023
rect 83 35632 93 35696
rect 157 35632 167 35696
rect 873 35632 883 35696
rect 947 35632 957 35696
rect 2240 35632 2398 35696
rect 93 35630 157 35632
rect 3427 35350 3491 36467
rect 6701 36087 6765 40449
rect 7082 39092 7200 43012
rect 7072 38974 7082 39092
rect 7200 38974 7210 39092
rect 11926 38974 11936 39092
rect 12054 38974 17164 39092
rect 7420 36971 7430 37035
rect 7494 36971 7504 37035
rect 5419 36023 5429 36087
rect 5493 36023 5503 36087
rect 6691 36023 6701 36087
rect 6765 36023 6775 36087
rect 5429 35345 5493 36023
rect 7430 35332 7494 36971
rect 9418 36467 9428 36531
rect 9492 36467 9502 36531
rect 9428 35340 9492 36467
rect -6999 34935 -6989 34999
rect -6925 34935 -6861 34999
rect -6989 31811 -6861 34935
rect 5420 34356 5430 34420
rect 5494 34356 5504 34420
rect 7418 34354 7428 34418
rect 7492 34354 7502 34418
rect 3866 34180 4878 34244
rect 7854 34181 8873 34245
rect -6999 31747 -6989 31811
rect -6861 31747 -6851 31811
rect -6989 31712 -6861 31747
rect 4354 30432 4418 34180
rect 8328 30437 8392 34181
rect 4344 30368 4354 30432
rect 4418 30368 4428 30432
rect 8318 30373 8328 30437
rect 8392 30373 8402 30437
rect -9398 29417 -9334 29481
rect -9270 29417 -9260 29481
rect -9398 29195 -9270 29417
rect -9407 29131 -9397 29195
rect -9269 29131 -9259 29195
rect -9398 29091 -9270 29131
rect 1941 28784 1951 28848
rect 2079 28784 2089 28848
rect -18326 27575 -18262 27600
rect -18336 27511 -18326 27575
rect -18262 27511 -18252 27575
rect -17635 27568 -17507 27644
rect 1951 27634 2079 28784
rect -12206 27598 2079 27634
rect -12206 27579 -6086 27598
rect -17635 27516 -17334 27568
rect -14546 27519 -14536 27571
rect -14484 27519 -13619 27571
rect -12491 27534 -6086 27579
rect -5958 27534 2079 27598
rect -12491 27515 2079 27534
rect -18326 27098 -18262 27511
rect -12206 27506 2079 27515
rect 3368 28595 3496 28627
rect 3368 28531 3399 28595
rect 3463 28531 3496 28595
rect -18336 27034 -18326 27098
rect -18262 27034 -18252 27098
rect -15239 27082 -14536 27083
rect -18891 26696 -18881 26760
rect -18817 26696 -18807 26760
rect -18881 25977 -18817 26696
rect -18892 25913 -18882 25977
rect -18818 25913 -18808 25977
rect -35142 24984 -27540 25112
rect -27412 24984 -24312 25112
rect -22964 24984 -22131 25112
rect -22259 21702 -22131 24984
rect -18881 24456 -18817 25913
rect -18891 24392 -18881 24456
rect -18817 24392 -18807 24456
rect -18326 24117 -18262 27034
rect -15242 27031 -14536 27082
rect -14484 27031 -14474 27083
rect -17266 26696 -17256 26760
rect -17192 26696 -17182 26760
rect -17635 26363 -17334 26415
rect -17635 26287 -17507 26363
rect -14546 25915 -14536 25967
rect -14484 25915 -13624 25967
rect -12478 25914 -10016 25978
rect -9888 25914 -9878 25978
rect 1952 25820 2080 25825
rect 1942 25756 1952 25820
rect 2080 25756 2090 25820
rect -17635 24926 -17507 25002
rect -17635 24874 -17339 24926
rect -15202 24389 -14538 24441
rect -14486 24389 -14480 24441
rect 1952 24408 2080 25756
rect -14538 24369 -14480 24389
rect -12198 24376 2080 24408
rect -12469 24374 2080 24376
rect -14538 24317 -13620 24369
rect -12469 24312 -3501 24374
rect -12198 24310 -3501 24312
rect -3373 24310 2080 24374
rect -12198 24280 2080 24310
rect -18336 24053 -18326 24117
rect -18262 24053 -18252 24117
rect -17265 24053 -17255 24117
rect -17191 24053 -17181 24117
rect -17635 23721 -17338 23773
rect -17635 23645 -17507 23721
rect 3368 23701 3496 28531
rect 9366 28592 9494 28632
rect 9366 28528 9399 28592
rect 9463 28528 9494 28592
rect 9366 23701 9494 28528
rect 3368 23637 3399 23701
rect 3463 23637 3496 23701
rect -14548 22719 -14538 22771
rect -14486 22719 -13614 22771
rect -12465 22712 -11601 22776
rect -11473 22712 -11463 22776
rect 3368 22535 3496 23637
rect 5633 23633 5643 23697
rect 5707 23633 5717 23697
rect 7007 23637 7017 23701
rect 7081 23637 7091 23701
rect 9366 23637 9399 23701
rect 9463 23637 9494 23701
rect 9366 22535 9494 23637
rect 13272 23295 27530 23423
rect -22259 21671 -5931 21702
rect -22259 21607 -6086 21671
rect -5958 21607 -5931 21671
rect -22259 21574 -5931 21607
rect 9394 21228 9458 21231
rect 3395 21221 3459 21226
rect -22293 20809 -3339 20842
rect -22293 20745 -3501 20809
rect -3373 20745 -3339 20809
rect -22293 20714 -3339 20745
rect -35142 17454 -25679 17582
rect -25551 17454 -24304 17582
rect -22293 17579 -22165 20714
rect -454 19981 -444 20109
rect -380 19981 -370 20109
rect -444 18993 -380 19981
rect 1674 19282 1684 19410
rect 1748 19282 1812 19410
rect -22986 17451 -22165 17579
rect -445 17221 -381 17690
rect 1684 17221 1812 19282
rect 3361 19346 3489 21221
rect 9363 20109 9491 21228
rect 5384 19981 5394 20109
rect 5458 19981 5468 20109
rect 9363 19981 9394 20109
rect 9458 19981 9491 20109
rect 3361 19282 3395 19346
rect 3459 19282 3489 19346
rect 3361 19072 3489 19282
rect 5394 19098 5458 19981
rect 7384 19282 7394 19410
rect 7458 19282 7468 19410
rect 7394 19103 7458 19282
rect 9363 19074 9491 19981
rect 13272 19716 13347 23295
rect 33170 22549 41297 22677
rect 13877 21996 13887 22124
rect 13951 21996 27510 22124
rect 13877 17983 13887 18047
rect 13951 17983 13961 18047
rect -455 17093 -445 17221
rect -381 17093 -371 17221
rect 1674 17093 1684 17221
rect 1748 17093 1812 17221
rect 3393 16866 3457 17769
rect 5393 16866 5457 17768
rect 7393 17359 7457 17775
rect 9396 17359 9460 17774
rect 7383 17231 7393 17359
rect 7457 17231 7467 17359
rect 9386 17231 9396 17359
rect 9460 17231 9470 17359
rect 13875 17231 13885 17359
rect 13949 17231 13959 17359
rect 3383 16738 3393 16866
rect 3457 16738 3467 16866
rect 5383 16738 5393 16866
rect 5457 16738 5467 16866
rect 13267 16738 13277 16866
rect 13341 16738 13351 16866
rect -3926 16288 -3862 16297
rect -3936 16224 -3926 16288
rect -3862 16224 -3852 16288
rect -3927 15083 -3914 15135
rect -3862 15083 -2971 15135
rect -1824 15084 -678 15136
rect -626 15084 -616 15136
rect -27550 13974 -27540 14102
rect -27412 13974 -24548 14102
rect -23154 14073 -15769 14105
rect -10703 14077 -10693 14141
rect -10629 14077 -5457 14141
rect -3963 14087 -3914 14139
rect -3862 14087 -3852 14139
rect -23385 14009 -15852 14073
rect -15788 14009 -15769 14073
rect -23154 13977 -15769 14009
rect -5633 12892 -5569 14077
rect -5633 12828 -4962 12892
rect -5026 12173 -4962 12828
rect -3914 12635 -3027 12636
rect -3924 12583 -3914 12635
rect -3862 12583 -3027 12635
rect -1725 12585 -279 12637
rect -227 12585 -217 12637
rect -3425 10982 -3415 11034
rect -3363 10982 -3032 11034
rect -1724 10983 -279 11035
rect -227 10983 -217 11035
rect -5025 10891 -5015 10943
rect -4963 10891 -4953 10943
rect 5662 10402 5714 11030
rect -4840 10401 -678 10402
rect -4840 10349 -4828 10401
rect -4776 10350 -678 10401
rect -626 10350 5714 10402
rect -4776 10349 5714 10350
rect 3748 9911 5265 9945
rect -4838 9404 -4828 9456
rect -4776 9404 -4766 9456
rect -3924 9385 -3914 9437
rect -3862 9385 -3040 9437
rect -1726 9383 -1149 9435
rect -1097 9383 -1087 9435
rect 5231 9418 5265 9911
rect 5213 9365 5223 9418
rect 5276 9365 5286 9418
rect 24534 9360 24544 9424
rect 24608 9360 24618 9424
rect -4837 7595 -4773 8191
rect -3425 7783 -3415 7835
rect -3363 7783 -3029 7835
rect -1726 7783 -1149 7835
rect -1097 7783 -1087 7835
rect 23198 7792 23208 7845
rect 23261 7792 23271 7845
rect -5594 7531 -4773 7595
rect -25689 6209 -25679 6337
rect -25551 6209 -24537 6337
rect -23167 6303 -15778 6336
rect -5594 6313 -5530 7531
rect -23396 6239 -15880 6303
rect -15816 6239 -15778 6303
rect -10714 6249 -10704 6313
rect -10640 6249 -5431 6313
rect -3976 6258 -3415 6310
rect -3363 6258 -3353 6310
rect -23167 6208 -15778 6239
rect -3425 5671 -3415 5723
rect -3363 5671 -2970 5723
rect -1832 5671 -678 5723
rect -626 5671 -616 5723
rect -1149 5129 899 5130
rect -1159 5077 -1149 5129
rect -1097 5077 899 5129
rect -3437 4983 -3427 5047
rect -3363 4983 -3353 5047
rect -3427 4973 -3363 4983
rect 23208 4916 23261 7792
rect 24544 6312 24608 9360
rect 27586 7587 27596 7651
rect 27660 7587 27670 7651
rect 24534 6248 24544 6312
rect 24608 6248 24618 6312
rect 27574 6248 27584 6312
rect 27648 6248 27658 6312
rect 34206 5616 41540 5744
rect 23198 4863 23208 4916
rect 23261 4863 23271 4916
rect 27582 4863 27592 4916
rect 27645 4863 27655 4916
rect -253 3789 867 3790
rect -289 3737 -279 3789
rect -227 3737 867 3789
rect -2131 3298 -2121 3416
rect -2003 3298 3361 3416
rect 23422 2354 23432 2407
rect 23485 2354 23495 2407
rect 22579 1044 22589 1097
rect 22642 1044 22652 1097
rect 22589 -2017 22642 1044
rect 23432 -640 23485 2354
rect 26001 716 26076 4397
rect 25991 641 26001 716
rect 26076 641 26086 716
rect 27570 641 27580 716
rect 27655 641 27665 716
rect 23422 -693 23432 -640
rect 23485 -693 23495 -640
rect 27581 -693 27591 -640
rect 27644 -693 27654 -640
rect 34216 -1324 41540 -1196
rect 22579 -2070 22589 -2017
rect 22643 -2070 22653 -2017
rect 27597 -2070 27607 -2017
rect 27660 -2070 27670 -2017
rect 22589 -2073 22642 -2070
rect -2131 -2631 -2121 -2513
rect -2003 -2631 -1993 -2513
rect -2121 -7531 -2003 -2631
<< via1 >>
rect -12553 53536 -12425 53600
rect -7550 53536 -7486 53600
rect -6989 53536 -6861 53600
rect -9398 52928 -9270 52992
rect -9398 49923 -9270 49987
rect -6989 49921 -6861 49985
rect -9398 39741 -9270 39805
rect -6989 39741 -6861 39805
rect -14172 33901 -14108 33965
rect -19353 32624 -19289 32688
rect -18522 31791 -18458 31855
rect -14240 30470 -14176 30534
rect 93 37382 157 37446
rect 1230 37382 1294 37446
rect 2626 37384 2690 37448
rect 5361 37384 5425 37448
rect 5361 36971 5425 37035
rect 93 36467 157 36531
rect 3427 36467 3491 36531
rect 2334 36023 2398 36087
rect 93 35632 157 35696
rect 883 35632 947 35696
rect 7082 38974 7200 39092
rect 11936 38974 12054 39092
rect 7430 36971 7494 37035
rect 5429 36023 5493 36087
rect 6701 36023 6765 36087
rect 9428 36467 9492 36531
rect -6989 34935 -6925 34999
rect 5430 34356 5494 34420
rect 7428 34354 7492 34418
rect -6989 31747 -6861 31811
rect 4354 30368 4418 30432
rect 8328 30373 8392 30437
rect -9334 29417 -9270 29481
rect -9397 29131 -9269 29195
rect 1951 28784 2079 28848
rect -18326 27511 -18262 27575
rect -14536 27519 -14484 27571
rect -6086 27534 -5958 27598
rect 3399 28531 3463 28595
rect -18326 27034 -18262 27098
rect -18881 26696 -18817 26760
rect -18882 25913 -18818 25977
rect -27540 24984 -27412 25112
rect -18881 24392 -18817 24456
rect -14536 27031 -14484 27083
rect -17256 26696 -17192 26760
rect -14536 25915 -14484 25967
rect -10016 25914 -9888 25978
rect 1952 25756 2080 25820
rect -14538 24389 -14486 24441
rect -3501 24310 -3373 24374
rect -18326 24053 -18262 24117
rect -17255 24053 -17191 24117
rect 9399 28528 9463 28592
rect 3399 23637 3463 23701
rect -14538 22719 -14486 22771
rect -11601 22712 -11473 22776
rect 5643 23633 5707 23697
rect 7017 23637 7081 23701
rect 9399 23637 9463 23701
rect -6086 21607 -5958 21671
rect -3501 20745 -3373 20809
rect -25679 17454 -25551 17582
rect -444 19981 -380 20109
rect 1684 19282 1748 19410
rect 5394 19981 5458 20109
rect 9394 19981 9458 20109
rect 3395 19282 3459 19346
rect 7394 19282 7458 19410
rect 13887 21996 13951 22124
rect 13887 17983 13951 18047
rect -445 17093 -381 17221
rect 1684 17093 1748 17221
rect 7393 17231 7457 17359
rect 9396 17231 9460 17359
rect 13885 17231 13949 17359
rect 3393 16738 3457 16866
rect 5393 16738 5457 16866
rect 13277 16738 13341 16866
rect -3926 16224 -3862 16288
rect -3914 15083 -3862 15135
rect -678 15084 -626 15136
rect -27540 13974 -27412 14102
rect -10693 14077 -10629 14141
rect -3914 14087 -3862 14139
rect -15852 14009 -15788 14073
rect -3914 12583 -3862 12635
rect -279 12585 -227 12637
rect -3415 10982 -3363 11034
rect -279 10983 -227 11035
rect -5015 10891 -4963 10943
rect -4828 10349 -4776 10401
rect -678 10350 -626 10402
rect -4828 9404 -4776 9456
rect -3914 9385 -3862 9437
rect -1149 9383 -1097 9435
rect 5223 9365 5276 9418
rect 24544 9360 24608 9424
rect -3415 7783 -3363 7835
rect -1149 7783 -1097 7835
rect 23208 7792 23261 7845
rect -25679 6209 -25551 6337
rect -15880 6239 -15816 6303
rect -10704 6249 -10640 6313
rect -3415 6258 -3363 6310
rect -3415 5671 -3363 5723
rect -678 5671 -626 5723
rect -1149 5077 -1097 5129
rect -3427 4983 -3363 5047
rect 27596 7587 27660 7651
rect 24544 6248 24608 6312
rect 27584 6248 27648 6312
rect 23208 4863 23261 4916
rect 27592 4863 27645 4916
rect -279 3737 -227 3789
rect -2121 3298 -2003 3416
rect 23432 2354 23485 2407
rect 22589 1044 22642 1097
rect 26001 641 26076 716
rect 27580 641 27655 716
rect 23432 -693 23485 -640
rect 27591 -693 27644 -640
rect 22589 -2070 22643 -2017
rect 27607 -2070 27660 -2017
rect -2121 -2631 -2003 -2513
<< metal2 >>
rect -12553 53600 -12425 53610
rect -7550 53600 -7486 53610
rect -12425 53536 -7550 53600
rect -12553 53526 -12425 53536
rect -7550 53526 -7486 53536
rect -6989 53600 -6861 53610
rect -9398 52992 -9270 53002
rect -9398 49987 -9270 52928
rect -9398 39805 -9270 49923
rect -9398 39728 -9270 39741
rect -6989 49985 -6861 53536
rect -6989 39805 -6861 49921
rect -6989 39731 -6861 39741
rect 7082 39092 7200 39102
rect 11936 39092 12054 39102
rect 7200 38974 11936 39092
rect 7082 38964 7200 38974
rect 11936 38964 12054 38974
rect 93 37446 157 37456
rect 1230 37446 1294 37456
rect 87 37382 93 37446
rect 157 37382 1230 37446
rect 93 37372 157 37382
rect 1230 37372 1294 37382
rect 2626 37448 2690 37458
rect 5361 37448 5425 37458
rect 2690 37384 5361 37448
rect 2626 37374 2690 37384
rect 5361 37374 5425 37384
rect 5361 37035 5425 37045
rect 7430 37035 7494 37045
rect 5425 36971 7430 37035
rect 5361 36961 5425 36971
rect 7430 36961 7494 36971
rect 93 36531 157 36541
rect 3427 36531 3491 36541
rect 9428 36531 9492 36541
rect 157 36467 3427 36531
rect 3491 36467 9428 36531
rect 93 36457 157 36467
rect 3427 36457 3491 36467
rect 9428 36457 9492 36467
rect 2334 36087 2398 36097
rect 5429 36087 5493 36097
rect 6701 36087 6765 36097
rect 2398 36023 5429 36087
rect 5493 36023 6701 36087
rect 2334 36013 2398 36023
rect 5429 36013 5493 36023
rect 6701 36013 6765 36023
rect 93 35696 157 35706
rect 883 35696 947 35706
rect 90 35632 93 35696
rect 157 35632 883 35696
rect 93 35622 157 35632
rect 883 35622 947 35632
rect -6989 34999 -6925 35009
rect -6989 34925 -6925 34935
rect 5430 34420 5494 34430
rect -14172 33965 -14108 33975
rect -12818 33965 -12754 33975
rect -14108 33901 -12818 33965
rect -14172 33891 -14108 33901
rect -12818 33891 -12754 33901
rect -19353 32688 -19289 32698
rect -19383 32624 -19353 32688
rect -19289 32624 -19254 32688
rect -19383 26015 -19254 32624
rect 5317 32345 5381 32355
rect 5430 32345 5494 34356
rect 7428 34418 7492 34428
rect 7428 32362 7492 34354
rect 5381 32281 5494 32345
rect 7364 32352 7492 32362
rect 7428 32288 7492 32352
rect 5317 32271 5381 32281
rect 7364 32278 7428 32288
rect -18522 31855 -18458 31865
rect -18523 31791 -18522 31855
rect -18458 31791 -18394 31855
rect -18523 27609 -18394 31791
rect -6989 31811 8057 31840
rect -6861 31747 7965 31811
rect 8029 31747 8057 31811
rect -6989 31712 8057 31747
rect -14240 30534 -14176 30544
rect -12813 30534 -12749 30544
rect -14176 30470 -12813 30534
rect -14240 30460 -14176 30470
rect -12813 30460 -12749 30470
rect 4354 30432 4418 30442
rect 4354 30358 4418 30368
rect 8328 30437 8392 30447
rect 8328 30363 8392 30373
rect -9334 29481 -9270 29491
rect -9334 29407 -9270 29417
rect -9347 29205 2453 29228
rect -9397 29195 2453 29205
rect 3326 29195 3390 29205
rect -9269 29131 3326 29195
rect -9397 29121 2453 29131
rect 3326 29121 3390 29131
rect -9347 29100 2453 29121
rect 1951 28848 2079 28858
rect 4701 28848 4765 28858
rect 2079 28784 4701 28848
rect 1951 28774 2079 28784
rect 4701 28774 4765 28784
rect 7960 28846 8024 28856
rect 3399 28595 3463 28605
rect 4328 28595 4392 28605
rect 3463 28531 4328 28595
rect 4392 28531 4398 28595
rect 3399 28521 3463 28531
rect 4328 28521 4392 28531
rect -18523 27575 -18246 27609
rect -6086 27598 -5958 27623
rect -18523 27511 -18326 27575
rect -18262 27511 -18246 27575
rect -18523 27480 -18246 27511
rect -14536 27571 -14484 27581
rect -18326 27098 -18262 27108
rect -18262 27034 -17257 27098
rect -14536 27083 -14484 27519
rect -18326 27024 -18262 27034
rect -18881 26760 -18817 26770
rect -17256 26760 -17192 26770
rect -18817 26696 -17256 26760
rect -18881 26686 -18817 26696
rect -17256 26686 -17192 26696
rect -19383 25977 -18816 26015
rect -19383 25913 -18882 25977
rect -18818 25913 -18816 25977
rect -19383 25886 -18816 25913
rect -14536 25967 -14484 27031
rect -14536 25905 -14484 25915
rect -10016 25978 -9888 25988
rect -27540 25112 -27412 25122
rect -27540 14102 -27412 24984
rect -18881 24456 -18817 24466
rect -18885 24392 -18881 24456
rect -18817 24392 -17231 24456
rect -14538 24441 -14486 24451
rect -18881 24382 -18817 24392
rect -18326 24117 -18262 24127
rect -17255 24117 -17191 24127
rect -18334 24053 -18326 24117
rect -18262 24053 -17255 24117
rect -18326 24043 -18262 24053
rect -17255 24043 -17191 24053
rect -14538 22771 -14486 24389
rect -14538 22713 -14486 22719
rect -11601 22776 -11473 22786
rect -27540 13964 -27412 13974
rect -25679 17582 -25551 17592
rect -25679 6337 -25551 17454
rect -15852 14073 -15788 14083
rect -15852 13999 -15788 14009
rect -11601 10181 -11473 22712
rect -10016 17968 -9888 25914
rect -6086 21671 -5958 27534
rect 1952 25820 2080 25830
rect 7960 25820 8024 28782
rect 8338 28592 8402 28602
rect 9399 28592 9463 28602
rect 8402 28528 9399 28592
rect 9463 28528 9473 28592
rect 8338 28518 8402 28528
rect 9399 28518 9463 28528
rect 2080 25756 8024 25820
rect 1952 25746 2080 25756
rect -6086 21597 -5958 21607
rect -3501 24374 -3373 24393
rect -3501 20809 -3373 24310
rect 3399 23701 3463 23709
rect 5643 23697 5707 23707
rect 3463 23637 5643 23697
rect 3399 23633 5643 23637
rect 3399 23627 3463 23633
rect 5643 23623 5707 23633
rect 7017 23701 7081 23711
rect 9399 23701 9463 23711
rect 7081 23637 9399 23701
rect 9463 23637 9467 23701
rect 7017 23627 7081 23637
rect 9399 23627 9463 23637
rect -3501 20735 -3373 20745
rect 13887 22124 13951 22134
rect -444 20109 -380 20119
rect 5394 20109 5458 20119
rect 9394 20109 9458 20119
rect -10016 17904 -9984 17968
rect -9920 17904 -9888 17968
rect -8599 19981 -444 20109
rect -380 19981 5394 20109
rect 5458 19981 9394 20109
rect 9458 19981 9474 20109
rect -9984 17894 -9920 17904
rect -10693 14141 -10629 14151
rect -10693 14067 -10629 14077
rect -11601 10117 -11570 10181
rect -11506 10117 -11473 10181
rect -8599 10223 -8471 19981
rect -444 19971 -380 19981
rect 5394 19971 5458 19981
rect 9394 19971 9458 19981
rect 1684 19410 1748 19420
rect 7394 19410 7458 19420
rect 1748 19346 7394 19410
rect 1748 19282 3395 19346
rect 3459 19282 7394 19346
rect 7458 19282 7468 19410
rect 1684 19272 1748 19282
rect 3395 19272 3459 19282
rect 7394 19272 7458 19282
rect 13887 18047 13951 21996
rect 13887 17973 13951 17983
rect 7393 17359 7457 17369
rect 9396 17359 9460 17369
rect 13885 17359 13949 17369
rect 7457 17231 9396 17359
rect 9460 17231 13885 17359
rect 13949 17231 13962 17359
rect -445 17221 -381 17231
rect 1684 17221 1748 17231
rect 7393 17221 7457 17231
rect 9396 17221 9460 17231
rect 13885 17221 13949 17231
rect -8108 17157 -445 17221
rect -8108 17093 -8045 17157
rect -7981 17093 -445 17157
rect -381 17093 1684 17221
rect -8108 17092 1748 17093
rect -8045 17083 -7981 17092
rect -445 17083 -381 17092
rect 1684 17083 1748 17092
rect 3393 16866 3457 16876
rect 5393 16866 5457 16876
rect 13277 16866 13341 16876
rect 3457 16738 5393 16866
rect 5457 16738 13277 16866
rect 13341 16738 13351 16866
rect 3393 16728 3457 16738
rect 5393 16728 5457 16738
rect 13277 16728 13341 16738
rect -8044 16288 -7980 16298
rect -3926 16288 -3862 16298
rect -7980 16224 -3926 16288
rect -8044 16214 -7980 16224
rect -3926 16214 -3862 16224
rect -3914 15135 -3862 16214
rect -3914 14139 -3862 15083
rect -3914 12635 -3862 14087
rect -5015 10943 -4963 10953
rect -5015 10401 -4963 10891
rect -4828 10401 -4776 10411
rect -5015 10349 -4828 10401
rect -8535 10159 -8471 10223
rect -8599 10139 -8471 10159
rect -11601 10113 -11473 10117
rect -11570 10107 -11506 10113
rect -4828 9456 -4776 10349
rect -4828 9394 -4776 9404
rect -3914 9437 -3862 12583
rect -678 15136 -626 15146
rect -3914 9375 -3862 9385
rect -3415 11034 -3363 11044
rect -3415 7835 -3363 10982
rect -678 10402 -626 15084
rect -10704 6313 -10640 6323
rect -15880 6303 -15816 6313
rect -10704 6239 -10640 6249
rect -3415 6310 -3363 7783
rect -15880 6229 -15816 6239
rect -25679 6199 -25551 6209
rect -3415 5723 -3363 6258
rect -3415 5057 -3363 5671
rect -1149 9435 -1097 9451
rect -1149 7835 -1097 9383
rect -1149 5129 -1097 7783
rect -678 5723 -626 10350
rect -678 5661 -626 5671
rect -279 12637 -227 12647
rect -279 11035 -227 12585
rect -1149 5067 -1097 5077
rect -8395 5047 -8331 5057
rect -3427 5047 -3363 5057
rect -8331 4983 -3427 5047
rect -8395 4973 -8331 4983
rect -3427 4973 -3363 4983
rect -279 3789 -227 10983
rect 5223 9418 5276 9428
rect 24544 9424 24608 9434
rect 5276 9365 24544 9418
rect 5223 9355 5276 9365
rect 24544 9350 24608 9360
rect 23208 7845 23261 7855
rect 17672 7792 23208 7845
rect 17672 7717 17725 7792
rect 23208 7782 23261 7792
rect 12920 7664 17725 7717
rect 25495 7651 25559 9116
rect 27596 7651 27660 7661
rect 25495 7587 27596 7651
rect 27596 7577 27660 7587
rect 24544 6312 24608 6322
rect 27584 6312 27648 6322
rect 24608 6248 27584 6312
rect 24544 6238 24608 6248
rect 27584 6238 27648 6248
rect 23208 4916 23261 4926
rect 27592 4916 27645 4926
rect 23261 4863 27592 4916
rect 23208 4853 23261 4863
rect 27592 4853 27645 4863
rect -279 3727 -227 3737
rect -2121 3416 -2003 3426
rect -2121 -2513 -2003 3298
rect 3670 2688 5404 2741
rect 5351 2407 5404 2688
rect 23432 2407 23485 2417
rect 5351 2354 23432 2407
rect 23432 2344 23485 2354
rect 22589 1097 22642 1107
rect 18808 1044 22589 1097
rect 22589 1034 22642 1044
rect 26001 716 26076 726
rect 27580 716 27655 726
rect 26076 641 27580 716
rect 26001 631 26076 641
rect 27580 631 27655 641
rect 23432 -640 23485 -630
rect 27591 -640 27644 -630
rect 23485 -693 27591 -640
rect 23432 -703 23485 -693
rect 27591 -703 27644 -693
rect 22589 -2017 22643 -2007
rect 27607 -2017 27660 -2007
rect 22643 -2070 27607 -2017
rect 22589 -2080 22643 -2070
rect 27607 -2080 27660 -2070
rect -2121 -2641 -2003 -2631
<< via2 >>
rect -6989 34935 -6925 34999
rect -12818 33901 -12754 33965
rect 5317 32281 5381 32345
rect 7364 32288 7428 32352
rect 7965 31747 8029 31811
rect -12813 30470 -12749 30534
rect 4354 30368 4418 30432
rect 8328 30373 8392 30437
rect -9334 29417 -9270 29481
rect 3326 29131 3390 29195
rect 4701 28784 4765 28848
rect 7960 28782 8024 28846
rect 4328 28531 4392 28595
rect -15852 14009 -15788 14073
rect 8338 28528 8402 28592
rect -9984 17904 -9920 17968
rect -10693 14077 -10629 14141
rect -11570 10117 -11506 10181
rect -8045 17093 -7981 17157
rect -8044 16224 -7980 16288
rect -8599 10159 -8535 10223
rect -15880 6239 -15816 6303
rect -10704 6249 -10640 6313
rect -8395 4983 -8331 5047
<< metal3 >>
rect -7018 34999 -6902 35031
rect -7018 34935 -6989 34999
rect -6925 34935 -6902 34999
rect -7018 34908 -6902 34935
rect -12840 33965 -12734 33991
rect -12840 33901 -12818 33965
rect -12754 33901 -12734 33965
rect -12840 33875 -12734 33901
rect -11166 31738 -11102 32675
rect 7354 32352 7438 32357
rect 5307 32345 5391 32350
rect 5121 32281 5317 32345
rect 5381 32281 5391 32345
rect 7354 32288 7364 32352
rect 7428 32288 7607 32352
rect 7354 32283 7438 32288
rect 5307 32276 5391 32281
rect 4964 31452 5028 32173
rect 7702 31452 7766 32173
rect 7942 31811 8053 31841
rect 7942 31747 7965 31811
rect 8029 31747 8053 31811
rect 7942 31723 8053 31747
rect 4964 31375 5028 31388
rect 7702 31375 7766 31388
rect 5702 31191 5766 31192
rect 3944 31123 4742 31187
rect 4941 31127 5766 31191
rect -12838 30534 -12729 30558
rect -12838 30470 -12813 30534
rect -12749 30470 -12729 30534
rect -12838 30442 -12729 30470
rect 3961 30389 4025 31123
rect 4325 30432 4440 30460
rect 4325 30368 4354 30432
rect 4418 30368 4440 30432
rect 5702 30394 5766 31127
rect 6964 31191 7028 31192
rect 6964 31127 7789 31191
rect 6964 30394 7028 31127
rect 7988 31123 8786 31187
rect 8300 30437 8415 30464
rect 4325 30342 4440 30368
rect 8300 30373 8328 30437
rect 8392 30373 8415 30437
rect 8705 30389 8769 31123
rect 8300 30348 8415 30373
rect -9361 29481 -9251 29512
rect -9361 29417 -9334 29481
rect -9270 29417 -9251 29481
rect -9361 29393 -9251 29417
rect 3961 29389 4025 30187
rect 4328 29982 4609 30046
rect 3298 29195 3418 29225
rect 3298 29131 3326 29195
rect 3390 29131 3418 29195
rect 3298 29102 3418 29131
rect 3961 28389 4025 29187
rect 4328 28600 4392 29982
rect 5702 29394 5766 30192
rect 6964 29394 7028 30192
rect 8121 29982 8402 30046
rect 4701 28853 4765 29012
rect 4691 28848 4775 28853
rect 4691 28784 4701 28848
rect 4765 28784 4775 28848
rect 4691 28779 4775 28784
rect 4318 28595 4402 28600
rect 4318 28531 4328 28595
rect 4392 28593 4402 28595
rect 4392 28531 4579 28593
rect 4318 28529 4579 28531
rect 4318 28526 4402 28529
rect 5702 28394 5766 29192
rect 6964 28394 7028 29192
rect 7960 28851 8024 29021
rect 7950 28846 8034 28851
rect 7950 28782 7960 28846
rect 8024 28782 8034 28846
rect 7950 28777 8034 28782
rect 8338 28597 8402 29982
rect 8705 29389 8769 30187
rect 8328 28593 8412 28597
rect 8151 28592 8412 28593
rect 8151 28529 8338 28592
rect 8328 28528 8338 28529
rect 8402 28528 8412 28592
rect 8328 28523 8412 28528
rect 8705 28389 8769 29187
rect 3961 27451 4025 28187
rect 5702 27451 5766 28192
rect 3961 27389 4764 27451
rect 3966 27387 4764 27389
rect 4966 27394 5766 27451
rect 6964 27451 7028 28192
rect 8705 27451 8769 28187
rect 6964 27394 7764 27451
rect 4966 27387 5764 27394
rect 6966 27387 7764 27394
rect 7966 27389 8769 27451
rect 7966 27387 8764 27389
rect 4966 26402 5030 27200
rect 7700 26402 7764 27200
rect -10016 17968 -9888 17999
rect -10016 17904 -9984 17968
rect -9920 17904 -9888 17968
rect -10016 17870 -9888 17904
rect -8074 17157 -7950 17194
rect -8074 17093 -8045 17157
rect -7981 17093 -7950 17157
rect -8074 17061 -7950 17093
rect -8054 16288 -7970 16293
rect -16348 16203 -15328 16267
rect -13748 16203 -12728 16267
rect -11148 16203 -10128 16267
rect -8414 16224 -8044 16288
rect -7980 16224 -7970 16288
rect -8054 16219 -7970 16224
rect -16700 14880 -16636 15900
rect -9826 14873 -9762 15893
rect -13594 14472 -12861 14536
rect -10703 14141 -10619 14146
rect -15869 14073 -15768 14097
rect -10960 14077 -10693 14141
rect -10629 14077 -10619 14141
rect -15869 14009 -15852 14073
rect -15788 14009 -15768 14073
rect -10703 14072 -10619 14077
rect -15869 13986 -15768 14009
rect -16700 12280 -16636 13300
rect -9826 12273 -9762 13293
rect -16351 11937 -15331 12001
rect -13751 11937 -12731 12001
rect -11151 11937 -10131 12001
rect -8628 10223 -8510 10250
rect -11598 10181 -11475 10211
rect -11598 10117 -11570 10181
rect -11506 10117 -11475 10181
rect -8628 10159 -8599 10223
rect -8535 10159 -8510 10223
rect -8628 10138 -8510 10159
rect -11598 10089 -11475 10117
rect -16348 8403 -15328 8467
rect -13748 8403 -12728 8467
rect -11148 8403 -10128 8467
rect -16700 7080 -16636 8100
rect -9826 7073 -9762 8093
rect -13594 6672 -12861 6736
rect -15900 6303 -15800 6328
rect -10714 6313 -10630 6318
rect -15900 6239 -15880 6303
rect -15816 6239 -15800 6303
rect -10955 6249 -10704 6313
rect -10640 6249 -10630 6313
rect -10714 6244 -10630 6249
rect -15900 6217 -15800 6239
rect -16700 4480 -16636 5500
rect -9826 4473 -9762 5493
rect -8395 5052 -8331 5314
rect -8405 5047 -8321 5052
rect -8405 4983 -8395 5047
rect -8331 4983 -8321 5047
rect -8405 4978 -8321 4983
rect -16351 4137 -15331 4201
rect -13751 4137 -12731 4201
rect -11151 4137 -10131 4201
<< via3 >>
rect -6989 34935 -6925 34999
rect -12818 33901 -12754 33965
rect 7965 31747 8029 31811
rect -12813 30470 -12749 30534
rect 4354 30368 4418 30432
rect 8328 30373 8392 30437
rect -9334 29417 -9270 29481
rect 3326 29131 3390 29195
rect -9984 17904 -9920 17968
rect -8045 17093 -7981 17157
rect -15852 14009 -15788 14073
rect -11570 10117 -11506 10181
rect -8599 10159 -8535 10223
rect -15880 6239 -15816 6303
<< metal4 >>
rect -6990 34999 -6924 35000
rect -10105 34935 -6989 34999
rect -6925 34935 -6924 34999
rect -6990 34934 -6924 34935
rect -12819 33965 -12753 33966
rect -12819 33901 -12818 33965
rect -12754 33901 -12298 33965
rect -12819 33900 -12753 33901
rect 4701 31450 4765 32172
rect 7965 31812 8029 32172
rect 7964 31811 8030 31812
rect 7964 31747 7965 31811
rect 8029 31747 8030 31811
rect 7964 31746 8030 31747
rect 3944 31386 4765 31450
rect 4941 31390 5739 31454
rect 6991 31390 7789 31454
rect 7965 31450 8029 31746
rect 4701 31372 4765 31386
rect 7965 31386 8786 31450
rect 7965 31372 8029 31386
rect -12814 30534 -12748 30535
rect -12814 30470 -12813 30534
rect -12749 30470 -12207 30534
rect -12814 30469 -12748 30470
rect 3698 30389 3762 31187
rect 4353 30432 4419 30433
rect 4353 30368 4354 30432
rect 4418 30368 4705 30432
rect 5965 30394 6029 31192
rect 6701 30394 6765 31192
rect 8327 30437 8393 30438
rect 8028 30373 8328 30437
rect 8392 30373 8393 30437
rect 8968 30389 9032 31187
rect 8327 30372 8393 30373
rect 4353 30367 4419 30368
rect -9335 29481 -9269 29482
rect -10091 29417 -9334 29481
rect -9270 29417 -9269 29481
rect -9335 29416 -9269 29417
rect 3698 29389 3762 30187
rect 4701 29396 4765 30194
rect 5965 29394 6029 30192
rect 6701 29394 6765 30192
rect 7965 29396 8029 30194
rect 8968 29389 9032 30187
rect 3325 29195 3391 29196
rect 3325 29131 3326 29195
rect 3390 29131 3762 29195
rect 3325 29130 3391 29131
rect 3698 28389 3762 29131
rect 4967 28378 5031 29176
rect 5965 28394 6029 29192
rect 6701 28394 6765 29192
rect 7699 28378 7763 29176
rect 8968 28389 9032 29187
rect 3698 27389 3762 28187
rect 5965 27394 6029 28192
rect 6701 27394 6765 28192
rect 8968 27389 9032 28187
rect 4703 27188 4767 27200
rect 7963 27188 8027 27200
rect 3966 27124 4767 27188
rect 4966 27124 5764 27188
rect 6966 27124 7764 27188
rect 7963 27124 8764 27188
rect 4703 26402 4767 27124
rect 7963 26402 8027 27124
rect -9985 17968 -9919 17969
rect -9985 17904 -9984 17968
rect -9920 17904 -9919 17968
rect -9985 17903 -9919 17904
rect -9984 17495 -9920 17903
rect -16348 17145 -15328 17209
rect -13748 17145 -12728 17209
rect -11148 17145 -10128 17209
rect -8046 17157 -7980 17158
rect -8541 17093 -8045 17157
rect -7981 17093 -7980 17157
rect -8046 17092 -7980 17093
rect -17642 14880 -17578 15900
rect -8884 14873 -8820 15893
rect -15853 14073 -15787 14074
rect -15853 14009 -15852 14073
rect -15788 14009 -15361 14073
rect -15853 14008 -15787 14009
rect -13753 13625 -12733 13689
rect -17642 12280 -17578 13300
rect -8884 12273 -8820 13293
rect -16351 10995 -15331 11059
rect -13751 10995 -12731 11059
rect -11151 10995 -10131 11059
rect -8600 10223 -8534 10224
rect -11571 10181 -11505 10182
rect -11571 10117 -11570 10181
rect -11506 10117 -11505 10181
rect -8600 10159 -8599 10223
rect -8535 10159 -8534 10223
rect -8600 10158 -8534 10159
rect -11571 10116 -11505 10117
rect -11570 9700 -11506 10116
rect -8599 9696 -8535 10158
rect -16348 9345 -15328 9409
rect -13748 9345 -12728 9409
rect -11148 9345 -10128 9409
rect -17642 7080 -17578 8100
rect -8884 7073 -8820 8093
rect -15881 6303 -15815 6304
rect -15881 6239 -15880 6303
rect -15816 6239 -15329 6303
rect -15881 6238 -15815 6239
rect -13753 5825 -12733 5889
rect -17642 4480 -17578 5500
rect -8884 4473 -8820 5493
rect -16351 3195 -15331 3259
rect -13751 3195 -12731 3259
rect -11151 3195 -10131 3259
use a_mux2_en  a_mux2_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/a_mux2_en
timestamp 1653911004
transform 1 0 29925 0 1 23897
box -2638 -2585 3429 115
use a_mux2_en  a_mux2_en_1
timestamp 1653911004
transform 0 -1 -14354 1 0 68726
box -2638 -2585 3429 115
use a_mux4_en  a_mux4_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/a_mux4_en
timestamp 1653911004
transform 1 0 30933 0 1 1386
box -3690 -5314 3456 148
use a_mux4_en  a_mux4_en_1
timestamp 1653911004
transform 1 0 30933 0 1 8326
box -3690 -5314 3456 148
use comparator  comparator_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/comparator
timestamp 1653911004
transform 0 -1 -12766 1 0 31540
box -171 198 1585 4870
use esd_cell  esd_cell_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/esd_cell
timestamp 1653911004
transform 1 0 -32809 0 1 16027
box -65 -65 3553 3095
use esd_cell  esd_cell_1
timestamp 1653911004
transform 1 0 -32809 0 1 23557
box -65 -65 3553 3095
use esd_cell  esd_cell_2
timestamp 1653911004
transform 1 0 12350 0 1 37546
box -65 -65 3553 3095
use esd_cell  esd_cell_3
timestamp 1653911004
transform 0 1 -3548 -1 0 -2736
box -65 -65 3553 3095
use esd_cell  esd_cell_4
timestamp 1653911004
transform 0 -1 -11568 1 0 73319
box -65 -65 3553 3095
use esd_cell  esd_cell_5
timestamp 1653911004
transform 1 0 36372 0 1 21122
box -65 -65 3553 3095
use esd_cell  esd_cell_6
timestamp 1653911004
transform 1 0 36372 0 1 -2751
box -65 -65 3553 3095
use esd_cell  esd_cell_7
timestamp 1653911004
transform 1 0 36372 0 1 4189
box -65 -65 3553 3095
use onebit_dac  onebit_dac_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/onebit_dac
timestamp 1653911004
transform 1 0 -17091 0 1 24436
box -313 -1154 1895 1114
use onebit_dac  onebit_dac_1
timestamp 1653911004
transform 1 0 -17086 0 1 27078
box -313 -1154 1895 1114
use ota  ota_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/ota
timestamp 1653911004
transform 1 0 7664 0 1 17642
box -7664 -17642 18422 2891
use ota  ota_1
timestamp 1653911004
transform 0 -1 -7144 1 0 47315
box -7664 -17642 18422 2891
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_0
timestamp 1653911004
transform 0 1 9865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_1
timestamp 1653911004
transform 0 1 9865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_2
timestamp 1653911004
transform 0 1 9865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_3
timestamp 1653911004
transform 0 1 9865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_4
timestamp 1653911004
transform 0 1 9865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_5
timestamp 1653911004
transform 0 1 9865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_6
timestamp 1653911004
transform 0 1 9865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_7
timestamp 1653911004
transform 0 1 9865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_8
timestamp 1653911004
transform 0 1 8865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_9
timestamp 1653911004
transform 0 1 8865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_10
timestamp 1653911004
transform 0 1 8865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_11
timestamp 1653911004
transform 0 1 8865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_12
timestamp 1653911004
transform 0 1 8865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_13
timestamp 1653911004
transform 0 1 8865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_14
timestamp 1653911004
transform 0 1 8865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_15
timestamp 1653911004
transform 0 1 8865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_16
timestamp 1653911004
transform 0 1 8865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_17
timestamp 1653911004
transform 0 1 7865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_18
timestamp 1653911004
transform 0 1 7865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_19
timestamp 1653911004
transform 0 1 7865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_20
timestamp 1653911004
transform 0 1 7865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_21
timestamp 1653911004
transform 0 1 7865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_22
timestamp 1653911004
transform 0 1 7865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_23
timestamp 1653911004
transform 0 1 7865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_24
timestamp 1653911004
transform 0 1 7865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_25
timestamp 1653911004
transform 0 1 7865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_26
timestamp 1653911004
transform 0 1 6865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_27
timestamp 1653911004
transform 0 1 6865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_28
timestamp 1653911004
transform 0 1 6865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_29
timestamp 1653911004
transform 0 1 6865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_30
timestamp 1653911004
transform 0 1 6865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_31
timestamp 1653911004
transform 0 1 6865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_32
timestamp 1653911004
transform 0 1 6865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_33
timestamp 1653911004
transform 0 1 6865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_34
timestamp 1653911004
transform 0 1 6865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_35
timestamp 1653911004
transform 0 -1 3865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_36
timestamp 1653911004
transform 0 -1 3865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_37
timestamp 1653911004
transform 0 -1 2865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_38
timestamp 1653911004
transform 0 -1 2865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_39
timestamp 1653911004
transform 0 -1 3865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_40
timestamp 1653911004
transform 0 -1 3865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_41
timestamp 1653911004
transform 0 -1 2865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_42
timestamp 1653911004
transform 0 -1 2865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_43
timestamp 1653911004
transform 0 -1 3865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_44
timestamp 1653911004
transform 0 -1 3865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_45
timestamp 1653911004
transform 0 -1 2865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_46
timestamp 1653911004
transform 0 -1 2865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_47
timestamp 1653911004
transform 0 -1 3865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_48
timestamp 1653911004
transform 0 -1 3865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_49
timestamp 1653911004
transform 0 -1 2865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_50
timestamp 1653911004
transform 0 -1 2865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_51
timestamp 1653911004
transform 0 -1 3865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_52
timestamp 1653911004
transform 0 -1 2865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_53
timestamp 1653911004
transform 0 -1 5865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_54
timestamp 1653911004
transform 0 -1 4865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_55
timestamp 1653911004
transform 0 -1 5865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_56
timestamp 1653911004
transform 0 -1 4865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_57
timestamp 1653911004
transform 0 -1 5865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_58
timestamp 1653911004
transform 0 -1 4865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_59
timestamp 1653911004
transform 0 -1 5865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_60
timestamp 1653911004
transform 0 -1 4865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_61
timestamp 1653911004
transform 0 -1 5865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_62
timestamp 1653911004
transform 0 -1 5865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_63
timestamp 1653911004
transform 0 -1 4865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_64
timestamp 1653911004
transform 0 -1 4865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_65
timestamp 1653911004
transform 0 -1 5865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_66
timestamp 1653911004
transform 0 -1 5865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_67
timestamp 1653911004
transform 0 -1 4865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_68
timestamp 1653911004
transform 0 -1 4865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_69
timestamp 1653911004
transform 0 -1 5865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_70
timestamp 1653911004
transform 0 1 9865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_71
timestamp 1653911004
transform 0 -1 4865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_0
timestamp 1653911004
transform 1 0 -6697 0 1 19276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_1
timestamp 1653911004
transform 1 0 -6697 0 1 16676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_2
timestamp 1653911004
transform 1 0 -6697 0 1 14076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_3
timestamp 1653911004
transform 1 0 -6697 0 1 11476
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_4
timestamp 1653911004
transform 1 0 -6697 0 1 8876
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_5
timestamp 1653911004
transform 1 0 -17097 0 1 3676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_6
timestamp 1653911004
transform 1 0 -9297 0 1 11476
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_7
timestamp 1653911004
transform 1 0 -9297 0 1 14076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_8
timestamp 1653911004
transform 1 0 -9297 0 1 16676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_9
timestamp 1653911004
transform 1 0 -9297 0 1 19276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_10
timestamp 1653911004
transform 1 0 -14497 0 1 3676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_11
timestamp 1653911004
transform 1 0 -11897 0 1 11476
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_12
timestamp 1653911004
transform 1 0 -11897 0 1 14076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_13
timestamp 1653911004
transform 1 0 -11897 0 1 16676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_14
timestamp 1653911004
transform 1 0 -11897 0 1 19276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_15
timestamp 1653911004
transform 1 0 -9297 0 1 3676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_16
timestamp 1653911004
transform 1 0 -14497 0 1 11476
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_17
timestamp 1653911004
transform 1 0 -14497 0 1 14076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_18
timestamp 1653911004
transform 1 0 -14497 0 1 16676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_19
timestamp 1653911004
transform 1 0 -14497 0 1 19276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_20
timestamp 1653911004
transform 1 0 -11897 0 1 3676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_21
timestamp 1653911004
transform 1 0 -17097 0 1 11476
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_22
timestamp 1653911004
transform 1 0 -17097 0 1 14076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_23
timestamp 1653911004
transform 1 0 -17097 0 1 16676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_24
timestamp 1653911004
transform 1 0 -17097 0 1 19276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_25
timestamp 1653911004
transform 1 0 -19697 0 1 8876
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_26
timestamp 1653911004
transform 1 0 -19697 0 1 11476
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_27
timestamp 1653911004
transform 1 0 -19697 0 1 14076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_28
timestamp 1653911004
transform 1 0 -19697 0 1 16676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_29
timestamp 1653911004
transform 1 0 -19697 0 1 19276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_30
timestamp 1653911004
transform 1 0 -14497 0 1 8876
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_31
timestamp 1653911004
transform 1 0 -17097 0 1 8876
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_32
timestamp 1653911004
transform 1 0 -14497 0 1 6276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_33
timestamp 1653911004
transform 1 0 -17097 0 1 6276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_34
timestamp 1653911004
transform 1 0 -9297 0 1 8876
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_35
timestamp 1653911004
transform 1 0 -11897 0 1 8876
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_36
timestamp 1653911004
transform 1 0 -9297 0 1 6276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_37
timestamp 1653911004
transform 1 0 -11897 0 1 6276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_38
timestamp 1653911004
transform 1 0 -19697 0 1 6276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_39
timestamp 1653911004
transform 1 0 -6697 0 1 6276
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_40
timestamp 1653911004
transform 1 0 -19697 0 1 3676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_41
timestamp 1653911004
transform 1 0 -6697 0 1 3676
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_42
timestamp 1653911004
transform 1 0 -19697 0 1 1076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_43
timestamp 1653911004
transform 1 0 -6697 0 1 1076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_44
timestamp 1653911004
transform 1 0 -17097 0 1 1076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_45
timestamp 1653911004
transform 1 0 -14497 0 1 1076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_46
timestamp 1653911004
transform 1 0 -11897 0 1 1076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_47
timestamp 1653911004
transform 1 0 -9297 0 1 1076
box -1030 -980 977 980
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_0
timestamp 1653911004
transform 1 0 -11147 0 -1 30508
box -1310 -1260 1210 1261
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_1
timestamp 1653911004
transform 1 0 -11147 0 -1 33918
box -1310 -1260 1210 1261
use sky130_fd_pr__nfet_01v8_CFEPS5  sky130_fd_pr__nfet_01v8_CFEPS5_0
timestamp 1653911004
transform 1 0 -20105 0 -1 33421
box -311 -275 311 275
use sky130_fd_pr__pfet_01v8_XAYTAL  sky130_fd_pr__pfet_01v8_XAYTAL_0
timestamp 1653911004
transform 1 0 -20105 0 -1 32821
box -311 -319 311 319
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/transmission_gate
timestamp 1653911004
transform 1 0 -24468 0 1 13627
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1653911004
transform 1 0 -5241 0 1 13700
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1653911004
transform 1 0 -24468 0 1 5859
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1653911004
transform 1 0 -2967 0 1 12195
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1653911004
transform 1 0 -2967 0 1 10595
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1653911004
transform 1 0 -2967 0 1 8995
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1653911004
transform 1 0 -2967 0 1 7395
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1653911004
transform 1 0 -5241 0 1 5869
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1653911004
transform 0 1 -5401 -1 0 11991
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1653911004
transform 0 -1 -4389 1 0 8354
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1653911004
transform -1 0 -1901 0 -1 15522
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1653911004
transform -1 0 -1903 0 -1 6110
box -216 -51 1283 1063
use transmission_gate  transmission_gate_12
timestamp 1653911004
transform 0 -1 3839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_13
timestamp 1653911004
transform 0 -1 5839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_14
timestamp 1653911004
transform 0 -1 7839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_15
timestamp 1653911004
transform 0 -1 9839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_16
timestamp 1653911004
transform 0 1 -826 -1 0 18922
box -216 -51 1283 1063
use transmission_gate  transmission_gate_17
timestamp 1653911004
transform 0 -1 3845 1 0 21294
box -216 -51 1283 1063
use transmission_gate  transmission_gate_18
timestamp 1653911004
transform 0 -1 9844 1 0 21294
box -216 -51 1283 1063
use transmission_gate  transmission_gate_19
timestamp 1653911004
transform -1 0 6948 0 -1 24081
box -216 -51 1283 1063
use transmission_gate  transmission_gate_20
timestamp 1653911004
transform 0 -1 3873 1 0 34268
box -216 -51 1283 1063
use transmission_gate  transmission_gate_21
timestamp 1653911004
transform 0 -1 5873 1 0 34268
box -216 -51 1283 1063
use transmission_gate  transmission_gate_22
timestamp 1653911004
transform 0 -1 7873 1 0 34268
box -216 -51 1283 1063
use transmission_gate  transmission_gate_23
timestamp 1653911004
transform 0 -1 9873 1 0 34268
box -216 -51 1283 1063
use transmission_gate  transmission_gate_24
timestamp 1653911004
transform 1 0 1359 0 -1 37827
box -216 -51 1283 1063
use transmission_gate  transmission_gate_25
timestamp 1653911004
transform 1 0 1007 0 -1 36077
box -216 -51 1283 1063
use transmission_gate  transmission_gate_26
timestamp 1653911004
transform -1 0 -7618 0 -1 50365
box -216 -51 1283 1063
use transmission_gate  transmission_gate_27
timestamp 1653911004
transform 1 0 -13548 0 1 27131
box -216 -51 1283 1063
use transmission_gate  transmission_gate_28
timestamp 1653911004
transform 1 0 -13548 0 1 25531
box -216 -51 1283 1063
use transmission_gate  transmission_gate_29
timestamp 1653911004
transform 1 0 -13548 0 1 23931
box -216 -51 1283 1063
use transmission_gate  transmission_gate_30
timestamp 1653911004
transform 1 0 -13548 0 1 22331
box -216 -51 1283 1063
use transmission_gate  transmission_gate_31
timestamp 1653911004
transform 1 0 -24236 0 1 24644
box -216 -51 1283 1063
use transmission_gate  transmission_gate_32
timestamp 1653911004
transform 1 0 -24236 0 1 17101
box -216 -51 1283 1063
<< labels >>
flabel metal1 34371 5685 34371 5685 1 FreeSans 400 0 0 0 out
<< end >>
