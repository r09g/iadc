magic
tech sky130A
magscale 1 2
timestamp 1654894248
<< error_p >>
rect -29 17 29 23
rect -29 -17 17 17
rect -29 -23 29 -17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -29 17 29 23
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -23 29 -17
<< properties >>
string GDS_END 504212
string GDS_FILE digital_filter_3a.gds
string GDS_START 504016
<< end >>
