magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< pwell >>
rect -455 -548 455 330
<< nmos >>
rect -255 -48 -225 52
rect -159 -48 -129 52
rect -63 -48 -33 52
rect 33 -48 63 52
rect 129 -48 159 52
rect 225 -48 255 52
rect -255 -270 -225 -170
rect -159 -270 -129 -170
rect -63 -270 -33 -170
rect 33 -270 63 -170
rect 129 -270 159 -170
rect 225 -270 255 -170
<< ndiff >>
rect -317 40 -255 52
rect -317 -36 -305 40
rect -271 -36 -255 40
rect -317 -48 -255 -36
rect -225 40 -159 52
rect -225 -36 -209 40
rect -175 -36 -159 40
rect -225 -48 -159 -36
rect -129 40 -63 52
rect -129 -36 -113 40
rect -79 -36 -63 40
rect -129 -48 -63 -36
rect -33 40 33 52
rect -33 -36 -17 40
rect 17 -36 33 40
rect -33 -48 33 -36
rect 63 40 129 52
rect 63 -36 79 40
rect 113 -36 129 40
rect 63 -48 129 -36
rect 159 40 225 52
rect 159 -36 175 40
rect 209 -36 225 40
rect 159 -48 225 -36
rect 255 40 317 52
rect 255 -36 271 40
rect 305 -36 317 40
rect 255 -48 317 -36
rect -317 -182 -255 -170
rect -317 -258 -305 -182
rect -271 -258 -255 -182
rect -317 -270 -255 -258
rect -225 -182 -159 -170
rect -225 -258 -209 -182
rect -175 -258 -159 -182
rect -225 -270 -159 -258
rect -129 -182 -63 -170
rect -129 -258 -113 -182
rect -79 -258 -63 -182
rect -129 -270 -63 -258
rect -33 -182 33 -170
rect -33 -258 -17 -182
rect 17 -258 33 -182
rect -33 -270 33 -258
rect 63 -182 129 -170
rect 63 -258 79 -182
rect 113 -258 129 -182
rect 63 -270 129 -258
rect 159 -182 225 -170
rect 159 -258 175 -182
rect 209 -258 225 -182
rect 159 -270 225 -258
rect 255 -182 317 -170
rect 255 -258 271 -182
rect 305 -258 317 -182
rect 255 -270 317 -258
<< ndiffc >>
rect -305 -36 -271 40
rect -209 -36 -175 40
rect -113 -36 -79 40
rect -17 -36 17 40
rect 79 -36 113 40
rect 175 -36 209 40
rect 271 -36 305 40
rect -305 -258 -271 -182
rect -209 -258 -175 -182
rect -113 -258 -79 -182
rect -17 -258 17 -182
rect 79 -258 113 -182
rect 175 -258 209 -182
rect 271 -258 305 -182
<< psubdiff >>
rect -419 260 -323 294
rect 323 260 419 294
rect -419 198 -385 260
rect 385 198 419 260
rect -419 -478 -385 -416
rect 385 -478 419 -416
rect -419 -512 -323 -478
rect 323 -512 419 -478
<< psubdiffcont >>
rect -323 260 323 294
rect -419 -416 -385 198
rect 385 -416 419 198
rect -323 -512 323 -478
<< poly >>
rect -63 192 63 208
rect -63 158 -17 192
rect 17 158 63 192
rect -63 142 63 158
rect -291 124 -225 140
rect -291 90 -275 124
rect -241 90 -225 124
rect -291 74 -225 90
rect -177 124 -111 140
rect -177 90 -161 124
rect -127 90 -111 124
rect -177 74 -111 90
rect -255 52 -225 74
rect -159 52 -129 74
rect -63 52 -33 142
rect 33 52 63 142
rect 111 124 177 140
rect 111 90 127 124
rect 161 90 177 124
rect 111 74 177 90
rect 225 124 291 140
rect 225 90 241 124
rect 275 90 291 124
rect 225 74 291 90
rect 129 52 159 74
rect 225 52 255 74
rect -255 -74 -225 -48
rect -159 -74 -129 -48
rect -63 -74 -33 -48
rect 33 -74 63 -48
rect 129 -74 159 -48
rect 225 -74 255 -48
rect -255 -170 -225 -144
rect -159 -170 -129 -144
rect -63 -170 -33 -144
rect 33 -170 63 -144
rect 129 -170 159 -144
rect 225 -170 255 -144
rect -255 -292 -225 -270
rect -159 -292 -129 -270
rect -291 -308 -225 -292
rect -291 -342 -275 -308
rect -241 -342 -225 -308
rect -291 -358 -225 -342
rect -177 -308 -111 -292
rect -177 -342 -161 -308
rect -127 -342 -111 -308
rect -177 -358 -111 -342
rect -63 -360 -33 -270
rect 33 -360 63 -270
rect 129 -292 159 -270
rect 225 -292 255 -270
rect 111 -308 177 -292
rect 111 -342 127 -308
rect 161 -342 177 -308
rect 111 -358 177 -342
rect 225 -308 291 -292
rect 225 -342 241 -308
rect 275 -342 291 -308
rect 225 -358 291 -342
rect -63 -376 63 -360
rect -63 -410 -17 -376
rect 17 -410 63 -376
rect -63 -426 63 -410
<< polycont >>
rect -17 158 17 192
rect -275 90 -241 124
rect -161 90 -127 124
rect 127 90 161 124
rect 241 90 275 124
rect -275 -342 -241 -308
rect -161 -342 -127 -308
rect 127 -342 161 -308
rect 241 -342 275 -308
rect -17 -410 17 -376
<< locali >>
rect -419 260 -323 294
rect 323 260 419 294
rect -419 198 -385 260
rect 385 198 419 260
rect -33 158 -17 192
rect 17 158 33 192
rect -385 90 -275 124
rect -241 90 -225 124
rect -177 90 -161 124
rect -127 90 -111 124
rect 111 90 127 124
rect 161 90 177 124
rect 225 90 241 124
rect 275 90 385 124
rect -305 40 -271 90
rect -305 -52 -271 -36
rect -209 48 -175 56
rect -209 -52 -175 -36
rect -113 40 -79 56
rect -113 -92 -79 -36
rect -17 40 17 56
rect 79 40 113 56
rect 79 -92 113 -36
rect 175 48 209 56
rect 175 -52 209 -36
rect 271 40 305 90
rect 271 -52 305 -36
rect -79 -126 79 -92
rect -305 -182 -271 -166
rect -305 -308 -271 -258
rect -209 -182 -175 -166
rect -209 -274 -175 -266
rect -113 -182 -79 -126
rect -113 -274 -79 -258
rect -17 -274 17 -258
rect 79 -182 113 -126
rect 79 -274 113 -258
rect 175 -182 209 -166
rect 175 -274 209 -266
rect 271 -182 305 -166
rect 271 -308 305 -258
rect -385 -342 -275 -308
rect -241 -342 -225 -308
rect -177 -342 -161 -308
rect -127 -342 -111 -308
rect 111 -342 127 -308
rect 161 -342 177 -308
rect 225 -342 241 -308
rect 275 -342 385 -308
rect -33 -410 -17 -376
rect 17 -410 33 -376
rect -419 -478 -385 -416
rect 385 -478 419 -416
rect -419 -512 -323 -478
rect 323 -512 419 -478
<< viali >>
rect -17 158 17 192
rect -161 90 -127 124
rect 127 90 161 124
rect -209 40 -175 48
rect -209 14 -175 40
rect -17 -36 17 -20
rect -17 -54 17 -36
rect 175 40 209 48
rect 175 14 209 40
rect -113 -126 -79 -92
rect 79 -126 113 -92
rect -209 -258 -175 -232
rect -209 -266 -175 -258
rect -17 -182 17 -164
rect -17 -198 17 -182
rect 175 -258 209 -232
rect 175 -266 209 -258
rect -161 -342 -127 -308
rect 127 -342 161 -308
rect -17 -410 17 -376
<< metal1 >>
rect -303 192 -293 210
rect -455 158 -293 192
rect -241 192 -231 210
rect -29 192 29 198
rect -241 158 -17 192
rect 17 158 63 192
rect -29 152 29 158
rect -173 124 -115 130
rect 115 124 173 130
rect 231 124 241 142
rect -177 90 -161 124
rect -127 90 127 124
rect 161 90 241 124
rect 293 124 303 142
rect 293 90 455 124
rect -173 84 -115 90
rect 115 84 173 90
rect -221 48 -163 54
rect 163 48 221 54
rect -221 14 -209 48
rect -175 14 175 48
rect 209 14 455 48
rect -221 8 -163 14
rect 163 8 221 14
rect -29 -20 29 -14
rect -455 -54 -17 -20
rect 17 -54 29 -20
rect -305 -232 -271 -54
rect -29 -60 29 -54
rect -133 -134 -123 -82
rect -71 -92 -61 -82
rect 61 -92 71 -82
rect -71 -126 71 -92
rect -71 -134 -61 -126
rect 61 -134 71 -126
rect 123 -134 133 -82
rect -29 -164 29 -158
rect 271 -164 305 14
rect -29 -198 -17 -164
rect 17 -198 305 -164
rect -29 -204 29 -198
rect -221 -232 -163 -226
rect 163 -232 221 -226
rect -305 -266 -209 -232
rect -175 -266 175 -232
rect 209 -266 271 -232
rect -221 -272 -163 -266
rect 163 -272 221 -266
rect -173 -308 -115 -302
rect 115 -308 173 -302
rect -303 -360 -293 -308
rect -241 -342 -161 -308
rect -127 -342 127 -308
rect 161 -342 177 -308
rect -241 -360 -231 -342
rect -173 -348 -115 -342
rect 115 -348 173 -342
rect -29 -376 29 -370
rect -63 -410 -17 -376
rect 17 -410 241 -376
rect -29 -416 29 -410
rect 231 -428 241 -410
rect 293 -428 303 -376
<< via1 >>
rect -293 158 -241 210
rect 241 90 293 142
rect -123 -92 -71 -82
rect 71 -92 123 -82
rect -123 -126 -113 -92
rect -113 -126 -79 -92
rect -79 -126 -71 -92
rect 71 -126 79 -92
rect 79 -126 113 -92
rect 113 -126 123 -92
rect -123 -134 -71 -126
rect 71 -134 123 -126
rect -293 -360 -241 -308
rect 241 -428 293 -376
<< metal2 >>
rect -293 210 -241 220
rect -293 -308 -241 158
rect 241 142 293 152
rect -129 -134 -123 -82
rect -71 -134 71 -82
rect 123 -134 129 -82
rect -293 -370 -241 -360
rect -27 -512 27 -134
rect 241 -376 293 90
rect 241 -438 293 -428
<< properties >>
string FIXED_BBOX -402 -206 402 206
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
