magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< nwell >>
rect -2112 -240 2112 240
<< pmos >>
rect -2018 -140 -1898 140
rect -1840 -140 -1720 140
rect -1662 -140 -1542 140
rect -1484 -140 -1364 140
rect -1306 -140 -1186 140
rect -1128 -140 -1008 140
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
rect 1008 -140 1128 140
rect 1186 -140 1306 140
rect 1364 -140 1484 140
rect 1542 -140 1662 140
rect 1720 -140 1840 140
rect 1898 -140 2018 140
<< pdiff >>
rect -2076 119 -2018 140
rect -2076 85 -2064 119
rect -2030 85 -2018 119
rect -2076 51 -2018 85
rect -2076 17 -2064 51
rect -2030 17 -2018 51
rect -2076 -17 -2018 17
rect -2076 -51 -2064 -17
rect -2030 -51 -2018 -17
rect -2076 -85 -2018 -51
rect -2076 -119 -2064 -85
rect -2030 -119 -2018 -85
rect -2076 -140 -2018 -119
rect -1898 119 -1840 140
rect -1898 85 -1886 119
rect -1852 85 -1840 119
rect -1898 51 -1840 85
rect -1898 17 -1886 51
rect -1852 17 -1840 51
rect -1898 -17 -1840 17
rect -1898 -51 -1886 -17
rect -1852 -51 -1840 -17
rect -1898 -85 -1840 -51
rect -1898 -119 -1886 -85
rect -1852 -119 -1840 -85
rect -1898 -140 -1840 -119
rect -1720 119 -1662 140
rect -1720 85 -1708 119
rect -1674 85 -1662 119
rect -1720 51 -1662 85
rect -1720 17 -1708 51
rect -1674 17 -1662 51
rect -1720 -17 -1662 17
rect -1720 -51 -1708 -17
rect -1674 -51 -1662 -17
rect -1720 -85 -1662 -51
rect -1720 -119 -1708 -85
rect -1674 -119 -1662 -85
rect -1720 -140 -1662 -119
rect -1542 119 -1484 140
rect -1542 85 -1530 119
rect -1496 85 -1484 119
rect -1542 51 -1484 85
rect -1542 17 -1530 51
rect -1496 17 -1484 51
rect -1542 -17 -1484 17
rect -1542 -51 -1530 -17
rect -1496 -51 -1484 -17
rect -1542 -85 -1484 -51
rect -1542 -119 -1530 -85
rect -1496 -119 -1484 -85
rect -1542 -140 -1484 -119
rect -1364 119 -1306 140
rect -1364 85 -1352 119
rect -1318 85 -1306 119
rect -1364 51 -1306 85
rect -1364 17 -1352 51
rect -1318 17 -1306 51
rect -1364 -17 -1306 17
rect -1364 -51 -1352 -17
rect -1318 -51 -1306 -17
rect -1364 -85 -1306 -51
rect -1364 -119 -1352 -85
rect -1318 -119 -1306 -85
rect -1364 -140 -1306 -119
rect -1186 119 -1128 140
rect -1186 85 -1174 119
rect -1140 85 -1128 119
rect -1186 51 -1128 85
rect -1186 17 -1174 51
rect -1140 17 -1128 51
rect -1186 -17 -1128 17
rect -1186 -51 -1174 -17
rect -1140 -51 -1128 -17
rect -1186 -85 -1128 -51
rect -1186 -119 -1174 -85
rect -1140 -119 -1128 -85
rect -1186 -140 -1128 -119
rect -1008 119 -950 140
rect -1008 85 -996 119
rect -962 85 -950 119
rect -1008 51 -950 85
rect -1008 17 -996 51
rect -962 17 -950 51
rect -1008 -17 -950 17
rect -1008 -51 -996 -17
rect -962 -51 -950 -17
rect -1008 -85 -950 -51
rect -1008 -119 -996 -85
rect -962 -119 -950 -85
rect -1008 -140 -950 -119
rect -830 119 -772 140
rect -830 85 -818 119
rect -784 85 -772 119
rect -830 51 -772 85
rect -830 17 -818 51
rect -784 17 -772 51
rect -830 -17 -772 17
rect -830 -51 -818 -17
rect -784 -51 -772 -17
rect -830 -85 -772 -51
rect -830 -119 -818 -85
rect -784 -119 -772 -85
rect -830 -140 -772 -119
rect -652 119 -594 140
rect -652 85 -640 119
rect -606 85 -594 119
rect -652 51 -594 85
rect -652 17 -640 51
rect -606 17 -594 51
rect -652 -17 -594 17
rect -652 -51 -640 -17
rect -606 -51 -594 -17
rect -652 -85 -594 -51
rect -652 -119 -640 -85
rect -606 -119 -594 -85
rect -652 -140 -594 -119
rect -474 119 -416 140
rect -474 85 -462 119
rect -428 85 -416 119
rect -474 51 -416 85
rect -474 17 -462 51
rect -428 17 -416 51
rect -474 -17 -416 17
rect -474 -51 -462 -17
rect -428 -51 -416 -17
rect -474 -85 -416 -51
rect -474 -119 -462 -85
rect -428 -119 -416 -85
rect -474 -140 -416 -119
rect -296 119 -238 140
rect -296 85 -284 119
rect -250 85 -238 119
rect -296 51 -238 85
rect -296 17 -284 51
rect -250 17 -238 51
rect -296 -17 -238 17
rect -296 -51 -284 -17
rect -250 -51 -238 -17
rect -296 -85 -238 -51
rect -296 -119 -284 -85
rect -250 -119 -238 -85
rect -296 -140 -238 -119
rect -118 119 -60 140
rect -118 85 -106 119
rect -72 85 -60 119
rect -118 51 -60 85
rect -118 17 -106 51
rect -72 17 -60 51
rect -118 -17 -60 17
rect -118 -51 -106 -17
rect -72 -51 -60 -17
rect -118 -85 -60 -51
rect -118 -119 -106 -85
rect -72 -119 -60 -85
rect -118 -140 -60 -119
rect 60 119 118 140
rect 60 85 72 119
rect 106 85 118 119
rect 60 51 118 85
rect 60 17 72 51
rect 106 17 118 51
rect 60 -17 118 17
rect 60 -51 72 -17
rect 106 -51 118 -17
rect 60 -85 118 -51
rect 60 -119 72 -85
rect 106 -119 118 -85
rect 60 -140 118 -119
rect 238 119 296 140
rect 238 85 250 119
rect 284 85 296 119
rect 238 51 296 85
rect 238 17 250 51
rect 284 17 296 51
rect 238 -17 296 17
rect 238 -51 250 -17
rect 284 -51 296 -17
rect 238 -85 296 -51
rect 238 -119 250 -85
rect 284 -119 296 -85
rect 238 -140 296 -119
rect 416 119 474 140
rect 416 85 428 119
rect 462 85 474 119
rect 416 51 474 85
rect 416 17 428 51
rect 462 17 474 51
rect 416 -17 474 17
rect 416 -51 428 -17
rect 462 -51 474 -17
rect 416 -85 474 -51
rect 416 -119 428 -85
rect 462 -119 474 -85
rect 416 -140 474 -119
rect 594 119 652 140
rect 594 85 606 119
rect 640 85 652 119
rect 594 51 652 85
rect 594 17 606 51
rect 640 17 652 51
rect 594 -17 652 17
rect 594 -51 606 -17
rect 640 -51 652 -17
rect 594 -85 652 -51
rect 594 -119 606 -85
rect 640 -119 652 -85
rect 594 -140 652 -119
rect 772 119 830 140
rect 772 85 784 119
rect 818 85 830 119
rect 772 51 830 85
rect 772 17 784 51
rect 818 17 830 51
rect 772 -17 830 17
rect 772 -51 784 -17
rect 818 -51 830 -17
rect 772 -85 830 -51
rect 772 -119 784 -85
rect 818 -119 830 -85
rect 772 -140 830 -119
rect 950 119 1008 140
rect 950 85 962 119
rect 996 85 1008 119
rect 950 51 1008 85
rect 950 17 962 51
rect 996 17 1008 51
rect 950 -17 1008 17
rect 950 -51 962 -17
rect 996 -51 1008 -17
rect 950 -85 1008 -51
rect 950 -119 962 -85
rect 996 -119 1008 -85
rect 950 -140 1008 -119
rect 1128 119 1186 140
rect 1128 85 1140 119
rect 1174 85 1186 119
rect 1128 51 1186 85
rect 1128 17 1140 51
rect 1174 17 1186 51
rect 1128 -17 1186 17
rect 1128 -51 1140 -17
rect 1174 -51 1186 -17
rect 1128 -85 1186 -51
rect 1128 -119 1140 -85
rect 1174 -119 1186 -85
rect 1128 -140 1186 -119
rect 1306 119 1364 140
rect 1306 85 1318 119
rect 1352 85 1364 119
rect 1306 51 1364 85
rect 1306 17 1318 51
rect 1352 17 1364 51
rect 1306 -17 1364 17
rect 1306 -51 1318 -17
rect 1352 -51 1364 -17
rect 1306 -85 1364 -51
rect 1306 -119 1318 -85
rect 1352 -119 1364 -85
rect 1306 -140 1364 -119
rect 1484 119 1542 140
rect 1484 85 1496 119
rect 1530 85 1542 119
rect 1484 51 1542 85
rect 1484 17 1496 51
rect 1530 17 1542 51
rect 1484 -17 1542 17
rect 1484 -51 1496 -17
rect 1530 -51 1542 -17
rect 1484 -85 1542 -51
rect 1484 -119 1496 -85
rect 1530 -119 1542 -85
rect 1484 -140 1542 -119
rect 1662 119 1720 140
rect 1662 85 1674 119
rect 1708 85 1720 119
rect 1662 51 1720 85
rect 1662 17 1674 51
rect 1708 17 1720 51
rect 1662 -17 1720 17
rect 1662 -51 1674 -17
rect 1708 -51 1720 -17
rect 1662 -85 1720 -51
rect 1662 -119 1674 -85
rect 1708 -119 1720 -85
rect 1662 -140 1720 -119
rect 1840 119 1898 140
rect 1840 85 1852 119
rect 1886 85 1898 119
rect 1840 51 1898 85
rect 1840 17 1852 51
rect 1886 17 1898 51
rect 1840 -17 1898 17
rect 1840 -51 1852 -17
rect 1886 -51 1898 -17
rect 1840 -85 1898 -51
rect 1840 -119 1852 -85
rect 1886 -119 1898 -85
rect 1840 -140 1898 -119
rect 2018 119 2076 140
rect 2018 85 2030 119
rect 2064 85 2076 119
rect 2018 51 2076 85
rect 2018 17 2030 51
rect 2064 17 2076 51
rect 2018 -17 2076 17
rect 2018 -51 2030 -17
rect 2064 -51 2076 -17
rect 2018 -85 2076 -51
rect 2018 -119 2030 -85
rect 2064 -119 2076 -85
rect 2018 -140 2076 -119
<< pdiffc >>
rect -2064 85 -2030 119
rect -2064 17 -2030 51
rect -2064 -51 -2030 -17
rect -2064 -119 -2030 -85
rect -1886 85 -1852 119
rect -1886 17 -1852 51
rect -1886 -51 -1852 -17
rect -1886 -119 -1852 -85
rect -1708 85 -1674 119
rect -1708 17 -1674 51
rect -1708 -51 -1674 -17
rect -1708 -119 -1674 -85
rect -1530 85 -1496 119
rect -1530 17 -1496 51
rect -1530 -51 -1496 -17
rect -1530 -119 -1496 -85
rect -1352 85 -1318 119
rect -1352 17 -1318 51
rect -1352 -51 -1318 -17
rect -1352 -119 -1318 -85
rect -1174 85 -1140 119
rect -1174 17 -1140 51
rect -1174 -51 -1140 -17
rect -1174 -119 -1140 -85
rect -996 85 -962 119
rect -996 17 -962 51
rect -996 -51 -962 -17
rect -996 -119 -962 -85
rect -818 85 -784 119
rect -818 17 -784 51
rect -818 -51 -784 -17
rect -818 -119 -784 -85
rect -640 85 -606 119
rect -640 17 -606 51
rect -640 -51 -606 -17
rect -640 -119 -606 -85
rect -462 85 -428 119
rect -462 17 -428 51
rect -462 -51 -428 -17
rect -462 -119 -428 -85
rect -284 85 -250 119
rect -284 17 -250 51
rect -284 -51 -250 -17
rect -284 -119 -250 -85
rect -106 85 -72 119
rect -106 17 -72 51
rect -106 -51 -72 -17
rect -106 -119 -72 -85
rect 72 85 106 119
rect 72 17 106 51
rect 72 -51 106 -17
rect 72 -119 106 -85
rect 250 85 284 119
rect 250 17 284 51
rect 250 -51 284 -17
rect 250 -119 284 -85
rect 428 85 462 119
rect 428 17 462 51
rect 428 -51 462 -17
rect 428 -119 462 -85
rect 606 85 640 119
rect 606 17 640 51
rect 606 -51 640 -17
rect 606 -119 640 -85
rect 784 85 818 119
rect 784 17 818 51
rect 784 -51 818 -17
rect 784 -119 818 -85
rect 962 85 996 119
rect 962 17 996 51
rect 962 -51 996 -17
rect 962 -119 996 -85
rect 1140 85 1174 119
rect 1140 17 1174 51
rect 1140 -51 1174 -17
rect 1140 -119 1174 -85
rect 1318 85 1352 119
rect 1318 17 1352 51
rect 1318 -51 1352 -17
rect 1318 -119 1352 -85
rect 1496 85 1530 119
rect 1496 17 1530 51
rect 1496 -51 1530 -17
rect 1496 -119 1530 -85
rect 1674 85 1708 119
rect 1674 17 1708 51
rect 1674 -51 1708 -17
rect 1674 -119 1708 -85
rect 1852 85 1886 119
rect 1852 17 1886 51
rect 1852 -51 1886 -17
rect 1852 -119 1886 -85
rect 2030 85 2064 119
rect 2030 17 2064 51
rect 2030 -51 2064 -17
rect 2030 -119 2064 -85
<< poly >>
rect -1996 221 -1920 237
rect -1996 205 -1975 221
rect -2018 187 -1975 205
rect -1941 205 -1920 221
rect -1818 221 -1742 237
rect -1818 205 -1797 221
rect -1941 187 -1898 205
rect -2018 140 -1898 187
rect -1840 187 -1797 205
rect -1763 205 -1742 221
rect -1640 221 -1564 237
rect -1640 205 -1619 221
rect -1763 187 -1720 205
rect -1840 140 -1720 187
rect -1662 187 -1619 205
rect -1585 205 -1564 221
rect -1462 221 -1386 237
rect -1462 205 -1441 221
rect -1585 187 -1542 205
rect -1662 140 -1542 187
rect -1484 187 -1441 205
rect -1407 205 -1386 221
rect -1284 221 -1208 237
rect -1284 205 -1263 221
rect -1407 187 -1364 205
rect -1484 140 -1364 187
rect -1306 187 -1263 205
rect -1229 205 -1208 221
rect -1106 221 -1030 237
rect -1106 205 -1085 221
rect -1229 187 -1186 205
rect -1306 140 -1186 187
rect -1128 187 -1085 205
rect -1051 205 -1030 221
rect -928 221 -852 237
rect -928 205 -907 221
rect -1051 187 -1008 205
rect -1128 140 -1008 187
rect -950 187 -907 205
rect -873 205 -852 221
rect -750 221 -674 237
rect -750 205 -729 221
rect -873 187 -830 205
rect -950 140 -830 187
rect -772 187 -729 205
rect -695 205 -674 221
rect -572 221 -496 237
rect -572 205 -551 221
rect -695 187 -652 205
rect -772 140 -652 187
rect -594 187 -551 205
rect -517 205 -496 221
rect -394 221 -318 237
rect -394 205 -373 221
rect -517 187 -474 205
rect -594 140 -474 187
rect -416 187 -373 205
rect -339 205 -318 221
rect -216 221 -140 237
rect -216 205 -195 221
rect -339 187 -296 205
rect -416 140 -296 187
rect -238 187 -195 205
rect -161 205 -140 221
rect -38 221 38 237
rect -38 205 -17 221
rect -161 187 -118 205
rect -238 140 -118 187
rect -60 187 -17 205
rect 17 205 38 221
rect 140 221 216 237
rect 140 205 161 221
rect 17 187 60 205
rect -60 140 60 187
rect 118 187 161 205
rect 195 205 216 221
rect 318 221 394 237
rect 318 205 339 221
rect 195 187 238 205
rect 118 140 238 187
rect 296 187 339 205
rect 373 205 394 221
rect 496 221 572 237
rect 496 205 517 221
rect 373 187 416 205
rect 296 140 416 187
rect 474 187 517 205
rect 551 205 572 221
rect 674 221 750 237
rect 674 205 695 221
rect 551 187 594 205
rect 474 140 594 187
rect 652 187 695 205
rect 729 205 750 221
rect 852 221 928 237
rect 852 205 873 221
rect 729 187 772 205
rect 652 140 772 187
rect 830 187 873 205
rect 907 205 928 221
rect 1030 221 1106 237
rect 1030 205 1051 221
rect 907 187 950 205
rect 830 140 950 187
rect 1008 187 1051 205
rect 1085 205 1106 221
rect 1208 221 1284 237
rect 1208 205 1229 221
rect 1085 187 1128 205
rect 1008 140 1128 187
rect 1186 187 1229 205
rect 1263 205 1284 221
rect 1386 221 1462 237
rect 1386 205 1407 221
rect 1263 187 1306 205
rect 1186 140 1306 187
rect 1364 187 1407 205
rect 1441 205 1462 221
rect 1564 221 1640 237
rect 1564 205 1585 221
rect 1441 187 1484 205
rect 1364 140 1484 187
rect 1542 187 1585 205
rect 1619 205 1640 221
rect 1742 221 1818 237
rect 1742 205 1763 221
rect 1619 187 1662 205
rect 1542 140 1662 187
rect 1720 187 1763 205
rect 1797 205 1818 221
rect 1920 221 1996 237
rect 1920 205 1941 221
rect 1797 187 1840 205
rect 1720 140 1840 187
rect 1898 187 1941 205
rect 1975 205 1996 221
rect 1975 187 2018 205
rect 1898 140 2018 187
rect -2018 -187 -1898 -140
rect -2018 -205 -1975 -187
rect -1996 -221 -1975 -205
rect -1941 -205 -1898 -187
rect -1840 -187 -1720 -140
rect -1840 -205 -1797 -187
rect -1941 -221 -1920 -205
rect -1996 -237 -1920 -221
rect -1818 -221 -1797 -205
rect -1763 -205 -1720 -187
rect -1662 -187 -1542 -140
rect -1662 -205 -1619 -187
rect -1763 -221 -1742 -205
rect -1818 -237 -1742 -221
rect -1640 -221 -1619 -205
rect -1585 -205 -1542 -187
rect -1484 -187 -1364 -140
rect -1484 -205 -1441 -187
rect -1585 -221 -1564 -205
rect -1640 -237 -1564 -221
rect -1462 -221 -1441 -205
rect -1407 -205 -1364 -187
rect -1306 -187 -1186 -140
rect -1306 -205 -1263 -187
rect -1407 -221 -1386 -205
rect -1462 -237 -1386 -221
rect -1284 -221 -1263 -205
rect -1229 -205 -1186 -187
rect -1128 -187 -1008 -140
rect -1128 -205 -1085 -187
rect -1229 -221 -1208 -205
rect -1284 -237 -1208 -221
rect -1106 -221 -1085 -205
rect -1051 -205 -1008 -187
rect -950 -187 -830 -140
rect -950 -205 -907 -187
rect -1051 -221 -1030 -205
rect -1106 -237 -1030 -221
rect -928 -221 -907 -205
rect -873 -205 -830 -187
rect -772 -187 -652 -140
rect -772 -205 -729 -187
rect -873 -221 -852 -205
rect -928 -237 -852 -221
rect -750 -221 -729 -205
rect -695 -205 -652 -187
rect -594 -187 -474 -140
rect -594 -205 -551 -187
rect -695 -221 -674 -205
rect -750 -237 -674 -221
rect -572 -221 -551 -205
rect -517 -205 -474 -187
rect -416 -187 -296 -140
rect -416 -205 -373 -187
rect -517 -221 -496 -205
rect -572 -237 -496 -221
rect -394 -221 -373 -205
rect -339 -205 -296 -187
rect -238 -187 -118 -140
rect -238 -205 -195 -187
rect -339 -221 -318 -205
rect -394 -237 -318 -221
rect -216 -221 -195 -205
rect -161 -205 -118 -187
rect -60 -187 60 -140
rect -60 -205 -17 -187
rect -161 -221 -140 -205
rect -216 -237 -140 -221
rect -38 -221 -17 -205
rect 17 -205 60 -187
rect 118 -187 238 -140
rect 118 -205 161 -187
rect 17 -221 38 -205
rect -38 -237 38 -221
rect 140 -221 161 -205
rect 195 -205 238 -187
rect 296 -187 416 -140
rect 296 -205 339 -187
rect 195 -221 216 -205
rect 140 -237 216 -221
rect 318 -221 339 -205
rect 373 -205 416 -187
rect 474 -187 594 -140
rect 474 -205 517 -187
rect 373 -221 394 -205
rect 318 -237 394 -221
rect 496 -221 517 -205
rect 551 -205 594 -187
rect 652 -187 772 -140
rect 652 -205 695 -187
rect 551 -221 572 -205
rect 496 -237 572 -221
rect 674 -221 695 -205
rect 729 -205 772 -187
rect 830 -187 950 -140
rect 830 -205 873 -187
rect 729 -221 750 -205
rect 674 -237 750 -221
rect 852 -221 873 -205
rect 907 -205 950 -187
rect 1008 -187 1128 -140
rect 1008 -205 1051 -187
rect 907 -221 928 -205
rect 852 -237 928 -221
rect 1030 -221 1051 -205
rect 1085 -205 1128 -187
rect 1186 -187 1306 -140
rect 1186 -205 1229 -187
rect 1085 -221 1106 -205
rect 1030 -237 1106 -221
rect 1208 -221 1229 -205
rect 1263 -205 1306 -187
rect 1364 -187 1484 -140
rect 1364 -205 1407 -187
rect 1263 -221 1284 -205
rect 1208 -237 1284 -221
rect 1386 -221 1407 -205
rect 1441 -205 1484 -187
rect 1542 -187 1662 -140
rect 1542 -205 1585 -187
rect 1441 -221 1462 -205
rect 1386 -237 1462 -221
rect 1564 -221 1585 -205
rect 1619 -205 1662 -187
rect 1720 -187 1840 -140
rect 1720 -205 1763 -187
rect 1619 -221 1640 -205
rect 1564 -237 1640 -221
rect 1742 -221 1763 -205
rect 1797 -205 1840 -187
rect 1898 -187 2018 -140
rect 1898 -205 1941 -187
rect 1797 -221 1818 -205
rect 1742 -237 1818 -221
rect 1920 -221 1941 -205
rect 1975 -205 2018 -187
rect 1975 -221 1996 -205
rect 1920 -237 1996 -221
<< polycont >>
rect -1975 187 -1941 221
rect -1797 187 -1763 221
rect -1619 187 -1585 221
rect -1441 187 -1407 221
rect -1263 187 -1229 221
rect -1085 187 -1051 221
rect -907 187 -873 221
rect -729 187 -695 221
rect -551 187 -517 221
rect -373 187 -339 221
rect -195 187 -161 221
rect -17 187 17 221
rect 161 187 195 221
rect 339 187 373 221
rect 517 187 551 221
rect 695 187 729 221
rect 873 187 907 221
rect 1051 187 1085 221
rect 1229 187 1263 221
rect 1407 187 1441 221
rect 1585 187 1619 221
rect 1763 187 1797 221
rect 1941 187 1975 221
rect -1975 -221 -1941 -187
rect -1797 -221 -1763 -187
rect -1619 -221 -1585 -187
rect -1441 -221 -1407 -187
rect -1263 -221 -1229 -187
rect -1085 -221 -1051 -187
rect -907 -221 -873 -187
rect -729 -221 -695 -187
rect -551 -221 -517 -187
rect -373 -221 -339 -187
rect -195 -221 -161 -187
rect -17 -221 17 -187
rect 161 -221 195 -187
rect 339 -221 373 -187
rect 517 -221 551 -187
rect 695 -221 729 -187
rect 873 -221 907 -187
rect 1051 -221 1085 -187
rect 1229 -221 1263 -187
rect 1407 -221 1441 -187
rect 1585 -221 1619 -187
rect 1763 -221 1797 -187
rect 1941 -221 1975 -187
<< locali >>
rect -1996 187 -1975 221
rect -1941 187 -1920 221
rect -1818 187 -1797 221
rect -1763 187 -1742 221
rect -1640 187 -1619 221
rect -1585 187 -1564 221
rect -1462 187 -1441 221
rect -1407 187 -1386 221
rect -1284 187 -1263 221
rect -1229 187 -1208 221
rect -1106 187 -1085 221
rect -1051 187 -1030 221
rect -928 187 -907 221
rect -873 187 -852 221
rect -750 187 -729 221
rect -695 187 -674 221
rect -572 187 -551 221
rect -517 187 -496 221
rect -394 187 -373 221
rect -339 187 -318 221
rect -216 187 -195 221
rect -161 187 -140 221
rect -38 187 -17 221
rect 17 187 38 221
rect 140 187 161 221
rect 195 187 216 221
rect 318 187 339 221
rect 373 187 394 221
rect 496 187 517 221
rect 551 187 572 221
rect 674 187 695 221
rect 729 187 750 221
rect 852 187 873 221
rect 907 187 928 221
rect 1030 187 1051 221
rect 1085 187 1106 221
rect 1208 187 1229 221
rect 1263 187 1284 221
rect 1386 187 1407 221
rect 1441 187 1462 221
rect 1564 187 1585 221
rect 1619 187 1640 221
rect 1742 187 1763 221
rect 1797 187 1818 221
rect 1920 187 1941 221
rect 1975 187 1996 221
rect -2064 125 -2030 144
rect -2064 53 -2030 85
rect -2064 -17 -2030 17
rect -2064 -85 -2030 -53
rect -2064 -144 -2030 -125
rect -1886 125 -1852 144
rect -1886 53 -1852 85
rect -1886 -17 -1852 17
rect -1886 -85 -1852 -53
rect -1886 -144 -1852 -125
rect -1708 125 -1674 144
rect -1708 53 -1674 85
rect -1708 -17 -1674 17
rect -1708 -85 -1674 -53
rect -1708 -144 -1674 -125
rect -1530 125 -1496 144
rect -1530 53 -1496 85
rect -1530 -17 -1496 17
rect -1530 -85 -1496 -53
rect -1530 -144 -1496 -125
rect -1352 125 -1318 144
rect -1352 53 -1318 85
rect -1352 -17 -1318 17
rect -1352 -85 -1318 -53
rect -1352 -144 -1318 -125
rect -1174 125 -1140 144
rect -1174 53 -1140 85
rect -1174 -17 -1140 17
rect -1174 -85 -1140 -53
rect -1174 -144 -1140 -125
rect -996 125 -962 144
rect -996 53 -962 85
rect -996 -17 -962 17
rect -996 -85 -962 -53
rect -996 -144 -962 -125
rect -818 125 -784 144
rect -818 53 -784 85
rect -818 -17 -784 17
rect -818 -85 -784 -53
rect -818 -144 -784 -125
rect -640 125 -606 144
rect -640 53 -606 85
rect -640 -17 -606 17
rect -640 -85 -606 -53
rect -640 -144 -606 -125
rect -462 125 -428 144
rect -462 53 -428 85
rect -462 -17 -428 17
rect -462 -85 -428 -53
rect -462 -144 -428 -125
rect -284 125 -250 144
rect -284 53 -250 85
rect -284 -17 -250 17
rect -284 -85 -250 -53
rect -284 -144 -250 -125
rect -106 125 -72 144
rect -106 53 -72 85
rect -106 -17 -72 17
rect -106 -85 -72 -53
rect -106 -144 -72 -125
rect 72 125 106 144
rect 72 53 106 85
rect 72 -17 106 17
rect 72 -85 106 -53
rect 72 -144 106 -125
rect 250 125 284 144
rect 250 53 284 85
rect 250 -17 284 17
rect 250 -85 284 -53
rect 250 -144 284 -125
rect 428 125 462 144
rect 428 53 462 85
rect 428 -17 462 17
rect 428 -85 462 -53
rect 428 -144 462 -125
rect 606 125 640 144
rect 606 53 640 85
rect 606 -17 640 17
rect 606 -85 640 -53
rect 606 -144 640 -125
rect 784 125 818 144
rect 784 53 818 85
rect 784 -17 818 17
rect 784 -85 818 -53
rect 784 -144 818 -125
rect 962 125 996 144
rect 962 53 996 85
rect 962 -17 996 17
rect 962 -85 996 -53
rect 962 -144 996 -125
rect 1140 125 1174 144
rect 1140 53 1174 85
rect 1140 -17 1174 17
rect 1140 -85 1174 -53
rect 1140 -144 1174 -125
rect 1318 125 1352 144
rect 1318 53 1352 85
rect 1318 -17 1352 17
rect 1318 -85 1352 -53
rect 1318 -144 1352 -125
rect 1496 125 1530 144
rect 1496 53 1530 85
rect 1496 -17 1530 17
rect 1496 -85 1530 -53
rect 1496 -144 1530 -125
rect 1674 125 1708 144
rect 1674 53 1708 85
rect 1674 -17 1708 17
rect 1674 -85 1708 -53
rect 1674 -144 1708 -125
rect 1852 125 1886 144
rect 1852 53 1886 85
rect 1852 -17 1886 17
rect 1852 -85 1886 -53
rect 1852 -144 1886 -125
rect 2030 125 2064 144
rect 2030 53 2064 85
rect 2030 -17 2064 17
rect 2030 -85 2064 -53
rect 2030 -144 2064 -125
rect -1996 -221 -1975 -187
rect -1941 -221 -1920 -187
rect -1818 -221 -1797 -187
rect -1763 -221 -1742 -187
rect -1640 -221 -1619 -187
rect -1585 -221 -1564 -187
rect -1462 -221 -1441 -187
rect -1407 -221 -1386 -187
rect -1284 -221 -1263 -187
rect -1229 -221 -1208 -187
rect -1106 -221 -1085 -187
rect -1051 -221 -1030 -187
rect -928 -221 -907 -187
rect -873 -221 -852 -187
rect -750 -221 -729 -187
rect -695 -221 -674 -187
rect -572 -221 -551 -187
rect -517 -221 -496 -187
rect -394 -221 -373 -187
rect -339 -221 -318 -187
rect -216 -221 -195 -187
rect -161 -221 -140 -187
rect -38 -221 -17 -187
rect 17 -221 38 -187
rect 140 -221 161 -187
rect 195 -221 216 -187
rect 318 -221 339 -187
rect 373 -221 394 -187
rect 496 -221 517 -187
rect 551 -221 572 -187
rect 674 -221 695 -187
rect 729 -221 750 -187
rect 852 -221 873 -187
rect 907 -221 928 -187
rect 1030 -221 1051 -187
rect 1085 -221 1106 -187
rect 1208 -221 1229 -187
rect 1263 -221 1284 -187
rect 1386 -221 1407 -187
rect 1441 -221 1462 -187
rect 1564 -221 1585 -187
rect 1619 -221 1640 -187
rect 1742 -221 1763 -187
rect 1797 -221 1818 -187
rect 1920 -221 1941 -187
rect 1975 -221 1996 -187
<< viali >>
rect -1975 187 -1941 221
rect -1797 187 -1763 221
rect -1619 187 -1585 221
rect -1441 187 -1407 221
rect -1263 187 -1229 221
rect -1085 187 -1051 221
rect -907 187 -873 221
rect -729 187 -695 221
rect -551 187 -517 221
rect -373 187 -339 221
rect -195 187 -161 221
rect -17 187 17 221
rect 161 187 195 221
rect 339 187 373 221
rect 517 187 551 221
rect 695 187 729 221
rect 873 187 907 221
rect 1051 187 1085 221
rect 1229 187 1263 221
rect 1407 187 1441 221
rect 1585 187 1619 221
rect 1763 187 1797 221
rect 1941 187 1975 221
rect -2064 119 -2030 125
rect -2064 91 -2030 119
rect -2064 51 -2030 53
rect -2064 19 -2030 51
rect -2064 -51 -2030 -19
rect -2064 -53 -2030 -51
rect -2064 -119 -2030 -91
rect -2064 -125 -2030 -119
rect -1886 119 -1852 125
rect -1886 91 -1852 119
rect -1886 51 -1852 53
rect -1886 19 -1852 51
rect -1886 -51 -1852 -19
rect -1886 -53 -1852 -51
rect -1886 -119 -1852 -91
rect -1886 -125 -1852 -119
rect -1708 119 -1674 125
rect -1708 91 -1674 119
rect -1708 51 -1674 53
rect -1708 19 -1674 51
rect -1708 -51 -1674 -19
rect -1708 -53 -1674 -51
rect -1708 -119 -1674 -91
rect -1708 -125 -1674 -119
rect -1530 119 -1496 125
rect -1530 91 -1496 119
rect -1530 51 -1496 53
rect -1530 19 -1496 51
rect -1530 -51 -1496 -19
rect -1530 -53 -1496 -51
rect -1530 -119 -1496 -91
rect -1530 -125 -1496 -119
rect -1352 119 -1318 125
rect -1352 91 -1318 119
rect -1352 51 -1318 53
rect -1352 19 -1318 51
rect -1352 -51 -1318 -19
rect -1352 -53 -1318 -51
rect -1352 -119 -1318 -91
rect -1352 -125 -1318 -119
rect -1174 119 -1140 125
rect -1174 91 -1140 119
rect -1174 51 -1140 53
rect -1174 19 -1140 51
rect -1174 -51 -1140 -19
rect -1174 -53 -1140 -51
rect -1174 -119 -1140 -91
rect -1174 -125 -1140 -119
rect -996 119 -962 125
rect -996 91 -962 119
rect -996 51 -962 53
rect -996 19 -962 51
rect -996 -51 -962 -19
rect -996 -53 -962 -51
rect -996 -119 -962 -91
rect -996 -125 -962 -119
rect -818 119 -784 125
rect -818 91 -784 119
rect -818 51 -784 53
rect -818 19 -784 51
rect -818 -51 -784 -19
rect -818 -53 -784 -51
rect -818 -119 -784 -91
rect -818 -125 -784 -119
rect -640 119 -606 125
rect -640 91 -606 119
rect -640 51 -606 53
rect -640 19 -606 51
rect -640 -51 -606 -19
rect -640 -53 -606 -51
rect -640 -119 -606 -91
rect -640 -125 -606 -119
rect -462 119 -428 125
rect -462 91 -428 119
rect -462 51 -428 53
rect -462 19 -428 51
rect -462 -51 -428 -19
rect -462 -53 -428 -51
rect -462 -119 -428 -91
rect -462 -125 -428 -119
rect -284 119 -250 125
rect -284 91 -250 119
rect -284 51 -250 53
rect -284 19 -250 51
rect -284 -51 -250 -19
rect -284 -53 -250 -51
rect -284 -119 -250 -91
rect -284 -125 -250 -119
rect -106 119 -72 125
rect -106 91 -72 119
rect -106 51 -72 53
rect -106 19 -72 51
rect -106 -51 -72 -19
rect -106 -53 -72 -51
rect -106 -119 -72 -91
rect -106 -125 -72 -119
rect 72 119 106 125
rect 72 91 106 119
rect 72 51 106 53
rect 72 19 106 51
rect 72 -51 106 -19
rect 72 -53 106 -51
rect 72 -119 106 -91
rect 72 -125 106 -119
rect 250 119 284 125
rect 250 91 284 119
rect 250 51 284 53
rect 250 19 284 51
rect 250 -51 284 -19
rect 250 -53 284 -51
rect 250 -119 284 -91
rect 250 -125 284 -119
rect 428 119 462 125
rect 428 91 462 119
rect 428 51 462 53
rect 428 19 462 51
rect 428 -51 462 -19
rect 428 -53 462 -51
rect 428 -119 462 -91
rect 428 -125 462 -119
rect 606 119 640 125
rect 606 91 640 119
rect 606 51 640 53
rect 606 19 640 51
rect 606 -51 640 -19
rect 606 -53 640 -51
rect 606 -119 640 -91
rect 606 -125 640 -119
rect 784 119 818 125
rect 784 91 818 119
rect 784 51 818 53
rect 784 19 818 51
rect 784 -51 818 -19
rect 784 -53 818 -51
rect 784 -119 818 -91
rect 784 -125 818 -119
rect 962 119 996 125
rect 962 91 996 119
rect 962 51 996 53
rect 962 19 996 51
rect 962 -51 996 -19
rect 962 -53 996 -51
rect 962 -119 996 -91
rect 962 -125 996 -119
rect 1140 119 1174 125
rect 1140 91 1174 119
rect 1140 51 1174 53
rect 1140 19 1174 51
rect 1140 -51 1174 -19
rect 1140 -53 1174 -51
rect 1140 -119 1174 -91
rect 1140 -125 1174 -119
rect 1318 119 1352 125
rect 1318 91 1352 119
rect 1318 51 1352 53
rect 1318 19 1352 51
rect 1318 -51 1352 -19
rect 1318 -53 1352 -51
rect 1318 -119 1352 -91
rect 1318 -125 1352 -119
rect 1496 119 1530 125
rect 1496 91 1530 119
rect 1496 51 1530 53
rect 1496 19 1530 51
rect 1496 -51 1530 -19
rect 1496 -53 1530 -51
rect 1496 -119 1530 -91
rect 1496 -125 1530 -119
rect 1674 119 1708 125
rect 1674 91 1708 119
rect 1674 51 1708 53
rect 1674 19 1708 51
rect 1674 -51 1708 -19
rect 1674 -53 1708 -51
rect 1674 -119 1708 -91
rect 1674 -125 1708 -119
rect 1852 119 1886 125
rect 1852 91 1886 119
rect 1852 51 1886 53
rect 1852 19 1886 51
rect 1852 -51 1886 -19
rect 1852 -53 1886 -51
rect 1852 -119 1886 -91
rect 1852 -125 1886 -119
rect 2030 119 2064 125
rect 2030 91 2064 119
rect 2030 51 2064 53
rect 2030 19 2064 51
rect 2030 -51 2064 -19
rect 2030 -53 2064 -51
rect 2030 -119 2064 -91
rect 2030 -125 2064 -119
rect -1975 -221 -1941 -187
rect -1797 -221 -1763 -187
rect -1619 -221 -1585 -187
rect -1441 -221 -1407 -187
rect -1263 -221 -1229 -187
rect -1085 -221 -1051 -187
rect -907 -221 -873 -187
rect -729 -221 -695 -187
rect -551 -221 -517 -187
rect -373 -221 -339 -187
rect -195 -221 -161 -187
rect -17 -221 17 -187
rect 161 -221 195 -187
rect 339 -221 373 -187
rect 517 -221 551 -187
rect 695 -221 729 -187
rect 873 -221 907 -187
rect 1051 -221 1085 -187
rect 1229 -221 1263 -187
rect 1407 -221 1441 -187
rect 1585 -221 1619 -187
rect 1763 -221 1797 -187
rect 1941 -221 1975 -187
<< metal1 >>
rect -1996 221 -1920 237
rect -1996 187 -1975 221
rect -1941 187 -1920 221
rect -1996 181 -1920 187
rect -1818 221 -1742 237
rect -1818 187 -1797 221
rect -1763 187 -1742 221
rect -1818 181 -1742 187
rect -1640 221 -1564 237
rect -1640 187 -1619 221
rect -1585 187 -1564 221
rect -1640 181 -1564 187
rect -1462 221 -1386 237
rect -1462 187 -1441 221
rect -1407 187 -1386 221
rect -1462 181 -1386 187
rect -1284 221 -1208 237
rect -1284 187 -1263 221
rect -1229 187 -1208 221
rect -1284 181 -1208 187
rect -1106 221 -1030 237
rect -1106 187 -1085 221
rect -1051 187 -1030 221
rect -1106 181 -1030 187
rect -928 221 -852 237
rect -928 187 -907 221
rect -873 187 -852 221
rect -928 181 -852 187
rect -750 221 -674 237
rect -750 187 -729 221
rect -695 187 -674 221
rect -750 181 -674 187
rect -572 221 -496 237
rect -572 187 -551 221
rect -517 187 -496 221
rect -572 181 -496 187
rect -394 221 -318 237
rect -394 187 -373 221
rect -339 187 -318 221
rect -394 181 -318 187
rect -216 221 -140 237
rect -216 187 -195 221
rect -161 187 -140 221
rect -216 181 -140 187
rect -38 221 38 237
rect -38 187 -17 221
rect 17 187 38 221
rect -38 181 38 187
rect 140 221 216 237
rect 140 187 161 221
rect 195 187 216 221
rect 140 181 216 187
rect 318 221 394 237
rect 318 187 339 221
rect 373 187 394 221
rect 318 181 394 187
rect 496 221 572 237
rect 496 187 517 221
rect 551 187 572 221
rect 496 181 572 187
rect 674 221 750 237
rect 674 187 695 221
rect 729 187 750 221
rect 674 181 750 187
rect 852 221 928 237
rect 852 187 873 221
rect 907 187 928 221
rect 852 181 928 187
rect 1030 221 1106 237
rect 1030 187 1051 221
rect 1085 187 1106 221
rect 1030 181 1106 187
rect 1208 221 1284 237
rect 1208 187 1229 221
rect 1263 187 1284 221
rect 1208 181 1284 187
rect 1386 221 1462 237
rect 1386 187 1407 221
rect 1441 187 1462 221
rect 1386 181 1462 187
rect 1564 221 1640 237
rect 1564 187 1585 221
rect 1619 187 1640 221
rect 1564 181 1640 187
rect 1742 221 1818 237
rect 1742 187 1763 221
rect 1797 187 1818 221
rect 1742 181 1818 187
rect 1920 221 1996 237
rect 1920 187 1941 221
rect 1975 187 1996 221
rect 1920 181 1996 187
rect -2070 125 -2024 140
rect -2070 91 -2064 125
rect -2030 91 -2024 125
rect -2070 53 -2024 91
rect -2070 19 -2064 53
rect -2030 19 -2024 53
rect -2070 -19 -2024 19
rect -2070 -53 -2064 -19
rect -2030 -53 -2024 -19
rect -2070 -91 -2024 -53
rect -2070 -125 -2064 -91
rect -2030 -125 -2024 -91
rect -2070 -140 -2024 -125
rect -1892 125 -1846 140
rect -1892 91 -1886 125
rect -1852 91 -1846 125
rect -1892 53 -1846 91
rect -1892 19 -1886 53
rect -1852 19 -1846 53
rect -1892 -19 -1846 19
rect -1892 -53 -1886 -19
rect -1852 -53 -1846 -19
rect -1892 -91 -1846 -53
rect -1892 -125 -1886 -91
rect -1852 -125 -1846 -91
rect -1892 -140 -1846 -125
rect -1714 125 -1668 140
rect -1714 91 -1708 125
rect -1674 91 -1668 125
rect -1714 53 -1668 91
rect -1714 19 -1708 53
rect -1674 19 -1668 53
rect -1714 -19 -1668 19
rect -1714 -53 -1708 -19
rect -1674 -53 -1668 -19
rect -1714 -91 -1668 -53
rect -1714 -125 -1708 -91
rect -1674 -125 -1668 -91
rect -1714 -140 -1668 -125
rect -1536 125 -1490 140
rect -1536 91 -1530 125
rect -1496 91 -1490 125
rect -1536 53 -1490 91
rect -1536 19 -1530 53
rect -1496 19 -1490 53
rect -1536 -19 -1490 19
rect -1536 -53 -1530 -19
rect -1496 -53 -1490 -19
rect -1536 -91 -1490 -53
rect -1536 -125 -1530 -91
rect -1496 -125 -1490 -91
rect -1536 -140 -1490 -125
rect -1358 125 -1312 140
rect -1358 91 -1352 125
rect -1318 91 -1312 125
rect -1358 53 -1312 91
rect -1358 19 -1352 53
rect -1318 19 -1312 53
rect -1358 -19 -1312 19
rect -1358 -53 -1352 -19
rect -1318 -53 -1312 -19
rect -1358 -91 -1312 -53
rect -1358 -125 -1352 -91
rect -1318 -125 -1312 -91
rect -1358 -140 -1312 -125
rect -1180 125 -1134 140
rect -1180 91 -1174 125
rect -1140 91 -1134 125
rect -1180 53 -1134 91
rect -1180 19 -1174 53
rect -1140 19 -1134 53
rect -1180 -19 -1134 19
rect -1180 -53 -1174 -19
rect -1140 -53 -1134 -19
rect -1180 -91 -1134 -53
rect -1180 -125 -1174 -91
rect -1140 -125 -1134 -91
rect -1180 -140 -1134 -125
rect -1002 125 -956 140
rect -1002 91 -996 125
rect -962 91 -956 125
rect -1002 53 -956 91
rect -1002 19 -996 53
rect -962 19 -956 53
rect -1002 -19 -956 19
rect -1002 -53 -996 -19
rect -962 -53 -956 -19
rect -1002 -91 -956 -53
rect -1002 -125 -996 -91
rect -962 -125 -956 -91
rect -1002 -140 -956 -125
rect -824 125 -778 140
rect -824 91 -818 125
rect -784 91 -778 125
rect -824 53 -778 91
rect -824 19 -818 53
rect -784 19 -778 53
rect -824 -19 -778 19
rect -824 -53 -818 -19
rect -784 -53 -778 -19
rect -824 -91 -778 -53
rect -824 -125 -818 -91
rect -784 -125 -778 -91
rect -824 -140 -778 -125
rect -646 125 -600 140
rect -646 91 -640 125
rect -606 91 -600 125
rect -646 53 -600 91
rect -646 19 -640 53
rect -606 19 -600 53
rect -646 -19 -600 19
rect -646 -53 -640 -19
rect -606 -53 -600 -19
rect -646 -91 -600 -53
rect -646 -125 -640 -91
rect -606 -125 -600 -91
rect -646 -140 -600 -125
rect -468 125 -422 140
rect -468 91 -462 125
rect -428 91 -422 125
rect -468 53 -422 91
rect -468 19 -462 53
rect -428 19 -422 53
rect -468 -19 -422 19
rect -468 -53 -462 -19
rect -428 -53 -422 -19
rect -468 -91 -422 -53
rect -468 -125 -462 -91
rect -428 -125 -422 -91
rect -468 -140 -422 -125
rect -290 125 -244 140
rect -290 91 -284 125
rect -250 91 -244 125
rect -290 53 -244 91
rect -290 19 -284 53
rect -250 19 -244 53
rect -290 -19 -244 19
rect -290 -53 -284 -19
rect -250 -53 -244 -19
rect -290 -91 -244 -53
rect -290 -125 -284 -91
rect -250 -125 -244 -91
rect -290 -140 -244 -125
rect -112 125 -66 140
rect -112 91 -106 125
rect -72 91 -66 125
rect -112 53 -66 91
rect -112 19 -106 53
rect -72 19 -66 53
rect -112 -19 -66 19
rect -112 -53 -106 -19
rect -72 -53 -66 -19
rect -112 -91 -66 -53
rect -112 -125 -106 -91
rect -72 -125 -66 -91
rect -112 -140 -66 -125
rect 66 125 112 140
rect 66 91 72 125
rect 106 91 112 125
rect 66 53 112 91
rect 66 19 72 53
rect 106 19 112 53
rect 66 -19 112 19
rect 66 -53 72 -19
rect 106 -53 112 -19
rect 66 -91 112 -53
rect 66 -125 72 -91
rect 106 -125 112 -91
rect 66 -140 112 -125
rect 244 125 290 140
rect 244 91 250 125
rect 284 91 290 125
rect 244 53 290 91
rect 244 19 250 53
rect 284 19 290 53
rect 244 -19 290 19
rect 244 -53 250 -19
rect 284 -53 290 -19
rect 244 -91 290 -53
rect 244 -125 250 -91
rect 284 -125 290 -91
rect 244 -140 290 -125
rect 422 125 468 140
rect 422 91 428 125
rect 462 91 468 125
rect 422 53 468 91
rect 422 19 428 53
rect 462 19 468 53
rect 422 -19 468 19
rect 422 -53 428 -19
rect 462 -53 468 -19
rect 422 -91 468 -53
rect 422 -125 428 -91
rect 462 -125 468 -91
rect 422 -140 468 -125
rect 600 125 646 140
rect 600 91 606 125
rect 640 91 646 125
rect 600 53 646 91
rect 600 19 606 53
rect 640 19 646 53
rect 600 -19 646 19
rect 600 -53 606 -19
rect 640 -53 646 -19
rect 600 -91 646 -53
rect 600 -125 606 -91
rect 640 -125 646 -91
rect 600 -140 646 -125
rect 778 125 824 140
rect 778 91 784 125
rect 818 91 824 125
rect 778 53 824 91
rect 778 19 784 53
rect 818 19 824 53
rect 778 -19 824 19
rect 778 -53 784 -19
rect 818 -53 824 -19
rect 778 -91 824 -53
rect 778 -125 784 -91
rect 818 -125 824 -91
rect 778 -140 824 -125
rect 956 125 1002 140
rect 956 91 962 125
rect 996 91 1002 125
rect 956 53 1002 91
rect 956 19 962 53
rect 996 19 1002 53
rect 956 -19 1002 19
rect 956 -53 962 -19
rect 996 -53 1002 -19
rect 956 -91 1002 -53
rect 956 -125 962 -91
rect 996 -125 1002 -91
rect 956 -140 1002 -125
rect 1134 125 1180 140
rect 1134 91 1140 125
rect 1174 91 1180 125
rect 1134 53 1180 91
rect 1134 19 1140 53
rect 1174 19 1180 53
rect 1134 -19 1180 19
rect 1134 -53 1140 -19
rect 1174 -53 1180 -19
rect 1134 -91 1180 -53
rect 1134 -125 1140 -91
rect 1174 -125 1180 -91
rect 1134 -140 1180 -125
rect 1312 125 1358 140
rect 1312 91 1318 125
rect 1352 91 1358 125
rect 1312 53 1358 91
rect 1312 19 1318 53
rect 1352 19 1358 53
rect 1312 -19 1358 19
rect 1312 -53 1318 -19
rect 1352 -53 1358 -19
rect 1312 -91 1358 -53
rect 1312 -125 1318 -91
rect 1352 -125 1358 -91
rect 1312 -140 1358 -125
rect 1490 125 1536 140
rect 1490 91 1496 125
rect 1530 91 1536 125
rect 1490 53 1536 91
rect 1490 19 1496 53
rect 1530 19 1536 53
rect 1490 -19 1536 19
rect 1490 -53 1496 -19
rect 1530 -53 1536 -19
rect 1490 -91 1536 -53
rect 1490 -125 1496 -91
rect 1530 -125 1536 -91
rect 1490 -140 1536 -125
rect 1668 125 1714 140
rect 1668 91 1674 125
rect 1708 91 1714 125
rect 1668 53 1714 91
rect 1668 19 1674 53
rect 1708 19 1714 53
rect 1668 -19 1714 19
rect 1668 -53 1674 -19
rect 1708 -53 1714 -19
rect 1668 -91 1714 -53
rect 1668 -125 1674 -91
rect 1708 -125 1714 -91
rect 1668 -140 1714 -125
rect 1846 125 1892 140
rect 1846 91 1852 125
rect 1886 91 1892 125
rect 1846 53 1892 91
rect 1846 19 1852 53
rect 1886 19 1892 53
rect 1846 -19 1892 19
rect 1846 -53 1852 -19
rect 1886 -53 1892 -19
rect 1846 -91 1892 -53
rect 1846 -125 1852 -91
rect 1886 -125 1892 -91
rect 1846 -140 1892 -125
rect 2024 125 2070 140
rect 2024 91 2030 125
rect 2064 91 2070 125
rect 2024 53 2070 91
rect 2024 19 2030 53
rect 2064 19 2070 53
rect 2024 -19 2070 19
rect 2024 -53 2030 -19
rect 2064 -53 2070 -19
rect 2024 -91 2070 -53
rect 2024 -125 2030 -91
rect 2064 -125 2070 -91
rect 2024 -140 2070 -125
rect -1996 -187 -1920 -181
rect -1996 -221 -1975 -187
rect -1941 -221 -1920 -187
rect -1996 -237 -1920 -221
rect -1818 -187 -1742 -181
rect -1818 -221 -1797 -187
rect -1763 -221 -1742 -187
rect -1818 -237 -1742 -221
rect -1640 -187 -1564 -181
rect -1640 -221 -1619 -187
rect -1585 -221 -1564 -187
rect -1640 -237 -1564 -221
rect -1462 -187 -1386 -181
rect -1462 -221 -1441 -187
rect -1407 -221 -1386 -187
rect -1462 -237 -1386 -221
rect -1284 -187 -1208 -181
rect -1284 -221 -1263 -187
rect -1229 -221 -1208 -187
rect -1284 -237 -1208 -221
rect -1106 -187 -1030 -181
rect -1106 -221 -1085 -187
rect -1051 -221 -1030 -187
rect -1106 -237 -1030 -221
rect -928 -187 -852 -181
rect -928 -221 -907 -187
rect -873 -221 -852 -187
rect -928 -237 -852 -221
rect -750 -187 -674 -181
rect -750 -221 -729 -187
rect -695 -221 -674 -187
rect -750 -237 -674 -221
rect -572 -187 -496 -181
rect -572 -221 -551 -187
rect -517 -221 -496 -187
rect -572 -237 -496 -221
rect -394 -187 -318 -181
rect -394 -221 -373 -187
rect -339 -221 -318 -187
rect -394 -237 -318 -221
rect -216 -187 -140 -181
rect -216 -221 -195 -187
rect -161 -221 -140 -187
rect -216 -237 -140 -221
rect -38 -187 38 -181
rect -38 -221 -17 -187
rect 17 -221 38 -187
rect -38 -237 38 -221
rect 140 -187 216 -181
rect 140 -221 161 -187
rect 195 -221 216 -187
rect 140 -237 216 -221
rect 318 -187 394 -181
rect 318 -221 339 -187
rect 373 -221 394 -187
rect 318 -237 394 -221
rect 496 -187 572 -181
rect 496 -221 517 -187
rect 551 -221 572 -187
rect 496 -237 572 -221
rect 674 -187 750 -181
rect 674 -221 695 -187
rect 729 -221 750 -187
rect 674 -237 750 -221
rect 852 -187 928 -181
rect 852 -221 873 -187
rect 907 -221 928 -187
rect 852 -237 928 -221
rect 1030 -187 1106 -181
rect 1030 -221 1051 -187
rect 1085 -221 1106 -187
rect 1030 -237 1106 -221
rect 1208 -187 1284 -181
rect 1208 -221 1229 -187
rect 1263 -221 1284 -187
rect 1208 -237 1284 -221
rect 1386 -187 1462 -181
rect 1386 -221 1407 -187
rect 1441 -221 1462 -187
rect 1386 -237 1462 -221
rect 1564 -187 1640 -181
rect 1564 -221 1585 -187
rect 1619 -221 1640 -187
rect 1564 -237 1640 -221
rect 1742 -187 1818 -181
rect 1742 -221 1763 -187
rect 1797 -221 1818 -187
rect 1742 -237 1818 -221
rect 1920 -187 1996 -181
rect 1920 -221 1941 -187
rect 1975 -221 1996 -187
rect 1920 -237 1996 -221
<< end >>
