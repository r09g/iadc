magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< error_p >>
rect -29 83 29 89
rect -29 49 -17 83
rect -29 43 29 49
<< nmos >>
rect -15 -89 15 11
<< ndiff >>
rect -73 -1 -15 11
rect -73 -77 -61 -1
rect -27 -77 -15 -1
rect -73 -89 -15 -77
rect 15 -1 73 11
rect 15 -77 27 -1
rect 61 -77 73 -1
rect 15 -89 73 -77
<< ndiffc >>
rect -61 -77 -27 -1
rect 27 -77 61 -1
<< poly >>
rect -33 83 33 99
rect -33 49 -17 83
rect 17 49 33 83
rect -33 33 33 49
rect -15 11 15 33
rect -15 -115 15 -89
<< polycont >>
rect -17 49 17 83
<< locali >>
rect -33 49 -17 83
rect 17 49 33 83
rect -61 -1 -27 15
rect -61 -93 -27 -77
rect 27 -1 61 15
rect 27 -93 61 -77
<< viali >>
rect -17 49 17 83
rect -61 -77 -27 -1
rect 27 -77 61 -1
<< metal1 >>
rect -29 83 29 89
rect -29 49 -17 83
rect 17 49 29 83
rect -29 43 29 49
rect -67 -1 -21 11
rect -67 -77 -61 -1
rect -27 -77 -21 -1
rect -67 -89 -21 -77
rect 21 -1 67 11
rect 21 -77 27 -1
rect 61 -77 67 -1
rect 21 -89 67 -77
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
