magic
tech sky130A
magscale 1 2
timestamp 1653627323
<< nwell >>
rect -2386 -1864 -1092 -530
rect -589 -1479 -145 -913
rect 285 -1180 3100 -530
rect 285 -2514 3100 -1864
<< pwell >>
rect -2386 -528 -1092 -66
rect 285 -528 3100 -66
rect 1553 -530 1809 -528
rect -430 -669 -396 -635
rect -417 -673 -396 -669
rect -548 -700 -462 -690
rect -417 -700 -231 -673
rect -548 -815 -231 -700
rect -548 -847 -462 -815
rect -417 -855 -231 -815
rect -548 -1692 -231 -1537
rect -548 -1702 -462 -1692
rect -417 -1719 -231 -1692
rect -417 -1723 -396 -1719
rect -430 -1757 -396 -1723
rect 285 -1862 3100 -1400
rect 1553 -1864 1809 -1862
rect -2386 -2328 -1092 -1866
<< nmos >>
rect -2186 -380 -2156 -276
rect -2090 -380 -2060 -276
rect -1994 -380 -1964 -276
rect -1898 -380 -1868 -276
rect -1802 -380 -1772 -276
rect -1706 -380 -1676 -276
rect -1610 -380 -1580 -276
rect -1514 -380 -1484 -276
rect -1418 -380 -1388 -276
rect -1322 -380 -1292 -276
rect 485 -380 515 -276
rect 581 -380 611 -276
rect 677 -380 707 -276
rect 773 -380 803 -276
rect 869 -380 899 -276
rect 965 -380 995 -276
rect 1061 -380 1091 -276
rect 1157 -380 1187 -276
rect 1253 -380 1283 -276
rect 1349 -380 1379 -276
rect 1661 -385 1691 -285
rect 2006 -380 2036 -276
rect 2102 -380 2132 -276
rect 2198 -380 2228 -276
rect 2294 -380 2324 -276
rect 2390 -380 2420 -276
rect 2486 -380 2516 -276
rect 2582 -380 2612 -276
rect 2678 -380 2708 -276
rect 2774 -380 2804 -276
rect 2870 -380 2900 -276
rect 485 -1714 515 -1610
rect 581 -1714 611 -1610
rect 677 -1714 707 -1610
rect 773 -1714 803 -1610
rect 869 -1714 899 -1610
rect 965 -1714 995 -1610
rect 1061 -1714 1091 -1610
rect 1157 -1714 1187 -1610
rect 1253 -1714 1283 -1610
rect 1349 -1714 1379 -1610
rect 1661 -1719 1691 -1619
rect 2006 -1714 2036 -1610
rect 2102 -1714 2132 -1610
rect 2198 -1714 2228 -1610
rect 2294 -1714 2324 -1610
rect 2390 -1714 2420 -1610
rect 2486 -1714 2516 -1610
rect 2582 -1714 2612 -1610
rect 2678 -1714 2708 -1610
rect 2774 -1714 2804 -1610
rect 2870 -1714 2900 -1610
rect -2186 -2118 -2156 -2014
rect -2090 -2118 -2060 -2014
rect -1994 -2118 -1964 -2014
rect -1898 -2118 -1868 -2014
rect -1802 -2118 -1772 -2014
rect -1706 -2118 -1676 -2014
rect -1610 -2118 -1580 -2014
rect -1514 -2118 -1484 -2014
rect -1418 -2118 -1388 -2014
rect -1322 -2118 -1292 -2014
<< scnmos >>
rect -339 -829 -309 -699
rect -339 -1693 -309 -1563
<< pmos >>
rect -2186 -960 -2156 -688
rect -2090 -960 -2060 -688
rect -1994 -960 -1964 -688
rect -1898 -960 -1868 -688
rect -1802 -960 -1772 -688
rect -1706 -960 -1676 -688
rect -1610 -960 -1580 -688
rect -1514 -960 -1484 -688
rect -1418 -960 -1388 -688
rect -1322 -960 -1292 -688
rect 485 -960 515 -688
rect 581 -960 611 -688
rect 677 -960 707 -688
rect 773 -960 803 -688
rect 869 -960 899 -688
rect 965 -960 995 -688
rect 1061 -960 1091 -688
rect 1157 -960 1187 -688
rect 1253 -960 1283 -688
rect 1349 -960 1379 -688
rect 2006 -960 2036 -688
rect 2102 -960 2132 -688
rect 2198 -960 2228 -688
rect 2294 -960 2324 -688
rect 2390 -960 2420 -688
rect 2486 -960 2516 -688
rect 2582 -960 2612 -688
rect 2678 -960 2708 -688
rect 2774 -960 2804 -688
rect 2870 -960 2900 -688
rect -2186 -1706 -2156 -1434
rect -2090 -1706 -2060 -1434
rect -1994 -1706 -1964 -1434
rect -1898 -1706 -1868 -1434
rect -1802 -1706 -1772 -1434
rect -1706 -1706 -1676 -1434
rect -1610 -1706 -1580 -1434
rect -1514 -1706 -1484 -1434
rect -1418 -1706 -1388 -1434
rect -1322 -1706 -1292 -1434
rect 485 -2294 515 -2022
rect 581 -2294 611 -2022
rect 677 -2294 707 -2022
rect 773 -2294 803 -2022
rect 869 -2294 899 -2022
rect 965 -2294 995 -2022
rect 1061 -2294 1091 -2022
rect 1157 -2294 1187 -2022
rect 1253 -2294 1283 -2022
rect 1349 -2294 1379 -2022
rect 2006 -2294 2036 -2022
rect 2102 -2294 2132 -2022
rect 2198 -2294 2228 -2022
rect 2294 -2294 2324 -2022
rect 2390 -2294 2420 -2022
rect 2486 -2294 2516 -2022
rect 2582 -2294 2612 -2022
rect 2678 -2294 2708 -2022
rect 2774 -2294 2804 -2022
rect 2870 -2294 2900 -2022
<< scpmoshvt >>
rect -339 -1149 -309 -949
rect -339 -1443 -309 -1243
<< ndiff >>
rect -2248 -288 -2186 -276
rect -2248 -368 -2236 -288
rect -2202 -368 -2186 -288
rect -2248 -380 -2186 -368
rect -2156 -288 -2090 -276
rect -2156 -368 -2140 -288
rect -2106 -368 -2090 -288
rect -2156 -380 -2090 -368
rect -2060 -288 -1994 -276
rect -2060 -368 -2044 -288
rect -2010 -368 -1994 -288
rect -2060 -380 -1994 -368
rect -1964 -288 -1898 -276
rect -1964 -368 -1948 -288
rect -1914 -368 -1898 -288
rect -1964 -380 -1898 -368
rect -1868 -288 -1802 -276
rect -1868 -368 -1852 -288
rect -1818 -368 -1802 -288
rect -1868 -380 -1802 -368
rect -1772 -288 -1706 -276
rect -1772 -368 -1756 -288
rect -1722 -368 -1706 -288
rect -1772 -380 -1706 -368
rect -1676 -288 -1610 -276
rect -1676 -368 -1660 -288
rect -1626 -368 -1610 -288
rect -1676 -380 -1610 -368
rect -1580 -288 -1514 -276
rect -1580 -368 -1564 -288
rect -1530 -368 -1514 -288
rect -1580 -380 -1514 -368
rect -1484 -288 -1418 -276
rect -1484 -368 -1468 -288
rect -1434 -368 -1418 -288
rect -1484 -380 -1418 -368
rect -1388 -288 -1322 -276
rect -1388 -368 -1372 -288
rect -1338 -368 -1322 -288
rect -1388 -380 -1322 -368
rect -1292 -288 -1230 -276
rect -1292 -368 -1276 -288
rect -1242 -368 -1230 -288
rect -1292 -380 -1230 -368
rect 423 -288 485 -276
rect 423 -368 435 -288
rect 469 -368 485 -288
rect 423 -380 485 -368
rect 515 -288 581 -276
rect 515 -368 531 -288
rect 565 -368 581 -288
rect 515 -380 581 -368
rect 611 -288 677 -276
rect 611 -368 627 -288
rect 661 -368 677 -288
rect 611 -380 677 -368
rect 707 -288 773 -276
rect 707 -368 723 -288
rect 757 -368 773 -288
rect 707 -380 773 -368
rect 803 -288 869 -276
rect 803 -368 819 -288
rect 853 -368 869 -288
rect 803 -380 869 -368
rect 899 -288 965 -276
rect 899 -368 915 -288
rect 949 -368 965 -288
rect 899 -380 965 -368
rect 995 -288 1061 -276
rect 995 -368 1011 -288
rect 1045 -368 1061 -288
rect 995 -380 1061 -368
rect 1091 -288 1157 -276
rect 1091 -368 1107 -288
rect 1141 -368 1157 -288
rect 1091 -380 1157 -368
rect 1187 -288 1253 -276
rect 1187 -368 1203 -288
rect 1237 -368 1253 -288
rect 1187 -380 1253 -368
rect 1283 -288 1349 -276
rect 1283 -368 1299 -288
rect 1333 -368 1349 -288
rect 1283 -380 1349 -368
rect 1379 -288 1441 -276
rect 1379 -368 1395 -288
rect 1429 -368 1441 -288
rect 1379 -380 1441 -368
rect 1603 -297 1661 -285
rect 1603 -373 1615 -297
rect 1649 -373 1661 -297
rect 1603 -385 1661 -373
rect 1691 -297 1749 -285
rect 1691 -373 1703 -297
rect 1737 -373 1749 -297
rect 1691 -385 1749 -373
rect 1944 -288 2006 -276
rect 1944 -368 1956 -288
rect 1990 -368 2006 -288
rect 1944 -380 2006 -368
rect 2036 -288 2102 -276
rect 2036 -368 2052 -288
rect 2086 -368 2102 -288
rect 2036 -380 2102 -368
rect 2132 -288 2198 -276
rect 2132 -368 2148 -288
rect 2182 -368 2198 -288
rect 2132 -380 2198 -368
rect 2228 -288 2294 -276
rect 2228 -368 2244 -288
rect 2278 -368 2294 -288
rect 2228 -380 2294 -368
rect 2324 -288 2390 -276
rect 2324 -368 2340 -288
rect 2374 -368 2390 -288
rect 2324 -380 2390 -368
rect 2420 -288 2486 -276
rect 2420 -368 2436 -288
rect 2470 -368 2486 -288
rect 2420 -380 2486 -368
rect 2516 -288 2582 -276
rect 2516 -368 2532 -288
rect 2566 -368 2582 -288
rect 2516 -380 2582 -368
rect 2612 -288 2678 -276
rect 2612 -368 2628 -288
rect 2662 -368 2678 -288
rect 2612 -380 2678 -368
rect 2708 -288 2774 -276
rect 2708 -368 2724 -288
rect 2758 -368 2774 -288
rect 2708 -380 2774 -368
rect 2804 -288 2870 -276
rect 2804 -368 2820 -288
rect 2854 -368 2870 -288
rect 2804 -380 2870 -368
rect 2900 -288 2962 -276
rect 2900 -368 2916 -288
rect 2950 -368 2962 -288
rect 2900 -380 2962 -368
rect -391 -715 -339 -699
rect -391 -749 -383 -715
rect -349 -749 -339 -715
rect -391 -783 -339 -749
rect -391 -817 -383 -783
rect -349 -817 -339 -783
rect -391 -829 -339 -817
rect -309 -715 -257 -699
rect -309 -749 -299 -715
rect -265 -749 -257 -715
rect -309 -783 -257 -749
rect -309 -817 -299 -783
rect -265 -817 -257 -783
rect -309 -829 -257 -817
rect -391 -1575 -339 -1563
rect -391 -1609 -383 -1575
rect -349 -1609 -339 -1575
rect -391 -1643 -339 -1609
rect -391 -1677 -383 -1643
rect -349 -1677 -339 -1643
rect -391 -1693 -339 -1677
rect -309 -1575 -257 -1563
rect -309 -1609 -299 -1575
rect -265 -1609 -257 -1575
rect -309 -1643 -257 -1609
rect -309 -1677 -299 -1643
rect -265 -1677 -257 -1643
rect -309 -1693 -257 -1677
rect 423 -1622 485 -1610
rect 423 -1702 435 -1622
rect 469 -1702 485 -1622
rect 423 -1714 485 -1702
rect 515 -1622 581 -1610
rect 515 -1702 531 -1622
rect 565 -1702 581 -1622
rect 515 -1714 581 -1702
rect 611 -1622 677 -1610
rect 611 -1702 627 -1622
rect 661 -1702 677 -1622
rect 611 -1714 677 -1702
rect 707 -1622 773 -1610
rect 707 -1702 723 -1622
rect 757 -1702 773 -1622
rect 707 -1714 773 -1702
rect 803 -1622 869 -1610
rect 803 -1702 819 -1622
rect 853 -1702 869 -1622
rect 803 -1714 869 -1702
rect 899 -1622 965 -1610
rect 899 -1702 915 -1622
rect 949 -1702 965 -1622
rect 899 -1714 965 -1702
rect 995 -1622 1061 -1610
rect 995 -1702 1011 -1622
rect 1045 -1702 1061 -1622
rect 995 -1714 1061 -1702
rect 1091 -1622 1157 -1610
rect 1091 -1702 1107 -1622
rect 1141 -1702 1157 -1622
rect 1091 -1714 1157 -1702
rect 1187 -1622 1253 -1610
rect 1187 -1702 1203 -1622
rect 1237 -1702 1253 -1622
rect 1187 -1714 1253 -1702
rect 1283 -1622 1349 -1610
rect 1283 -1702 1299 -1622
rect 1333 -1702 1349 -1622
rect 1283 -1714 1349 -1702
rect 1379 -1622 1441 -1610
rect 1379 -1702 1395 -1622
rect 1429 -1702 1441 -1622
rect 1379 -1714 1441 -1702
rect 1603 -1631 1661 -1619
rect 1603 -1707 1615 -1631
rect 1649 -1707 1661 -1631
rect 1603 -1719 1661 -1707
rect 1691 -1631 1749 -1619
rect 1691 -1707 1703 -1631
rect 1737 -1707 1749 -1631
rect 1691 -1719 1749 -1707
rect 1944 -1622 2006 -1610
rect 1944 -1702 1956 -1622
rect 1990 -1702 2006 -1622
rect 1944 -1714 2006 -1702
rect 2036 -1622 2102 -1610
rect 2036 -1702 2052 -1622
rect 2086 -1702 2102 -1622
rect 2036 -1714 2102 -1702
rect 2132 -1622 2198 -1610
rect 2132 -1702 2148 -1622
rect 2182 -1702 2198 -1622
rect 2132 -1714 2198 -1702
rect 2228 -1622 2294 -1610
rect 2228 -1702 2244 -1622
rect 2278 -1702 2294 -1622
rect 2228 -1714 2294 -1702
rect 2324 -1622 2390 -1610
rect 2324 -1702 2340 -1622
rect 2374 -1702 2390 -1622
rect 2324 -1714 2390 -1702
rect 2420 -1622 2486 -1610
rect 2420 -1702 2436 -1622
rect 2470 -1702 2486 -1622
rect 2420 -1714 2486 -1702
rect 2516 -1622 2582 -1610
rect 2516 -1702 2532 -1622
rect 2566 -1702 2582 -1622
rect 2516 -1714 2582 -1702
rect 2612 -1622 2678 -1610
rect 2612 -1702 2628 -1622
rect 2662 -1702 2678 -1622
rect 2612 -1714 2678 -1702
rect 2708 -1622 2774 -1610
rect 2708 -1702 2724 -1622
rect 2758 -1702 2774 -1622
rect 2708 -1714 2774 -1702
rect 2804 -1622 2870 -1610
rect 2804 -1702 2820 -1622
rect 2854 -1702 2870 -1622
rect 2804 -1714 2870 -1702
rect 2900 -1622 2962 -1610
rect 2900 -1702 2916 -1622
rect 2950 -1702 2962 -1622
rect 2900 -1714 2962 -1702
rect -2248 -2026 -2186 -2014
rect -2248 -2106 -2236 -2026
rect -2202 -2106 -2186 -2026
rect -2248 -2118 -2186 -2106
rect -2156 -2026 -2090 -2014
rect -2156 -2106 -2140 -2026
rect -2106 -2106 -2090 -2026
rect -2156 -2118 -2090 -2106
rect -2060 -2026 -1994 -2014
rect -2060 -2106 -2044 -2026
rect -2010 -2106 -1994 -2026
rect -2060 -2118 -1994 -2106
rect -1964 -2026 -1898 -2014
rect -1964 -2106 -1948 -2026
rect -1914 -2106 -1898 -2026
rect -1964 -2118 -1898 -2106
rect -1868 -2026 -1802 -2014
rect -1868 -2106 -1852 -2026
rect -1818 -2106 -1802 -2026
rect -1868 -2118 -1802 -2106
rect -1772 -2026 -1706 -2014
rect -1772 -2106 -1756 -2026
rect -1722 -2106 -1706 -2026
rect -1772 -2118 -1706 -2106
rect -1676 -2026 -1610 -2014
rect -1676 -2106 -1660 -2026
rect -1626 -2106 -1610 -2026
rect -1676 -2118 -1610 -2106
rect -1580 -2026 -1514 -2014
rect -1580 -2106 -1564 -2026
rect -1530 -2106 -1514 -2026
rect -1580 -2118 -1514 -2106
rect -1484 -2026 -1418 -2014
rect -1484 -2106 -1468 -2026
rect -1434 -2106 -1418 -2026
rect -1484 -2118 -1418 -2106
rect -1388 -2026 -1322 -2014
rect -1388 -2106 -1372 -2026
rect -1338 -2106 -1322 -2026
rect -1388 -2118 -1322 -2106
rect -1292 -2026 -1230 -2014
rect -1292 -2106 -1276 -2026
rect -1242 -2106 -1230 -2026
rect -1292 -2118 -1230 -2106
<< pdiff >>
rect -2248 -700 -2186 -688
rect -2248 -948 -2236 -700
rect -2202 -948 -2186 -700
rect -2248 -960 -2186 -948
rect -2156 -700 -2090 -688
rect -2156 -948 -2140 -700
rect -2106 -948 -2090 -700
rect -2156 -960 -2090 -948
rect -2060 -700 -1994 -688
rect -2060 -948 -2044 -700
rect -2010 -948 -1994 -700
rect -2060 -960 -1994 -948
rect -1964 -700 -1898 -688
rect -1964 -948 -1948 -700
rect -1914 -948 -1898 -700
rect -1964 -960 -1898 -948
rect -1868 -700 -1802 -688
rect -1868 -948 -1852 -700
rect -1818 -948 -1802 -700
rect -1868 -960 -1802 -948
rect -1772 -700 -1706 -688
rect -1772 -948 -1756 -700
rect -1722 -948 -1706 -700
rect -1772 -960 -1706 -948
rect -1676 -700 -1610 -688
rect -1676 -948 -1660 -700
rect -1626 -948 -1610 -700
rect -1676 -960 -1610 -948
rect -1580 -700 -1514 -688
rect -1580 -948 -1564 -700
rect -1530 -948 -1514 -700
rect -1580 -960 -1514 -948
rect -1484 -700 -1418 -688
rect -1484 -948 -1468 -700
rect -1434 -948 -1418 -700
rect -1484 -960 -1418 -948
rect -1388 -700 -1322 -688
rect -1388 -948 -1372 -700
rect -1338 -948 -1322 -700
rect -1388 -960 -1322 -948
rect -1292 -700 -1230 -688
rect -1292 -948 -1276 -700
rect -1242 -948 -1230 -700
rect -1292 -960 -1230 -948
rect -391 -967 -339 -949
rect -391 -1001 -383 -967
rect -349 -1001 -339 -967
rect -391 -1035 -339 -1001
rect -391 -1069 -383 -1035
rect -349 -1069 -339 -1035
rect -391 -1103 -339 -1069
rect -391 -1137 -383 -1103
rect -349 -1137 -339 -1103
rect -391 -1149 -339 -1137
rect -309 -967 -257 -949
rect -309 -1001 -299 -967
rect -265 -1001 -257 -967
rect -309 -1035 -257 -1001
rect -309 -1069 -299 -1035
rect -265 -1069 -257 -1035
rect -309 -1103 -257 -1069
rect -309 -1137 -299 -1103
rect -265 -1137 -257 -1103
rect -309 -1149 -257 -1137
rect 423 -700 485 -688
rect 423 -948 435 -700
rect 469 -948 485 -700
rect 423 -960 485 -948
rect 515 -700 581 -688
rect 515 -948 531 -700
rect 565 -948 581 -700
rect 515 -960 581 -948
rect 611 -700 677 -688
rect 611 -948 627 -700
rect 661 -948 677 -700
rect 611 -960 677 -948
rect 707 -700 773 -688
rect 707 -948 723 -700
rect 757 -948 773 -700
rect 707 -960 773 -948
rect 803 -700 869 -688
rect 803 -948 819 -700
rect 853 -948 869 -700
rect 803 -960 869 -948
rect 899 -700 965 -688
rect 899 -948 915 -700
rect 949 -948 965 -700
rect 899 -960 965 -948
rect 995 -700 1061 -688
rect 995 -948 1011 -700
rect 1045 -948 1061 -700
rect 995 -960 1061 -948
rect 1091 -700 1157 -688
rect 1091 -948 1107 -700
rect 1141 -948 1157 -700
rect 1091 -960 1157 -948
rect 1187 -700 1253 -688
rect 1187 -948 1203 -700
rect 1237 -948 1253 -700
rect 1187 -960 1253 -948
rect 1283 -700 1349 -688
rect 1283 -948 1299 -700
rect 1333 -948 1349 -700
rect 1283 -960 1349 -948
rect 1379 -700 1441 -688
rect 1379 -948 1395 -700
rect 1429 -948 1441 -700
rect 1379 -960 1441 -948
rect 1944 -700 2006 -688
rect 1944 -948 1956 -700
rect 1990 -948 2006 -700
rect 1944 -960 2006 -948
rect 2036 -700 2102 -688
rect 2036 -948 2052 -700
rect 2086 -948 2102 -700
rect 2036 -960 2102 -948
rect 2132 -700 2198 -688
rect 2132 -948 2148 -700
rect 2182 -948 2198 -700
rect 2132 -960 2198 -948
rect 2228 -700 2294 -688
rect 2228 -948 2244 -700
rect 2278 -948 2294 -700
rect 2228 -960 2294 -948
rect 2324 -700 2390 -688
rect 2324 -948 2340 -700
rect 2374 -948 2390 -700
rect 2324 -960 2390 -948
rect 2420 -700 2486 -688
rect 2420 -948 2436 -700
rect 2470 -948 2486 -700
rect 2420 -960 2486 -948
rect 2516 -700 2582 -688
rect 2516 -948 2532 -700
rect 2566 -948 2582 -700
rect 2516 -960 2582 -948
rect 2612 -700 2678 -688
rect 2612 -948 2628 -700
rect 2662 -948 2678 -700
rect 2612 -960 2678 -948
rect 2708 -700 2774 -688
rect 2708 -948 2724 -700
rect 2758 -948 2774 -700
rect 2708 -960 2774 -948
rect 2804 -700 2870 -688
rect 2804 -948 2820 -700
rect 2854 -948 2870 -700
rect 2804 -960 2870 -948
rect 2900 -700 2962 -688
rect 2900 -948 2916 -700
rect 2950 -948 2962 -700
rect 2900 -960 2962 -948
rect -391 -1255 -339 -1243
rect -2248 -1446 -2186 -1434
rect -2248 -1694 -2236 -1446
rect -2202 -1694 -2186 -1446
rect -2248 -1706 -2186 -1694
rect -2156 -1446 -2090 -1434
rect -2156 -1694 -2140 -1446
rect -2106 -1694 -2090 -1446
rect -2156 -1706 -2090 -1694
rect -2060 -1446 -1994 -1434
rect -2060 -1694 -2044 -1446
rect -2010 -1694 -1994 -1446
rect -2060 -1706 -1994 -1694
rect -1964 -1446 -1898 -1434
rect -1964 -1694 -1948 -1446
rect -1914 -1694 -1898 -1446
rect -1964 -1706 -1898 -1694
rect -1868 -1446 -1802 -1434
rect -1868 -1694 -1852 -1446
rect -1818 -1694 -1802 -1446
rect -1868 -1706 -1802 -1694
rect -1772 -1446 -1706 -1434
rect -1772 -1694 -1756 -1446
rect -1722 -1694 -1706 -1446
rect -1772 -1706 -1706 -1694
rect -1676 -1446 -1610 -1434
rect -1676 -1694 -1660 -1446
rect -1626 -1694 -1610 -1446
rect -1676 -1706 -1610 -1694
rect -1580 -1446 -1514 -1434
rect -1580 -1694 -1564 -1446
rect -1530 -1694 -1514 -1446
rect -1580 -1706 -1514 -1694
rect -1484 -1446 -1418 -1434
rect -1484 -1694 -1468 -1446
rect -1434 -1694 -1418 -1446
rect -1484 -1706 -1418 -1694
rect -1388 -1446 -1322 -1434
rect -1388 -1694 -1372 -1446
rect -1338 -1694 -1322 -1446
rect -1388 -1706 -1322 -1694
rect -1292 -1446 -1230 -1434
rect -1292 -1694 -1276 -1446
rect -1242 -1694 -1230 -1446
rect -1292 -1706 -1230 -1694
rect -391 -1289 -383 -1255
rect -349 -1289 -339 -1255
rect -391 -1323 -339 -1289
rect -391 -1357 -383 -1323
rect -349 -1357 -339 -1323
rect -391 -1391 -339 -1357
rect -391 -1425 -383 -1391
rect -349 -1425 -339 -1391
rect -391 -1443 -339 -1425
rect -309 -1255 -257 -1243
rect -309 -1289 -299 -1255
rect -265 -1289 -257 -1255
rect -309 -1323 -257 -1289
rect -309 -1357 -299 -1323
rect -265 -1357 -257 -1323
rect -309 -1391 -257 -1357
rect -309 -1425 -299 -1391
rect -265 -1425 -257 -1391
rect -309 -1443 -257 -1425
rect 423 -2034 485 -2022
rect 423 -2282 435 -2034
rect 469 -2282 485 -2034
rect 423 -2294 485 -2282
rect 515 -2034 581 -2022
rect 515 -2282 531 -2034
rect 565 -2282 581 -2034
rect 515 -2294 581 -2282
rect 611 -2034 677 -2022
rect 611 -2282 627 -2034
rect 661 -2282 677 -2034
rect 611 -2294 677 -2282
rect 707 -2034 773 -2022
rect 707 -2282 723 -2034
rect 757 -2282 773 -2034
rect 707 -2294 773 -2282
rect 803 -2034 869 -2022
rect 803 -2282 819 -2034
rect 853 -2282 869 -2034
rect 803 -2294 869 -2282
rect 899 -2034 965 -2022
rect 899 -2282 915 -2034
rect 949 -2282 965 -2034
rect 899 -2294 965 -2282
rect 995 -2034 1061 -2022
rect 995 -2282 1011 -2034
rect 1045 -2282 1061 -2034
rect 995 -2294 1061 -2282
rect 1091 -2034 1157 -2022
rect 1091 -2282 1107 -2034
rect 1141 -2282 1157 -2034
rect 1091 -2294 1157 -2282
rect 1187 -2034 1253 -2022
rect 1187 -2282 1203 -2034
rect 1237 -2282 1253 -2034
rect 1187 -2294 1253 -2282
rect 1283 -2034 1349 -2022
rect 1283 -2282 1299 -2034
rect 1333 -2282 1349 -2034
rect 1283 -2294 1349 -2282
rect 1379 -2034 1441 -2022
rect 1379 -2282 1395 -2034
rect 1429 -2282 1441 -2034
rect 1379 -2294 1441 -2282
rect 1944 -2034 2006 -2022
rect 1944 -2282 1956 -2034
rect 1990 -2282 2006 -2034
rect 1944 -2294 2006 -2282
rect 2036 -2034 2102 -2022
rect 2036 -2282 2052 -2034
rect 2086 -2282 2102 -2034
rect 2036 -2294 2102 -2282
rect 2132 -2034 2198 -2022
rect 2132 -2282 2148 -2034
rect 2182 -2282 2198 -2034
rect 2132 -2294 2198 -2282
rect 2228 -2034 2294 -2022
rect 2228 -2282 2244 -2034
rect 2278 -2282 2294 -2034
rect 2228 -2294 2294 -2282
rect 2324 -2034 2390 -2022
rect 2324 -2282 2340 -2034
rect 2374 -2282 2390 -2034
rect 2324 -2294 2390 -2282
rect 2420 -2034 2486 -2022
rect 2420 -2282 2436 -2034
rect 2470 -2282 2486 -2034
rect 2420 -2294 2486 -2282
rect 2516 -2034 2582 -2022
rect 2516 -2282 2532 -2034
rect 2566 -2282 2582 -2034
rect 2516 -2294 2582 -2282
rect 2612 -2034 2678 -2022
rect 2612 -2282 2628 -2034
rect 2662 -2282 2678 -2034
rect 2612 -2294 2678 -2282
rect 2708 -2034 2774 -2022
rect 2708 -2282 2724 -2034
rect 2758 -2282 2774 -2034
rect 2708 -2294 2774 -2282
rect 2804 -2034 2870 -2022
rect 2804 -2282 2820 -2034
rect 2854 -2282 2870 -2034
rect 2804 -2294 2870 -2282
rect 2900 -2034 2962 -2022
rect 2900 -2282 2916 -2034
rect 2950 -2282 2962 -2034
rect 2900 -2294 2962 -2282
<< ndiffc >>
rect -2236 -368 -2202 -288
rect -2140 -368 -2106 -288
rect -2044 -368 -2010 -288
rect -1948 -368 -1914 -288
rect -1852 -368 -1818 -288
rect -1756 -368 -1722 -288
rect -1660 -368 -1626 -288
rect -1564 -368 -1530 -288
rect -1468 -368 -1434 -288
rect -1372 -368 -1338 -288
rect -1276 -368 -1242 -288
rect 435 -368 469 -288
rect 531 -368 565 -288
rect 627 -368 661 -288
rect 723 -368 757 -288
rect 819 -368 853 -288
rect 915 -368 949 -288
rect 1011 -368 1045 -288
rect 1107 -368 1141 -288
rect 1203 -368 1237 -288
rect 1299 -368 1333 -288
rect 1395 -368 1429 -288
rect 1615 -373 1649 -297
rect 1703 -373 1737 -297
rect 1956 -368 1990 -288
rect 2052 -368 2086 -288
rect 2148 -368 2182 -288
rect 2244 -368 2278 -288
rect 2340 -368 2374 -288
rect 2436 -368 2470 -288
rect 2532 -368 2566 -288
rect 2628 -368 2662 -288
rect 2724 -368 2758 -288
rect 2820 -368 2854 -288
rect 2916 -368 2950 -288
rect -383 -749 -349 -715
rect -383 -817 -349 -783
rect -299 -749 -265 -715
rect -299 -817 -265 -783
rect -383 -1609 -349 -1575
rect -383 -1677 -349 -1643
rect -299 -1609 -265 -1575
rect -299 -1677 -265 -1643
rect 435 -1702 469 -1622
rect 531 -1702 565 -1622
rect 627 -1702 661 -1622
rect 723 -1702 757 -1622
rect 819 -1702 853 -1622
rect 915 -1702 949 -1622
rect 1011 -1702 1045 -1622
rect 1107 -1702 1141 -1622
rect 1203 -1702 1237 -1622
rect 1299 -1702 1333 -1622
rect 1395 -1702 1429 -1622
rect 1615 -1707 1649 -1631
rect 1703 -1707 1737 -1631
rect 1956 -1702 1990 -1622
rect 2052 -1702 2086 -1622
rect 2148 -1702 2182 -1622
rect 2244 -1702 2278 -1622
rect 2340 -1702 2374 -1622
rect 2436 -1702 2470 -1622
rect 2532 -1702 2566 -1622
rect 2628 -1702 2662 -1622
rect 2724 -1702 2758 -1622
rect 2820 -1702 2854 -1622
rect 2916 -1702 2950 -1622
rect -2236 -2106 -2202 -2026
rect -2140 -2106 -2106 -2026
rect -2044 -2106 -2010 -2026
rect -1948 -2106 -1914 -2026
rect -1852 -2106 -1818 -2026
rect -1756 -2106 -1722 -2026
rect -1660 -2106 -1626 -2026
rect -1564 -2106 -1530 -2026
rect -1468 -2106 -1434 -2026
rect -1372 -2106 -1338 -2026
rect -1276 -2106 -1242 -2026
<< pdiffc >>
rect -2236 -948 -2202 -700
rect -2140 -948 -2106 -700
rect -2044 -948 -2010 -700
rect -1948 -948 -1914 -700
rect -1852 -948 -1818 -700
rect -1756 -948 -1722 -700
rect -1660 -948 -1626 -700
rect -1564 -948 -1530 -700
rect -1468 -948 -1434 -700
rect -1372 -948 -1338 -700
rect -1276 -948 -1242 -700
rect -383 -1001 -349 -967
rect -383 -1069 -349 -1035
rect -383 -1137 -349 -1103
rect -299 -1001 -265 -967
rect -299 -1069 -265 -1035
rect -299 -1137 -265 -1103
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect -2236 -1694 -2202 -1446
rect -2140 -1694 -2106 -1446
rect -2044 -1694 -2010 -1446
rect -1948 -1694 -1914 -1446
rect -1852 -1694 -1818 -1446
rect -1756 -1694 -1722 -1446
rect -1660 -1694 -1626 -1446
rect -1564 -1694 -1530 -1446
rect -1468 -1694 -1434 -1446
rect -1372 -1694 -1338 -1446
rect -1276 -1694 -1242 -1446
rect -383 -1289 -349 -1255
rect -383 -1357 -349 -1323
rect -383 -1425 -349 -1391
rect -299 -1289 -265 -1255
rect -299 -1357 -265 -1323
rect -299 -1425 -265 -1391
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
<< psubdiff >>
rect -2350 -136 -2254 -102
rect -1224 -136 -1128 -102
rect -2350 -198 -2316 -136
rect -1162 -198 -1128 -136
rect -2350 -458 -2316 -396
rect -1162 -458 -1128 -396
rect -2350 -492 -2254 -458
rect -1224 -492 -1128 -458
rect 321 -136 417 -102
rect 1447 -136 1543 -102
rect 321 -198 355 -136
rect 1509 -198 1543 -136
rect 321 -458 355 -396
rect 1842 -136 1938 -102
rect 2968 -136 3064 -102
rect 1842 -198 1876 -136
rect 1509 -458 1543 -396
rect 3030 -198 3064 -136
rect 321 -492 417 -458
rect 1447 -492 1543 -458
rect 1842 -458 1876 -396
rect 3030 -458 3064 -396
rect 1842 -492 1938 -458
rect 2968 -492 3064 -458
rect -522 -763 -488 -716
rect -522 -821 -488 -797
rect 321 -1470 417 -1436
rect 1447 -1470 1543 -1436
rect 321 -1532 355 -1470
rect -522 -1595 -488 -1571
rect -522 -1676 -488 -1629
rect 1509 -1532 1543 -1470
rect 321 -1792 355 -1730
rect 1842 -1470 1938 -1436
rect 2968 -1470 3064 -1436
rect 1842 -1532 1876 -1470
rect 1509 -1792 1543 -1730
rect 3030 -1532 3064 -1470
rect 321 -1826 417 -1792
rect 1447 -1826 1543 -1792
rect 1842 -1792 1876 -1730
rect 3030 -1792 3064 -1730
rect 1842 -1826 1938 -1792
rect 2968 -1826 3064 -1792
rect -2350 -1936 -2254 -1902
rect -1224 -1936 -1128 -1902
rect -2350 -1998 -2316 -1936
rect -1162 -1998 -1128 -1936
rect -2350 -2258 -2316 -2196
rect -1162 -2258 -1128 -2196
rect -2350 -2292 -2254 -2258
rect -1224 -2292 -1128 -2258
<< nsubdiff >>
rect -2350 -600 -2254 -566
rect -1224 -600 -1128 -566
rect -2350 -662 -2316 -600
rect -1162 -662 -1128 -600
rect -2350 -1110 -2316 -1048
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect 1509 -662 1543 -600
rect -1162 -1110 -1128 -1048
rect -2350 -1144 -2254 -1110
rect -1224 -1144 -1128 -1110
rect -522 -981 -488 -957
rect -522 -1074 -488 -1015
rect -522 -1132 -488 -1108
rect 321 -1110 355 -1048
rect 1509 -1110 1543 -1048
rect 321 -1144 417 -1110
rect 1447 -1144 1543 -1110
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1842 -1110 1876 -1048
rect 3030 -1110 3064 -1048
rect 1842 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect -2350 -1284 -2254 -1250
rect -1224 -1284 -1128 -1250
rect -2350 -1346 -2316 -1284
rect -1162 -1346 -1128 -1284
rect -522 -1284 -488 -1260
rect -522 -1377 -488 -1318
rect -522 -1435 -488 -1411
rect -2350 -1794 -2316 -1732
rect -1162 -1794 -1128 -1732
rect -2350 -1828 -2254 -1794
rect -1224 -1828 -1128 -1794
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect 321 -2444 355 -2382
rect 1509 -2444 1543 -2382
rect 321 -2478 417 -2444
rect 1447 -2478 1543 -2444
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1842 -2444 1876 -2382
rect 3030 -2444 3064 -2382
rect 1842 -2478 1938 -2444
rect 2968 -2478 3064 -2444
<< psubdiffcont >>
rect -2254 -136 -1224 -102
rect -2350 -396 -2316 -198
rect -1162 -396 -1128 -198
rect -2254 -492 -1224 -458
rect 417 -136 1447 -102
rect 321 -396 355 -198
rect 1509 -396 1543 -198
rect 1938 -136 2968 -102
rect 1842 -396 1876 -198
rect 417 -492 1447 -458
rect 3030 -396 3064 -198
rect 1938 -492 2968 -458
rect -522 -797 -488 -763
rect 417 -1470 1447 -1436
rect -522 -1629 -488 -1595
rect 321 -1730 355 -1532
rect 1509 -1730 1543 -1532
rect 1938 -1470 2968 -1436
rect 1842 -1730 1876 -1532
rect 417 -1826 1447 -1792
rect 3030 -1730 3064 -1532
rect 1938 -1826 2968 -1792
rect -2254 -1936 -1224 -1902
rect -2350 -2196 -2316 -1998
rect -1162 -2196 -1128 -1998
rect -2254 -2292 -1224 -2258
<< nsubdiffcont >>
rect -2254 -600 -1224 -566
rect -2350 -1048 -2316 -662
rect -1162 -1048 -1128 -662
rect 417 -600 1447 -566
rect -2254 -1144 -1224 -1110
rect -522 -1015 -488 -981
rect -522 -1108 -488 -1074
rect 321 -1048 355 -662
rect 1509 -1048 1543 -662
rect 417 -1144 1447 -1110
rect 1938 -600 2968 -566
rect 1842 -1048 1876 -662
rect 3030 -1048 3064 -662
rect 1938 -1144 2968 -1110
rect -2254 -1284 -1224 -1250
rect -2350 -1732 -2316 -1346
rect -1162 -1732 -1128 -1346
rect -522 -1318 -488 -1284
rect -522 -1411 -488 -1377
rect -2254 -1828 -1224 -1794
rect 417 -1934 1447 -1900
rect 321 -2382 355 -1996
rect 1509 -2382 1543 -1996
rect 417 -2478 1447 -2444
rect 1938 -1934 2968 -1900
rect 1842 -2382 1876 -1996
rect 3030 -2382 3064 -1996
rect 1938 -2478 2968 -2444
<< poly >>
rect -2252 -200 -1226 -188
rect -2252 -234 -2236 -200
rect -2202 -234 -2044 -200
rect -2010 -234 -1852 -200
rect -1818 -234 -1660 -200
rect -1626 -234 -1468 -200
rect -1434 -234 -1276 -200
rect -1242 -234 -1226 -200
rect -2252 -254 -1226 -234
rect -2186 -276 -2156 -254
rect -2090 -276 -2060 -254
rect -1994 -276 -1964 -254
rect -1898 -276 -1868 -254
rect -1802 -276 -1772 -254
rect -1706 -276 -1676 -254
rect -1610 -276 -1580 -254
rect -1514 -276 -1484 -254
rect -1418 -276 -1388 -254
rect -1322 -276 -1292 -254
rect -2186 -406 -2156 -380
rect -2090 -406 -2060 -380
rect -1994 -406 -1964 -380
rect -1898 -406 -1868 -380
rect -1802 -406 -1772 -380
rect -1706 -406 -1676 -380
rect -1610 -406 -1580 -380
rect -1514 -406 -1484 -380
rect -1418 -406 -1388 -380
rect -1322 -406 -1292 -380
rect 419 -200 1445 -188
rect 419 -234 435 -200
rect 469 -234 627 -200
rect 661 -234 819 -200
rect 853 -234 1011 -200
rect 1045 -234 1203 -200
rect 1237 -234 1395 -200
rect 1429 -234 1445 -200
rect 419 -254 1445 -234
rect 485 -276 515 -254
rect 581 -276 611 -254
rect 677 -276 707 -254
rect 773 -276 803 -254
rect 869 -276 899 -254
rect 965 -276 995 -254
rect 1061 -276 1091 -254
rect 1157 -276 1187 -254
rect 1253 -276 1283 -254
rect 1349 -276 1379 -254
rect 485 -406 515 -380
rect 581 -406 611 -380
rect 677 -406 707 -380
rect 773 -406 803 -380
rect 869 -406 899 -380
rect 965 -406 995 -380
rect 1061 -406 1091 -380
rect 1157 -406 1187 -380
rect 1253 -406 1283 -380
rect 1349 -406 1379 -380
rect 1661 -285 1691 -259
rect 1661 -407 1691 -385
rect 1940 -200 2966 -188
rect 1940 -234 1956 -200
rect 1990 -234 2148 -200
rect 2182 -234 2340 -200
rect 2374 -234 2532 -200
rect 2566 -234 2724 -200
rect 2758 -234 2916 -200
rect 2950 -234 2966 -200
rect 1940 -254 2966 -234
rect 2006 -276 2036 -254
rect 2102 -276 2132 -254
rect 2198 -276 2228 -254
rect 2294 -276 2324 -254
rect 2390 -276 2420 -254
rect 2486 -276 2516 -254
rect 2582 -276 2612 -254
rect 2678 -276 2708 -254
rect 2774 -276 2804 -254
rect 2870 -276 2900 -254
rect 1643 -423 1709 -407
rect 1643 -457 1659 -423
rect 1693 -457 1709 -423
rect 1643 -473 1709 -457
rect 2006 -406 2036 -380
rect 2102 -406 2132 -380
rect 2198 -406 2228 -380
rect 2294 -406 2324 -380
rect 2390 -406 2420 -380
rect 2486 -406 2516 -380
rect 2582 -406 2612 -380
rect 2678 -406 2708 -380
rect 2774 -406 2804 -380
rect 2870 -406 2900 -380
rect -2186 -688 -2156 -662
rect -2090 -688 -2060 -662
rect -1994 -688 -1964 -662
rect -1898 -688 -1868 -662
rect -1802 -688 -1772 -662
rect -1706 -688 -1676 -662
rect -1610 -688 -1580 -662
rect -1514 -688 -1484 -662
rect -1418 -688 -1388 -662
rect -1322 -688 -1292 -662
rect -2186 -992 -2156 -960
rect -2090 -992 -2060 -960
rect -1994 -992 -1964 -960
rect -1898 -992 -1868 -960
rect -1802 -992 -1772 -960
rect -1706 -992 -1676 -960
rect -1610 -992 -1580 -960
rect -1514 -992 -1484 -960
rect -1418 -992 -1388 -960
rect -1322 -992 -1292 -960
rect -2252 -1008 -1226 -992
rect -2252 -1042 -2236 -1008
rect -2202 -1042 -2044 -1008
rect -2010 -1042 -1852 -1008
rect -1818 -1042 -1660 -1008
rect -1626 -1042 -1468 -1008
rect -1434 -1042 -1276 -1008
rect -1242 -1042 -1226 -1008
rect -2252 -1058 -1226 -1042
rect -339 -699 -309 -673
rect -339 -851 -309 -829
rect -395 -867 -309 -851
rect -395 -901 -379 -867
rect -345 -901 -309 -867
rect -395 -917 -309 -901
rect -339 -949 -309 -917
rect 485 -688 515 -662
rect 581 -688 611 -662
rect 677 -688 707 -662
rect 773 -688 803 -662
rect 869 -688 899 -662
rect 965 -688 995 -662
rect 1061 -688 1091 -662
rect 1157 -688 1187 -662
rect 1253 -688 1283 -662
rect 1349 -688 1379 -662
rect 485 -992 515 -960
rect 581 -992 611 -960
rect 677 -992 707 -960
rect 773 -992 803 -960
rect 869 -992 899 -960
rect 965 -992 995 -960
rect 1061 -992 1091 -960
rect 1157 -992 1187 -960
rect 1253 -992 1283 -960
rect 1349 -992 1379 -960
rect 419 -1008 1445 -992
rect 419 -1042 435 -1008
rect 469 -1042 627 -1008
rect 661 -1042 819 -1008
rect 853 -1042 1011 -1008
rect 1045 -1042 1203 -1008
rect 1237 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 419 -1058 1445 -1042
rect 2006 -688 2036 -662
rect 2102 -688 2132 -662
rect 2198 -688 2228 -662
rect 2294 -688 2324 -662
rect 2390 -688 2420 -662
rect 2486 -688 2516 -662
rect 2582 -688 2612 -662
rect 2678 -688 2708 -662
rect 2774 -688 2804 -662
rect 2870 -688 2900 -662
rect 2006 -992 2036 -960
rect 2102 -992 2132 -960
rect 2198 -992 2228 -960
rect 2294 -992 2324 -960
rect 2390 -992 2420 -960
rect 2486 -992 2516 -960
rect 2582 -992 2612 -960
rect 2678 -992 2708 -960
rect 2774 -992 2804 -960
rect 2870 -992 2900 -960
rect 1940 -1008 2966 -992
rect 1940 -1042 1956 -1008
rect 1990 -1042 2148 -1008
rect 2182 -1042 2340 -1008
rect 2374 -1042 2532 -1008
rect 2566 -1042 2724 -1008
rect 2758 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1940 -1058 2966 -1042
rect -339 -1175 -309 -1149
rect -339 -1243 -309 -1217
rect -2252 -1352 -1226 -1336
rect -2252 -1386 -2236 -1352
rect -2202 -1386 -2044 -1352
rect -2010 -1386 -1852 -1352
rect -1818 -1386 -1660 -1352
rect -1626 -1386 -1468 -1352
rect -1434 -1386 -1276 -1352
rect -1242 -1386 -1226 -1352
rect -2252 -1402 -1226 -1386
rect -2186 -1434 -2156 -1402
rect -2090 -1434 -2060 -1402
rect -1994 -1434 -1964 -1402
rect -1898 -1434 -1868 -1402
rect -1802 -1434 -1772 -1402
rect -1706 -1434 -1676 -1402
rect -1610 -1434 -1580 -1402
rect -1514 -1434 -1484 -1402
rect -1418 -1434 -1388 -1402
rect -1322 -1434 -1292 -1402
rect -2186 -1732 -2156 -1706
rect -2090 -1732 -2060 -1706
rect -1994 -1732 -1964 -1706
rect -1898 -1732 -1868 -1706
rect -1802 -1732 -1772 -1706
rect -1706 -1732 -1676 -1706
rect -1610 -1732 -1580 -1706
rect -1514 -1732 -1484 -1706
rect -1418 -1732 -1388 -1706
rect -1322 -1732 -1292 -1706
rect -339 -1475 -309 -1443
rect -395 -1491 -309 -1475
rect -395 -1525 -379 -1491
rect -345 -1525 -309 -1491
rect -395 -1541 -309 -1525
rect -339 -1563 -309 -1541
rect -339 -1719 -309 -1693
rect 419 -1534 1445 -1522
rect 419 -1568 435 -1534
rect 469 -1568 627 -1534
rect 661 -1568 819 -1534
rect 853 -1568 1011 -1534
rect 1045 -1568 1203 -1534
rect 1237 -1568 1395 -1534
rect 1429 -1568 1445 -1534
rect 419 -1588 1445 -1568
rect 485 -1610 515 -1588
rect 581 -1610 611 -1588
rect 677 -1610 707 -1588
rect 773 -1610 803 -1588
rect 869 -1610 899 -1588
rect 965 -1610 995 -1588
rect 1061 -1610 1091 -1588
rect 1157 -1610 1187 -1588
rect 1253 -1610 1283 -1588
rect 1349 -1610 1379 -1588
rect 485 -1740 515 -1714
rect 581 -1740 611 -1714
rect 677 -1740 707 -1714
rect 773 -1740 803 -1714
rect 869 -1740 899 -1714
rect 965 -1740 995 -1714
rect 1061 -1740 1091 -1714
rect 1157 -1740 1187 -1714
rect 1253 -1740 1283 -1714
rect 1349 -1740 1379 -1714
rect 1661 -1619 1691 -1593
rect 1661 -1741 1691 -1719
rect 1940 -1534 2966 -1522
rect 1940 -1568 1956 -1534
rect 1990 -1568 2148 -1534
rect 2182 -1568 2340 -1534
rect 2374 -1568 2532 -1534
rect 2566 -1568 2724 -1534
rect 2758 -1568 2916 -1534
rect 2950 -1568 2966 -1534
rect 1940 -1588 2966 -1568
rect 2006 -1610 2036 -1588
rect 2102 -1610 2132 -1588
rect 2198 -1610 2228 -1588
rect 2294 -1610 2324 -1588
rect 2390 -1610 2420 -1588
rect 2486 -1610 2516 -1588
rect 2582 -1610 2612 -1588
rect 2678 -1610 2708 -1588
rect 2774 -1610 2804 -1588
rect 2870 -1610 2900 -1588
rect 1643 -1757 1709 -1741
rect 1643 -1791 1659 -1757
rect 1693 -1791 1709 -1757
rect 1643 -1807 1709 -1791
rect 2006 -1740 2036 -1714
rect 2102 -1740 2132 -1714
rect 2198 -1740 2228 -1714
rect 2294 -1740 2324 -1714
rect 2390 -1740 2420 -1714
rect 2486 -1740 2516 -1714
rect 2582 -1740 2612 -1714
rect 2678 -1740 2708 -1714
rect 2774 -1740 2804 -1714
rect 2870 -1740 2900 -1714
rect -2186 -2014 -2156 -1988
rect -2090 -2014 -2060 -1988
rect -1994 -2014 -1964 -1988
rect -1898 -2014 -1868 -1988
rect -1802 -2014 -1772 -1988
rect -1706 -2014 -1676 -1988
rect -1610 -2014 -1580 -1988
rect -1514 -2014 -1484 -1988
rect -1418 -2014 -1388 -1988
rect -1322 -2014 -1292 -1988
rect -2186 -2140 -2156 -2118
rect -2090 -2140 -2060 -2118
rect -1994 -2140 -1964 -2118
rect -1898 -2140 -1868 -2118
rect -1802 -2140 -1772 -2118
rect -1706 -2140 -1676 -2118
rect -1610 -2140 -1580 -2118
rect -1514 -2140 -1484 -2118
rect -1418 -2140 -1388 -2118
rect -1322 -2140 -1292 -2118
rect -2252 -2160 -1226 -2140
rect -2252 -2194 -2236 -2160
rect -2202 -2194 -2044 -2160
rect -2010 -2194 -1852 -2160
rect -1818 -2194 -1660 -2160
rect -1626 -2194 -1468 -2160
rect -1434 -2194 -1276 -2160
rect -1242 -2194 -1226 -2160
rect -2252 -2206 -1226 -2194
rect 485 -2022 515 -1996
rect 581 -2022 611 -1996
rect 677 -2022 707 -1996
rect 773 -2022 803 -1996
rect 869 -2022 899 -1996
rect 965 -2022 995 -1996
rect 1061 -2022 1091 -1996
rect 1157 -2022 1187 -1996
rect 1253 -2022 1283 -1996
rect 1349 -2022 1379 -1996
rect 485 -2326 515 -2294
rect 581 -2326 611 -2294
rect 677 -2326 707 -2294
rect 773 -2326 803 -2294
rect 869 -2326 899 -2294
rect 965 -2326 995 -2294
rect 1061 -2326 1091 -2294
rect 1157 -2326 1187 -2294
rect 1253 -2326 1283 -2294
rect 1349 -2326 1379 -2294
rect 419 -2342 1445 -2326
rect 419 -2376 435 -2342
rect 469 -2376 627 -2342
rect 661 -2376 819 -2342
rect 853 -2376 1011 -2342
rect 1045 -2376 1203 -2342
rect 1237 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 419 -2392 1445 -2376
rect 2006 -2022 2036 -1996
rect 2102 -2022 2132 -1996
rect 2198 -2022 2228 -1996
rect 2294 -2022 2324 -1996
rect 2390 -2022 2420 -1996
rect 2486 -2022 2516 -1996
rect 2582 -2022 2612 -1996
rect 2678 -2022 2708 -1996
rect 2774 -2022 2804 -1996
rect 2870 -2022 2900 -1996
rect 2006 -2326 2036 -2294
rect 2102 -2326 2132 -2294
rect 2198 -2326 2228 -2294
rect 2294 -2326 2324 -2294
rect 2390 -2326 2420 -2294
rect 2486 -2326 2516 -2294
rect 2582 -2326 2612 -2294
rect 2678 -2326 2708 -2294
rect 2774 -2326 2804 -2294
rect 2870 -2326 2900 -2294
rect 1940 -2342 2966 -2326
rect 1940 -2376 1956 -2342
rect 1990 -2376 2148 -2342
rect 2182 -2376 2340 -2342
rect 2374 -2376 2532 -2342
rect 2566 -2376 2724 -2342
rect 2758 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1940 -2392 2966 -2376
<< polycont >>
rect -2236 -234 -2202 -200
rect -2044 -234 -2010 -200
rect -1852 -234 -1818 -200
rect -1660 -234 -1626 -200
rect -1468 -234 -1434 -200
rect -1276 -234 -1242 -200
rect 435 -234 469 -200
rect 627 -234 661 -200
rect 819 -234 853 -200
rect 1011 -234 1045 -200
rect 1203 -234 1237 -200
rect 1395 -234 1429 -200
rect 1956 -234 1990 -200
rect 2148 -234 2182 -200
rect 2340 -234 2374 -200
rect 2532 -234 2566 -200
rect 2724 -234 2758 -200
rect 2916 -234 2950 -200
rect 1659 -457 1693 -423
rect -2236 -1042 -2202 -1008
rect -2044 -1042 -2010 -1008
rect -1852 -1042 -1818 -1008
rect -1660 -1042 -1626 -1008
rect -1468 -1042 -1434 -1008
rect -1276 -1042 -1242 -1008
rect -379 -901 -345 -867
rect 435 -1042 469 -1008
rect 627 -1042 661 -1008
rect 819 -1042 853 -1008
rect 1011 -1042 1045 -1008
rect 1203 -1042 1237 -1008
rect 1395 -1042 1429 -1008
rect 1956 -1042 1990 -1008
rect 2148 -1042 2182 -1008
rect 2340 -1042 2374 -1008
rect 2532 -1042 2566 -1008
rect 2724 -1042 2758 -1008
rect 2916 -1042 2950 -1008
rect -2236 -1386 -2202 -1352
rect -2044 -1386 -2010 -1352
rect -1852 -1386 -1818 -1352
rect -1660 -1386 -1626 -1352
rect -1468 -1386 -1434 -1352
rect -1276 -1386 -1242 -1352
rect -379 -1525 -345 -1491
rect 435 -1568 469 -1534
rect 627 -1568 661 -1534
rect 819 -1568 853 -1534
rect 1011 -1568 1045 -1534
rect 1203 -1568 1237 -1534
rect 1395 -1568 1429 -1534
rect 1956 -1568 1990 -1534
rect 2148 -1568 2182 -1534
rect 2340 -1568 2374 -1534
rect 2532 -1568 2566 -1534
rect 2724 -1568 2758 -1534
rect 2916 -1568 2950 -1534
rect 1659 -1791 1693 -1757
rect -2236 -2194 -2202 -2160
rect -2044 -2194 -2010 -2160
rect -1852 -2194 -1818 -2160
rect -1660 -2194 -1626 -2160
rect -1468 -2194 -1434 -2160
rect -1276 -2194 -1242 -2160
rect 435 -2376 469 -2342
rect 627 -2376 661 -2342
rect 819 -2376 853 -2342
rect 1011 -2376 1045 -2342
rect 1203 -2376 1237 -2342
rect 1395 -2376 1429 -2342
rect 1956 -2376 1990 -2342
rect 2148 -2376 2182 -2342
rect 2340 -2376 2374 -2342
rect 2532 -2376 2566 -2342
rect 2724 -2376 2758 -2342
rect 2916 -2376 2950 -2342
<< locali >>
rect -2350 -136 -2254 -102
rect -1224 -136 -1128 -102
rect -2350 -198 -2316 -136
rect -1162 -198 -1128 -136
rect -2252 -234 -2236 -200
rect -2202 -234 -2186 -200
rect -2060 -234 -2044 -200
rect -2010 -234 -1994 -200
rect -1868 -234 -1852 -200
rect -1818 -234 -1802 -200
rect -1676 -234 -1660 -200
rect -1626 -234 -1610 -200
rect -1484 -234 -1468 -200
rect -1434 -234 -1418 -200
rect -1292 -234 -1276 -200
rect -1242 -234 -1226 -200
rect -2236 -288 -2202 -272
rect -2236 -384 -2202 -368
rect -2140 -288 -2106 -272
rect -2140 -384 -2106 -368
rect -2044 -288 -2010 -272
rect -2044 -384 -2010 -368
rect -1948 -288 -1914 -272
rect -1948 -384 -1914 -368
rect -1852 -288 -1818 -272
rect -1852 -384 -1818 -368
rect -1756 -288 -1722 -272
rect -1756 -384 -1722 -368
rect -1660 -288 -1626 -272
rect -1660 -384 -1626 -368
rect -1564 -288 -1530 -272
rect -1564 -384 -1530 -368
rect -1468 -288 -1434 -272
rect -1468 -384 -1434 -368
rect -1372 -288 -1338 -272
rect -1372 -384 -1338 -368
rect -1276 -288 -1242 -272
rect -1276 -384 -1242 -368
rect -2350 -458 -2316 -396
rect -1162 -458 -1128 -398
rect -2350 -492 -2254 -458
rect -1224 -492 -1128 -458
rect 321 -136 417 -102
rect 1447 -136 1543 -102
rect 321 -198 355 -136
rect 1509 -198 1543 -136
rect 419 -234 435 -200
rect 469 -234 485 -200
rect 611 -234 627 -200
rect 661 -234 677 -200
rect 803 -234 819 -200
rect 853 -234 869 -200
rect 995 -234 1011 -200
rect 1045 -234 1061 -200
rect 1187 -234 1203 -200
rect 1237 -234 1253 -200
rect 1379 -234 1395 -200
rect 1429 -234 1445 -200
rect 435 -288 469 -272
rect 435 -384 469 -368
rect 531 -288 565 -272
rect 531 -384 565 -368
rect 627 -288 661 -272
rect 627 -384 661 -368
rect 723 -288 757 -272
rect 723 -384 757 -368
rect 819 -288 853 -272
rect 819 -384 853 -368
rect 915 -288 949 -272
rect 915 -384 949 -368
rect 1011 -288 1045 -272
rect 1011 -384 1045 -368
rect 1107 -288 1141 -272
rect 1107 -384 1141 -368
rect 1203 -288 1237 -272
rect 1203 -384 1237 -368
rect 1299 -288 1333 -272
rect 1299 -384 1333 -368
rect 1395 -288 1429 -272
rect 1395 -384 1429 -368
rect 321 -458 355 -396
rect 1842 -136 1938 -102
rect 2968 -136 3064 -102
rect 1842 -198 1876 -136
rect 1615 -297 1649 -281
rect 1615 -389 1649 -373
rect 1703 -297 1737 -281
rect 1703 -389 1737 -373
rect 1509 -458 1543 -398
rect 3030 -198 3064 -136
rect 1940 -234 1956 -200
rect 1990 -234 2006 -200
rect 2132 -234 2148 -200
rect 2182 -234 2198 -200
rect 2324 -234 2340 -200
rect 2374 -234 2390 -200
rect 2516 -234 2532 -200
rect 2566 -234 2582 -200
rect 2708 -234 2724 -200
rect 2758 -234 2774 -200
rect 2900 -234 2916 -200
rect 2950 -234 2966 -200
rect 1956 -288 1990 -272
rect 1956 -384 1990 -368
rect 2052 -288 2086 -272
rect 2052 -384 2086 -368
rect 2148 -288 2182 -272
rect 2148 -384 2182 -368
rect 2244 -288 2278 -272
rect 2244 -384 2278 -368
rect 2340 -288 2374 -272
rect 2340 -384 2374 -368
rect 2436 -288 2470 -272
rect 2436 -384 2470 -368
rect 2532 -288 2566 -272
rect 2532 -384 2566 -368
rect 2628 -288 2662 -272
rect 2628 -384 2662 -368
rect 2724 -288 2758 -272
rect 2724 -384 2758 -368
rect 2820 -288 2854 -272
rect 2820 -384 2854 -368
rect 2916 -288 2950 -272
rect 2916 -384 2950 -368
rect 1643 -457 1659 -423
rect 1693 -457 1709 -423
rect 321 -492 417 -458
rect 1447 -492 1543 -458
rect 1842 -458 1876 -396
rect 3030 -458 3064 -398
rect 1842 -492 1938 -458
rect 2968 -492 3064 -458
rect -2350 -600 -2254 -566
rect -1224 -600 -1128 -566
rect -2350 -662 -2316 -600
rect -1162 -662 -1128 -600
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect -2236 -700 -2202 -684
rect -2236 -964 -2202 -948
rect -2140 -700 -2106 -684
rect -2140 -964 -2106 -948
rect -2044 -700 -2010 -684
rect -2044 -964 -2010 -948
rect -1948 -700 -1914 -684
rect -1948 -964 -1914 -948
rect -1852 -700 -1818 -684
rect -1852 -964 -1818 -948
rect -1756 -700 -1722 -684
rect -1756 -964 -1722 -948
rect -1660 -700 -1626 -684
rect -1660 -964 -1626 -948
rect -1564 -700 -1530 -684
rect -1564 -964 -1530 -948
rect -1468 -700 -1434 -684
rect -1468 -964 -1434 -948
rect -1372 -700 -1338 -684
rect -1372 -964 -1338 -948
rect -1276 -700 -1242 -684
rect -1276 -964 -1242 -948
rect -2252 -1042 -2236 -1008
rect -2202 -1042 -2186 -1008
rect -2060 -1042 -2044 -1008
rect -2010 -1042 -1994 -1008
rect -1868 -1042 -1852 -1008
rect -1818 -1042 -1802 -1008
rect -1676 -1042 -1660 -1008
rect -1626 -1042 -1610 -1008
rect -1484 -1042 -1468 -1008
rect -1434 -1042 -1418 -1008
rect -1292 -1042 -1276 -1008
rect -1242 -1042 -1226 -1008
rect -2350 -1110 -2316 -1048
rect -551 -669 -522 -635
rect -488 -669 -430 -635
rect -396 -669 -338 -635
rect -304 -669 -246 -635
rect -212 -669 -183 -635
rect 321 -662 355 -600
rect -534 -763 -476 -669
rect -534 -797 -522 -763
rect -488 -797 -476 -763
rect -534 -814 -476 -797
rect -395 -715 -349 -669
rect -395 -749 -383 -715
rect -395 -783 -349 -749
rect -395 -817 -383 -783
rect -395 -833 -349 -817
rect -315 -715 -249 -703
rect -315 -749 -299 -715
rect -265 -749 -249 -715
rect -315 -778 -249 -749
rect -315 -783 -298 -778
rect -315 -817 -299 -783
rect -264 -812 -249 -778
rect -265 -817 -249 -812
rect -315 -829 -249 -817
rect -395 -873 -379 -867
rect -395 -907 -381 -873
rect -345 -901 -329 -867
rect -347 -907 -329 -901
rect -395 -915 -329 -907
rect -1162 -1110 -1128 -1048
rect -2350 -1144 -2254 -1110
rect -1224 -1144 -1128 -1110
rect -534 -981 -476 -946
rect -295 -949 -249 -829
rect -534 -1015 -522 -981
rect -488 -1015 -476 -981
rect -534 -1074 -476 -1015
rect -534 -1108 -522 -1074
rect -488 -1108 -476 -1074
rect -534 -1179 -476 -1108
rect -391 -967 -349 -951
rect -391 -1001 -383 -967
rect -391 -1035 -349 -1001
rect -391 -1069 -383 -1035
rect -391 -1103 -349 -1069
rect -391 -1137 -383 -1103
rect -391 -1179 -349 -1137
rect -315 -967 -249 -949
rect -315 -1001 -299 -967
rect -265 -1001 -249 -967
rect -315 -1035 -249 -1001
rect -315 -1069 -299 -1035
rect -265 -1069 -249 -1035
rect -315 -1103 -249 -1069
rect -315 -1137 -299 -1103
rect -265 -1137 -249 -1103
rect -315 -1145 -249 -1137
rect 1509 -662 1543 -600
rect 435 -700 469 -684
rect 435 -964 469 -948
rect 531 -700 565 -684
rect 531 -964 565 -948
rect 627 -700 661 -684
rect 627 -964 661 -948
rect 723 -700 757 -684
rect 723 -964 757 -948
rect 819 -700 853 -684
rect 819 -964 853 -948
rect 915 -700 949 -684
rect 915 -964 949 -948
rect 1011 -700 1045 -684
rect 1011 -964 1045 -948
rect 1107 -700 1141 -684
rect 1107 -964 1141 -948
rect 1203 -700 1237 -684
rect 1203 -964 1237 -948
rect 1299 -700 1333 -684
rect 1299 -964 1333 -948
rect 1395 -700 1429 -684
rect 1395 -964 1429 -948
rect 419 -1042 435 -1008
rect 469 -1042 485 -1008
rect 611 -1042 627 -1008
rect 661 -1042 677 -1008
rect 803 -1042 819 -1008
rect 853 -1042 869 -1008
rect 995 -1042 1011 -1008
rect 1045 -1042 1061 -1008
rect 1187 -1042 1203 -1008
rect 1237 -1042 1253 -1008
rect 1379 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 321 -1110 355 -1048
rect 1509 -1110 1543 -1048
rect 321 -1144 417 -1110
rect 1447 -1144 1543 -1110
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1956 -700 1990 -684
rect 1956 -964 1990 -948
rect 2052 -700 2086 -684
rect 2052 -964 2086 -948
rect 2148 -700 2182 -684
rect 2148 -964 2182 -948
rect 2244 -700 2278 -684
rect 2244 -964 2278 -948
rect 2340 -700 2374 -684
rect 2340 -964 2374 -948
rect 2436 -700 2470 -684
rect 2436 -964 2470 -948
rect 2532 -700 2566 -684
rect 2532 -964 2566 -948
rect 2628 -700 2662 -684
rect 2628 -964 2662 -948
rect 2724 -700 2758 -684
rect 2724 -964 2758 -948
rect 2820 -700 2854 -684
rect 2820 -964 2854 -948
rect 2916 -700 2950 -684
rect 2916 -964 2950 -948
rect 1940 -1042 1956 -1008
rect 1990 -1042 2006 -1008
rect 2132 -1042 2148 -1008
rect 2182 -1042 2198 -1008
rect 2324 -1042 2340 -1008
rect 2374 -1042 2390 -1008
rect 2516 -1042 2532 -1008
rect 2566 -1042 2582 -1008
rect 2708 -1042 2724 -1008
rect 2758 -1042 2774 -1008
rect 2900 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1842 -1110 1876 -1048
rect 3030 -1110 3064 -1048
rect 1842 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect -551 -1213 -522 -1179
rect -488 -1213 -430 -1179
rect -396 -1213 -338 -1179
rect -304 -1213 -246 -1179
rect -212 -1213 -183 -1179
rect -2350 -1284 -2254 -1250
rect -1224 -1284 -1128 -1250
rect -2350 -1346 -2316 -1284
rect -1162 -1346 -1128 -1284
rect -2252 -1386 -2236 -1352
rect -2202 -1386 -2186 -1352
rect -2060 -1386 -2044 -1352
rect -2010 -1386 -1994 -1352
rect -1868 -1386 -1852 -1352
rect -1818 -1386 -1802 -1352
rect -1676 -1386 -1660 -1352
rect -1626 -1386 -1610 -1352
rect -1484 -1386 -1468 -1352
rect -1434 -1386 -1418 -1352
rect -1292 -1386 -1276 -1352
rect -1242 -1386 -1226 -1352
rect -2236 -1446 -2202 -1430
rect -2236 -1710 -2202 -1694
rect -2140 -1446 -2106 -1430
rect -2140 -1710 -2106 -1694
rect -2044 -1446 -2010 -1430
rect -2044 -1710 -2010 -1694
rect -1948 -1446 -1914 -1430
rect -1948 -1710 -1914 -1694
rect -1852 -1446 -1818 -1430
rect -1852 -1710 -1818 -1694
rect -1756 -1446 -1722 -1430
rect -1756 -1710 -1722 -1694
rect -1660 -1446 -1626 -1430
rect -1660 -1710 -1626 -1694
rect -1564 -1446 -1530 -1430
rect -1564 -1710 -1530 -1694
rect -1468 -1446 -1434 -1430
rect -1468 -1710 -1434 -1694
rect -1372 -1446 -1338 -1430
rect -1372 -1710 -1338 -1694
rect -1276 -1446 -1242 -1430
rect -1276 -1710 -1242 -1694
rect -2350 -1794 -2316 -1732
rect -534 -1284 -476 -1213
rect -534 -1318 -522 -1284
rect -488 -1318 -476 -1284
rect -534 -1377 -476 -1318
rect -534 -1411 -522 -1377
rect -488 -1411 -476 -1377
rect -534 -1446 -476 -1411
rect -391 -1255 -349 -1213
rect -391 -1289 -383 -1255
rect -391 -1323 -349 -1289
rect -391 -1357 -383 -1323
rect -391 -1391 -349 -1357
rect -391 -1425 -383 -1391
rect -391 -1441 -349 -1425
rect -315 -1255 -249 -1247
rect -315 -1289 -299 -1255
rect -265 -1289 -249 -1255
rect -315 -1323 -249 -1289
rect -315 -1382 -299 -1323
rect -265 -1382 -249 -1323
rect -315 -1391 -249 -1382
rect -315 -1425 -299 -1391
rect -265 -1425 -249 -1391
rect -315 -1443 -249 -1425
rect -395 -1486 -329 -1477
rect -395 -1520 -382 -1486
rect -348 -1491 -329 -1486
rect -395 -1525 -379 -1520
rect -345 -1525 -329 -1491
rect -395 -1575 -349 -1559
rect -295 -1563 -249 -1443
rect -534 -1595 -476 -1578
rect -534 -1629 -522 -1595
rect -488 -1629 -476 -1595
rect -534 -1723 -476 -1629
rect -395 -1609 -383 -1575
rect -395 -1643 -349 -1609
rect -395 -1677 -383 -1643
rect -395 -1723 -349 -1677
rect -315 -1575 -249 -1563
rect -315 -1609 -299 -1575
rect -265 -1609 -249 -1575
rect -315 -1643 -249 -1609
rect -315 -1677 -299 -1643
rect -265 -1677 -249 -1643
rect -315 -1689 -249 -1677
rect 321 -1470 417 -1436
rect 1447 -1470 1543 -1436
rect 321 -1532 355 -1470
rect -1162 -1794 -1128 -1732
rect -551 -1757 -522 -1723
rect -488 -1757 -430 -1723
rect -396 -1757 -338 -1723
rect -304 -1757 -246 -1723
rect -212 -1757 -183 -1723
rect 1509 -1532 1543 -1470
rect 419 -1568 435 -1534
rect 469 -1568 485 -1534
rect 611 -1568 627 -1534
rect 661 -1568 677 -1534
rect 803 -1568 819 -1534
rect 853 -1568 869 -1534
rect 995 -1568 1011 -1534
rect 1045 -1568 1061 -1534
rect 1187 -1568 1203 -1534
rect 1237 -1568 1253 -1534
rect 1379 -1568 1395 -1534
rect 1429 -1568 1445 -1534
rect 435 -1622 469 -1606
rect 435 -1718 469 -1702
rect 531 -1622 565 -1606
rect 531 -1718 565 -1702
rect 627 -1622 661 -1606
rect 627 -1718 661 -1702
rect 723 -1622 757 -1606
rect 723 -1718 757 -1702
rect 819 -1622 853 -1606
rect 819 -1718 853 -1702
rect 915 -1622 949 -1606
rect 915 -1718 949 -1702
rect 1011 -1622 1045 -1606
rect 1011 -1718 1045 -1702
rect 1107 -1622 1141 -1606
rect 1107 -1718 1141 -1702
rect 1203 -1622 1237 -1606
rect 1203 -1718 1237 -1702
rect 1299 -1622 1333 -1606
rect 1299 -1718 1333 -1702
rect 1395 -1622 1429 -1606
rect 1395 -1718 1429 -1702
rect -2350 -1828 -2254 -1794
rect -1224 -1828 -1128 -1794
rect 321 -1792 355 -1730
rect 1842 -1470 1938 -1436
rect 2968 -1470 3064 -1436
rect 1842 -1532 1876 -1470
rect 1615 -1631 1649 -1615
rect 1615 -1723 1649 -1707
rect 1703 -1631 1737 -1615
rect 1703 -1723 1737 -1707
rect 1509 -1792 1543 -1732
rect 3030 -1532 3064 -1470
rect 1940 -1568 1956 -1534
rect 1990 -1568 2006 -1534
rect 2132 -1568 2148 -1534
rect 2182 -1568 2198 -1534
rect 2324 -1568 2340 -1534
rect 2374 -1568 2390 -1534
rect 2516 -1568 2532 -1534
rect 2566 -1568 2582 -1534
rect 2708 -1568 2724 -1534
rect 2758 -1568 2774 -1534
rect 2900 -1568 2916 -1534
rect 2950 -1568 2966 -1534
rect 1956 -1622 1990 -1606
rect 1956 -1718 1990 -1702
rect 2052 -1622 2086 -1606
rect 2052 -1718 2086 -1702
rect 2148 -1622 2182 -1606
rect 2148 -1718 2182 -1702
rect 2244 -1622 2278 -1606
rect 2244 -1718 2278 -1702
rect 2340 -1622 2374 -1606
rect 2340 -1718 2374 -1702
rect 2436 -1622 2470 -1606
rect 2436 -1718 2470 -1702
rect 2532 -1622 2566 -1606
rect 2532 -1718 2566 -1702
rect 2628 -1622 2662 -1606
rect 2628 -1718 2662 -1702
rect 2724 -1622 2758 -1606
rect 2724 -1718 2758 -1702
rect 2820 -1622 2854 -1606
rect 2820 -1718 2854 -1702
rect 2916 -1622 2950 -1606
rect 2916 -1718 2950 -1702
rect 1643 -1791 1659 -1757
rect 1693 -1791 1709 -1757
rect 321 -1826 417 -1792
rect 1447 -1826 1543 -1792
rect 1842 -1792 1876 -1730
rect 3030 -1792 3064 -1732
rect 1842 -1826 1938 -1792
rect 2968 -1826 3064 -1792
rect -2350 -1936 -2254 -1902
rect -1224 -1936 -1128 -1902
rect -2350 -1998 -2316 -1936
rect -1162 -1996 -1128 -1936
rect -2236 -2026 -2202 -2010
rect -2236 -2122 -2202 -2106
rect -2140 -2026 -2106 -2010
rect -2140 -2122 -2106 -2106
rect -2044 -2026 -2010 -2010
rect -2044 -2122 -2010 -2106
rect -1948 -2026 -1914 -2010
rect -1948 -2122 -1914 -2106
rect -1852 -2026 -1818 -2010
rect -1852 -2122 -1818 -2106
rect -1756 -2026 -1722 -2010
rect -1756 -2122 -1722 -2106
rect -1660 -2026 -1626 -2010
rect -1660 -2122 -1626 -2106
rect -1564 -2026 -1530 -2010
rect -1564 -2122 -1530 -2106
rect -1468 -2026 -1434 -2010
rect -1468 -2122 -1434 -2106
rect -1372 -2026 -1338 -2010
rect -1372 -2122 -1338 -2106
rect -1276 -2026 -1242 -2010
rect -1276 -2122 -1242 -2106
rect -2252 -2194 -2236 -2160
rect -2202 -2194 -2186 -2160
rect -2060 -2194 -2044 -2160
rect -2010 -2194 -1994 -2160
rect -1868 -2194 -1852 -2160
rect -1818 -2194 -1802 -2160
rect -1676 -2194 -1660 -2160
rect -1626 -2194 -1610 -2160
rect -1484 -2194 -1468 -2160
rect -1434 -2194 -1418 -2160
rect -1292 -2194 -1276 -2160
rect -1242 -2194 -1226 -2160
rect -2350 -2258 -2316 -2196
rect -1162 -2258 -1128 -2196
rect -2350 -2292 -2254 -2258
rect -1224 -2292 -1128 -2258
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect 435 -2034 469 -2018
rect 435 -2298 469 -2282
rect 531 -2034 565 -2018
rect 531 -2298 565 -2282
rect 627 -2034 661 -2018
rect 627 -2298 661 -2282
rect 723 -2034 757 -2018
rect 723 -2298 757 -2282
rect 819 -2034 853 -2018
rect 819 -2298 853 -2282
rect 915 -2034 949 -2018
rect 915 -2298 949 -2282
rect 1011 -2034 1045 -2018
rect 1011 -2298 1045 -2282
rect 1107 -2034 1141 -2018
rect 1107 -2298 1141 -2282
rect 1203 -2034 1237 -2018
rect 1203 -2298 1237 -2282
rect 1299 -2034 1333 -2018
rect 1299 -2298 1333 -2282
rect 1395 -2034 1429 -2018
rect 1395 -2298 1429 -2282
rect 419 -2376 435 -2342
rect 469 -2376 485 -2342
rect 611 -2376 627 -2342
rect 661 -2376 677 -2342
rect 803 -2376 819 -2342
rect 853 -2376 869 -2342
rect 995 -2376 1011 -2342
rect 1045 -2376 1061 -2342
rect 1187 -2376 1203 -2342
rect 1237 -2376 1253 -2342
rect 1379 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 321 -2444 355 -2382
rect 1509 -2444 1543 -2382
rect 321 -2478 417 -2444
rect 1447 -2478 1543 -2444
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1956 -2034 1990 -2018
rect 1956 -2298 1990 -2282
rect 2052 -2034 2086 -2018
rect 2052 -2298 2086 -2282
rect 2148 -2034 2182 -2018
rect 2148 -2298 2182 -2282
rect 2244 -2034 2278 -2018
rect 2244 -2298 2278 -2282
rect 2340 -2034 2374 -2018
rect 2340 -2298 2374 -2282
rect 2436 -2034 2470 -2018
rect 2436 -2298 2470 -2282
rect 2532 -2034 2566 -2018
rect 2532 -2298 2566 -2282
rect 2628 -2034 2662 -2018
rect 2628 -2298 2662 -2282
rect 2724 -2034 2758 -2018
rect 2724 -2298 2758 -2282
rect 2820 -2034 2854 -2018
rect 2820 -2298 2854 -2282
rect 2916 -2034 2950 -2018
rect 2916 -2298 2950 -2282
rect 1940 -2376 1956 -2342
rect 1990 -2376 2006 -2342
rect 2132 -2376 2148 -2342
rect 2182 -2376 2198 -2342
rect 2324 -2376 2340 -2342
rect 2374 -2376 2390 -2342
rect 2516 -2376 2532 -2342
rect 2566 -2376 2582 -2342
rect 2708 -2376 2724 -2342
rect 2758 -2376 2774 -2342
rect 2900 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1842 -2444 1876 -2382
rect 3030 -2444 3064 -2382
rect 1842 -2478 1938 -2444
rect 2968 -2478 3064 -2444
<< viali >>
rect -2236 -234 -2202 -200
rect -2044 -234 -2010 -200
rect -1852 -234 -1818 -200
rect -1660 -234 -1626 -200
rect -1468 -234 -1434 -200
rect -1276 -234 -1242 -200
rect -2236 -368 -2202 -288
rect -2140 -368 -2106 -288
rect -2044 -368 -2010 -288
rect -1948 -368 -1914 -288
rect -1852 -368 -1818 -288
rect -1756 -368 -1722 -288
rect -1660 -368 -1626 -288
rect -1564 -368 -1530 -288
rect -1468 -368 -1434 -288
rect -1372 -368 -1338 -288
rect -1276 -368 -1242 -288
rect -1162 -396 -1128 -198
rect -1162 -398 -1128 -396
rect 435 -234 469 -200
rect 627 -234 661 -200
rect 819 -234 853 -200
rect 1011 -234 1045 -200
rect 1203 -234 1237 -200
rect 1395 -234 1429 -200
rect 435 -368 469 -288
rect 531 -368 565 -288
rect 627 -368 661 -288
rect 723 -368 757 -288
rect 819 -368 853 -288
rect 915 -368 949 -288
rect 1011 -368 1045 -288
rect 1107 -368 1141 -288
rect 1203 -368 1237 -288
rect 1299 -368 1333 -288
rect 1395 -368 1429 -288
rect 1509 -396 1543 -198
rect 1615 -373 1649 -297
rect 1703 -373 1737 -297
rect 1509 -398 1543 -396
rect 1956 -234 1990 -200
rect 2148 -234 2182 -200
rect 2340 -234 2374 -200
rect 2532 -234 2566 -200
rect 2724 -234 2758 -200
rect 2916 -234 2950 -200
rect 1956 -368 1990 -288
rect 2052 -368 2086 -288
rect 2148 -368 2182 -288
rect 2244 -368 2278 -288
rect 2340 -368 2374 -288
rect 2436 -368 2470 -288
rect 2532 -368 2566 -288
rect 2628 -368 2662 -288
rect 2724 -368 2758 -288
rect 2820 -368 2854 -288
rect 2916 -368 2950 -288
rect 1659 -457 1693 -423
rect 3030 -396 3064 -198
rect 3030 -398 3064 -396
rect -2236 -948 -2202 -700
rect -2140 -948 -2106 -700
rect -2044 -948 -2010 -700
rect -1948 -948 -1914 -700
rect -1852 -948 -1818 -700
rect -1756 -948 -1722 -700
rect -1660 -948 -1626 -700
rect -1564 -948 -1530 -700
rect -1468 -948 -1434 -700
rect -1372 -948 -1338 -700
rect -1276 -948 -1242 -700
rect -2236 -1042 -2202 -1008
rect -2044 -1042 -2010 -1008
rect -1852 -1042 -1818 -1008
rect -1660 -1042 -1626 -1008
rect -1468 -1042 -1434 -1008
rect -1276 -1042 -1242 -1008
rect -1162 -1048 -1128 -662
rect -522 -669 -488 -635
rect -430 -669 -396 -635
rect -338 -669 -304 -635
rect -246 -669 -212 -635
rect -298 -783 -264 -778
rect -298 -812 -265 -783
rect -265 -812 -264 -783
rect -381 -901 -379 -873
rect -379 -901 -347 -873
rect -381 -907 -347 -901
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect 435 -1042 469 -1008
rect 627 -1042 661 -1008
rect 819 -1042 853 -1008
rect 1011 -1042 1045 -1008
rect 1203 -1042 1237 -1008
rect 1395 -1042 1429 -1008
rect 1509 -1048 1543 -662
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect 1956 -1042 1990 -1008
rect 2148 -1042 2182 -1008
rect 2340 -1042 2374 -1008
rect 2532 -1042 2566 -1008
rect 2724 -1042 2758 -1008
rect 2916 -1042 2950 -1008
rect 3030 -1048 3064 -662
rect -522 -1213 -488 -1179
rect -430 -1213 -396 -1179
rect -338 -1213 -304 -1179
rect -246 -1213 -212 -1179
rect -2236 -1386 -2202 -1352
rect -2044 -1386 -2010 -1352
rect -1852 -1386 -1818 -1352
rect -1660 -1386 -1626 -1352
rect -1468 -1386 -1434 -1352
rect -1276 -1386 -1242 -1352
rect -2236 -1694 -2202 -1446
rect -2140 -1694 -2106 -1446
rect -2044 -1694 -2010 -1446
rect -1948 -1694 -1914 -1446
rect -1852 -1694 -1818 -1446
rect -1756 -1694 -1722 -1446
rect -1660 -1694 -1626 -1446
rect -1564 -1694 -1530 -1446
rect -1468 -1694 -1434 -1446
rect -1372 -1694 -1338 -1446
rect -1276 -1694 -1242 -1446
rect -1162 -1732 -1128 -1346
rect -299 -1357 -265 -1348
rect -299 -1382 -265 -1357
rect -382 -1491 -348 -1486
rect -382 -1520 -379 -1491
rect -379 -1520 -348 -1491
rect -522 -1757 -488 -1723
rect -430 -1757 -396 -1723
rect -338 -1757 -304 -1723
rect -246 -1757 -212 -1723
rect 435 -1568 469 -1534
rect 627 -1568 661 -1534
rect 819 -1568 853 -1534
rect 1011 -1568 1045 -1534
rect 1203 -1568 1237 -1534
rect 1395 -1568 1429 -1534
rect 435 -1702 469 -1622
rect 531 -1702 565 -1622
rect 627 -1702 661 -1622
rect 723 -1702 757 -1622
rect 819 -1702 853 -1622
rect 915 -1702 949 -1622
rect 1011 -1702 1045 -1622
rect 1107 -1702 1141 -1622
rect 1203 -1702 1237 -1622
rect 1299 -1702 1333 -1622
rect 1395 -1702 1429 -1622
rect 1509 -1730 1543 -1532
rect 1615 -1707 1649 -1631
rect 1703 -1707 1737 -1631
rect 1509 -1732 1543 -1730
rect 1956 -1568 1990 -1534
rect 2148 -1568 2182 -1534
rect 2340 -1568 2374 -1534
rect 2532 -1568 2566 -1534
rect 2724 -1568 2758 -1534
rect 2916 -1568 2950 -1534
rect 1956 -1702 1990 -1622
rect 2052 -1702 2086 -1622
rect 2148 -1702 2182 -1622
rect 2244 -1702 2278 -1622
rect 2340 -1702 2374 -1622
rect 2436 -1702 2470 -1622
rect 2532 -1702 2566 -1622
rect 2628 -1702 2662 -1622
rect 2724 -1702 2758 -1622
rect 2820 -1702 2854 -1622
rect 2916 -1702 2950 -1622
rect 1659 -1791 1693 -1757
rect 3030 -1730 3064 -1532
rect 3030 -1732 3064 -1730
rect -1162 -1998 -1128 -1996
rect -2236 -2106 -2202 -2026
rect -2140 -2106 -2106 -2026
rect -2044 -2106 -2010 -2026
rect -1948 -2106 -1914 -2026
rect -1852 -2106 -1818 -2026
rect -1756 -2106 -1722 -2026
rect -1660 -2106 -1626 -2026
rect -1564 -2106 -1530 -2026
rect -1468 -2106 -1434 -2026
rect -1372 -2106 -1338 -2026
rect -1276 -2106 -1242 -2026
rect -2236 -2194 -2202 -2160
rect -2044 -2194 -2010 -2160
rect -1852 -2194 -1818 -2160
rect -1660 -2194 -1626 -2160
rect -1468 -2194 -1434 -2160
rect -1276 -2194 -1242 -2160
rect -1162 -2196 -1128 -1998
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 435 -2376 469 -2342
rect 627 -2376 661 -2342
rect 819 -2376 853 -2342
rect 1011 -2376 1045 -2342
rect 1203 -2376 1237 -2342
rect 1395 -2376 1429 -2342
rect 1509 -2382 1543 -1996
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
rect 1956 -2376 1990 -2342
rect 2148 -2376 2182 -2342
rect 2340 -2376 2374 -2342
rect 2532 -2376 2566 -2342
rect 2724 -2376 2758 -2342
rect 2916 -2376 2950 -2342
rect 3030 -2382 3064 -1996
<< metal1 >>
rect -2420 -136 -1338 -102
rect -2549 -245 -2522 -193
rect -2470 -245 -2460 -193
rect -2420 -513 -2386 -136
rect -2252 -193 -2186 -188
rect -2255 -245 -2245 -193
rect -2193 -245 -2183 -193
rect -2252 -248 -2186 -245
rect -2140 -276 -2106 -136
rect -2060 -193 -1994 -188
rect -2064 -245 -2054 -193
rect -2002 -245 -1992 -193
rect -2060 -248 -1994 -245
rect -1948 -276 -1914 -136
rect -1868 -193 -1802 -188
rect -1872 -245 -1862 -193
rect -1810 -245 -1800 -193
rect -1868 -248 -1802 -245
rect -1756 -276 -1722 -136
rect -1676 -193 -1610 -188
rect -1680 -245 -1670 -193
rect -1618 -245 -1608 -193
rect -1676 -248 -1610 -245
rect -1564 -276 -1530 -136
rect -1484 -192 -1418 -188
rect -1487 -244 -1477 -192
rect -1425 -244 -1415 -192
rect -1484 -248 -1418 -244
rect -1372 -276 -1338 -136
rect -1292 -192 -1226 -188
rect -1295 -244 -1285 -192
rect -1233 -244 -1223 -192
rect -1168 -198 -1122 -24
rect 251 -136 1333 -102
rect -1292 -248 -1226 -244
rect -2242 -288 -2196 -276
rect -2242 -368 -2236 -288
rect -2202 -368 -2196 -288
rect -2242 -380 -2196 -368
rect -2146 -288 -2100 -276
rect -2146 -368 -2140 -288
rect -2106 -368 -2100 -288
rect -2146 -380 -2100 -368
rect -2050 -288 -2004 -276
rect -2050 -368 -2044 -288
rect -2010 -368 -2004 -288
rect -2050 -380 -2004 -368
rect -1954 -288 -1908 -276
rect -1954 -368 -1948 -288
rect -1914 -368 -1908 -288
rect -1954 -380 -1908 -368
rect -1858 -288 -1812 -276
rect -1858 -368 -1852 -288
rect -1818 -368 -1812 -288
rect -1858 -380 -1812 -368
rect -1762 -288 -1716 -276
rect -1762 -368 -1756 -288
rect -1722 -368 -1716 -288
rect -1762 -380 -1716 -368
rect -1666 -288 -1620 -276
rect -1666 -368 -1660 -288
rect -1626 -368 -1620 -288
rect -1666 -380 -1620 -368
rect -1570 -288 -1524 -276
rect -1570 -368 -1564 -288
rect -1530 -368 -1524 -288
rect -1570 -380 -1524 -368
rect -1474 -288 -1428 -276
rect -1474 -368 -1468 -288
rect -1434 -368 -1428 -288
rect -1474 -380 -1428 -368
rect -1378 -288 -1332 -276
rect -1378 -368 -1372 -288
rect -1338 -368 -1332 -288
rect -1378 -380 -1332 -368
rect -1282 -288 -1236 -276
rect -1282 -368 -1276 -288
rect -1242 -368 -1236 -288
rect -1282 -380 -1236 -368
rect -2638 -547 -2386 -513
rect -2549 -1052 -2522 -1000
rect -2470 -1052 -2460 -1000
rect -2420 -1110 -2386 -547
rect -2236 -513 -2202 -380
rect -2044 -513 -2010 -380
rect -1852 -513 -1818 -380
rect -1660 -513 -1626 -380
rect -1468 -513 -1434 -380
rect -1276 -513 -1242 -380
rect -1168 -398 -1162 -198
rect -1128 -398 -1122 -198
rect 70 -245 149 -193
rect 201 -245 211 -193
rect -1168 -410 -1122 -398
rect -1046 -479 104 -445
rect -1046 -513 -1012 -479
rect -2236 -547 -1012 -513
rect 70 -513 104 -479
rect 251 -513 285 -136
rect 419 -193 485 -188
rect 416 -245 426 -193
rect 478 -245 488 -193
rect 419 -248 485 -245
rect 531 -276 565 -136
rect 611 -193 677 -188
rect 607 -245 617 -193
rect 669 -245 679 -193
rect 611 -248 677 -245
rect 723 -276 757 -136
rect 803 -193 869 -188
rect 799 -245 809 -193
rect 861 -245 871 -193
rect 803 -248 869 -245
rect 915 -276 949 -136
rect 995 -193 1061 -188
rect 991 -245 1001 -193
rect 1053 -245 1063 -193
rect 995 -248 1061 -245
rect 1107 -276 1141 -136
rect 1187 -192 1253 -188
rect 1184 -244 1194 -192
rect 1246 -244 1256 -192
rect 1187 -248 1253 -244
rect 1299 -276 1333 -136
rect 1379 -192 1445 -188
rect 1376 -244 1386 -192
rect 1438 -244 1448 -192
rect 1503 -198 1549 8
rect 1772 -136 2854 -102
rect 1379 -248 1445 -244
rect 429 -288 475 -276
rect 429 -368 435 -288
rect 469 -368 475 -288
rect 429 -380 475 -368
rect 525 -288 571 -276
rect 525 -368 531 -288
rect 565 -368 571 -288
rect 525 -380 571 -368
rect 621 -288 667 -276
rect 621 -368 627 -288
rect 661 -368 667 -288
rect 621 -380 667 -368
rect 717 -288 763 -276
rect 717 -368 723 -288
rect 757 -368 763 -288
rect 717 -380 763 -368
rect 813 -288 859 -276
rect 813 -368 819 -288
rect 853 -368 859 -288
rect 813 -380 859 -368
rect 909 -288 955 -276
rect 909 -368 915 -288
rect 949 -368 955 -288
rect 909 -380 955 -368
rect 1005 -288 1051 -276
rect 1005 -368 1011 -288
rect 1045 -368 1051 -288
rect 1005 -380 1051 -368
rect 1101 -288 1147 -276
rect 1101 -368 1107 -288
rect 1141 -368 1147 -288
rect 1101 -380 1147 -368
rect 1197 -288 1243 -276
rect 1197 -368 1203 -288
rect 1237 -368 1243 -288
rect 1197 -380 1243 -368
rect 1293 -288 1339 -276
rect 1293 -368 1299 -288
rect 1333 -368 1339 -288
rect 1293 -380 1339 -368
rect 1389 -288 1435 -276
rect 1389 -368 1395 -288
rect 1429 -368 1435 -288
rect 1389 -380 1435 -368
rect 70 -547 285 -513
rect -2236 -688 -2202 -547
rect -2044 -688 -2010 -547
rect -1852 -688 -1818 -547
rect -1660 -688 -1626 -547
rect -1468 -688 -1434 -547
rect -1276 -688 -1242 -547
rect -624 -635 -183 -604
rect -1168 -662 -1122 -650
rect -2242 -700 -2196 -688
rect -2242 -948 -2236 -700
rect -2202 -948 -2196 -700
rect -2242 -960 -2196 -948
rect -2146 -700 -2100 -688
rect -2146 -948 -2140 -700
rect -2106 -948 -2100 -700
rect -2146 -960 -2100 -948
rect -2050 -700 -2004 -688
rect -2050 -948 -2044 -700
rect -2010 -948 -2004 -700
rect -2050 -960 -2004 -948
rect -1954 -700 -1908 -688
rect -1954 -948 -1948 -700
rect -1914 -948 -1908 -700
rect -1954 -960 -1908 -948
rect -1858 -700 -1812 -688
rect -1858 -948 -1852 -700
rect -1818 -948 -1812 -700
rect -1858 -960 -1812 -948
rect -1762 -700 -1716 -688
rect -1762 -948 -1756 -700
rect -1722 -948 -1716 -700
rect -1762 -960 -1716 -948
rect -1666 -700 -1620 -688
rect -1666 -948 -1660 -700
rect -1626 -948 -1620 -700
rect -1666 -960 -1620 -948
rect -1570 -700 -1524 -688
rect -1570 -948 -1564 -700
rect -1530 -948 -1524 -700
rect -1570 -960 -1524 -948
rect -1474 -700 -1428 -688
rect -1474 -948 -1468 -700
rect -1434 -948 -1428 -700
rect -1474 -960 -1428 -948
rect -1378 -700 -1332 -688
rect -1378 -948 -1372 -700
rect -1338 -948 -1332 -700
rect -1378 -960 -1332 -948
rect -1282 -700 -1236 -688
rect -1282 -948 -1276 -700
rect -1242 -948 -1236 -700
rect -1282 -960 -1236 -948
rect -2255 -1052 -2245 -1000
rect -2193 -1052 -2183 -1000
rect -2140 -1110 -2106 -960
rect -2062 -1052 -2052 -1000
rect -2000 -1052 -1990 -1000
rect -1948 -1110 -1914 -960
rect -1871 -1052 -1861 -1000
rect -1809 -1052 -1799 -1000
rect -1756 -1110 -1722 -960
rect -1679 -1052 -1669 -1000
rect -1617 -1052 -1607 -1000
rect -1564 -1110 -1530 -960
rect -1487 -1052 -1477 -1000
rect -1425 -1052 -1415 -1000
rect -1372 -1110 -1338 -960
rect -1295 -1052 -1285 -1000
rect -1233 -1052 -1223 -1000
rect -1168 -1048 -1162 -662
rect -1128 -1048 -1122 -662
rect -624 -669 -522 -635
rect -488 -669 -430 -635
rect -396 -669 -338 -635
rect -304 -669 -246 -635
rect -212 -669 -183 -635
rect -624 -700 -183 -669
rect -43 -772 -33 -769
rect -310 -778 -33 -772
rect -310 -812 -298 -778
rect -264 -812 -33 -778
rect -310 -818 -33 -812
rect -43 -821 -33 -818
rect 19 -821 29 -769
rect -401 -917 -391 -865
rect -339 -917 -329 -865
rect -2420 -1144 -1338 -1110
rect -1168 -1174 -1122 -1048
rect -176 -1052 -166 -1000
rect -114 -1052 149 -1000
rect 201 -1052 211 -1000
rect 251 -1110 285 -547
rect 435 -513 469 -380
rect 627 -513 661 -380
rect 819 -513 853 -380
rect 1011 -513 1045 -380
rect 1203 -513 1237 -380
rect 1395 -513 1429 -380
rect 1503 -398 1509 -198
rect 1543 -285 1549 -198
rect 1643 -245 1670 -193
rect 1722 -245 1732 -193
rect 1772 -285 1806 -136
rect 1940 -193 2006 -188
rect 1937 -245 1947 -193
rect 1999 -245 2009 -193
rect 1940 -248 2006 -245
rect 2052 -276 2086 -136
rect 2132 -193 2198 -188
rect 2128 -245 2138 -193
rect 2190 -245 2200 -193
rect 2132 -248 2198 -245
rect 2244 -276 2278 -136
rect 2324 -193 2390 -188
rect 2320 -245 2330 -193
rect 2382 -245 2392 -193
rect 2324 -248 2390 -245
rect 2436 -276 2470 -136
rect 2516 -193 2582 -188
rect 2512 -245 2522 -193
rect 2574 -245 2584 -193
rect 2516 -248 2582 -245
rect 2628 -276 2662 -136
rect 2708 -192 2774 -188
rect 2705 -244 2715 -192
rect 2767 -244 2777 -192
rect 2708 -248 2774 -244
rect 2820 -276 2854 -136
rect 2900 -192 2966 -188
rect 2897 -244 2907 -192
rect 2959 -244 2969 -192
rect 3024 -198 3070 15
rect 2900 -248 2966 -244
rect 1543 -297 1655 -285
rect 1543 -373 1615 -297
rect 1649 -373 1655 -297
rect 1543 -385 1655 -373
rect 1697 -297 1806 -285
rect 1697 -373 1703 -297
rect 1737 -373 1806 -297
rect 1697 -385 1806 -373
rect 1950 -288 1996 -276
rect 1950 -368 1956 -288
rect 1990 -368 1996 -288
rect 1950 -380 1996 -368
rect 2046 -288 2092 -276
rect 2046 -368 2052 -288
rect 2086 -368 2092 -288
rect 2046 -380 2092 -368
rect 2142 -288 2188 -276
rect 2142 -368 2148 -288
rect 2182 -368 2188 -288
rect 2142 -380 2188 -368
rect 2238 -288 2284 -276
rect 2238 -368 2244 -288
rect 2278 -368 2284 -288
rect 2238 -380 2284 -368
rect 2334 -288 2380 -276
rect 2334 -368 2340 -288
rect 2374 -368 2380 -288
rect 2334 -380 2380 -368
rect 2430 -288 2476 -276
rect 2430 -368 2436 -288
rect 2470 -368 2476 -288
rect 2430 -380 2476 -368
rect 2526 -288 2572 -276
rect 2526 -368 2532 -288
rect 2566 -368 2572 -288
rect 2526 -380 2572 -368
rect 2622 -288 2668 -276
rect 2622 -368 2628 -288
rect 2662 -368 2668 -288
rect 2622 -380 2668 -368
rect 2718 -288 2764 -276
rect 2718 -368 2724 -288
rect 2758 -368 2764 -288
rect 2718 -380 2764 -368
rect 2814 -288 2860 -276
rect 2814 -368 2820 -288
rect 2854 -368 2860 -288
rect 2814 -380 2860 -368
rect 2910 -288 2956 -276
rect 2910 -368 2916 -288
rect 2950 -368 2956 -288
rect 2910 -380 2956 -368
rect 1543 -398 1549 -385
rect 1503 -410 1549 -398
rect 1647 -423 1705 -417
rect 1640 -475 1650 -423
rect 1702 -475 1712 -423
rect 1772 -513 1806 -385
rect 435 -547 1806 -513
rect 435 -688 469 -547
rect 627 -688 661 -547
rect 819 -688 853 -547
rect 1011 -688 1045 -547
rect 1203 -688 1237 -547
rect 1395 -688 1429 -547
rect 1503 -662 1549 -650
rect 429 -700 475 -688
rect 429 -948 435 -700
rect 469 -948 475 -700
rect 429 -960 475 -948
rect 525 -700 571 -688
rect 525 -948 531 -700
rect 565 -948 571 -700
rect 525 -960 571 -948
rect 621 -700 667 -688
rect 621 -948 627 -700
rect 661 -948 667 -700
rect 621 -960 667 -948
rect 717 -700 763 -688
rect 717 -948 723 -700
rect 757 -948 763 -700
rect 717 -960 763 -948
rect 813 -700 859 -688
rect 813 -948 819 -700
rect 853 -948 859 -700
rect 813 -960 859 -948
rect 909 -700 955 -688
rect 909 -948 915 -700
rect 949 -948 955 -700
rect 909 -960 955 -948
rect 1005 -700 1051 -688
rect 1005 -948 1011 -700
rect 1045 -948 1051 -700
rect 1005 -960 1051 -948
rect 1101 -700 1147 -688
rect 1101 -948 1107 -700
rect 1141 -948 1147 -700
rect 1101 -960 1147 -948
rect 1197 -700 1243 -688
rect 1197 -948 1203 -700
rect 1237 -948 1243 -700
rect 1197 -960 1243 -948
rect 1293 -700 1339 -688
rect 1293 -948 1299 -700
rect 1333 -948 1339 -700
rect 1293 -960 1339 -948
rect 1389 -700 1435 -688
rect 1389 -948 1395 -700
rect 1429 -948 1435 -700
rect 1389 -960 1435 -948
rect 416 -1052 426 -1000
rect 478 -1052 488 -1000
rect 531 -1110 565 -960
rect 609 -1052 619 -1000
rect 671 -1052 681 -1000
rect 723 -1110 757 -960
rect 800 -1052 810 -1000
rect 862 -1052 872 -1000
rect 915 -1110 949 -960
rect 992 -1052 1002 -1000
rect 1054 -1052 1064 -1000
rect 1107 -1110 1141 -960
rect 1184 -1052 1194 -1000
rect 1246 -1052 1256 -1000
rect 1299 -1110 1333 -960
rect 1376 -1052 1386 -1000
rect 1438 -1052 1448 -1000
rect 1503 -1048 1509 -662
rect 1543 -1048 1549 -662
rect 251 -1144 1333 -1110
rect -1168 -1220 -1045 -1174
rect -624 -1179 -183 -1148
rect -624 -1213 -522 -1179
rect -488 -1213 -430 -1179
rect -396 -1213 -338 -1179
rect -304 -1213 -246 -1179
rect -212 -1213 -183 -1179
rect -2420 -1284 -1338 -1250
rect -2549 -1394 -2522 -1342
rect -2470 -1394 -2460 -1342
rect -2420 -1847 -2386 -1284
rect -2255 -1394 -2245 -1342
rect -2193 -1394 -2183 -1342
rect -2140 -1434 -2106 -1284
rect -2062 -1394 -2052 -1342
rect -2000 -1394 -1990 -1342
rect -1948 -1434 -1914 -1284
rect -1871 -1394 -1861 -1342
rect -1809 -1394 -1799 -1342
rect -1756 -1434 -1722 -1284
rect -1679 -1394 -1669 -1342
rect -1617 -1394 -1607 -1342
rect -1564 -1434 -1530 -1284
rect -1487 -1394 -1477 -1342
rect -1425 -1394 -1415 -1342
rect -1372 -1434 -1338 -1284
rect -1295 -1394 -1285 -1342
rect -1233 -1394 -1223 -1342
rect -1168 -1346 -1122 -1220
rect -624 -1244 -183 -1213
rect 1503 -1248 1549 -1048
rect 1643 -1052 1670 -1000
rect 1722 -1052 1732 -1000
rect 1772 -1110 1806 -547
rect 1956 -513 1990 -380
rect 2148 -513 2182 -380
rect 2340 -513 2374 -380
rect 2532 -513 2566 -380
rect 2724 -513 2758 -380
rect 2916 -513 2950 -380
rect 3024 -398 3030 -198
rect 3064 -398 3070 -198
rect 3024 -410 3070 -398
rect 1956 -547 3258 -513
rect 1956 -688 1990 -547
rect 2148 -688 2182 -547
rect 2340 -688 2374 -547
rect 2532 -688 2566 -547
rect 2724 -688 2758 -547
rect 2916 -688 2950 -547
rect 3024 -662 3070 -650
rect 1950 -700 1996 -688
rect 1950 -948 1956 -700
rect 1990 -948 1996 -700
rect 1950 -960 1996 -948
rect 2046 -700 2092 -688
rect 2046 -948 2052 -700
rect 2086 -948 2092 -700
rect 2046 -960 2092 -948
rect 2142 -700 2188 -688
rect 2142 -948 2148 -700
rect 2182 -948 2188 -700
rect 2142 -960 2188 -948
rect 2238 -700 2284 -688
rect 2238 -948 2244 -700
rect 2278 -948 2284 -700
rect 2238 -960 2284 -948
rect 2334 -700 2380 -688
rect 2334 -948 2340 -700
rect 2374 -948 2380 -700
rect 2334 -960 2380 -948
rect 2430 -700 2476 -688
rect 2430 -948 2436 -700
rect 2470 -948 2476 -700
rect 2430 -960 2476 -948
rect 2526 -700 2572 -688
rect 2526 -948 2532 -700
rect 2566 -948 2572 -700
rect 2526 -960 2572 -948
rect 2622 -700 2668 -688
rect 2622 -948 2628 -700
rect 2662 -948 2668 -700
rect 2622 -960 2668 -948
rect 2718 -700 2764 -688
rect 2718 -948 2724 -700
rect 2758 -948 2764 -700
rect 2718 -960 2764 -948
rect 2814 -700 2860 -688
rect 2814 -948 2820 -700
rect 2854 -948 2860 -700
rect 2814 -960 2860 -948
rect 2910 -700 2956 -688
rect 2910 -948 2916 -700
rect 2950 -948 2956 -700
rect 2910 -960 2956 -948
rect 1937 -1052 1947 -1000
rect 1999 -1052 2009 -1000
rect 2052 -1110 2086 -960
rect 2130 -1052 2140 -1000
rect 2192 -1052 2202 -1000
rect 2244 -1110 2278 -960
rect 2321 -1052 2331 -1000
rect 2383 -1052 2393 -1000
rect 2436 -1110 2470 -960
rect 2513 -1052 2523 -1000
rect 2575 -1052 2585 -1000
rect 2628 -1110 2662 -960
rect 2705 -1052 2715 -1000
rect 2767 -1052 2777 -1000
rect 2820 -1110 2854 -960
rect 2897 -1052 2907 -1000
rect 2959 -1052 2969 -1000
rect 3024 -1048 3030 -662
rect 3064 -1048 3070 -662
rect 1772 -1144 2854 -1110
rect 3024 -1246 3070 -1048
rect 3224 -1270 3258 -547
rect 3224 -1304 3429 -1270
rect -2242 -1446 -2196 -1434
rect -2242 -1694 -2236 -1446
rect -2202 -1694 -2196 -1446
rect -2242 -1706 -2196 -1694
rect -2146 -1446 -2100 -1434
rect -2146 -1694 -2140 -1446
rect -2106 -1694 -2100 -1446
rect -2146 -1706 -2100 -1694
rect -2050 -1446 -2004 -1434
rect -2050 -1694 -2044 -1446
rect -2010 -1694 -2004 -1446
rect -2050 -1706 -2004 -1694
rect -1954 -1446 -1908 -1434
rect -1954 -1694 -1948 -1446
rect -1914 -1694 -1908 -1446
rect -1954 -1706 -1908 -1694
rect -1858 -1446 -1812 -1434
rect -1858 -1694 -1852 -1446
rect -1818 -1694 -1812 -1446
rect -1858 -1706 -1812 -1694
rect -1762 -1446 -1716 -1434
rect -1762 -1694 -1756 -1446
rect -1722 -1694 -1716 -1446
rect -1762 -1706 -1716 -1694
rect -1666 -1446 -1620 -1434
rect -1666 -1694 -1660 -1446
rect -1626 -1694 -1620 -1446
rect -1666 -1706 -1620 -1694
rect -1570 -1446 -1524 -1434
rect -1570 -1694 -1564 -1446
rect -1530 -1694 -1524 -1446
rect -1570 -1706 -1524 -1694
rect -1474 -1446 -1428 -1434
rect -1474 -1694 -1468 -1446
rect -1434 -1694 -1428 -1446
rect -1474 -1706 -1428 -1694
rect -1378 -1446 -1332 -1434
rect -1378 -1694 -1372 -1446
rect -1338 -1694 -1332 -1446
rect -1378 -1706 -1332 -1694
rect -1282 -1446 -1236 -1434
rect -1282 -1694 -1276 -1446
rect -1242 -1694 -1236 -1446
rect -1282 -1706 -1236 -1694
rect -2638 -1881 -2386 -1847
rect -2549 -2201 -2522 -2149
rect -2470 -2201 -2460 -2149
rect -2420 -2258 -2386 -1881
rect -2236 -1847 -2202 -1706
rect -2044 -1847 -2010 -1706
rect -1852 -1847 -1818 -1706
rect -1660 -1847 -1626 -1706
rect -1468 -1847 -1434 -1706
rect -1276 -1847 -1242 -1706
rect -1168 -1732 -1162 -1346
rect -1128 -1732 -1122 -1346
rect -965 -1394 -955 -1342
rect -903 -1348 -253 -1342
rect -903 -1382 -299 -1348
rect -265 -1382 -253 -1348
rect -903 -1388 -253 -1382
rect -903 -1394 -893 -1388
rect 251 -1470 1333 -1436
rect -401 -1530 -391 -1478
rect -339 -1530 -329 -1478
rect 70 -1579 149 -1527
rect 201 -1579 211 -1527
rect -1168 -1744 -1122 -1732
rect -624 -1723 -183 -1692
rect -624 -1757 -522 -1723
rect -488 -1757 -430 -1723
rect -396 -1757 -338 -1723
rect -304 -1757 -246 -1723
rect -212 -1757 -183 -1723
rect -624 -1788 -183 -1757
rect 251 -1847 285 -1470
rect 419 -1527 485 -1522
rect 416 -1579 426 -1527
rect 478 -1579 488 -1527
rect 419 -1582 485 -1579
rect 531 -1610 565 -1470
rect 611 -1527 677 -1522
rect 607 -1579 617 -1527
rect 669 -1579 679 -1527
rect 611 -1582 677 -1579
rect 723 -1610 757 -1470
rect 803 -1527 869 -1522
rect 799 -1579 809 -1527
rect 861 -1579 871 -1527
rect 803 -1582 869 -1579
rect 915 -1610 949 -1470
rect 995 -1527 1061 -1522
rect 991 -1579 1001 -1527
rect 1053 -1579 1063 -1527
rect 995 -1582 1061 -1579
rect 1107 -1610 1141 -1470
rect 1187 -1526 1253 -1522
rect 1184 -1578 1194 -1526
rect 1246 -1578 1256 -1526
rect 1187 -1582 1253 -1578
rect 1299 -1610 1333 -1470
rect 1379 -1526 1445 -1522
rect 1376 -1578 1386 -1526
rect 1438 -1578 1448 -1526
rect 1503 -1532 1549 -1334
rect 1772 -1470 2854 -1436
rect 1379 -1582 1445 -1578
rect 429 -1622 475 -1610
rect 429 -1702 435 -1622
rect 469 -1702 475 -1622
rect 429 -1714 475 -1702
rect 525 -1622 571 -1610
rect 525 -1702 531 -1622
rect 565 -1702 571 -1622
rect 525 -1714 571 -1702
rect 621 -1622 667 -1610
rect 621 -1702 627 -1622
rect 661 -1702 667 -1622
rect 621 -1714 667 -1702
rect 717 -1622 763 -1610
rect 717 -1702 723 -1622
rect 757 -1702 763 -1622
rect 717 -1714 763 -1702
rect 813 -1622 859 -1610
rect 813 -1702 819 -1622
rect 853 -1702 859 -1622
rect 813 -1714 859 -1702
rect 909 -1622 955 -1610
rect 909 -1702 915 -1622
rect 949 -1702 955 -1622
rect 909 -1714 955 -1702
rect 1005 -1622 1051 -1610
rect 1005 -1702 1011 -1622
rect 1045 -1702 1051 -1622
rect 1005 -1714 1051 -1702
rect 1101 -1622 1147 -1610
rect 1101 -1702 1107 -1622
rect 1141 -1702 1147 -1622
rect 1101 -1714 1147 -1702
rect 1197 -1622 1243 -1610
rect 1197 -1702 1203 -1622
rect 1237 -1702 1243 -1622
rect 1197 -1714 1243 -1702
rect 1293 -1622 1339 -1610
rect 1293 -1702 1299 -1622
rect 1333 -1702 1339 -1622
rect 1293 -1714 1339 -1702
rect 1389 -1622 1435 -1610
rect 1389 -1702 1395 -1622
rect 1429 -1702 1435 -1622
rect 1389 -1714 1435 -1702
rect -2236 -1881 -989 -1847
rect -2236 -2014 -2202 -1881
rect -2044 -2014 -2010 -1881
rect -1852 -2014 -1818 -1881
rect -1660 -2014 -1626 -1881
rect -1468 -2014 -1434 -1881
rect -1276 -2014 -1242 -1881
rect -1168 -1996 -1122 -1984
rect -2242 -2026 -2196 -2014
rect -2242 -2106 -2236 -2026
rect -2202 -2106 -2196 -2026
rect -2242 -2118 -2196 -2106
rect -2146 -2026 -2100 -2014
rect -2146 -2106 -2140 -2026
rect -2106 -2106 -2100 -2026
rect -2146 -2118 -2100 -2106
rect -2050 -2026 -2004 -2014
rect -2050 -2106 -2044 -2026
rect -2010 -2106 -2004 -2026
rect -2050 -2118 -2004 -2106
rect -1954 -2026 -1908 -2014
rect -1954 -2106 -1948 -2026
rect -1914 -2106 -1908 -2026
rect -1954 -2118 -1908 -2106
rect -1858 -2026 -1812 -2014
rect -1858 -2106 -1852 -2026
rect -1818 -2106 -1812 -2026
rect -1858 -2118 -1812 -2106
rect -1762 -2026 -1716 -2014
rect -1762 -2106 -1756 -2026
rect -1722 -2106 -1716 -2026
rect -1762 -2118 -1716 -2106
rect -1666 -2026 -1620 -2014
rect -1666 -2106 -1660 -2026
rect -1626 -2106 -1620 -2026
rect -1666 -2118 -1620 -2106
rect -1570 -2026 -1524 -2014
rect -1570 -2106 -1564 -2026
rect -1530 -2106 -1524 -2026
rect -1570 -2118 -1524 -2106
rect -1474 -2026 -1428 -2014
rect -1474 -2106 -1468 -2026
rect -1434 -2106 -1428 -2026
rect -1474 -2118 -1428 -2106
rect -1378 -2026 -1332 -2014
rect -1378 -2106 -1372 -2026
rect -1338 -2106 -1332 -2026
rect -1378 -2118 -1332 -2106
rect -1282 -2026 -1236 -2014
rect -1282 -2106 -1276 -2026
rect -1242 -2106 -1236 -2026
rect -1282 -2118 -1236 -2106
rect -2252 -2149 -2186 -2146
rect -2255 -2201 -2245 -2149
rect -2193 -2201 -2183 -2149
rect -2252 -2206 -2186 -2201
rect -2140 -2258 -2106 -2118
rect -2060 -2149 -1994 -2146
rect -2064 -2201 -2054 -2149
rect -2002 -2201 -1992 -2149
rect -2060 -2206 -1994 -2201
rect -1948 -2258 -1914 -2118
rect -1868 -2149 -1802 -2146
rect -1872 -2201 -1862 -2149
rect -1810 -2201 -1800 -2149
rect -1868 -2206 -1802 -2201
rect -1756 -2258 -1722 -2118
rect -1676 -2149 -1610 -2146
rect -1680 -2201 -1670 -2149
rect -1618 -2201 -1608 -2149
rect -1676 -2206 -1610 -2201
rect -1564 -2258 -1530 -2118
rect -1484 -2150 -1418 -2146
rect -1487 -2202 -1477 -2150
rect -1425 -2202 -1415 -2150
rect -1484 -2206 -1418 -2202
rect -1372 -2258 -1338 -2118
rect -1292 -2150 -1226 -2146
rect -1295 -2202 -1285 -2150
rect -1233 -2202 -1223 -2150
rect -1168 -2196 -1162 -1996
rect -1128 -2196 -1122 -1996
rect -1023 -2007 -989 -1881
rect 69 -1881 285 -1847
rect 69 -2007 103 -1881
rect -1023 -2041 103 -2007
rect -1292 -2206 -1226 -2202
rect -2420 -2292 -1338 -2258
rect -1168 -2371 -1122 -2196
rect 70 -2386 149 -2334
rect 201 -2386 211 -2334
rect 251 -2444 285 -1881
rect 435 -1847 469 -1714
rect 627 -1847 661 -1714
rect 819 -1847 853 -1714
rect 1011 -1847 1045 -1714
rect 1203 -1847 1237 -1714
rect 1395 -1847 1429 -1714
rect 1503 -1732 1509 -1532
rect 1543 -1619 1549 -1532
rect 1643 -1579 1670 -1527
rect 1722 -1579 1732 -1527
rect 1772 -1619 1806 -1470
rect 1940 -1527 2006 -1522
rect 1937 -1579 1947 -1527
rect 1999 -1579 2009 -1527
rect 1940 -1582 2006 -1579
rect 2052 -1610 2086 -1470
rect 2132 -1527 2198 -1522
rect 2128 -1579 2138 -1527
rect 2190 -1579 2200 -1527
rect 2132 -1582 2198 -1579
rect 2244 -1610 2278 -1470
rect 2324 -1527 2390 -1522
rect 2320 -1579 2330 -1527
rect 2382 -1579 2392 -1527
rect 2324 -1582 2390 -1579
rect 2436 -1610 2470 -1470
rect 2516 -1527 2582 -1522
rect 2512 -1579 2522 -1527
rect 2574 -1579 2584 -1527
rect 2516 -1582 2582 -1579
rect 2628 -1610 2662 -1470
rect 2708 -1526 2774 -1522
rect 2705 -1578 2715 -1526
rect 2767 -1578 2777 -1526
rect 2708 -1582 2774 -1578
rect 2820 -1610 2854 -1470
rect 2900 -1526 2966 -1522
rect 2897 -1578 2907 -1526
rect 2959 -1578 2969 -1526
rect 3024 -1532 3070 -1336
rect 2900 -1582 2966 -1578
rect 1543 -1631 1655 -1619
rect 1543 -1707 1615 -1631
rect 1649 -1707 1655 -1631
rect 1543 -1719 1655 -1707
rect 1697 -1631 1806 -1619
rect 1697 -1707 1703 -1631
rect 1737 -1707 1806 -1631
rect 1697 -1719 1806 -1707
rect 1950 -1622 1996 -1610
rect 1950 -1702 1956 -1622
rect 1990 -1702 1996 -1622
rect 1950 -1714 1996 -1702
rect 2046 -1622 2092 -1610
rect 2046 -1702 2052 -1622
rect 2086 -1702 2092 -1622
rect 2046 -1714 2092 -1702
rect 2142 -1622 2188 -1610
rect 2142 -1702 2148 -1622
rect 2182 -1702 2188 -1622
rect 2142 -1714 2188 -1702
rect 2238 -1622 2284 -1610
rect 2238 -1702 2244 -1622
rect 2278 -1702 2284 -1622
rect 2238 -1714 2284 -1702
rect 2334 -1622 2380 -1610
rect 2334 -1702 2340 -1622
rect 2374 -1702 2380 -1622
rect 2334 -1714 2380 -1702
rect 2430 -1622 2476 -1610
rect 2430 -1702 2436 -1622
rect 2470 -1702 2476 -1622
rect 2430 -1714 2476 -1702
rect 2526 -1622 2572 -1610
rect 2526 -1702 2532 -1622
rect 2566 -1702 2572 -1622
rect 2526 -1714 2572 -1702
rect 2622 -1622 2668 -1610
rect 2622 -1702 2628 -1622
rect 2662 -1702 2668 -1622
rect 2622 -1714 2668 -1702
rect 2718 -1622 2764 -1610
rect 2718 -1702 2724 -1622
rect 2758 -1702 2764 -1622
rect 2718 -1714 2764 -1702
rect 2814 -1622 2860 -1610
rect 2814 -1702 2820 -1622
rect 2854 -1702 2860 -1622
rect 2814 -1714 2860 -1702
rect 2910 -1622 2956 -1610
rect 2910 -1702 2916 -1622
rect 2950 -1702 2956 -1622
rect 2910 -1714 2956 -1702
rect 1543 -1732 1549 -1719
rect 1503 -1744 1549 -1732
rect 1647 -1757 1705 -1751
rect 1640 -1809 1650 -1757
rect 1702 -1809 1712 -1757
rect 1772 -1847 1806 -1719
rect 435 -1881 1806 -1847
rect 435 -2022 469 -1881
rect 627 -2022 661 -1881
rect 819 -2022 853 -1881
rect 1011 -2022 1045 -1881
rect 1203 -2022 1237 -1881
rect 1395 -2022 1429 -1881
rect 1503 -1996 1549 -1984
rect 429 -2034 475 -2022
rect 429 -2282 435 -2034
rect 469 -2282 475 -2034
rect 429 -2294 475 -2282
rect 525 -2034 571 -2022
rect 525 -2282 531 -2034
rect 565 -2282 571 -2034
rect 525 -2294 571 -2282
rect 621 -2034 667 -2022
rect 621 -2282 627 -2034
rect 661 -2282 667 -2034
rect 621 -2294 667 -2282
rect 717 -2034 763 -2022
rect 717 -2282 723 -2034
rect 757 -2282 763 -2034
rect 717 -2294 763 -2282
rect 813 -2034 859 -2022
rect 813 -2282 819 -2034
rect 853 -2282 859 -2034
rect 813 -2294 859 -2282
rect 909 -2034 955 -2022
rect 909 -2282 915 -2034
rect 949 -2282 955 -2034
rect 909 -2294 955 -2282
rect 1005 -2034 1051 -2022
rect 1005 -2282 1011 -2034
rect 1045 -2282 1051 -2034
rect 1005 -2294 1051 -2282
rect 1101 -2034 1147 -2022
rect 1101 -2282 1107 -2034
rect 1141 -2282 1147 -2034
rect 1101 -2294 1147 -2282
rect 1197 -2034 1243 -2022
rect 1197 -2282 1203 -2034
rect 1237 -2282 1243 -2034
rect 1197 -2294 1243 -2282
rect 1293 -2034 1339 -2022
rect 1293 -2282 1299 -2034
rect 1333 -2282 1339 -2034
rect 1293 -2294 1339 -2282
rect 1389 -2034 1435 -2022
rect 1389 -2282 1395 -2034
rect 1429 -2282 1435 -2034
rect 1389 -2294 1435 -2282
rect 416 -2386 426 -2334
rect 478 -2386 488 -2334
rect 531 -2444 565 -2294
rect 609 -2386 619 -2334
rect 671 -2386 681 -2334
rect 723 -2444 757 -2294
rect 800 -2386 810 -2334
rect 862 -2386 872 -2334
rect 915 -2444 949 -2294
rect 992 -2386 1002 -2334
rect 1054 -2386 1064 -2334
rect 1107 -2444 1141 -2294
rect 1184 -2386 1194 -2334
rect 1246 -2386 1256 -2334
rect 1299 -2444 1333 -2294
rect 1376 -2386 1386 -2334
rect 1438 -2386 1448 -2334
rect 1503 -2382 1509 -1996
rect 1543 -2382 1549 -1996
rect 251 -2478 1333 -2444
rect 1503 -2585 1549 -2382
rect 1643 -2386 1670 -2334
rect 1722 -2386 1732 -2334
rect 1772 -2444 1806 -1881
rect 1956 -1847 1990 -1714
rect 2148 -1847 2182 -1714
rect 2340 -1847 2374 -1714
rect 2532 -1847 2566 -1714
rect 2724 -1847 2758 -1714
rect 2916 -1847 2950 -1714
rect 3024 -1732 3030 -1532
rect 3064 -1732 3070 -1532
rect 3024 -1744 3070 -1732
rect 3224 -1847 3258 -1304
rect 1956 -1881 3258 -1847
rect 1956 -2022 1990 -1881
rect 2148 -2022 2182 -1881
rect 2340 -2022 2374 -1881
rect 2532 -2022 2566 -1881
rect 2724 -2022 2758 -1881
rect 2916 -2022 2950 -1881
rect 3024 -1996 3070 -1984
rect 1950 -2034 1996 -2022
rect 1950 -2282 1956 -2034
rect 1990 -2282 1996 -2034
rect 1950 -2294 1996 -2282
rect 2046 -2034 2092 -2022
rect 2046 -2282 2052 -2034
rect 2086 -2282 2092 -2034
rect 2046 -2294 2092 -2282
rect 2142 -2034 2188 -2022
rect 2142 -2282 2148 -2034
rect 2182 -2282 2188 -2034
rect 2142 -2294 2188 -2282
rect 2238 -2034 2284 -2022
rect 2238 -2282 2244 -2034
rect 2278 -2282 2284 -2034
rect 2238 -2294 2284 -2282
rect 2334 -2034 2380 -2022
rect 2334 -2282 2340 -2034
rect 2374 -2282 2380 -2034
rect 2334 -2294 2380 -2282
rect 2430 -2034 2476 -2022
rect 2430 -2282 2436 -2034
rect 2470 -2282 2476 -2034
rect 2430 -2294 2476 -2282
rect 2526 -2034 2572 -2022
rect 2526 -2282 2532 -2034
rect 2566 -2282 2572 -2034
rect 2526 -2294 2572 -2282
rect 2622 -2034 2668 -2022
rect 2622 -2282 2628 -2034
rect 2662 -2282 2668 -2034
rect 2622 -2294 2668 -2282
rect 2718 -2034 2764 -2022
rect 2718 -2282 2724 -2034
rect 2758 -2282 2764 -2034
rect 2718 -2294 2764 -2282
rect 2814 -2034 2860 -2022
rect 2814 -2282 2820 -2034
rect 2854 -2282 2860 -2034
rect 2814 -2294 2860 -2282
rect 2910 -2034 2956 -2022
rect 2910 -2282 2916 -2034
rect 2950 -2282 2956 -2034
rect 2910 -2294 2956 -2282
rect 1937 -2386 1947 -2334
rect 1999 -2386 2009 -2334
rect 2052 -2444 2086 -2294
rect 2130 -2386 2140 -2334
rect 2192 -2386 2202 -2334
rect 2244 -2444 2278 -2294
rect 2321 -2386 2331 -2334
rect 2383 -2386 2393 -2334
rect 2436 -2444 2470 -2294
rect 2513 -2386 2523 -2334
rect 2575 -2386 2585 -2334
rect 2628 -2444 2662 -2294
rect 2705 -2386 2715 -2334
rect 2767 -2386 2777 -2334
rect 2820 -2444 2854 -2294
rect 2897 -2386 2907 -2334
rect 2959 -2386 2969 -2334
rect 3024 -2382 3030 -1996
rect 3064 -2382 3070 -1996
rect 1772 -2478 2854 -2444
rect 3024 -2580 3070 -2382
<< via1 >>
rect -2522 -245 -2470 -193
rect -2245 -200 -2193 -193
rect -2245 -234 -2236 -200
rect -2236 -234 -2202 -200
rect -2202 -234 -2193 -200
rect -2245 -245 -2193 -234
rect -2054 -200 -2002 -193
rect -2054 -234 -2044 -200
rect -2044 -234 -2010 -200
rect -2010 -234 -2002 -200
rect -2054 -245 -2002 -234
rect -1862 -200 -1810 -193
rect -1862 -234 -1852 -200
rect -1852 -234 -1818 -200
rect -1818 -234 -1810 -200
rect -1862 -245 -1810 -234
rect -1670 -200 -1618 -193
rect -1670 -234 -1660 -200
rect -1660 -234 -1626 -200
rect -1626 -234 -1618 -200
rect -1670 -245 -1618 -234
rect -1477 -200 -1425 -192
rect -1477 -234 -1468 -200
rect -1468 -234 -1434 -200
rect -1434 -234 -1425 -200
rect -1477 -244 -1425 -234
rect -1285 -200 -1233 -192
rect -1285 -234 -1276 -200
rect -1276 -234 -1242 -200
rect -1242 -234 -1233 -200
rect -1285 -244 -1233 -234
rect -2522 -1052 -2470 -1000
rect 149 -245 201 -193
rect 426 -200 478 -193
rect 426 -234 435 -200
rect 435 -234 469 -200
rect 469 -234 478 -200
rect 426 -245 478 -234
rect 617 -200 669 -193
rect 617 -234 627 -200
rect 627 -234 661 -200
rect 661 -234 669 -200
rect 617 -245 669 -234
rect 809 -200 861 -193
rect 809 -234 819 -200
rect 819 -234 853 -200
rect 853 -234 861 -200
rect 809 -245 861 -234
rect 1001 -200 1053 -193
rect 1001 -234 1011 -200
rect 1011 -234 1045 -200
rect 1045 -234 1053 -200
rect 1001 -245 1053 -234
rect 1194 -200 1246 -192
rect 1194 -234 1203 -200
rect 1203 -234 1237 -200
rect 1237 -234 1246 -200
rect 1194 -244 1246 -234
rect 1386 -200 1438 -192
rect 1386 -234 1395 -200
rect 1395 -234 1429 -200
rect 1429 -234 1438 -200
rect 1386 -244 1438 -234
rect -2245 -1008 -2193 -1000
rect -2245 -1042 -2236 -1008
rect -2236 -1042 -2202 -1008
rect -2202 -1042 -2193 -1008
rect -2245 -1052 -2193 -1042
rect -2052 -1008 -2000 -1000
rect -2052 -1042 -2044 -1008
rect -2044 -1042 -2010 -1008
rect -2010 -1042 -2000 -1008
rect -2052 -1052 -2000 -1042
rect -1861 -1008 -1809 -1000
rect -1861 -1042 -1852 -1008
rect -1852 -1042 -1818 -1008
rect -1818 -1042 -1809 -1008
rect -1861 -1052 -1809 -1042
rect -1669 -1008 -1617 -1000
rect -1669 -1042 -1660 -1008
rect -1660 -1042 -1626 -1008
rect -1626 -1042 -1617 -1008
rect -1669 -1052 -1617 -1042
rect -1477 -1008 -1425 -1000
rect -1477 -1042 -1468 -1008
rect -1468 -1042 -1434 -1008
rect -1434 -1042 -1425 -1008
rect -1477 -1052 -1425 -1042
rect -1285 -1008 -1233 -1000
rect -1285 -1042 -1276 -1008
rect -1276 -1042 -1242 -1008
rect -1242 -1042 -1233 -1008
rect -1285 -1052 -1233 -1042
rect -33 -821 19 -769
rect -391 -873 -339 -865
rect -391 -907 -381 -873
rect -381 -907 -347 -873
rect -347 -907 -339 -873
rect -391 -917 -339 -907
rect -166 -1052 -114 -1000
rect 149 -1052 201 -1000
rect 1670 -245 1722 -193
rect 1947 -200 1999 -193
rect 1947 -234 1956 -200
rect 1956 -234 1990 -200
rect 1990 -234 1999 -200
rect 1947 -245 1999 -234
rect 2138 -200 2190 -193
rect 2138 -234 2148 -200
rect 2148 -234 2182 -200
rect 2182 -234 2190 -200
rect 2138 -245 2190 -234
rect 2330 -200 2382 -193
rect 2330 -234 2340 -200
rect 2340 -234 2374 -200
rect 2374 -234 2382 -200
rect 2330 -245 2382 -234
rect 2522 -200 2574 -193
rect 2522 -234 2532 -200
rect 2532 -234 2566 -200
rect 2566 -234 2574 -200
rect 2522 -245 2574 -234
rect 2715 -200 2767 -192
rect 2715 -234 2724 -200
rect 2724 -234 2758 -200
rect 2758 -234 2767 -200
rect 2715 -244 2767 -234
rect 2907 -200 2959 -192
rect 2907 -234 2916 -200
rect 2916 -234 2950 -200
rect 2950 -234 2959 -200
rect 2907 -244 2959 -234
rect 1650 -457 1659 -423
rect 1659 -457 1693 -423
rect 1693 -457 1702 -423
rect 1650 -475 1702 -457
rect 426 -1008 478 -1000
rect 426 -1042 435 -1008
rect 435 -1042 469 -1008
rect 469 -1042 478 -1008
rect 426 -1052 478 -1042
rect 619 -1008 671 -1000
rect 619 -1042 627 -1008
rect 627 -1042 661 -1008
rect 661 -1042 671 -1008
rect 619 -1052 671 -1042
rect 810 -1008 862 -1000
rect 810 -1042 819 -1008
rect 819 -1042 853 -1008
rect 853 -1042 862 -1008
rect 810 -1052 862 -1042
rect 1002 -1008 1054 -1000
rect 1002 -1042 1011 -1008
rect 1011 -1042 1045 -1008
rect 1045 -1042 1054 -1008
rect 1002 -1052 1054 -1042
rect 1194 -1008 1246 -1000
rect 1194 -1042 1203 -1008
rect 1203 -1042 1237 -1008
rect 1237 -1042 1246 -1008
rect 1194 -1052 1246 -1042
rect 1386 -1008 1438 -1000
rect 1386 -1042 1395 -1008
rect 1395 -1042 1429 -1008
rect 1429 -1042 1438 -1008
rect 1386 -1052 1438 -1042
rect -2522 -1394 -2470 -1342
rect -2245 -1352 -2193 -1342
rect -2245 -1386 -2236 -1352
rect -2236 -1386 -2202 -1352
rect -2202 -1386 -2193 -1352
rect -2245 -1394 -2193 -1386
rect -2052 -1352 -2000 -1342
rect -2052 -1386 -2044 -1352
rect -2044 -1386 -2010 -1352
rect -2010 -1386 -2000 -1352
rect -2052 -1394 -2000 -1386
rect -1861 -1352 -1809 -1342
rect -1861 -1386 -1852 -1352
rect -1852 -1386 -1818 -1352
rect -1818 -1386 -1809 -1352
rect -1861 -1394 -1809 -1386
rect -1669 -1352 -1617 -1342
rect -1669 -1386 -1660 -1352
rect -1660 -1386 -1626 -1352
rect -1626 -1386 -1617 -1352
rect -1669 -1394 -1617 -1386
rect -1477 -1352 -1425 -1342
rect -1477 -1386 -1468 -1352
rect -1468 -1386 -1434 -1352
rect -1434 -1386 -1425 -1352
rect -1477 -1394 -1425 -1386
rect -1285 -1352 -1233 -1342
rect -1285 -1386 -1276 -1352
rect -1276 -1386 -1242 -1352
rect -1242 -1386 -1233 -1352
rect -1285 -1394 -1233 -1386
rect 1670 -1052 1722 -1000
rect 1947 -1008 1999 -1000
rect 1947 -1042 1956 -1008
rect 1956 -1042 1990 -1008
rect 1990 -1042 1999 -1008
rect 1947 -1052 1999 -1042
rect 2140 -1008 2192 -1000
rect 2140 -1042 2148 -1008
rect 2148 -1042 2182 -1008
rect 2182 -1042 2192 -1008
rect 2140 -1052 2192 -1042
rect 2331 -1008 2383 -1000
rect 2331 -1042 2340 -1008
rect 2340 -1042 2374 -1008
rect 2374 -1042 2383 -1008
rect 2331 -1052 2383 -1042
rect 2523 -1008 2575 -1000
rect 2523 -1042 2532 -1008
rect 2532 -1042 2566 -1008
rect 2566 -1042 2575 -1008
rect 2523 -1052 2575 -1042
rect 2715 -1008 2767 -1000
rect 2715 -1042 2724 -1008
rect 2724 -1042 2758 -1008
rect 2758 -1042 2767 -1008
rect 2715 -1052 2767 -1042
rect 2907 -1008 2959 -1000
rect 2907 -1042 2916 -1008
rect 2916 -1042 2950 -1008
rect 2950 -1042 2959 -1008
rect 2907 -1052 2959 -1042
rect -2522 -2201 -2470 -2149
rect -955 -1394 -903 -1342
rect -391 -1486 -339 -1478
rect -391 -1520 -382 -1486
rect -382 -1520 -348 -1486
rect -348 -1520 -339 -1486
rect -391 -1530 -339 -1520
rect 149 -1579 201 -1527
rect 426 -1534 478 -1527
rect 426 -1568 435 -1534
rect 435 -1568 469 -1534
rect 469 -1568 478 -1534
rect 426 -1579 478 -1568
rect 617 -1534 669 -1527
rect 617 -1568 627 -1534
rect 627 -1568 661 -1534
rect 661 -1568 669 -1534
rect 617 -1579 669 -1568
rect 809 -1534 861 -1527
rect 809 -1568 819 -1534
rect 819 -1568 853 -1534
rect 853 -1568 861 -1534
rect 809 -1579 861 -1568
rect 1001 -1534 1053 -1527
rect 1001 -1568 1011 -1534
rect 1011 -1568 1045 -1534
rect 1045 -1568 1053 -1534
rect 1001 -1579 1053 -1568
rect 1194 -1534 1246 -1526
rect 1194 -1568 1203 -1534
rect 1203 -1568 1237 -1534
rect 1237 -1568 1246 -1534
rect 1194 -1578 1246 -1568
rect 1386 -1534 1438 -1526
rect 1386 -1568 1395 -1534
rect 1395 -1568 1429 -1534
rect 1429 -1568 1438 -1534
rect 1386 -1578 1438 -1568
rect -2245 -2160 -2193 -2149
rect -2245 -2194 -2236 -2160
rect -2236 -2194 -2202 -2160
rect -2202 -2194 -2193 -2160
rect -2245 -2201 -2193 -2194
rect -2054 -2160 -2002 -2149
rect -2054 -2194 -2044 -2160
rect -2044 -2194 -2010 -2160
rect -2010 -2194 -2002 -2160
rect -2054 -2201 -2002 -2194
rect -1862 -2160 -1810 -2149
rect -1862 -2194 -1852 -2160
rect -1852 -2194 -1818 -2160
rect -1818 -2194 -1810 -2160
rect -1862 -2201 -1810 -2194
rect -1670 -2160 -1618 -2149
rect -1670 -2194 -1660 -2160
rect -1660 -2194 -1626 -2160
rect -1626 -2194 -1618 -2160
rect -1670 -2201 -1618 -2194
rect -1477 -2160 -1425 -2150
rect -1477 -2194 -1468 -2160
rect -1468 -2194 -1434 -2160
rect -1434 -2194 -1425 -2160
rect -1477 -2202 -1425 -2194
rect -1285 -2160 -1233 -2150
rect -1285 -2194 -1276 -2160
rect -1276 -2194 -1242 -2160
rect -1242 -2194 -1233 -2160
rect -1285 -2202 -1233 -2194
rect 149 -2386 201 -2334
rect 1670 -1579 1722 -1527
rect 1947 -1534 1999 -1527
rect 1947 -1568 1956 -1534
rect 1956 -1568 1990 -1534
rect 1990 -1568 1999 -1534
rect 1947 -1579 1999 -1568
rect 2138 -1534 2190 -1527
rect 2138 -1568 2148 -1534
rect 2148 -1568 2182 -1534
rect 2182 -1568 2190 -1534
rect 2138 -1579 2190 -1568
rect 2330 -1534 2382 -1527
rect 2330 -1568 2340 -1534
rect 2340 -1568 2374 -1534
rect 2374 -1568 2382 -1534
rect 2330 -1579 2382 -1568
rect 2522 -1534 2574 -1527
rect 2522 -1568 2532 -1534
rect 2532 -1568 2566 -1534
rect 2566 -1568 2574 -1534
rect 2522 -1579 2574 -1568
rect 2715 -1534 2767 -1526
rect 2715 -1568 2724 -1534
rect 2724 -1568 2758 -1534
rect 2758 -1568 2767 -1534
rect 2715 -1578 2767 -1568
rect 2907 -1534 2959 -1526
rect 2907 -1568 2916 -1534
rect 2916 -1568 2950 -1534
rect 2950 -1568 2959 -1534
rect 2907 -1578 2959 -1568
rect 1650 -1791 1659 -1757
rect 1659 -1791 1693 -1757
rect 1693 -1791 1702 -1757
rect 1650 -1809 1702 -1791
rect 426 -2342 478 -2334
rect 426 -2376 435 -2342
rect 435 -2376 469 -2342
rect 469 -2376 478 -2342
rect 426 -2386 478 -2376
rect 619 -2342 671 -2334
rect 619 -2376 627 -2342
rect 627 -2376 661 -2342
rect 661 -2376 671 -2342
rect 619 -2386 671 -2376
rect 810 -2342 862 -2334
rect 810 -2376 819 -2342
rect 819 -2376 853 -2342
rect 853 -2376 862 -2342
rect 810 -2386 862 -2376
rect 1002 -2342 1054 -2334
rect 1002 -2376 1011 -2342
rect 1011 -2376 1045 -2342
rect 1045 -2376 1054 -2342
rect 1002 -2386 1054 -2376
rect 1194 -2342 1246 -2334
rect 1194 -2376 1203 -2342
rect 1203 -2376 1237 -2342
rect 1237 -2376 1246 -2342
rect 1194 -2386 1246 -2376
rect 1386 -2342 1438 -2334
rect 1386 -2376 1395 -2342
rect 1395 -2376 1429 -2342
rect 1429 -2376 1438 -2342
rect 1386 -2386 1438 -2376
rect 1670 -2386 1722 -2334
rect 1947 -2342 1999 -2334
rect 1947 -2376 1956 -2342
rect 1956 -2376 1990 -2342
rect 1990 -2376 1999 -2342
rect 1947 -2386 1999 -2376
rect 2140 -2342 2192 -2334
rect 2140 -2376 2148 -2342
rect 2148 -2376 2182 -2342
rect 2182 -2376 2192 -2342
rect 2140 -2386 2192 -2376
rect 2331 -2342 2383 -2334
rect 2331 -2376 2340 -2342
rect 2340 -2376 2374 -2342
rect 2374 -2376 2383 -2342
rect 2331 -2386 2383 -2376
rect 2523 -2342 2575 -2334
rect 2523 -2376 2532 -2342
rect 2532 -2376 2566 -2342
rect 2566 -2376 2575 -2342
rect 2523 -2386 2575 -2376
rect 2715 -2342 2767 -2334
rect 2715 -2376 2724 -2342
rect 2724 -2376 2758 -2342
rect 2758 -2376 2767 -2342
rect 2715 -2386 2767 -2376
rect 2907 -2342 2959 -2334
rect 2907 -2376 2916 -2342
rect 2916 -2376 2950 -2342
rect 2950 -2376 2959 -2342
rect 2907 -2386 2959 -2376
<< metal2 >>
rect -2522 -193 -2470 -183
rect -2245 -193 -2193 -183
rect -2054 -193 -2002 -183
rect -1862 -193 -1810 -183
rect -1670 -193 -1618 -183
rect -1477 -192 -1425 -182
rect -1285 -192 -1233 -182
rect -2470 -245 -2245 -193
rect -2193 -245 -2054 -193
rect -2002 -245 -1862 -193
rect -1810 -245 -1670 -193
rect -1618 -244 -1477 -193
rect -1425 -244 -1285 -192
rect -1233 -244 -723 -192
rect -1618 -245 -1226 -244
rect -2522 -255 -2470 -245
rect -2245 -255 -2193 -245
rect -2054 -255 -2002 -245
rect -1862 -255 -1810 -245
rect -1670 -255 -1618 -245
rect -1477 -254 -1425 -245
rect -1285 -254 -1233 -245
rect -2522 -1000 -2470 -990
rect -2245 -1000 -2193 -990
rect -2052 -1000 -2000 -990
rect -1861 -1000 -1809 -990
rect -1669 -1000 -1617 -990
rect -1477 -1000 -1425 -990
rect -1285 -1000 -1233 -990
rect -2470 -1052 -2245 -1000
rect -2193 -1052 -2052 -1000
rect -2000 -1052 -1861 -1000
rect -1809 -1052 -1669 -1000
rect -1617 -1052 -1477 -1000
rect -1425 -1052 -1285 -1000
rect -1233 -1052 -903 -1000
rect -2522 -1062 -2470 -1052
rect -2245 -1062 -2193 -1052
rect -2052 -1062 -2000 -1052
rect -1861 -1062 -1809 -1052
rect -1669 -1062 -1617 -1052
rect -1477 -1062 -1425 -1052
rect -1285 -1062 -1233 -1052
rect -2522 -1342 -2470 -1332
rect -2245 -1342 -2193 -1332
rect -2052 -1342 -2000 -1332
rect -1861 -1342 -1809 -1332
rect -1669 -1342 -1617 -1332
rect -1477 -1342 -1425 -1332
rect -1285 -1342 -1233 -1332
rect -955 -1342 -903 -1052
rect -2470 -1394 -2245 -1342
rect -2193 -1394 -2052 -1342
rect -2000 -1394 -1861 -1342
rect -1809 -1394 -1669 -1342
rect -1617 -1394 -1477 -1342
rect -1425 -1394 -1285 -1342
rect -1233 -1394 -955 -1342
rect -2522 -1404 -2470 -1394
rect -2245 -1404 -2193 -1394
rect -2052 -1404 -2000 -1394
rect -1861 -1404 -1809 -1394
rect -1669 -1404 -1617 -1394
rect -1477 -1404 -1425 -1394
rect -1285 -1404 -1233 -1394
rect -955 -1404 -903 -1394
rect -775 -1927 -723 -244
rect -391 -865 -339 115
rect 149 -193 201 -183
rect 426 -193 478 -183
rect 617 -193 669 -183
rect 809 -193 861 -183
rect 1001 -193 1053 -183
rect 1194 -192 1246 -182
rect -391 -1000 -339 -917
rect -33 -245 149 -193
rect 201 -245 426 -193
rect 478 -245 617 -193
rect 669 -245 809 -193
rect 861 -245 1001 -193
rect 1053 -244 1194 -193
rect 1386 -192 1438 -182
rect 1246 -244 1386 -193
rect 1670 -193 1722 -183
rect 1947 -193 1999 -183
rect 2138 -193 2190 -183
rect 2330 -193 2382 -183
rect 2522 -193 2574 -183
rect 2715 -192 2767 -182
rect 1438 -244 1670 -193
rect 1053 -245 1670 -244
rect 1722 -245 1947 -193
rect 1999 -245 2138 -193
rect 2190 -245 2330 -193
rect 2382 -245 2522 -193
rect 2574 -244 2715 -193
rect 2907 -192 2959 -182
rect 2767 -244 2907 -193
rect 2959 -244 2966 -193
rect 2574 -245 2966 -244
rect -33 -769 19 -245
rect 149 -255 201 -245
rect 426 -255 478 -245
rect 617 -255 669 -245
rect 809 -255 861 -245
rect 1001 -255 1053 -245
rect 1194 -254 1246 -245
rect 1386 -254 1438 -245
rect 1670 -255 1722 -245
rect 1947 -255 1999 -245
rect 2138 -255 2190 -245
rect 2330 -255 2382 -245
rect 2522 -255 2574 -245
rect 2715 -254 2767 -245
rect 2907 -254 2959 -245
rect -166 -1000 -114 -990
rect -391 -1052 -166 -1000
rect -166 -1062 -114 -1052
rect -391 -1478 -339 -1468
rect -391 -1927 -339 -1530
rect -775 -1979 -339 -1927
rect -2522 -2149 -2470 -2139
rect -2245 -2149 -2193 -2139
rect -2054 -2149 -2002 -2139
rect -1862 -2149 -1810 -2139
rect -1670 -2149 -1618 -2139
rect -1477 -2149 -1425 -2140
rect -1285 -2149 -1233 -2140
rect -775 -2149 -723 -1979
rect -2470 -2201 -2245 -2149
rect -2193 -2201 -2054 -2149
rect -2002 -2201 -1862 -2149
rect -1810 -2201 -1670 -2149
rect -1618 -2150 -723 -2149
rect -1618 -2201 -1477 -2150
rect -2522 -2211 -2470 -2201
rect -2245 -2211 -2193 -2201
rect -2054 -2211 -2002 -2201
rect -1862 -2211 -1810 -2201
rect -1670 -2211 -1618 -2201
rect -1425 -2201 -1285 -2150
rect -1477 -2212 -1425 -2202
rect -1233 -2201 -723 -2150
rect -1285 -2212 -1233 -2202
rect -391 -2457 -339 -1979
rect -33 -2334 19 -821
rect 1650 -423 1702 -413
rect 1650 -990 1702 -475
rect 149 -1000 201 -990
rect 426 -1000 478 -990
rect 619 -1000 671 -990
rect 810 -1000 862 -990
rect 1002 -1000 1054 -990
rect 1194 -1000 1246 -990
rect 1386 -1000 1438 -990
rect 1650 -1000 1722 -990
rect 1947 -1000 1999 -990
rect 2140 -1000 2192 -990
rect 2331 -1000 2383 -990
rect 2523 -1000 2575 -990
rect 2715 -1000 2767 -990
rect 2907 -1000 2959 -990
rect 201 -1052 426 -1000
rect 478 -1052 619 -1000
rect 671 -1052 810 -1000
rect 862 -1052 1002 -1000
rect 1054 -1052 1194 -1000
rect 1246 -1052 1386 -1000
rect 1438 -1052 1670 -1000
rect 1722 -1052 1947 -1000
rect 1999 -1052 2140 -1000
rect 2192 -1052 2331 -1000
rect 2383 -1052 2523 -1000
rect 2575 -1052 2715 -1000
rect 2767 -1052 2907 -1000
rect 2959 -1052 2966 -1000
rect 149 -1527 201 -1052
rect 426 -1062 478 -1052
rect 619 -1062 671 -1052
rect 810 -1062 862 -1052
rect 1002 -1062 1054 -1052
rect 1194 -1062 1246 -1052
rect 1386 -1062 1438 -1052
rect 1670 -1062 1722 -1052
rect 1947 -1062 1999 -1052
rect 2140 -1062 2192 -1052
rect 2331 -1062 2383 -1052
rect 2523 -1062 2575 -1052
rect 2715 -1062 2767 -1052
rect 2907 -1062 2959 -1052
rect 426 -1527 478 -1517
rect 617 -1527 669 -1517
rect 809 -1527 861 -1517
rect 1001 -1527 1053 -1517
rect 1194 -1526 1246 -1516
rect 201 -1579 426 -1527
rect 478 -1579 617 -1527
rect 669 -1579 809 -1527
rect 861 -1579 1001 -1527
rect 1053 -1578 1194 -1527
rect 1386 -1526 1438 -1516
rect 1246 -1578 1386 -1527
rect 1670 -1527 1722 -1517
rect 1947 -1527 1999 -1517
rect 2138 -1527 2190 -1517
rect 2330 -1527 2382 -1517
rect 2522 -1527 2574 -1517
rect 2715 -1526 2767 -1516
rect 1438 -1578 1670 -1527
rect 1053 -1579 1670 -1578
rect 1722 -1579 1947 -1527
rect 1999 -1579 2138 -1527
rect 2190 -1579 2330 -1527
rect 2382 -1579 2522 -1527
rect 2574 -1578 2715 -1527
rect 2907 -1526 2959 -1516
rect 2767 -1578 2907 -1527
rect 2959 -1578 2966 -1527
rect 2574 -1579 2966 -1578
rect 149 -1589 201 -1579
rect 426 -1589 478 -1579
rect 617 -1589 669 -1579
rect 809 -1589 861 -1579
rect 1001 -1589 1053 -1579
rect 1194 -1588 1246 -1579
rect 1386 -1588 1438 -1579
rect 1670 -1589 1722 -1579
rect 1947 -1589 1999 -1579
rect 2138 -1589 2190 -1579
rect 2330 -1589 2382 -1579
rect 2522 -1589 2574 -1579
rect 2715 -1588 2767 -1579
rect 2907 -1588 2959 -1579
rect 1650 -1757 1702 -1747
rect 1650 -2324 1702 -1809
rect 149 -2334 201 -2324
rect 426 -2334 478 -2324
rect 619 -2334 671 -2324
rect 810 -2334 862 -2324
rect 1002 -2334 1054 -2324
rect 1194 -2334 1246 -2324
rect 1386 -2334 1438 -2324
rect 1650 -2334 1722 -2324
rect 1947 -2334 1999 -2324
rect 2140 -2334 2192 -2324
rect 2331 -2334 2383 -2324
rect 2523 -2334 2575 -2324
rect 2715 -2334 2767 -2324
rect 2907 -2334 2959 -2324
rect -33 -2386 149 -2334
rect 201 -2386 426 -2334
rect 478 -2386 619 -2334
rect 671 -2386 810 -2334
rect 862 -2386 1002 -2334
rect 1054 -2386 1194 -2334
rect 1246 -2386 1386 -2334
rect 1438 -2386 1670 -2334
rect 1722 -2386 1947 -2334
rect 1999 -2386 2140 -2334
rect 2192 -2386 2331 -2334
rect 2383 -2386 2523 -2334
rect 2575 -2386 2715 -2334
rect 2767 -2386 2907 -2334
rect 2959 -2386 2966 -2334
rect 149 -2396 201 -2386
rect 426 -2396 478 -2386
rect 619 -2396 671 -2386
rect 810 -2396 862 -2386
rect 1002 -2396 1054 -2386
rect 1194 -2396 1246 -2386
rect 1386 -2396 1438 -2386
rect 1670 -2396 1722 -2386
rect 1947 -2396 1999 -2386
rect 2140 -2396 2192 -2386
rect 2331 -2396 2383 -2386
rect 2523 -2396 2575 -2386
rect 2715 -2396 2767 -2386
rect 2907 -2396 2959 -2386
<< labels >>
flabel metal1 -2635 -530 -2635 -530 3 FreeSans 400 0 0 0 in0
port 3 e
flabel metal1 -2634 -1864 -2634 -1864 3 FreeSans 400 0 0 0 in1
port 4 e
flabel metal1 -1144 -2365 -1144 -2365 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 -1051 -1198 -1051 -1198 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 -1145 -35 -1145 -35 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal2 -366 110 -366 110 5 FreeSans 400 0 0 0 s0
port 2 s
flabel metal2 -365 -2445 -365 -2445 1 FreeSans 400 0 0 0 en
port 1 n
flabel metal1 -615 -1743 -615 -1743 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 -617 -1196 -617 -1196 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 -616 -652 -616 -652 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 1526 -1 1526 -1 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 3048 4 3048 4 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 1526 -1242 1526 -1242 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 3048 -1239 3048 -1239 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 3047 -1344 3047 -1344 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 1526 -1342 1526 -1342 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal1 1527 -2577 1527 -2577 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 3048 -2574 3048 -2574 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 3423 -1288 3423 -1288 1 FreeSans 400 0 0 0 out
port 5 n
flabel metal1 -2544 -1368 -2544 -1368 3 FreeSans 400 0 0 0 transmission_gate_1/en_b
flabel metal1 -2545 -1864 -2545 -1864 3 FreeSans 400 0 0 0 transmission_gate_1/in
flabel metal1 -2545 -2175 -2545 -2175 3 FreeSans 400 0 0 0 transmission_gate_1/en
flabel metal1 -1054 -1865 -1054 -1865 7 FreeSans 400 0 0 0 transmission_gate_1/out
flabel metal1 -1145 -1219 -1145 -1219 5 FreeSans 400 0 0 0 transmission_gate_1/VDD
flabel metal1 -1145 -2325 -1145 -2325 1 FreeSans 400 0 0 0 transmission_gate_1/VSS
flabel metal1 -2544 -1026 -2544 -1026 3 FreeSans 400 0 0 0 transmission_gate_0/en_b
flabel metal1 -2545 -530 -2545 -530 3 FreeSans 400 0 0 0 transmission_gate_0/in
flabel metal1 -2545 -219 -2545 -219 3 FreeSans 400 0 0 0 transmission_gate_0/en
flabel metal1 -1054 -529 -1054 -529 7 FreeSans 400 0 0 0 transmission_gate_0/out
flabel metal1 -1145 -1175 -1145 -1175 1 FreeSans 400 0 0 0 transmission_gate_0/VDD
flabel metal1 -1145 -69 -1145 -69 5 FreeSans 400 0 0 0 transmission_gate_0/VSS
flabel metal1 1526 -1215 1526 -1215 5 FreeSans 400 0 0 0 switch_5t_1/VDD
flabel metal1 1526 -33 1526 -33 5 FreeSans 400 0 0 0 switch_5t_1/VSS
flabel metal1 80 -1025 80 -1025 5 FreeSans 400 0 0 0 switch_5t_1/en_b
flabel metal1 78 -219 78 -219 5 FreeSans 400 0 0 0 switch_5t_1/en
flabel metal1 79 -530 79 -530 5 FreeSans 400 0 0 0 switch_5t_1/in
flabel metal1 3174 -529 3174 -529 7 FreeSans 400 0 0 0 switch_5t_1/out
flabel metal1 3047 -1216 3047 -1216 5 FreeSans 400 0 0 0 switch_5t_1/VDD
flabel metal1 3047 -34 3047 -34 5 FreeSans 400 0 0 0 switch_5t_1/VSS
flabel metal1 1648 -1026 1648 -1026 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/en_b
flabel metal1 1647 -530 1647 -530 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/in
flabel metal1 1647 -219 1647 -219 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/en
flabel metal1 3138 -529 3138 -529 7 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/out
flabel metal1 3047 -1175 3047 -1175 1 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/VDD
flabel metal1 3047 -69 3047 -69 5 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/VSS
flabel metal1 127 -1026 127 -1026 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/en_b
flabel metal1 126 -530 126 -530 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/in
flabel metal1 126 -219 126 -219 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/en
flabel metal1 1617 -529 1617 -529 7 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/out
flabel metal1 1526 -1175 1526 -1175 1 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/VDD
flabel metal1 1526 -69 1526 -69 5 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/VSS
flabel metal1 1526 -2549 1526 -2549 5 FreeSans 400 0 0 0 switch_5t_0/VDD
flabel metal1 1526 -1367 1526 -1367 5 FreeSans 400 0 0 0 switch_5t_0/VSS
flabel metal1 80 -2359 80 -2359 5 FreeSans 400 0 0 0 switch_5t_0/en_b
flabel metal1 78 -1553 78 -1553 5 FreeSans 400 0 0 0 switch_5t_0/en
flabel metal1 79 -1864 79 -1864 5 FreeSans 400 0 0 0 switch_5t_0/in
flabel metal1 3174 -1863 3174 -1863 7 FreeSans 400 0 0 0 switch_5t_0/out
flabel metal1 3047 -2550 3047 -2550 5 FreeSans 400 0 0 0 switch_5t_0/VDD
flabel metal1 3047 -1368 3047 -1368 5 FreeSans 400 0 0 0 switch_5t_0/VSS
flabel metal1 1648 -2360 1648 -2360 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/en_b
flabel metal1 1647 -1864 1647 -1864 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/in
flabel metal1 1647 -1553 1647 -1553 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/en
flabel metal1 3138 -1863 3138 -1863 7 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/out
flabel metal1 3047 -2509 3047 -2509 1 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/VDD
flabel metal1 3047 -1403 3047 -1403 5 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/VSS
flabel metal1 127 -2360 127 -2360 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/en_b
flabel metal1 126 -1864 126 -1864 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/in
flabel metal1 126 -1553 126 -1553 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/en
flabel metal1 1617 -1863 1617 -1863 7 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/out
flabel metal1 1526 -2509 1526 -2509 1 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/VDD
flabel metal1 1526 -1403 1526 -1403 5 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/VSS
flabel metal1 -534 -1205 -481 -1176 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -531 -672 -480 -634 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment -459 -652 -459 -652 8 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
rlabel metal1 -551 -700 -459 -604 5 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel metal1 -551 -1244 -459 -1148 5 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -529 -1216 -476 -1187 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -530 -1758 -479 -1720 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment -551 -1740 -551 -1740 4 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
rlabel metal1 -551 -1788 -459 -1692 1 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel metal1 -551 -1244 -459 -1148 1 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel locali -295 -975 -261 -941 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali -295 -907 -261 -873 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali -387 -907 -353 -873 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/A
flabel nwell -430 -1213 -396 -1179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell -430 -669 -396 -635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 -430 -669 -396 -635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 -430 -1213 -396 -1179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment -459 -652 -459 -652 2 sky130_fd_sc_hd__inv_1_1/inv_1
rlabel metal1 -459 -700 -183 -604 5 sky130_fd_sc_hd__inv_1_1/VGND
rlabel metal1 -459 -1244 -183 -1148 5 sky130_fd_sc_hd__inv_1_1/VPWR
flabel locali -295 -1451 -261 -1417 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -295 -1519 -261 -1485 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -387 -1519 -353 -1485 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell -430 -1213 -396 -1179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -430 -1757 -396 -1723 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -430 -1757 -396 -1723 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -430 -1213 -396 -1179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -459 -1740 -459 -1740 4 sky130_fd_sc_hd__inv_1_0/inv_1
rlabel metal1 -459 -1788 -183 -1692 1 sky130_fd_sc_hd__inv_1_0/VGND
rlabel metal1 -459 -1244 -183 -1148 1 sky130_fd_sc_hd__inv_1_0/VPWR
<< end >>
