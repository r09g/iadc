* NGSPICE file created from analog_top_v2.ext - technology: sky130A

.subckt esd_cell_flat esd VDD VSS
X0 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+13p pd=1.058e+08u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=500000u
X1 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.595e+13p pd=1.1638e+08u as=1.45e+13p ps=1.058e+08u w=5e+06u l=500000u
X2 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X3 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X4 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X5 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X6 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X7 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X8 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X9 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X10 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X11 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X12 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X13 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X14 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X20 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X21 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X22 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X23 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X24 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X25 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X26 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X27 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X28 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X29 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X30 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X31 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X32 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X33 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X34 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X35 VSS VSS esd VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X36 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X37 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X38 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X39 VDD VDD esd VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 esd VDD 24.78fF
C1 esd VSS 25.63fF
C2 VDD VSS 19.27fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CEWQ64 c1_n260_n210# m3_n360_n310# VSUBS
X0 c1_n260_n210# m3_n360_n310# sky130_fd_pr__cap_mim_m3_1 l=2.1e+06u w=2.1e+06u
C0 m3_n360_n310# c1_n260_n210# 0.73fF
C1 m3_n360_n310# VSUBS 0.63fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CGPBWM m3_n1030_n980# c1_n930_n880# VSUBS
X0 c1_n930_n880# m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1 l=8.8e+06u w=8.79e+06u
C0 c1_n930_n880# m3_n1030_n980# 8.31fF
C1 m3_n1030_n980# VSUBS 2.79fF
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
C0 VPB VPWR 0.47fF
C1 VPB VGND 0.87fF
C2 VPWR VGND 3.03fF
C3 VPWR VNB 1.33fF
C4 VGND VNB 0.77fF
C5 VPB VNB 1.14fF
.ends

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_352_n136# a_256_n136# 0.33fF
C1 a_n416_n136# a_256_n136# 0.03fF
C2 a_n128_n136# w_n646_n356# 0.05fF
C3 a_352_n136# a_n224_n136# 0.03fF
C4 a_n224_n136# a_n416_n136# 0.12fF
C5 a_n32_n136# a_448_n136# 0.04fF
C6 a_n128_n136# a_64_n136# 0.12fF
C7 a_352_n136# a_n32_n136# 0.05fF
C8 a_n32_n136# a_n416_n136# 0.05fF
C9 a_160_n136# a_n128_n136# 0.07fF
C10 w_n646_n356# a_64_n136# 0.05fF
C11 a_160_n136# w_n646_n356# 0.06fF
C12 a_n512_n234# a_n320_n136# 0.03fF
C13 a_n508_n136# a_n128_n136# 0.05fF
C14 a_160_n136# a_64_n136# 0.33fF
C15 a_n320_n136# a_448_n136# 0.02fF
C16 a_n128_n136# a_256_n136# 0.05fF
C17 a_n508_n136# w_n646_n356# 0.13fF
C18 a_n224_n136# a_n128_n136# 0.33fF
C19 a_352_n136# a_n320_n136# 0.03fF
C20 a_n416_n136# a_n320_n136# 0.33fF
C21 a_256_n136# w_n646_n356# 0.06fF
C22 a_n508_n136# a_64_n136# 0.03fF
C23 a_n224_n136# w_n646_n356# 0.06fF
C24 a_n512_n234# a_448_n136# 0.03fF
C25 a_n32_n136# a_n128_n136# 0.33fF
C26 a_n508_n136# a_160_n136# 0.03fF
C27 a_256_n136# a_64_n136# 0.12fF
C28 a_352_n136# a_n512_n234# 0.03fF
C29 a_160_n136# a_256_n136# 0.33fF
C30 a_n512_n234# a_n416_n136# 0.03fF
C31 a_n32_n136# w_n646_n356# 0.05fF
C32 a_n224_n136# a_64_n136# 0.07fF
C33 a_n224_n136# a_160_n136# 0.05fF
C34 a_352_n136# a_448_n136# 0.33fF
C35 a_n416_n136# a_448_n136# 0.02fF
C36 a_n32_n136# a_64_n136# 0.33fF
C37 a_n508_n136# a_256_n136# 0.02fF
C38 a_n32_n136# a_160_n136# 0.12fF
C39 a_352_n136# a_n416_n136# 0.02fF
C40 a_n508_n136# a_n224_n136# 0.07fF
C41 a_n320_n136# a_n128_n136# 0.12fF
C42 a_n224_n136# a_256_n136# 0.04fF
C43 a_n508_n136# a_n32_n136# 0.04fF
C44 a_n320_n136# w_n646_n356# 0.06fF
C45 a_n32_n136# a_256_n136# 0.07fF
C46 a_n512_n234# a_n128_n136# 0.03fF
C47 a_n224_n136# a_n32_n136# 0.12fF
C48 a_n320_n136# a_64_n136# 0.05fF
C49 a_n320_n136# a_160_n136# 0.04fF
C50 a_448_n136# a_n128_n136# 0.03fF
C51 a_n512_n234# w_n646_n356# 1.47fF
C52 a_352_n136# a_n128_n136# 0.04fF
C53 a_448_n136# w_n646_n356# 0.13fF
C54 a_n416_n136# a_n128_n136# 0.07fF
C55 a_n512_n234# a_64_n136# 0.03fF
C56 a_n508_n136# a_n320_n136# 0.12fF
C57 a_n512_n234# a_160_n136# 0.03fF
C58 a_352_n136# w_n646_n356# 0.08fF
C59 a_n416_n136# w_n646_n356# 0.08fF
C60 a_448_n136# a_64_n136# 0.05fF
C61 a_n320_n136# a_256_n136# 0.03fF
C62 a_160_n136# a_448_n136# 0.07fF
C63 a_n224_n136# a_n320_n136# 0.33fF
C64 a_352_n136# a_64_n136# 0.07fF
C65 a_n416_n136# a_64_n136# 0.04fF
C66 a_n508_n136# a_n512_n234# 0.03fF
C67 a_352_n136# a_160_n136# 0.12fF
C68 a_n416_n136# a_160_n136# 0.03fF
C69 a_n32_n136# a_n320_n136# 0.07fF
C70 a_n512_n234# a_256_n136# 0.03fF
C71 a_n508_n136# a_448_n136# 0.02fF
C72 a_n512_n234# a_n224_n136# 0.03fF
C73 a_448_n136# a_256_n136# 0.12fF
C74 a_352_n136# a_n508_n136# 0.02fF
C75 a_n508_n136# a_n416_n136# 0.33fF
C76 a_n224_n136# a_448_n136# 0.03fF
C77 a_n512_n234# a_n32_n136# 0.03fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# w_n646_n262# a_448_n52# a_n416_n52#
+ a_160_n52# a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149#
+ a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_352_n52# a_160_n52# 0.05fF
C1 a_n416_n52# a_160_n52# 0.01fF
C2 a_n128_n52# a_n512_n149# 0.03fF
C3 a_352_n52# a_n320_n52# 0.01fF
C4 a_n320_n52# a_n416_n52# 0.13fF
C5 a_n32_n52# a_448_n52# 0.02fF
C6 a_n128_n52# a_64_n52# 0.05fF
C7 a_352_n52# a_n32_n52# 0.02fF
C8 a_n32_n52# a_n416_n52# 0.02fF
C9 a_256_n52# a_n128_n52# 0.02fF
C10 a_n512_n149# a_64_n52# 0.03fF
C11 a_256_n52# a_n512_n149# 0.03fF
C12 a_n508_n52# a_n224_n52# 0.03fF
C13 a_256_n52# a_64_n52# 0.05fF
C14 a_n224_n52# a_448_n52# 0.01fF
C15 a_n128_n52# a_160_n52# 0.03fF
C16 a_n320_n52# a_n128_n52# 0.05fF
C17 a_352_n52# a_n224_n52# 0.01fF
C18 a_n416_n52# a_n224_n52# 0.05fF
C19 a_160_n52# a_n512_n149# 0.03fF
C20 a_n320_n52# a_n512_n149# 0.03fF
C21 a_n508_n52# a_448_n52# 0.01fF
C22 a_n32_n52# a_n128_n52# 0.13fF
C23 a_160_n52# a_64_n52# 0.13fF
C24 a_352_n52# a_n508_n52# 0.01fF
C25 a_256_n52# a_160_n52# 0.13fF
C26 a_n32_n52# a_n512_n149# 0.03fF
C27 a_n508_n52# a_n416_n52# 0.13fF
C28 a_n320_n52# a_64_n52# 0.02fF
C29 a_n320_n52# a_256_n52# 0.01fF
C30 a_352_n52# a_448_n52# 0.13fF
C31 a_n416_n52# a_448_n52# 0.01fF
C32 a_n32_n52# a_64_n52# 0.13fF
C33 a_n32_n52# a_256_n52# 0.03fF
C34 a_352_n52# a_n416_n52# 0.01fF
C35 a_n224_n52# a_n128_n52# 0.13fF
C36 a_n320_n52# a_160_n52# 0.02fF
C37 a_n224_n52# a_n512_n149# 0.03fF
C38 a_n32_n52# a_160_n52# 0.05fF
C39 a_n508_n52# a_n128_n52# 0.02fF
C40 a_n320_n52# a_n32_n52# 0.03fF
C41 a_n224_n52# a_64_n52# 0.03fF
C42 a_n224_n52# a_256_n52# 0.02fF
C43 a_448_n52# a_n128_n52# 0.01fF
C44 a_n508_n52# a_n512_n149# 0.03fF
C45 a_352_n52# a_n128_n52# 0.02fF
C46 a_448_n52# a_n512_n149# 0.03fF
C47 a_n416_n52# a_n128_n52# 0.03fF
C48 a_n508_n52# a_64_n52# 0.01fF
C49 a_n508_n52# a_256_n52# 0.01fF
C50 a_352_n52# a_n512_n149# 0.03fF
C51 a_n416_n52# a_n512_n149# 0.03fF
C52 a_448_n52# a_64_n52# 0.02fF
C53 a_n224_n52# a_160_n52# 0.02fF
C54 a_256_n52# a_448_n52# 0.05fF
C55 a_n320_n52# a_n224_n52# 0.13fF
C56 a_352_n52# a_64_n52# 0.03fF
C57 a_n416_n52# a_64_n52# 0.02fF
C58 a_352_n52# a_256_n52# 0.13fF
C59 a_n416_n52# a_256_n52# 0.01fF
C60 a_n32_n52# a_n224_n52# 0.05fF
C61 a_n508_n52# a_160_n52# 0.01fF
C62 a_n508_n52# a_n320_n52# 0.05fF
C63 a_448_n52# a_160_n52# 0.03fF
C64 a_n320_n52# a_448_n52# 0.01fF
C65 a_n508_n52# a_n32_n52# 0.02fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate en VDD nmos_tgate_0/w_n646_n262# in out en_b VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in nmos_tgate_0/w_n646_n262# out in in VSS out in out out en
+ out nmos_tgate
C0 en_b en 0.07fF
C1 en_b VDD -0.11fF
C2 in out 0.77fF
C3 en out 0.01fF
C4 in en 0.13fF
C5 out VDD 0.29fF
C6 in VDD 0.70fF
C7 en_b out 0.01fF
C8 en VDD 0.12fF
C9 in en_b 0.15fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

.subckt sky130_fd_sc_hd__clkinv_16 A VGND VPWR Y VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.0605e+12p pd=1.261e+07u as=1.0059e+12p ps=1.151e+07u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.515e+12p pd=3.103e+07u as=3.655e+12p ps=3.331e+07u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VPB A 1.26fF
C1 VPWR A 0.64fF
C2 A Y 1.32fF
C3 VPB VPWR 0.89fF
C4 VGND A 0.66fF
C5 VPB Y 0.09fF
C6 VPWR Y 4.41fF
C7 VPWR VGND 0.34fF
C8 VGND Y 1.58fF
C9 VGND VNB 1.26fF
C10 Y VNB 0.13fF
C11 VPWR VNB 0.47fF
C12 A VNB 1.70fF
C13 VPB VNB 2.20fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_YVTR7C a_n207_n140# a_n1039_n205# a_29_n205# a_327_n140#
+ a_n683_n205# a_n1275_n140# a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_1097_n205#
+ a_n505_n205# a_n741_n140# a_563_n205# a_861_n140# w_n1311_n241# a_919_n205# a_n327_n205#
+ a_n563_n140# a_385_n205# a_683_n140# a_n919_n140# a_n149_n205# a_1039_n140# a_n385_n140#
+ a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_327_n140# a_207_n205# a_149_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_149_n140# a_29_n205# a_n29_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_861_n140# a_741_n205# a_683_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_n140# a_n327_n205# a_n385_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1097_n205# a_1097_n205# a_1039_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n741_n140# a_n861_n205# a_n919_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n1097_n140# a_n1275_n140# a_n1275_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_683_n140# a_563_n205# a_505_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1039_n140# a_919_n205# a_861_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n29_n140# a_n149_n205# a_n207_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n563_n140# a_n683_n205# a_n741_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n207_n140# a_327_n140# 0.02fF
C1 a_1039_n140# a_683_n140# 0.03fF
C2 a_n919_n140# a_683_n140# 0.01fF
C3 a_919_n205# a_741_n205# 0.10fF
C4 a_1097_n205# a_861_n140# 0.03fF
C5 a_n505_n205# a_n149_n205# 0.03fF
C6 a_1097_n205# a_n149_n205# 0.00fF
C7 a_29_n205# a_741_n205# 0.01fF
C8 a_n207_n140# a_505_n140# 0.01fF
C9 w_n1311_n241# a_327_n140# 0.02fF
C10 a_n741_n140# a_n919_n140# 0.06fF
C11 a_149_n140# a_861_n140# 0.01fF
C12 a_n683_n205# a_n861_n205# 0.10fF
C13 a_n1275_n140# a_385_n205# 0.00fF
C14 w_n1311_n241# a_505_n140# 0.02fF
C15 a_1039_n140# a_1097_n205# 0.06fF
C16 a_n29_n140# a_683_n140# 0.01fF
C17 a_n741_n140# a_n1275_n140# 0.02fF
C18 a_n1039_n205# a_n861_n205# 0.10fF
C19 a_n385_n140# a_327_n140# 0.01fF
C20 a_1039_n140# a_149_n140# 0.01fF
C21 a_n505_n205# a_n1275_n140# 0.01fF
C22 a_n683_n205# a_919_n205# 0.01fF
C23 a_n29_n140# a_n741_n140# 0.01fF
C24 a_n861_n205# a_n327_n205# 0.02fF
C25 a_149_n140# a_n919_n140# 0.01fF
C26 a_n683_n205# a_29_n205# 0.01fF
C27 a_n563_n140# a_n1097_n140# 0.02fF
C28 a_505_n140# a_n385_n140# 0.01fF
C29 w_n1311_n241# a_207_n205# 0.18fF
C30 a_149_n140# a_n1275_n140# 0.01fF
C31 a_n29_n140# a_1097_n205# 0.01fF
C32 a_919_n205# a_n327_n205# 0.01fF
C33 a_n683_n205# a_741_n205# 0.01fF
C34 a_n1039_n205# a_29_n205# 0.01fF
C35 a_n861_n205# a_n149_n205# 0.01fF
C36 a_29_n205# a_n327_n205# 0.03fF
C37 a_563_n205# w_n1311_n241# 0.16fF
C38 a_n29_n140# a_149_n140# 0.06fF
C39 a_n207_n140# a_683_n140# 0.01fF
C40 a_n327_n205# a_741_n205# 0.01fF
C41 a_919_n205# a_n149_n205# 0.01fF
C42 a_n207_n140# a_n741_n140# 0.02fF
C43 w_n1311_n241# a_683_n140# 0.02fF
C44 a_n149_n205# a_29_n205# 0.10fF
C45 w_n1311_n241# a_385_n205# 0.17fF
C46 a_n149_n205# a_741_n205# 0.01fF
C47 a_n207_n140# a_1097_n205# 0.01fF
C48 w_n1311_n241# a_n741_n140# 0.02fF
C49 a_n861_n205# a_n1275_n140# 0.02fF
C50 a_505_n140# a_327_n140# 0.06fF
C51 a_n563_n140# a_861_n140# 0.01fF
C52 a_n385_n140# a_683_n140# 0.01fF
C53 a_n207_n140# a_149_n140# 0.03fF
C54 a_n683_n205# a_n1039_n205# 0.03fF
C55 w_n1311_n241# a_n505_n205# 0.20fF
C56 w_n1311_n241# a_1097_n205# 0.28fF
C57 a_n683_n205# a_n327_n205# 0.03fF
C58 a_n741_n140# a_n385_n140# 0.03fF
C59 a_29_n205# a_n1275_n140# 0.00fF
C60 w_n1311_n241# a_149_n140# 0.02fF
C61 a_n1039_n205# a_n327_n205# 0.01fF
C62 a_1039_n140# a_n563_n140# 0.01fF
C63 a_n919_n140# a_n563_n140# 0.03fF
C64 a_1097_n205# a_n385_n140# 0.01fF
C65 a_n683_n205# a_n149_n205# 0.02fF
C66 a_n919_n140# a_n1097_n140# 0.06fF
C67 a_n563_n140# a_n1275_n140# 0.01fF
C68 a_n1039_n205# a_n149_n205# 0.01fF
C69 a_149_n140# a_n385_n140# 0.02fF
C70 a_n149_n205# a_n327_n205# 0.10fF
C71 a_n1097_n140# a_n1275_n140# 0.06fF
C72 a_n29_n140# a_n563_n140# 0.02fF
C73 a_683_n140# a_327_n140# 0.03fF
C74 a_n29_n140# a_n1097_n140# 0.01fF
C75 w_n1311_n241# a_n861_n205# 0.20fF
C76 a_505_n140# a_683_n140# 0.06fF
C77 a_n683_n205# a_n1275_n140# 0.01fF
C78 a_n741_n140# a_327_n140# 0.01fF
C79 a_563_n205# a_207_n205# 0.03fF
C80 a_n1039_n205# a_n1275_n140# 0.07fF
C81 a_n741_n140# a_505_n140# 0.01fF
C82 a_919_n205# w_n1311_n241# 0.14fF
C83 a_1097_n205# a_327_n140# 0.01fF
C84 a_n1275_n140# a_n327_n205# 0.01fF
C85 w_n1311_n241# a_29_n205# 0.19fF
C86 a_1039_n140# a_861_n140# 0.06fF
C87 a_n207_n140# a_n563_n140# 0.03fF
C88 a_1097_n205# a_505_n140# 0.01fF
C89 a_149_n140# a_327_n140# 0.06fF
C90 w_n1311_n241# a_741_n205# 0.15fF
C91 a_n207_n140# a_n1097_n140# 0.01fF
C92 a_n149_n205# a_n1275_n140# 0.01fF
C93 a_207_n205# a_385_n205# 0.10fF
C94 a_149_n140# a_505_n140# 0.03fF
C95 w_n1311_n241# a_n563_n140# 0.02fF
C96 a_n29_n140# a_861_n140# 0.01fF
C97 a_563_n205# a_385_n205# 0.10fF
C98 w_n1311_n241# a_n1097_n140# 0.02fF
C99 a_n505_n205# a_207_n205# 0.01fF
C100 a_207_n205# a_1097_n205# 0.01fF
C101 a_n919_n140# a_n1275_n140# 0.03fF
C102 a_n563_n140# a_n385_n140# 0.06fF
C103 a_563_n205# a_n505_n205# 0.01fF
C104 a_563_n205# a_1097_n205# 0.01fF
C105 a_n683_n205# w_n1311_n241# 0.20fF
C106 a_n741_n140# a_683_n140# 0.01fF
C107 a_n1097_n140# a_n385_n140# 0.01fF
C108 a_1039_n140# a_n29_n140# 0.01fF
C109 a_n29_n140# a_n919_n140# 0.01fF
C110 a_n1039_n205# w_n1311_n241# 0.20fF
C111 a_1097_n205# a_683_n140# 0.02fF
C112 w_n1311_n241# a_n327_n205# 0.20fF
C113 a_n29_n140# a_n1275_n140# 0.01fF
C114 a_n207_n140# a_861_n140# 0.01fF
C115 a_n505_n205# a_385_n205# 0.01fF
C116 a_1097_n205# a_385_n205# 0.01fF
C117 a_149_n140# a_683_n140# 0.02fF
C118 w_n1311_n241# a_861_n140# 0.01fF
C119 w_n1311_n241# a_n149_n205# 0.19fF
C120 a_n741_n140# a_149_n140# 0.01fF
C121 a_207_n205# a_n861_n205# 0.01fF
C122 a_n505_n205# a_1097_n205# 0.00fF
C123 a_1039_n140# a_n207_n140# 0.01fF
C124 a_n563_n140# a_327_n140# 0.01fF
C125 a_n207_n140# a_n919_n140# 0.01fF
C126 a_563_n205# a_n861_n205# 0.01fF
C127 a_n1097_n140# a_327_n140# 0.01fF
C128 a_1097_n205# a_149_n140# 0.01fF
C129 a_n563_n140# a_505_n140# 0.01fF
C130 a_n207_n140# a_n1275_n140# 0.01fF
C131 a_861_n140# a_n385_n140# 0.01fF
C132 a_919_n205# a_207_n205# 0.01fF
C133 a_1039_n140# w_n1311_n241# 0.01fF
C134 w_n1311_n241# a_n919_n140# 0.02fF
C135 a_207_n205# a_29_n205# 0.10fF
C136 a_505_n140# a_n1097_n140# 0.01fF
C137 a_563_n205# a_919_n205# 0.03fF
C138 a_n29_n140# a_n207_n140# 0.06fF
C139 w_n1311_n241# a_n1275_n140# 0.33fF
C140 a_563_n205# a_29_n205# 0.02fF
C141 a_207_n205# a_741_n205# 0.02fF
C142 a_1039_n140# a_n385_n140# 0.01fF
C143 a_n861_n205# a_385_n205# 0.01fF
C144 a_n919_n140# a_n385_n140# 0.02fF
C145 a_563_n205# a_741_n205# 0.10fF
C146 w_n1311_n241# a_n29_n140# 0.02fF
C147 a_n385_n140# a_n1275_n140# 0.01fF
C148 a_n505_n205# a_n861_n205# 0.03fF
C149 a_919_n205# a_385_n205# 0.02fF
C150 a_29_n205# a_385_n205# 0.03fF
C151 a_n29_n140# a_n385_n140# 0.03fF
C152 a_861_n140# a_327_n140# 0.02fF
C153 a_919_n205# a_n505_n205# 0.01fF
C154 a_n683_n205# a_207_n205# 0.01fF
C155 a_n563_n140# a_683_n140# 0.01fF
C156 a_919_n205# a_1097_n205# 0.07fF
C157 a_741_n205# a_385_n205# 0.03fF
C158 a_n505_n205# a_29_n205# 0.02fF
C159 a_1097_n205# a_29_n205# 0.01fF
C160 a_505_n140# a_861_n140# 0.03fF
C161 a_563_n205# a_n683_n205# 0.01fF
C162 a_n1039_n205# a_207_n205# 0.01fF
C163 w_n1311_n241# a_n207_n140# 0.02fF
C164 a_n741_n140# a_n563_n140# 0.06fF
C165 a_n505_n205# a_741_n205# 0.01fF
C166 a_207_n205# a_n327_n205# 0.02fF
C167 a_1097_n205# a_741_n205# 0.02fF
C168 a_1039_n140# a_327_n140# 0.01fF
C169 a_n919_n140# a_327_n140# 0.01fF
C170 a_563_n205# a_n1039_n205# 0.01fF
C171 a_n741_n140# a_n1097_n140# 0.03fF
C172 a_563_n205# a_n327_n205# 0.01fF
C173 a_1039_n140# a_505_n140# 0.02fF
C174 a_327_n140# a_n1275_n140# 0.01fF
C175 a_n919_n140# a_505_n140# 0.01fF
C176 a_n207_n140# a_n385_n140# 0.06fF
C177 a_207_n205# a_n149_n205# 0.03fF
C178 a_n683_n205# a_385_n205# 0.01fF
C179 a_149_n140# a_n563_n140# 0.01fF
C180 a_n29_n140# a_327_n140# 0.03fF
C181 a_563_n205# a_n149_n205# 0.01fF
C182 a_149_n140# a_n1097_n140# 0.01fF
C183 w_n1311_n241# a_n385_n140# 0.02fF
C184 a_n1039_n205# a_385_n205# 0.01fF
C185 a_n683_n205# a_n505_n205# 0.10fF
C186 a_n327_n205# a_385_n205# 0.01fF
C187 a_n29_n140# a_505_n140# 0.02fF
C188 a_n861_n205# a_29_n205# 0.01fF
C189 a_861_n140# a_683_n140# 0.06fF
C190 a_n1039_n205# a_n505_n205# 0.02fF
C191 a_207_n205# a_n1275_n140# 0.00fF
C192 a_n505_n205# a_n327_n205# 0.10fF
C193 a_n861_n205# a_741_n205# 0.01fF
C194 a_1097_n205# a_n327_n205# 0.00fF
C195 a_n149_n205# a_385_n205# 0.02fF
C196 a_n741_n140# a_861_n140# 0.01fF
C197 a_919_n205# a_29_n205# 0.01fF
C198 w_n1311_n241# VSUBS 3.79fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AKSJZW a_n149_n195# a_n207_n140# a_207_n195# a_327_n140#
+ a_n1275_n140# a_n861_n195# a_n29_n140# a_149_n140# a_n1097_n140# a_n1039_n195# a_29_n195#
+ a_n683_n195# a_n741_n140# a_741_n195# a_861_n140# a_1097_n195# a_n563_n140# a_n505_n195#
+ a_563_n195# a_683_n140# a_n919_n140# a_919_n195# a_1039_n140# a_n385_n140# a_n327_n195#
+ a_385_n195# a_505_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n195# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n195# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n195# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n195# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_327_n140# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_861_n140# a_741_n195# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n207_n140# a_n327_n195# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_1097_n195# a_1097_n195# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n195# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1275_n140# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n195# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n195# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n505_n195# a_n149_n195# 0.03fF
C1 a_n327_n195# a_n1039_n195# 0.01fF
C2 a_n207_n140# a_149_n140# 0.03fF
C3 a_29_n195# a_n1275_n140# 0.00fF
C4 a_327_n140# a_n1275_n140# 0.01fF
C5 a_327_n140# a_n1097_n140# 0.01fF
C6 a_n919_n140# a_149_n140# 0.01fF
C7 a_861_n140# a_1097_n195# 0.03fF
C8 a_n207_n140# a_505_n140# 0.01fF
C9 a_919_n195# a_n683_n195# 0.01fF
C10 a_n505_n195# a_n1275_n140# 0.01fF
C11 a_505_n140# a_n919_n140# 0.01fF
C12 a_n207_n140# a_n741_n140# 0.02fF
C13 a_207_n195# a_385_n195# 0.10fF
C14 a_n741_n140# a_n919_n140# 0.06fF
C15 a_505_n140# a_149_n140# 0.03fF
C16 a_29_n195# a_n327_n195# 0.03fF
C17 a_563_n195# a_385_n195# 0.10fF
C18 a_1039_n140# a_n29_n140# 0.01fF
C19 a_n741_n140# a_149_n140# 0.01fF
C20 a_29_n195# a_741_n195# 0.01fF
C21 a_385_n195# a_n149_n195# 0.02fF
C22 a_n505_n195# a_n327_n195# 0.10fF
C23 a_505_n140# a_n741_n140# 0.01fF
C24 a_n385_n140# a_1039_n140# 0.01fF
C25 a_n505_n195# a_741_n195# 0.01fF
C26 a_385_n195# a_n1275_n140# 0.00fF
C27 a_n207_n140# a_n1275_n140# 0.01fF
C28 a_n29_n140# a_861_n140# 0.01fF
C29 a_n207_n140# a_n1097_n140# 0.01fF
C30 a_1039_n140# a_n563_n140# 0.01fF
C31 a_1039_n140# a_683_n140# 0.03fF
C32 a_n1275_n140# a_n919_n140# 0.03fF
C33 a_n1097_n140# a_n919_n140# 0.06fF
C34 a_385_n195# a_n327_n195# 0.01fF
C35 a_n385_n140# a_861_n140# 0.01fF
C36 a_n1275_n140# a_149_n140# 0.01fF
C37 a_n1097_n140# a_149_n140# 0.01fF
C38 a_1039_n140# a_327_n140# 0.01fF
C39 a_385_n195# a_741_n195# 0.03fF
C40 a_n861_n195# a_n683_n195# 0.10fF
C41 a_n29_n140# a_1097_n195# 0.01fF
C42 a_505_n140# a_n1097_n140# 0.01fF
C43 a_207_n195# a_563_n195# 0.03fF
C44 a_919_n195# a_29_n195# 0.01fF
C45 a_n385_n140# a_1097_n195# 0.01fF
C46 a_n741_n140# a_n1275_n140# 0.02fF
C47 a_207_n195# a_n149_n195# 0.03fF
C48 a_n1097_n140# a_n741_n140# 0.03fF
C49 a_861_n140# a_n563_n140# 0.01fF
C50 a_683_n140# a_861_n140# 0.06fF
C51 a_919_n195# a_n505_n195# 0.01fF
C52 a_563_n195# a_n149_n195# 0.01fF
C53 a_207_n195# a_n1275_n140# 0.00fF
C54 a_327_n140# a_861_n140# 0.02fF
C55 a_683_n140# a_1097_n195# 0.02fF
C56 a_n1275_n140# a_n149_n195# 0.01fF
C57 a_29_n195# a_1097_n195# 0.01fF
C58 a_n1039_n195# a_n683_n195# 0.03fF
C59 a_327_n140# a_1097_n195# 0.01fF
C60 a_207_n195# a_n327_n195# 0.02fF
C61 a_919_n195# a_385_n195# 0.02fF
C62 a_n207_n140# a_1039_n140# 0.01fF
C63 a_n861_n195# a_n1039_n195# 0.10fF
C64 a_n1097_n140# a_n1275_n140# 0.06fF
C65 a_207_n195# a_741_n195# 0.02fF
C66 a_563_n195# a_n327_n195# 0.01fF
C67 a_n505_n195# a_1097_n195# 0.00fF
C68 a_n327_n195# a_n149_n195# 0.10fF
C69 a_n385_n140# a_n29_n140# 0.03fF
C70 a_563_n195# a_741_n195# 0.10fF
C71 a_29_n195# a_n683_n195# 0.01fF
C72 a_1039_n140# a_149_n140# 0.01fF
C73 a_741_n195# a_n149_n195# 0.01fF
C74 a_n327_n195# a_n1275_n140# 0.01fF
C75 a_1039_n140# a_505_n140# 0.02fF
C76 a_29_n195# a_n861_n195# 0.01fF
C77 a_n505_n195# a_n683_n195# 0.10fF
C78 a_n207_n140# a_861_n140# 0.01fF
C79 a_n29_n140# a_n563_n140# 0.02fF
C80 a_n505_n195# a_n861_n195# 0.03fF
C81 a_n29_n140# a_683_n140# 0.01fF
C82 a_385_n195# a_1097_n195# 0.01fF
C83 a_n385_n140# a_n563_n140# 0.06fF
C84 a_n385_n140# a_683_n140# 0.01fF
C85 a_861_n140# a_149_n140# 0.01fF
C86 a_n29_n140# a_327_n140# 0.03fF
C87 a_n207_n140# a_1097_n195# 0.01fF
C88 a_n327_n195# a_741_n195# 0.01fF
C89 a_505_n140# a_861_n140# 0.03fF
C90 a_n385_n140# a_327_n140# 0.01fF
C91 a_207_n195# a_919_n195# 0.01fF
C92 a_385_n195# a_n683_n195# 0.01fF
C93 a_n741_n140# a_861_n140# 0.01fF
C94 a_1097_n195# a_149_n140# 0.01fF
C95 a_563_n195# a_919_n195# 0.03fF
C96 a_683_n140# a_n563_n140# 0.01fF
C97 a_385_n195# a_n861_n195# 0.01fF
C98 a_29_n195# a_n1039_n195# 0.01fF
C99 a_505_n140# a_1097_n195# 0.01fF
C100 a_919_n195# a_n149_n195# 0.01fF
C101 a_327_n140# a_n563_n140# 0.01fF
C102 a_n505_n195# a_n1039_n195# 0.02fF
C103 a_683_n140# a_327_n140# 0.03fF
C104 a_207_n195# a_1097_n195# 0.01fF
C105 a_29_n195# a_n505_n195# 0.02fF
C106 a_563_n195# a_1097_n195# 0.01fF
C107 a_n207_n140# a_n29_n140# 0.06fF
C108 a_919_n195# a_n327_n195# 0.01fF
C109 a_1097_n195# a_n149_n195# 0.00fF
C110 a_n29_n140# a_n919_n140# 0.01fF
C111 a_n385_n140# a_n207_n140# 0.06fF
C112 a_385_n195# a_n1039_n195# 0.01fF
C113 a_919_n195# a_741_n195# 0.10fF
C114 a_207_n195# a_n683_n195# 0.01fF
C115 a_n385_n140# a_n919_n140# 0.02fF
C116 a_n29_n140# a_149_n140# 0.06fF
C117 a_n29_n140# a_505_n140# 0.02fF
C118 a_207_n195# a_n861_n195# 0.01fF
C119 a_563_n195# a_n683_n195# 0.01fF
C120 a_n385_n140# a_149_n140# 0.02fF
C121 a_n683_n195# a_n149_n195# 0.02fF
C122 a_n29_n140# a_n741_n140# 0.01fF
C123 a_n385_n140# a_505_n140# 0.01fF
C124 a_563_n195# a_n861_n195# 0.01fF
C125 a_29_n195# a_385_n195# 0.03fF
C126 a_n207_n140# a_n563_n140# 0.03fF
C127 a_n207_n140# a_683_n140# 0.01fF
C128 a_n861_n195# a_n149_n195# 0.01fF
C129 a_n919_n140# a_n563_n140# 0.03fF
C130 a_n385_n140# a_n741_n140# 0.03fF
C131 a_n327_n195# a_1097_n195# 0.00fF
C132 a_683_n140# a_n919_n140# 0.01fF
C133 a_n1275_n140# a_n683_n195# 0.01fF
C134 a_385_n195# a_n505_n195# 0.01fF
C135 a_n207_n140# a_327_n140# 0.02fF
C136 a_149_n140# a_n563_n140# 0.01fF
C137 a_683_n140# a_149_n140# 0.02fF
C138 a_1097_n195# a_741_n195# 0.02fF
C139 a_327_n140# a_n919_n140# 0.01fF
C140 a_n861_n195# a_n1275_n140# 0.02fF
C141 a_505_n140# a_n563_n140# 0.01fF
C142 a_683_n140# a_505_n140# 0.06fF
C143 a_327_n140# a_149_n140# 0.06fF
C144 a_n741_n140# a_n563_n140# 0.06fF
C145 a_n327_n195# a_n683_n195# 0.03fF
C146 a_683_n140# a_n741_n140# 0.01fF
C147 a_327_n140# a_505_n140# 0.06fF
C148 a_207_n195# a_n1039_n195# 0.01fF
C149 a_n683_n195# a_741_n195# 0.01fF
C150 a_n327_n195# a_n861_n195# 0.02fF
C151 a_1039_n140# a_861_n140# 0.06fF
C152 a_n29_n140# a_n1275_n140# 0.01fF
C153 a_n29_n140# a_n1097_n140# 0.01fF
C154 a_327_n140# a_n741_n140# 0.01fF
C155 a_563_n195# a_n1039_n195# 0.01fF
C156 a_n861_n195# a_741_n195# 0.01fF
C157 a_n385_n140# a_n1275_n140# 0.01fF
C158 a_n1039_n195# a_n149_n195# 0.01fF
C159 a_n385_n140# a_n1097_n140# 0.01fF
C160 a_207_n195# a_29_n195# 0.10fF
C161 a_1039_n140# a_1097_n195# 0.06fF
C162 a_n1275_n140# a_n1039_n195# 0.06fF
C163 a_563_n195# a_29_n195# 0.02fF
C164 a_207_n195# a_n505_n195# 0.01fF
C165 a_29_n195# a_n149_n195# 0.10fF
C166 a_919_n195# a_1097_n195# 0.06fF
C167 a_n1275_n140# a_n563_n140# 0.01fF
C168 a_n1097_n140# a_n563_n140# 0.02fF
C169 a_n207_n140# a_n919_n140# 0.01fF
C170 a_563_n195# a_n505_n195# 0.01fF
C171 a_1039_n140# VSUBS 0.01fF
C172 a_861_n140# VSUBS 0.01fF
C173 a_683_n140# VSUBS 0.02fF
C174 a_505_n140# VSUBS 0.02fF
C175 a_327_n140# VSUBS 0.02fF
C176 a_149_n140# VSUBS 0.02fF
C177 a_n29_n140# VSUBS 0.02fF
C178 a_n207_n140# VSUBS 0.02fF
C179 a_n385_n140# VSUBS 0.02fF
C180 a_n563_n140# VSUBS 0.02fF
C181 a_n741_n140# VSUBS 0.02fF
C182 a_n919_n140# VSUBS 0.02fF
C183 a_n1097_n140# VSUBS 0.02fF
C184 a_1097_n195# VSUBS 0.31fF
C185 a_919_n195# VSUBS 0.19fF
C186 a_741_n195# VSUBS 0.20fF
C187 a_563_n195# VSUBS 0.21fF
C188 a_385_n195# VSUBS 0.22fF
C189 a_207_n195# VSUBS 0.23fF
C190 a_29_n195# VSUBS 0.23fF
C191 a_n149_n195# VSUBS 0.24fF
C192 a_n327_n195# VSUBS 0.24fF
C193 a_n505_n195# VSUBS 0.24fF
C194 a_n683_n195# VSUBS 0.24fF
C195 a_n861_n195# VSUBS 0.24fF
C196 a_n1039_n195# VSUBS 0.24fF
C197 a_n1275_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_K7HVMB a_664_n120# a_n608_n120# a_n86_n120# a_72_n208#
+ a_240_n120# a_n184_n120# a_n562_142# a_n510_n120# a_28_n120# a_n298_n120# a_126_n120#
+ a_452_n120# a_n396_n120# a_284_142# a_n138_142# a_550_n120# a_496_n208# a_338_n120#
+ a_n350_n208# a_n820_n120# VSUBS
X0 a_n820_n120# a_n820_n120# a_n820_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X1 a_n510_n120# a_n562_142# a_n608_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X2 a_664_n120# a_664_n120# a_664_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X3 a_n298_n120# a_n350_n208# a_n396_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X4 a_550_n120# a_496_n208# a_452_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X5 a_126_n120# a_72_n208# a_28_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X6 a_n86_n120# a_n138_142# a_n184_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X7 a_338_n120# a_284_142# a_240_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
C0 a_n184_n120# a_n396_n120# 0.04fF
C1 a_338_n120# a_126_n120# 0.04fF
C2 a_n298_n120# a_126_n120# 0.02fF
C3 a_n510_n120# a_240_n120# 0.01fF
C4 a_n510_n120# a_452_n120# 0.01fF
C5 a_496_n208# a_n138_142# 0.00fF
C6 a_n184_n120# a_240_n120# 0.02fF
C7 a_n184_n120# a_452_n120# 0.01fF
C8 a_338_n120# a_n510_n120# 0.01fF
C9 a_n510_n120# a_n298_n120# 0.04fF
C10 a_664_n120# a_496_n208# 0.01fF
C11 a_338_n120# a_n184_n120# 0.01fF
C12 a_n184_n120# a_n298_n120# 0.09fF
C13 a_n608_n120# a_550_n120# 0.01fF
C14 a_284_142# a_n562_142# 0.01fF
C15 a_664_n120# a_550_n120# 0.13fF
C16 a_496_n208# a_452_n120# 0.00fF
C17 a_550_n120# a_n396_n120# 0.01fF
C18 a_n820_n120# a_284_142# 0.00fF
C19 a_240_n120# a_550_n120# 0.03fF
C20 a_452_n120# a_550_n120# 0.11fF
C21 a_664_n120# a_n138_142# 0.00fF
C22 a_496_n208# a_72_n208# 0.01fF
C23 a_28_n120# a_n86_n120# 0.09fF
C24 a_n562_142# a_n350_n208# 0.01fF
C25 a_338_n120# a_550_n120# 0.04fF
C26 a_n298_n120# a_550_n120# 0.01fF
C27 a_n608_n120# a_664_n120# 0.01fF
C28 a_n820_n120# a_n350_n208# 0.01fF
C29 a_n608_n120# a_n396_n120# 0.04fF
C30 a_664_n120# a_n396_n120# 0.01fF
C31 a_n608_n120# a_240_n120# 0.01fF
C32 a_n608_n120# a_452_n120# 0.01fF
C33 a_n820_n120# a_n86_n120# 0.02fF
C34 a_664_n120# a_240_n120# 0.03fF
C35 a_664_n120# a_452_n120# 0.06fF
C36 a_240_n120# a_n396_n120# 0.01fF
C37 a_452_n120# a_n396_n120# 0.01fF
C38 a_n138_142# a_72_n208# 0.01fF
C39 a_n820_n120# a_28_n120# 0.02fF
C40 a_338_n120# a_n608_n120# 0.01fF
C41 a_126_n120# a_n86_n120# 0.04fF
C42 a_n608_n120# a_n298_n120# 0.03fF
C43 a_284_142# a_496_n208# 0.01fF
C44 a_338_n120# a_664_n120# 0.04fF
C45 a_452_n120# a_240_n120# 0.04fF
C46 a_28_n120# a_126_n120# 0.11fF
C47 a_664_n120# a_n298_n120# 0.01fF
C48 a_338_n120# a_n396_n120# 0.01fF
C49 a_n298_n120# a_n396_n120# 0.11fF
C50 a_n820_n120# a_n562_142# 0.01fF
C51 a_664_n120# a_72_n208# 0.00fF
C52 a_n510_n120# a_n86_n120# 0.02fF
C53 a_338_n120# a_240_n120# 0.11fF
C54 a_338_n120# a_452_n120# 0.09fF
C55 a_n298_n120# a_240_n120# 0.01fF
C56 a_n298_n120# a_452_n120# 0.01fF
C57 a_n510_n120# a_28_n120# 0.01fF
C58 a_n184_n120# a_n86_n120# 0.11fF
C59 a_n820_n120# a_126_n120# 0.02fF
C60 a_n184_n120# a_28_n120# 0.04fF
C61 a_496_n208# a_n350_n208# 0.01fF
C62 a_338_n120# a_n298_n120# 0.01fF
C63 a_284_142# a_n138_142# 0.01fF
C64 a_n510_n120# a_n562_142# 0.00fF
C65 a_n820_n120# a_n510_n120# 0.06fF
C66 a_n820_n120# a_n184_n120# 0.03fF
C67 a_664_n120# a_284_142# 0.01fF
C68 a_n510_n120# a_126_n120# 0.01fF
C69 a_550_n120# a_n86_n120# 0.01fF
C70 a_n138_142# a_n350_n208# 0.01fF
C71 a_n184_n120# a_126_n120# 0.03fF
C72 a_284_142# a_240_n120# 0.00fF
C73 a_28_n120# a_550_n120# 0.01fF
C74 a_n562_142# a_496_n208# 0.00fF
C75 a_n820_n120# a_496_n208# 0.00fF
C76 a_n510_n120# a_n184_n120# 0.02fF
C77 a_n138_142# a_n86_n120# 0.00fF
C78 a_664_n120# a_n350_n208# 0.00fF
C79 a_284_142# a_72_n208# 0.01fF
C80 a_n608_n120# a_n86_n120# 0.01fF
C81 a_n820_n120# a_550_n120# 0.01fF
C82 a_n608_n120# a_28_n120# 0.01fF
C83 a_664_n120# a_n86_n120# 0.02fF
C84 a_n86_n120# a_n396_n120# 0.03fF
C85 a_550_n120# a_126_n120# 0.02fF
C86 a_n562_142# a_n138_142# 0.01fF
C87 a_664_n120# a_28_n120# 0.02fF
C88 a_28_n120# a_n396_n120# 0.02fF
C89 a_n820_n120# a_n138_142# 0.00fF
C90 a_n298_n120# a_n350_n208# 0.00fF
C91 a_240_n120# a_n86_n120# 0.02fF
C92 a_452_n120# a_n86_n120# 0.01fF
C93 a_n350_n208# a_72_n208# 0.01fF
C94 a_n510_n120# a_550_n120# 0.01fF
C95 a_28_n120# a_240_n120# 0.04fF
C96 a_28_n120# a_452_n120# 0.02fF
C97 a_n820_n120# a_n608_n120# 0.13fF
C98 a_664_n120# a_n562_142# 0.00fF
C99 a_338_n120# a_n86_n120# 0.02fF
C100 a_n184_n120# a_550_n120# 0.01fF
C101 a_n298_n120# a_n86_n120# 0.04fF
C102 a_n820_n120# a_664_n120# 0.02fF
C103 a_n820_n120# a_n396_n120# 0.04fF
C104 a_n608_n120# a_126_n120# 0.01fF
C105 a_338_n120# a_28_n120# 0.03fF
C106 a_n298_n120# a_28_n120# 0.02fF
C107 a_664_n120# a_126_n120# 0.03fF
C108 a_28_n120# a_72_n208# 0.00fF
C109 a_n820_n120# a_240_n120# 0.01fF
C110 a_126_n120# a_n396_n120# 0.01fF
C111 a_n820_n120# a_452_n120# 0.01fF
C112 a_n608_n120# a_n510_n120# 0.11fF
C113 a_240_n120# a_126_n120# 0.09fF
C114 a_452_n120# a_126_n120# 0.02fF
C115 a_664_n120# a_n510_n120# 0.01fF
C116 a_n608_n120# a_n184_n120# 0.02fF
C117 a_338_n120# a_n820_n120# 0.01fF
C118 a_n820_n120# a_n298_n120# 0.03fF
C119 a_n562_142# a_72_n208# 0.00fF
C120 a_n510_n120# a_n396_n120# 0.09fF
C121 a_284_142# a_n350_n208# 0.00fF
C122 a_664_n120# a_n184_n120# 0.02fF
C123 a_n820_n120# a_72_n208# 0.00fF
C124 a_550_n120# VSUBS 0.01fF
C125 a_452_n120# VSUBS 0.01fF
C126 a_338_n120# VSUBS 0.01fF
C127 a_240_n120# VSUBS 0.01fF
C128 a_126_n120# VSUBS 0.02fF
C129 a_28_n120# VSUBS 0.01fF
C130 a_n86_n120# VSUBS 0.01fF
C131 a_n184_n120# VSUBS 0.02fF
C132 a_n298_n120# VSUBS 0.02fF
C133 a_n396_n120# VSUBS 0.02fF
C134 a_n510_n120# VSUBS 0.02fF
C135 a_n608_n120# VSUBS 0.02fF
C136 a_496_n208# VSUBS 0.11fF
C137 a_664_n120# VSUBS 0.17fF
C138 a_72_n208# VSUBS 0.10fF
C139 a_284_142# VSUBS 0.10fF
C140 a_n350_n208# VSUBS 0.12fF
C141 a_n138_142# VSUBS 0.11fF
C142 a_n820_n120# VSUBS 0.20fF
C143 a_n562_142# VSUBS 0.14fF
.ends

.subckt sky130_fd_pr__nfet_01v8_S6RQQZ a_n149_n194# a_n207_n140# a_207_n194# a_1453_n194#
+ a_n1217_n194# a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140#
+ a_n1097_n140# a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194#
+ a_861_n140# a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140#
+ a_n919_n140# a_919_n194# a_n1631_n140# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194#
+ a_n1395_n194# a_505_n140# a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n1453_n140# a_n1631_n140# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1453_n194# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n861_n194# a_n505_n194# 0.03fF
C1 a_n919_n140# a_n1097_n140# 0.06fF
C2 a_n683_n194# a_n1395_n194# 0.01fF
C3 a_n327_n194# a_n1631_n140# 0.00fF
C4 a_1453_n194# a_1217_n140# 0.03fF
C5 a_29_n194# a_919_n194# 0.01fF
C6 a_n1275_n140# a_n1097_n140# 0.06fF
C7 a_505_n140# a_149_n140# 0.03fF
C8 a_1217_n140# a_1395_n140# 0.06fF
C9 a_n919_n140# a_n563_n140# 0.03fF
C10 a_563_n194# a_n1039_n194# 0.01fF
C11 a_683_n140# a_n563_n140# 0.01fF
C12 a_505_n140# a_1039_n140# 0.02fF
C13 a_n861_n194# a_n1631_n140# 0.01fF
C14 a_n563_n140# a_n1275_n140# 0.01fF
C15 a_n149_n194# a_29_n194# 0.10fF
C16 a_n563_n140# a_n1097_n140# 0.02fF
C17 a_n327_n194# a_n683_n194# 0.03fF
C18 a_207_n194# a_29_n194# 0.10fF
C19 a_n207_n140# a_n741_n140# 0.02fF
C20 a_n327_n194# a_385_n194# 0.01fF
C21 a_n207_n140# a_n385_n140# 0.06fF
C22 a_29_n194# a_n505_n194# 0.02fF
C23 a_1453_n194# a_385_n194# 0.01fF
C24 a_n861_n194# a_n683_n194# 0.10fF
C25 a_563_n194# a_1275_n194# 0.01fF
C26 a_n861_n194# a_385_n194# 0.01fF
C27 a_29_n194# a_n1631_n140# 0.00fF
C28 a_n207_n140# a_1395_n140# 0.01fF
C29 a_1097_n194# a_563_n194# 0.02fF
C30 a_n919_n140# a_n1631_n140# 0.01fF
C31 a_n149_n194# a_919_n194# 0.01fF
C32 a_n919_n140# a_n1453_n140# 0.02fF
C33 a_n29_n140# a_n741_n140# 0.01fF
C34 a_683_n140# a_1217_n140# 0.02fF
C35 a_n29_n140# a_n385_n140# 0.03fF
C36 a_n1631_n140# a_n1275_n140# 0.03fF
C37 a_n1453_n140# a_n1275_n140# 0.06fF
C38 a_861_n140# a_n741_n140# 0.01fF
C39 a_29_n194# a_n683_n194# 0.01fF
C40 a_327_n140# a_n741_n140# 0.01fF
C41 a_861_n140# a_n385_n140# 0.01fF
C42 a_327_n140# a_n385_n140# 0.01fF
C43 a_207_n194# a_919_n194# 0.01fF
C44 a_n1631_n140# a_n1097_n140# 0.02fF
C45 a_919_n194# a_n505_n194# 0.01fF
C46 a_n1453_n140# a_n1097_n140# 0.03fF
C47 a_n29_n140# a_1453_n194# 0.01fF
C48 a_29_n194# a_385_n194# 0.03fF
C49 a_n1217_n194# a_n1039_n194# 0.10fF
C50 a_1275_n194# a_741_n194# 0.02fF
C51 a_861_n140# a_1453_n194# 0.01fF
C52 a_327_n140# a_1453_n194# 0.01fF
C53 a_n29_n140# a_1395_n140# 0.01fF
C54 a_n563_n140# a_n1631_n140# 0.01fF
C55 a_n563_n140# a_n1453_n140# 0.01fF
C56 a_861_n140# a_1395_n140# 0.02fF
C57 a_n149_n194# a_207_n194# 0.03fF
C58 a_327_n140# a_1395_n140# 0.01fF
C59 a_563_n194# a_n327_n194# 0.01fF
C60 a_563_n194# a_1453_n194# 0.01fF
C61 a_1097_n194# a_741_n194# 0.03fF
C62 a_n149_n194# a_n505_n194# 0.03fF
C63 a_149_n140# a_n741_n140# 0.01fF
C64 a_n385_n140# a_149_n140# 0.02fF
C65 a_563_n194# a_n861_n194# 0.01fF
C66 a_207_n194# a_n505_n194# 0.01fF
C67 a_1039_n140# a_n385_n140# 0.01fF
C68 a_n919_n140# a_n207_n140# 0.01fF
C69 a_n207_n140# a_683_n140# 0.01fF
C70 a_n149_n194# a_n1631_n140# 0.00fF
C71 a_n207_n140# a_n1275_n140# 0.01fF
C72 a_1453_n194# a_149_n140# 0.01fF
C73 a_n683_n194# a_919_n194# 0.01fF
C74 a_505_n140# a_n741_n140# 0.01fF
C75 a_1039_n140# a_1453_n194# 0.02fF
C76 a_1395_n140# a_149_n140# 0.01fF
C77 a_505_n140# a_n385_n140# 0.01fF
C78 a_n207_n140# a_n1097_n140# 0.01fF
C79 a_1039_n140# a_1395_n140# 0.03fF
C80 a_n1631_n140# a_n505_n194# 0.01fF
C81 a_919_n194# a_385_n194# 0.02fF
C82 a_n207_n140# a_n563_n140# 0.03fF
C83 a_n327_n194# a_741_n194# 0.01fF
C84 a_505_n140# a_1453_n194# 0.01fF
C85 a_1453_n194# a_741_n194# 0.01fF
C86 a_n1395_n194# a_n1039_n194# 0.03fF
C87 a_n149_n194# a_n683_n194# 0.02fF
C88 a_505_n140# a_1395_n140# 0.01fF
C89 a_563_n194# a_29_n194# 0.02fF
C90 a_n919_n140# a_n29_n140# 0.01fF
C91 a_n1453_n140# a_n1631_n140# 0.06fF
C92 a_n1217_n194# a_n1395_n194# 0.10fF
C93 a_207_n194# a_n683_n194# 0.01fF
C94 a_n149_n194# a_385_n194# 0.02fF
C95 a_n861_n194# a_741_n194# 0.01fF
C96 a_n29_n140# a_683_n140# 0.01fF
C97 a_n29_n140# a_n1275_n140# 0.01fF
C98 a_327_n140# a_n919_n140# 0.01fF
C99 a_n683_n194# a_n505_n194# 0.10fF
C100 a_861_n140# a_683_n140# 0.06fF
C101 a_327_n140# a_683_n140# 0.03fF
C102 a_1097_n194# a_1275_n194# 0.10fF
C103 a_327_n140# a_n1275_n140# 0.01fF
C104 a_207_n194# a_385_n194# 0.10fF
C105 a_n327_n194# a_n1039_n194# 0.01fF
C106 a_n29_n140# a_n1097_n140# 0.01fF
C107 a_385_n194# a_n505_n194# 0.01fF
C108 a_327_n140# a_n1097_n140# 0.01fF
C109 a_n683_n194# a_n1631_n140# 0.01fF
C110 a_n29_n140# a_n563_n140# 0.02fF
C111 a_n327_n194# a_n1217_n194# 0.01fF
C112 a_n861_n194# a_n1039_n194# 0.10fF
C113 a_861_n140# a_n563_n140# 0.01fF
C114 a_327_n140# a_n563_n140# 0.01fF
C115 a_n919_n140# a_149_n140# 0.01fF
C116 a_n861_n194# a_n1217_n194# 0.03fF
C117 a_683_n140# a_149_n140# 0.02fF
C118 a_149_n140# a_n1275_n140# 0.01fF
C119 a_29_n194# a_741_n194# 0.01fF
C120 a_1039_n140# a_683_n140# 0.03fF
C121 a_n207_n140# a_1217_n140# 0.01fF
C122 a_n207_n140# a_n1631_n140# 0.01fF
C123 a_563_n194# a_919_n194# 0.03fF
C124 a_n207_n140# a_n1453_n140# 0.01fF
C125 a_149_n140# a_n1097_n140# 0.01fF
C126 a_n327_n194# a_1275_n194# 0.01fF
C127 a_1275_n194# a_1453_n194# 0.06fF
C128 a_n919_n140# a_505_n140# 0.01fF
C129 a_n683_n194# a_385_n194# 0.01fF
C130 a_n563_n140# a_149_n140# 0.01fF
C131 a_505_n140# a_683_n140# 0.06fF
C132 a_1097_n194# a_n327_n194# 0.01fF
C133 a_1097_n194# a_1453_n194# 0.02fF
C134 a_n149_n194# a_563_n194# 0.01fF
C135 a_1039_n140# a_n563_n140# 0.01fF
C136 a_29_n194# a_n1039_n194# 0.01fF
C137 a_505_n140# a_n1097_n140# 0.01fF
C138 a_207_n194# a_563_n194# 0.03fF
C139 a_n385_n140# a_n741_n140# 0.03fF
C140 a_29_n194# a_n1217_n194# 0.01fF
C141 a_n327_n194# a_n1395_n194# 0.01fF
C142 a_505_n140# a_n563_n140# 0.01fF
C143 a_563_n194# a_n505_n194# 0.01fF
C144 a_n29_n140# a_1217_n140# 0.01fF
C145 a_n29_n140# a_n1631_n140# 0.01fF
C146 a_n29_n140# a_n1453_n140# 0.01fF
C147 a_861_n140# a_1217_n140# 0.03fF
C148 a_327_n140# a_1217_n140# 0.01fF
C149 a_919_n194# a_741_n194# 0.10fF
C150 a_n861_n194# a_n1395_n194# 0.02fF
C151 a_1275_n194# a_29_n194# 0.01fF
C152 a_n149_n194# a_741_n194# 0.01fF
C153 a_1453_n194# a_1395_n140# 0.06fF
C154 a_1097_n194# a_29_n194# 0.01fF
C155 a_n327_n194# a_n861_n194# 0.02fF
C156 a_1217_n140# a_149_n140# 0.01fF
C157 a_207_n194# a_741_n194# 0.02fF
C158 a_n1453_n140# a_149_n140# 0.01fF
C159 a_563_n194# a_n683_n194# 0.01fF
C160 a_741_n194# a_n505_n194# 0.01fF
C161 a_1039_n140# a_1217_n140# 0.06fF
C162 a_n207_n140# a_n29_n140# 0.06fF
C163 a_29_n194# a_n1395_n194# 0.01fF
C164 a_563_n194# a_385_n194# 0.10fF
C165 a_n149_n194# a_n1039_n194# 0.01fF
C166 a_n207_n140# a_861_n140# 0.01fF
C167 a_327_n140# a_n207_n140# 0.02fF
C168 a_505_n140# a_1217_n140# 0.01fF
C169 a_n149_n194# a_n1217_n194# 0.01fF
C170 a_207_n194# a_n1039_n194# 0.01fF
C171 a_n1039_n194# a_n505_n194# 0.02fF
C172 a_1275_n194# a_919_n194# 0.03fF
C173 a_207_n194# a_n1217_n194# 0.01fF
C174 a_n327_n194# a_29_n194# 0.03fF
C175 a_n919_n140# a_n741_n140# 0.06fF
C176 a_29_n194# a_1453_n194# 0.00fF
C177 a_n919_n140# a_n385_n140# 0.02fF
C178 a_683_n140# a_n741_n140# 0.01fF
C179 a_n1217_n194# a_n505_n194# 0.01fF
C180 a_n1275_n140# a_n741_n140# 0.02fF
C181 a_n385_n140# a_683_n140# 0.01fF
C182 a_1097_n194# a_919_n194# 0.10fF
C183 a_n683_n194# a_741_n194# 0.01fF
C184 a_n385_n140# a_n1275_n140# 0.01fF
C185 a_n207_n140# a_149_n140# 0.03fF
C186 a_n1631_n140# a_n1039_n194# 0.01fF
C187 a_29_n194# a_n861_n194# 0.01fF
C188 a_n149_n194# a_1275_n194# 0.01fF
C189 a_n1097_n140# a_n741_n140# 0.03fF
C190 a_n29_n140# a_861_n140# 0.01fF
C191 a_n207_n140# a_1039_n140# 0.01fF
C192 a_327_n140# a_n29_n140# 0.03fF
C193 a_n385_n140# a_n1097_n140# 0.01fF
C194 a_683_n140# a_1453_n194# 0.01fF
C195 a_741_n194# a_385_n194# 0.03fF
C196 a_n1217_n194# a_n1631_n140# 0.02fF
C197 a_327_n140# a_861_n140# 0.02fF
C198 a_1097_n194# a_n149_n194# 0.01fF
C199 a_n563_n140# a_n741_n140# 0.06fF
C200 a_207_n194# a_1275_n194# 0.01fF
C201 a_683_n140# a_1395_n140# 0.01fF
C202 a_n385_n140# a_n563_n140# 0.06fF
C203 a_n207_n140# a_505_n140# 0.01fF
C204 a_n683_n194# a_n1039_n194# 0.03fF
C205 a_1097_n194# a_207_n194# 0.01fF
C206 a_1097_n194# a_n505_n194# 0.01fF
C207 a_n149_n194# a_n1395_n194# 0.01fF
C208 a_n1039_n194# a_385_n194# 0.01fF
C209 a_n683_n194# a_n1217_n194# 0.02fF
C210 a_n29_n140# a_149_n140# 0.06fF
C211 a_n327_n194# a_919_n194# 0.01fF
C212 a_1453_n194# a_919_n194# 0.01fF
C213 a_861_n140# a_149_n140# 0.01fF
C214 a_207_n194# a_n1395_n194# 0.01fF
C215 a_327_n140# a_149_n140# 0.06fF
C216 a_n29_n140# a_1039_n140# 0.01fF
C217 a_n1217_n194# a_385_n194# 0.01fF
C218 a_n1395_n194# a_n505_n194# 0.01fF
C219 a_861_n140# a_1039_n140# 0.06fF
C220 a_327_n140# a_1039_n140# 0.01fF
C221 a_n149_n194# a_n327_n194# 0.10fF
C222 a_n149_n194# a_1453_n194# 0.00fF
C223 a_n29_n140# a_505_n140# 0.02fF
C224 a_505_n140# a_861_n140# 0.03fF
C225 a_n1631_n140# a_n1395_n194# 0.06fF
C226 a_327_n140# a_505_n140# 0.06fF
C227 a_207_n194# a_n327_n194# 0.02fF
C228 a_207_n194# a_1453_n194# 0.00fF
C229 a_n149_n194# a_n861_n194# 0.01fF
C230 a_n327_n194# a_n505_n194# 0.10fF
C231 a_1275_n194# a_385_n194# 0.01fF
C232 a_563_n194# a_741_n194# 0.10fF
C233 a_n1631_n140# a_n741_n140# 0.01fF
C234 a_n919_n140# a_683_n140# 0.01fF
C235 a_n1453_n140# a_n741_n140# 0.01fF
C236 a_n385_n140# a_1217_n140# 0.01fF
C237 a_n385_n140# a_n1631_n140# 0.01fF
C238 a_n919_n140# a_n1275_n140# 0.03fF
C239 a_n385_n140# a_n1453_n140# 0.01fF
C240 a_1039_n140# a_149_n140# 0.01fF
C241 a_207_n194# a_n861_n194# 0.01fF
C242 a_1097_n194# a_385_n194# 0.01fF
C243 a_1395_n140# VSUBS 0.01fF
C244 a_1217_n140# VSUBS 0.01fF
C245 a_1039_n140# VSUBS 0.02fF
C246 a_861_n140# VSUBS 0.02fF
C247 a_683_n140# VSUBS 0.02fF
C248 a_505_n140# VSUBS 0.02fF
C249 a_327_n140# VSUBS 0.02fF
C250 a_149_n140# VSUBS 0.02fF
C251 a_n29_n140# VSUBS 0.02fF
C252 a_n207_n140# VSUBS 0.02fF
C253 a_n385_n140# VSUBS 0.02fF
C254 a_n563_n140# VSUBS 0.02fF
C255 a_n741_n140# VSUBS 0.02fF
C256 a_n919_n140# VSUBS 0.02fF
C257 a_n1097_n140# VSUBS 0.02fF
C258 a_n1275_n140# VSUBS 0.02fF
C259 a_n1453_n140# VSUBS 0.02fF
C260 a_1453_n194# VSUBS 0.31fF
C261 a_1275_n194# VSUBS 0.19fF
C262 a_1097_n194# VSUBS 0.20fF
C263 a_919_n194# VSUBS 0.21fF
C264 a_741_n194# VSUBS 0.22fF
C265 a_563_n194# VSUBS 0.23fF
C266 a_385_n194# VSUBS 0.23fF
C267 a_207_n194# VSUBS 0.24fF
C268 a_29_n194# VSUBS 0.24fF
C269 a_n149_n194# VSUBS 0.24fF
C270 a_n327_n194# VSUBS 0.24fF
C271 a_n505_n194# VSUBS 0.24fF
C272 a_n683_n194# VSUBS 0.24fF
C273 a_n861_n194# VSUBS 0.24fF
C274 a_n1039_n194# VSUBS 0.24fF
C275 a_n1217_n194# VSUBS 0.24fF
C276 a_n1395_n194# VSUBS 0.24fF
C277 a_n1631_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6RUDQZ a_n594_n195# a_n1008_n140# a_n652_n140# a_652_n195#
+ a_772_n140# a_n60_n195# a_n474_n140# a_n416_n195# a_474_n195# a_594_n140# a_n296_n140#
+ a_n238_n195# a_60_n140# a_296_n195# a_416_n140# a_n118_n140# a_118_n195# a_238_n140#
+ a_n772_n195# a_n830_n140# a_830_n195# VSUBS
X0 a_772_n140# a_652_n195# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n195# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n195# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n195# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n195# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_830_n195# a_830_n195# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n1008_n140# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n195# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n195# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n195# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n195# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_594_n140# a_238_n140# 0.03fF
C1 a_n594_n195# a_n238_n195# 0.03fF
C2 a_n238_n195# a_830_n195# 0.01fF
C3 a_n830_n140# a_772_n140# 0.01fF
C4 a_n60_n195# a_652_n195# 0.01fF
C5 a_n118_n140# a_n296_n140# 0.06fF
C6 a_n772_n195# a_652_n195# 0.01fF
C7 a_60_n140# a_416_n140# 0.03fF
C8 a_n594_n195# a_830_n195# 0.00fF
C9 a_n474_n140# a_n296_n140# 0.06fF
C10 a_60_n140# a_n652_n140# 0.01fF
C11 a_n296_n140# a_238_n140# 0.02fF
C12 a_594_n140# a_416_n140# 0.06fF
C13 a_296_n195# a_n1008_n140# 0.00fF
C14 a_n416_n195# a_296_n195# 0.01fF
C15 a_594_n140# a_n652_n140# 0.01fF
C16 a_474_n195# a_n1008_n140# 0.00fF
C17 a_474_n195# a_n416_n195# 0.01fF
C18 a_830_n195# a_772_n140# 0.06fF
C19 a_296_n195# a_n238_n195# 0.02fF
C20 a_n296_n140# a_416_n140# 0.01fF
C21 a_474_n195# a_n238_n195# 0.01fF
C22 a_n296_n140# a_n652_n140# 0.03fF
C23 a_60_n140# a_n1008_n140# 0.01fF
C24 a_296_n195# a_830_n195# 0.01fF
C25 a_n1008_n140# a_118_n195# 0.01fF
C26 a_n594_n195# a_296_n195# 0.01fF
C27 a_n416_n195# a_118_n195# 0.02fF
C28 a_n118_n140# a_n474_n140# 0.03fF
C29 a_n830_n140# a_60_n140# 0.01fF
C30 a_474_n195# a_830_n195# 0.02fF
C31 a_474_n195# a_n594_n195# 0.01fF
C32 a_n1008_n140# a_594_n140# 0.01fF
C33 a_n118_n140# a_238_n140# 0.03fF
C34 a_n830_n140# a_594_n140# 0.01fF
C35 a_n474_n140# a_238_n140# 0.01fF
C36 a_118_n195# a_n238_n195# 0.03fF
C37 a_n1008_n140# a_n296_n140# 0.01fF
C38 a_60_n140# a_830_n195# 0.01fF
C39 a_n594_n195# a_118_n195# 0.01fF
C40 a_118_n195# a_830_n195# 0.01fF
C41 a_n118_n140# a_416_n140# 0.02fF
C42 a_n830_n140# a_n296_n140# 0.02fF
C43 a_n474_n140# a_416_n140# 0.01fF
C44 a_n118_n140# a_n652_n140# 0.02fF
C45 a_594_n140# a_830_n195# 0.03fF
C46 a_n60_n195# a_n1008_n140# 0.01fF
C47 a_n416_n195# a_n60_n195# 0.03fF
C48 a_416_n140# a_238_n140# 0.06fF
C49 a_n1008_n140# a_n772_n195# 0.06fF
C50 a_n416_n195# a_n772_n195# 0.03fF
C51 a_474_n195# a_296_n195# 0.10fF
C52 a_n474_n140# a_n652_n140# 0.06fF
C53 a_60_n140# a_772_n140# 0.01fF
C54 a_n652_n140# a_238_n140# 0.01fF
C55 a_594_n140# a_772_n140# 0.06fF
C56 a_n60_n195# a_n238_n195# 0.10fF
C57 a_n1008_n140# a_652_n195# 0.00fF
C58 a_n772_n195# a_n238_n195# 0.02fF
C59 a_n416_n195# a_652_n195# 0.01fF
C60 a_n296_n140# a_830_n195# 0.01fF
C61 a_296_n195# a_118_n195# 0.10fF
C62 a_n118_n140# a_n1008_n140# 0.01fF
C63 a_n60_n195# a_830_n195# 0.01fF
C64 a_n60_n195# a_n594_n195# 0.02fF
C65 a_416_n140# a_n652_n140# 0.01fF
C66 a_n772_n195# a_830_n195# 0.00fF
C67 a_n594_n195# a_n772_n195# 0.10fF
C68 a_474_n195# a_118_n195# 0.03fF
C69 a_n118_n140# a_n830_n140# 0.01fF
C70 a_n474_n140# a_n1008_n140# 0.02fF
C71 a_n296_n140# a_772_n140# 0.01fF
C72 a_652_n195# a_n238_n195# 0.01fF
C73 a_n1008_n140# a_238_n140# 0.01fF
C74 a_n474_n140# a_n830_n140# 0.03fF
C75 a_n830_n140# a_238_n140# 0.01fF
C76 a_652_n195# a_830_n195# 0.06fF
C77 a_n594_n195# a_652_n195# 0.01fF
C78 a_n118_n140# a_830_n195# 0.01fF
C79 a_n1008_n140# a_416_n140# 0.01fF
C80 a_60_n140# a_594_n140# 0.02fF
C81 a_n60_n195# a_296_n195# 0.03fF
C82 a_n474_n140# a_830_n195# 0.01fF
C83 a_n830_n140# a_416_n140# 0.01fF
C84 a_296_n195# a_n772_n195# 0.01fF
C85 a_n1008_n140# a_n652_n140# 0.03fF
C86 a_830_n195# a_238_n140# 0.01fF
C87 a_474_n195# a_n60_n195# 0.02fF
C88 a_n830_n140# a_n652_n140# 0.06fF
C89 a_474_n195# a_n772_n195# 0.01fF
C90 a_n118_n140# a_772_n140# 0.01fF
C91 a_n474_n140# a_772_n140# 0.01fF
C92 a_772_n140# a_238_n140# 0.02fF
C93 a_296_n195# a_652_n195# 0.03fF
C94 a_60_n140# a_n296_n140# 0.03fF
C95 a_474_n195# a_652_n195# 0.10fF
C96 a_416_n140# a_830_n195# 0.02fF
C97 a_n296_n140# a_594_n140# 0.01fF
C98 a_n60_n195# a_118_n195# 0.10fF
C99 a_n772_n195# a_118_n195# 0.01fF
C100 a_830_n195# a_n652_n140# 0.01fF
C101 a_n416_n195# a_n1008_n140# 0.01fF
C102 a_n830_n140# a_n1008_n140# 0.06fF
C103 a_416_n140# a_772_n140# 0.03fF
C104 a_772_n140# a_n652_n140# 0.01fF
C105 a_118_n195# a_652_n195# 0.02fF
C106 a_n1008_n140# a_n238_n195# 0.01fF
C107 a_n416_n195# a_n238_n195# 0.10fF
C108 a_n118_n140# a_60_n140# 0.06fF
C109 a_n594_n195# a_n1008_n140# 0.02fF
C110 a_n416_n195# a_830_n195# 0.00fF
C111 a_n416_n195# a_n594_n195# 0.10fF
C112 a_n474_n140# a_60_n140# 0.02fF
C113 a_n118_n140# a_594_n140# 0.01fF
C114 a_60_n140# a_238_n140# 0.06fF
C115 a_n60_n195# a_n772_n195# 0.01fF
C116 a_n474_n140# a_594_n140# 0.01fF
C117 a_772_n140# VSUBS 0.01fF
C118 a_594_n140# VSUBS 0.01fF
C119 a_416_n140# VSUBS 0.02fF
C120 a_238_n140# VSUBS 0.02fF
C121 a_60_n140# VSUBS 0.02fF
C122 a_n118_n140# VSUBS 0.02fF
C123 a_n296_n140# VSUBS 0.02fF
C124 a_n474_n140# VSUBS 0.02fF
C125 a_n652_n140# VSUBS 0.02fF
C126 a_n830_n140# VSUBS 0.02fF
C127 a_830_n195# VSUBS 0.31fF
C128 a_652_n195# VSUBS 0.19fF
C129 a_474_n195# VSUBS 0.20fF
C130 a_296_n195# VSUBS 0.21fF
C131 a_118_n195# VSUBS 0.22fF
C132 a_n60_n195# VSUBS 0.23fF
C133 a_n238_n195# VSUBS 0.23fF
C134 a_n416_n195# VSUBS 0.24fF
C135 a_n594_n195# VSUBS 0.24fF
C136 a_n772_n195# VSUBS 0.24fF
C137 a_n1008_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_SD55Q9 a_352_607# a_644_607# a_174_607# a_60_607#
+ a_232_553# a_n232_n389# a_466_607# a_n524_n389# a_524_553# a_n410_n887# a_n702_n887#
+ a_n994_n887# a_644_n389# a_352_n389# a_60_n389# a_524_55# a_n60_55# a_n352_55# a_n232_n887#
+ a_n524_n887# a_174_n389# a_n352_n445# a_466_n389# a_n60_n445# a_n644_n445# a_644_n887#
+ a_352_n887# a_n118_n389# a_60_n887# a_174_n887# a_n352_n943# a_466_n887# a_n118_n887#
+ a_n60_n943# a_n644_n943# a_232_n445# a_n118_109# a_n410_109# a_758_n887# a_524_n445#
+ a_n232_109# a_n702_109# a_n644_55# a_n524_109# a_352_109# a_232_55# a_n352_553#
+ a_644_109# a_174_109# a_60_109# a_n644_553# a_n60_553# a_466_109# a_n410_607# a_524_n943#
+ a_232_n943# a_n410_n389# a_n118_607# a_n702_n389# a_n232_607# a_n702_607# a_n524_607#
+ VSUBS
X0 a_60_n389# a_n60_n445# a_n118_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_644_n887# a_524_n943# a_466_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_644_607# a_524_553# a_466_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n524_607# a_n644_553# a_n702_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_352_n389# a_232_n445# a_174_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_644_n389# a_524_n445# a_466_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n232_n887# a_n352_n943# a_n410_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_644_109# a_524_55# a_466_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n524_n887# a_n644_n943# a_n702_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_352_607# a_232_553# a_174_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n524_109# a_n644_55# a_n702_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n232_607# a_n352_553# a_n410_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n232_n389# a_n352_n445# a_n410_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n524_n389# a_n644_n445# a_n702_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_60_607# a_n60_553# a_n118_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_352_109# a_232_55# a_174_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n232_109# a_n352_55# a_n410_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_60_n887# a_n60_n943# a_n118_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_60_109# a_n60_55# a_n118_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_352_n887# a_232_n943# a_174_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_232_n445# a_232_553# 0.03fF
C1 a_n352_553# a_n994_n887# 0.02fF
C2 a_174_n389# a_n994_n887# 0.04fF
C3 a_758_n887# a_n994_n887# 0.07fF
C4 a_n410_607# a_n410_n389# 0.00fF
C5 a_n60_553# a_232_553# 0.04fF
C6 a_174_n887# a_n994_n887# 0.04fF
C7 a_n232_607# a_466_607# 0.03fF
C8 a_n524_109# a_352_109# 0.02fF
C9 a_60_109# a_352_109# 0.07fF
C10 a_174_n389# a_174_109# 0.01fF
C11 a_758_n887# a_174_109# 0.06fF
C12 a_n352_553# a_n352_n445# 0.03fF
C13 a_n994_n887# a_60_607# 0.04fF
C14 a_n524_109# a_644_109# 0.02fF
C15 a_174_n887# a_174_109# 0.00fF
C16 a_n352_n445# a_758_n887# 0.01fF
C17 a_524_553# a_n644_553# 0.01fF
C18 a_524_n445# a_n994_n887# 0.01fF
C19 a_524_n943# a_n994_n887# 0.01fF
C20 a_644_109# a_60_109# 0.03fF
C21 a_n118_n887# a_644_n887# 0.03fF
C22 a_n702_109# a_466_109# 0.02fF
C23 a_644_n887# a_644_n389# 0.01fF
C24 a_n410_n389# a_60_n389# 0.04fF
C25 a_n702_n389# a_352_n389# 0.02fF
C26 a_n644_n445# a_n644_553# 0.03fF
C27 a_n410_607# a_n232_607# 0.13fF
C28 a_n352_553# a_n352_55# 0.15fF
C29 a_n60_n445# a_n994_n887# 0.01fF
C30 a_644_109# a_352_109# 0.07fF
C31 a_n524_607# a_758_n887# 0.03fF
C32 a_n352_55# a_758_n887# 0.01fF
C33 a_524_n445# a_n352_n445# 0.01fF
C34 a_n524_n887# a_60_n887# 0.03fF
C35 a_n702_n389# a_n524_n389# 0.13fF
C36 a_n60_n943# a_n60_55# 0.03fF
C37 a_n118_607# a_n232_607# 0.25fF
C38 a_232_55# a_232_553# 0.15fF
C39 a_n702_n887# a_n702_n389# 0.01fF
C40 a_n352_553# a_524_553# 0.01fF
C41 a_n524_607# a_60_607# 0.03fF
C42 a_n60_n445# a_n352_n445# 0.04fF
C43 a_352_n389# a_n994_n887# 0.03fF
C44 a_n232_607# a_n702_607# 0.04fF
C45 a_524_553# a_758_n887# 0.05fF
C46 a_352_n887# a_n994_n887# 0.03fF
C47 a_524_55# a_n644_55# 0.01fF
C48 a_n118_n389# a_n118_607# 0.00fF
C49 a_n644_n445# a_758_n887# 0.01fF
C50 a_n524_n389# a_n994_n887# 0.12fF
C51 a_n118_n389# a_60_n389# 0.13fF
C52 a_n644_n943# a_n60_n943# 0.02fF
C53 a_524_n445# a_524_553# 0.03fF
C54 a_524_n943# a_524_553# 0.01fF
C55 a_n702_n887# a_n994_n887# 0.33fF
C56 a_n232_607# a_n232_109# 0.01fF
C57 a_n232_n887# a_60_n887# 0.07fF
C58 a_n410_n389# a_174_n389# 0.03fF
C59 a_n702_n389# a_466_n389# 0.02fF
C60 a_524_n445# a_n644_n445# 0.01fF
C61 a_n410_n389# a_758_n887# 0.03fF
C62 a_644_607# a_174_607# 0.04fF
C63 a_n702_n389# a_n232_n389# 0.04fF
C64 a_60_n389# a_60_109# 0.01fF
C65 a_232_n445# a_n994_n887# 0.01fF
C66 a_n524_n887# a_758_n887# 0.03fF
C67 a_60_n887# a_60_109# 0.00fF
C68 a_n118_n389# a_n118_109# 0.01fF
C69 a_n524_n887# a_174_n887# 0.03fF
C70 a_n410_109# a_n994_n887# 0.08fF
C71 a_n60_553# a_n994_n887# 0.01fF
C72 a_n232_n887# a_n232_109# 0.00fF
C73 a_524_55# a_n994_n887# 0.01fF
C74 a_n60_n445# a_n644_n445# 0.02fF
C75 a_n644_55# a_232_55# 0.01fF
C76 a_n410_607# a_466_607# 0.02fF
C77 a_n524_n389# a_n524_607# 0.00fF
C78 a_n524_109# a_n232_109# 0.07fF
C79 a_232_n445# a_n352_n445# 0.02fF
C80 a_466_n389# a_n994_n887# 0.03fF
C81 a_n524_109# a_n118_109# 0.05fF
C82 a_n232_109# a_60_109# 0.07fF
C83 a_174_607# a_n994_n887# 0.04fF
C84 a_n410_109# a_174_109# 0.03fF
C85 a_n118_109# a_60_109# 0.13fF
C86 a_n232_n389# a_n994_n887# 0.06fF
C87 a_466_n887# a_n994_n887# 0.03fF
C88 a_n232_607# a_758_n887# 0.04fF
C89 a_n410_n887# a_n994_n887# 0.08fF
C90 a_n118_607# a_466_607# 0.03fF
C91 a_n232_109# a_352_109# 0.03fF
C92 a_n118_n389# a_174_n389# 0.07fF
C93 a_174_607# a_174_109# 0.01fF
C94 a_466_607# a_n702_607# 0.02fF
C95 a_n118_109# a_352_109# 0.04fF
C96 a_n118_n389# a_758_n887# 0.04fF
C97 a_n644_n943# a_232_n943# 0.01fF
C98 a_n644_n943# a_n644_553# 0.01fF
C99 a_n232_607# a_60_607# 0.07fF
C100 a_n232_n887# a_758_n887# 0.04fF
C101 a_n232_n887# a_174_n887# 0.05fF
C102 a_n60_55# a_758_n887# 0.01fF
C103 a_524_55# a_n352_55# 0.01fF
C104 a_644_109# a_n232_109# 0.02fF
C105 a_n410_n389# a_352_n389# 0.03fF
C106 a_n702_n389# a_644_n389# 0.01fF
C107 a_644_607# a_644_n389# 0.00fF
C108 a_644_109# a_n118_109# 0.03fF
C109 a_n524_109# a_758_n887# 0.03fF
C110 a_232_55# a_n994_n887# 0.01fF
C111 a_644_607# a_644_n887# 0.00fF
C112 a_n410_607# a_n118_607# 0.07fF
C113 a_758_n887# a_60_109# 0.05fF
C114 a_174_607# a_n524_607# 0.03fF
C115 a_n524_n887# a_352_n887# 0.02fF
C116 a_n702_n389# a_n702_109# 0.01fF
C117 a_644_607# a_352_607# 0.07fF
C118 a_n410_607# a_n702_607# 0.07fF
C119 a_n60_553# a_524_553# 0.02fF
C120 a_524_55# a_524_553# 0.15fF
C121 a_n524_n389# a_n410_n389# 0.25fF
C122 a_232_n445# a_n644_n445# 0.01fF
C123 a_466_109# a_n994_n887# 0.03fF
C124 a_n118_n887# a_n994_n887# 0.05fF
C125 a_758_n887# a_352_109# 0.08fF
C126 a_n524_n887# a_n524_n389# 0.01fF
C127 a_60_109# a_60_607# 0.01fF
C128 a_644_n389# a_n994_n887# 0.02fF
C129 a_n644_n943# a_758_n887# 0.01fF
C130 a_n702_n887# a_n524_n887# 0.13fF
C131 a_644_n887# a_n994_n887# 0.02fF
C132 a_n118_607# a_n702_607# 0.03fF
C133 a_n60_n943# a_232_n943# 0.04fF
C134 a_466_109# a_174_109# 0.07fF
C135 a_n60_55# a_n60_n445# 0.15fF
C136 a_758_n887# a_644_109# 0.33fF
C137 a_n994_n887# a_352_607# 0.03fF
C138 a_n702_109# a_n994_n887# 0.33fF
C139 a_n352_55# a_232_55# 0.02fF
C140 a_n118_n389# a_352_n389# 0.04fF
C141 a_n410_n389# a_n410_109# 0.01fF
C142 a_n644_n943# a_524_n943# 0.01fF
C143 a_758_n887# a_466_607# 0.12fF
C144 a_60_n887# a_60_n389# 0.01fF
C145 a_n702_109# a_174_109# 0.02fF
C146 a_n352_n943# a_n994_n887# 0.02fF
C147 a_n232_n887# a_352_n887# 0.03fF
C148 a_n410_n389# a_466_n389# 0.02fF
C149 a_n118_607# a_n118_109# 0.01fF
C150 a_n524_n389# a_n118_n389# 0.05fF
C151 a_n410_n389# a_n232_n389# 0.13fF
C152 a_n410_n887# a_n410_n389# 0.01fF
C153 a_466_607# a_60_607# 0.05fF
C154 a_n524_n887# a_466_n887# 0.02fF
C155 a_n60_n943# a_758_n887# 0.01fF
C156 a_n524_n887# a_n410_n887# 0.25fF
C157 a_n702_n887# a_n232_n887# 0.04fF
C158 a_n352_n943# a_n352_n445# 0.15fF
C159 a_n524_n389# a_n524_109# 0.01fF
C160 a_n524_607# a_352_607# 0.02fF
C161 a_n994_n887# a_232_553# 0.01fF
C162 a_n410_607# a_758_n887# 0.03fF
C163 a_352_n389# a_352_109# 0.01fF
C164 a_352_n887# a_352_109# 0.00fF
C165 a_n60_n943# a_524_n943# 0.02fF
C166 a_174_607# a_n232_607# 0.05fF
C167 a_n232_n389# a_n232_607# 0.00fF
C168 a_n232_109# a_n118_109# 0.25fF
C169 a_n352_n943# a_n352_55# 0.03fF
C170 a_n410_607# a_60_607# 0.04fF
C171 a_n118_607# a_758_n887# 0.04fF
C172 a_n60_55# a_n60_553# 0.15fF
C173 a_524_55# a_n60_55# 0.02fF
C174 a_n118_n389# a_466_n389# 0.03fF
C175 a_758_n887# a_n702_607# 0.02fF
C176 a_60_n389# a_174_n389# 0.25fF
C177 a_n410_109# a_n524_109# 0.25fF
C178 a_n232_n389# a_n118_n389# 0.25fF
C179 a_758_n887# a_60_n389# 0.05fF
C180 a_n60_n943# a_n60_n445# 0.15fF
C181 a_n410_109# a_60_109# 0.04fF
C182 a_60_n887# a_758_n887# 0.05fF
C183 a_n232_n887# a_n232_n389# 0.01fF
C184 a_n118_607# a_60_607# 0.13fF
C185 a_n232_n887# a_466_n887# 0.03fF
C186 a_60_n887# a_174_n887# 0.25fF
C187 a_n410_n389# a_644_n389# 0.02fF
C188 a_n524_n887# a_n118_n887# 0.05fF
C189 a_n410_n887# a_n232_n887# 0.13fF
C190 a_60_607# a_n702_607# 0.03fF
C191 a_60_n389# a_60_607# 0.00fF
C192 a_n410_109# a_352_109# 0.03fF
C193 a_n352_553# a_n644_553# 0.04fF
C194 a_n524_n887# a_644_n887# 0.02fF
C195 a_758_n887# a_n232_109# 0.04fF
C196 a_60_n887# a_60_607# 0.00fF
C197 a_758_n887# a_n644_553# 0.01fF
C198 a_232_n943# a_758_n887# 0.02fF
C199 a_758_n887# a_n118_109# 0.04fF
C200 a_524_553# a_232_553# 0.04fF
C201 a_n644_55# a_n994_n887# 0.05fF
C202 a_n410_109# a_644_109# 0.02fF
C203 a_n60_55# a_232_55# 0.04fF
C204 a_232_n943# a_524_n943# 0.04fF
C205 a_n702_n389# a_n994_n887# 0.33fF
C206 a_644_607# a_n994_n887# 0.02fF
C207 a_n118_n887# a_n118_n389# 0.01fF
C208 a_n232_607# a_352_607# 0.03fF
C209 a_n118_n389# a_644_n389# 0.03fF
C210 a_60_n389# a_352_n389# 0.07fF
C211 a_n352_553# a_758_n887# 0.01fF
C212 a_n232_n887# a_n118_n887# 0.25fF
C213 a_758_n887# a_174_n389# 0.06fF
C214 a_466_n389# a_466_607# 0.00fF
C215 a_n524_109# a_466_109# 0.02fF
C216 a_174_n887# a_174_n389# 0.01fF
C217 a_174_607# a_466_607# 0.07fF
C218 a_174_n887# a_758_n887# 0.06fF
C219 a_466_n887# a_466_607# 0.00fF
C220 a_466_109# a_60_109# 0.05fF
C221 a_n232_n887# a_644_n887# 0.02fF
C222 a_60_n887# a_352_n887# 0.07fF
C223 a_n60_n943# a_n60_553# 0.01fF
C224 a_n644_55# a_n352_55# 0.04fF
C225 a_n524_n389# a_60_n389# 0.03fF
C226 a_n410_607# a_n410_109# 0.01fF
C227 a_n702_n887# a_n702_607# 0.00fF
C228 a_758_n887# a_60_607# 0.05fF
C229 a_466_109# a_352_109# 0.25fF
C230 a_n702_109# a_n524_109# 0.13fF
C231 a_524_n943# a_758_n887# 0.05fF
C232 a_524_n445# a_758_n887# 0.06fF
C233 a_644_607# a_n524_607# 0.02fF
C234 a_n702_109# a_60_109# 0.03fF
C235 a_n702_n887# a_60_n887# 0.03fF
C236 a_n994_n887# a_174_109# 0.04fF
C237 a_n410_607# a_174_607# 0.03fF
C238 a_n352_n445# a_n994_n887# 0.02fF
C239 a_644_109# a_466_109# 0.13fF
C240 a_n410_n887# a_n410_607# 0.00fF
C241 a_n60_n445# a_758_n887# 0.01fF
C242 a_n644_55# a_n644_n445# 0.15fF
C243 a_352_607# a_352_109# 0.01fF
C244 a_n702_109# a_352_109# 0.02fF
C245 a_524_n943# a_524_n445# 0.15fF
C246 a_644_109# a_644_n389# 0.01fF
C247 a_n118_607# a_174_607# 0.07fF
C248 a_644_n887# a_644_109# 0.00fF
C249 a_466_109# a_466_607# 0.01fF
C250 a_n524_607# a_n994_n887# 0.12fF
C251 a_n352_55# a_n994_n887# 0.02fF
C252 a_n702_109# a_644_109# 0.01fF
C253 a_174_607# a_n702_607# 0.02fF
C254 a_174_n389# a_352_n389# 0.13fF
C255 a_60_n389# a_466_n389# 0.05fF
C256 a_758_n887# a_352_n389# 0.08fF
C257 a_232_n943# a_232_n445# 0.15fF
C258 a_n60_n445# a_524_n445# 0.02fF
C259 a_n232_n389# a_60_n389# 0.07fF
C260 a_n644_n943# a_n352_n943# 0.04fF
C261 a_352_n887# a_758_n887# 0.08fF
C262 a_174_n887# a_352_n887# 0.13fF
C263 a_n410_109# a_n232_109# 0.13fF
C264 a_60_n887# a_466_n887# 0.05fF
C265 a_n60_553# a_n644_553# 0.02fF
C266 a_n410_109# a_n118_109# 0.07fF
C267 a_466_607# a_352_607# 0.25fF
C268 a_524_553# a_n994_n887# 0.01fF
C269 a_n410_n887# a_60_n887# 0.04fF
C270 a_n352_n445# a_n352_55# 0.15fF
C271 a_n524_n389# a_174_n389# 0.03fF
C272 a_n524_n389# a_758_n887# 0.03fF
C273 a_n702_n389# a_n410_n389# 0.07fF
C274 a_n702_n887# a_758_n887# 0.02fF
C275 a_n644_n445# a_n994_n887# 0.05fF
C276 a_n232_n389# a_n232_109# 0.01fF
C277 a_n702_n887# a_174_n887# 0.02fF
C278 a_232_n445# a_758_n887# 0.02fF
C279 a_n410_607# a_352_607# 0.03fF
C280 a_n118_n887# a_n118_607# 0.00fF
C281 a_n352_n445# a_n644_n445# 0.04fF
C282 a_n352_553# a_n60_553# 0.04fF
C283 a_n410_n389# a_n994_n887# 0.08fF
C284 a_n410_109# a_758_n887# 0.03fF
C285 a_n60_553# a_758_n887# 0.01fF
C286 a_524_55# a_758_n887# 0.05fF
C287 a_n352_n943# a_n60_n943# 0.04fF
C288 a_644_607# a_n232_607# 0.02fF
C289 a_n524_n887# a_n994_n887# 0.12fF
C290 a_232_n943# a_232_55# 0.03fF
C291 a_60_n389# a_644_n389# 0.03fF
C292 a_174_n389# a_466_n389# 0.07fF
C293 a_n118_607# a_352_607# 0.04fF
C294 a_n60_55# a_n644_55# 0.02fF
C295 a_n118_n887# a_60_n887# 0.13fF
C296 a_174_607# a_174_n389# 0.00fF
C297 a_758_n887# a_466_n389# 0.12fF
C298 a_n232_n389# a_174_n389# 0.05fF
C299 a_232_n445# a_524_n445# 0.04fF
C300 a_174_607# a_758_n887# 0.06fF
C301 a_352_n887# a_352_n389# 0.01fF
C302 a_n232_n389# a_758_n887# 0.04fF
C303 a_n702_n389# a_n118_n389# 0.03fF
C304 a_466_n887# a_758_n887# 0.12fF
C305 a_174_n887# a_174_607# 0.00fF
C306 a_352_607# a_n702_607# 0.02fF
C307 a_n702_109# a_n702_607# 0.01fF
C308 a_174_n887# a_466_n887# 0.07fF
C309 a_60_n887# a_644_n887# 0.03fF
C310 a_n410_n887# a_758_n887# 0.03fF
C311 a_524_55# a_524_n445# 0.15fF
C312 a_524_55# a_524_n943# 0.03fF
C313 a_n232_109# a_466_109# 0.03fF
C314 a_n410_n887# a_174_n887# 0.03fF
C315 a_466_109# a_n118_109# 0.03fF
C316 a_n524_n389# a_352_n389# 0.02fF
C317 a_n60_n445# a_232_n445# 0.04fF
C318 a_n232_607# a_n994_n887# 0.06fF
C319 a_n118_n887# a_n118_109# 0.00fF
C320 a_174_607# a_60_607# 0.25fF
C321 a_n60_n445# a_n60_553# 0.03fF
C322 a_n702_n887# a_352_n887# 0.02fF
C323 a_n644_n943# a_n644_55# 0.03fF
C324 a_n118_n389# a_n994_n887# 0.05fF
C325 a_n524_n887# a_n524_607# 0.00fF
C326 a_n702_109# a_n232_109# 0.04fF
C327 a_n702_109# a_n118_109# 0.03fF
C328 a_758_n887# a_232_55# 0.02fF
C329 a_n232_n887# a_n994_n887# 0.06fF
C330 a_n60_55# a_n994_n887# 0.01fF
C331 a_n524_109# a_n994_n887# 0.12fF
C332 a_n352_n943# a_232_n943# 0.02fF
C333 a_758_n887# a_466_109# 0.12fF
C334 a_60_109# a_n994_n887# 0.04fF
C335 a_644_607# a_644_109# 0.01fF
C336 a_n118_n887# a_758_n887# 0.04fF
C337 a_n524_607# a_n232_607# 0.07fF
C338 a_174_n389# a_644_n389# 0.04fF
C339 a_352_n389# a_466_n389# 0.25fF
C340 a_n118_n887# a_174_n887# 0.07fF
C341 a_758_n887# a_644_n389# 0.33fF
C342 a_n232_n389# a_352_n389# 0.03fF
C343 a_n524_109# a_174_109# 0.03fF
C344 a_644_n887# a_758_n887# 0.33fF
C345 a_n994_n887# a_352_109# 0.03fF
C346 a_60_109# a_174_109# 0.25fF
C347 a_352_n887# a_466_n887# 0.25fF
C348 a_174_n887# a_644_n887# 0.04fF
C349 a_644_607# a_466_607# 0.13fF
C350 a_758_n887# a_352_607# 0.08fF
C351 a_n644_n943# a_n994_n887# 0.05fF
C352 a_n702_109# a_758_n887# 0.02fF
C353 a_n410_n887# a_352_n887# 0.03fF
C354 a_232_n943# a_232_553# 0.01fF
C355 a_n644_553# a_232_553# 0.01fF
C356 a_n524_n389# a_466_n389# 0.02fF
C357 a_n524_n389# a_n232_n389# 0.07fF
C358 a_644_109# a_n994_n887# 0.02fF
C359 a_n60_55# a_n352_55# 0.04fF
C360 a_352_109# a_174_109# 0.13fF
C361 a_n352_553# a_n352_n943# 0.01fF
C362 a_n702_n887# a_466_n887# 0.02fF
C363 a_n524_607# a_n524_109# 0.01fF
C364 a_n352_n943# a_758_n887# 0.01fF
C365 a_352_607# a_60_607# 0.07fF
C366 a_n702_n887# a_n410_n887# 0.07fF
C367 a_466_607# a_n994_n887# 0.03fF
C368 a_644_607# a_n410_607# 0.02fF
C369 a_644_109# a_174_109# 0.04fF
C370 a_n352_553# a_232_553# 0.02fF
C371 a_n352_n943# a_524_n943# 0.01fF
C372 a_758_n887# a_232_553# 0.02fF
C373 a_644_607# a_n118_607# 0.03fF
C374 a_n410_n887# a_n410_109# 0.00fF
C375 a_n60_n943# a_n994_n887# 0.01fF
C376 a_352_n389# a_644_n389# 0.07fF
C377 a_n118_n887# a_352_n887# 0.04fF
C378 a_n232_n389# a_466_n389# 0.03fF
C379 a_n702_n389# a_n702_607# 0.00fF
C380 a_466_n887# a_466_n389# 0.01fF
C381 a_644_607# a_n702_607# 0.01fF
C382 a_n410_n389# a_n118_n389# 0.07fF
C383 a_n410_607# a_n994_n887# 0.08fF
C384 a_n702_n389# a_60_n389# 0.03fF
C385 a_352_n887# a_644_n887# 0.07fF
C386 a_352_n389# a_352_607# 0.00fF
C387 a_n410_n887# a_466_n887# 0.02fF
C388 a_232_n445# a_232_55# 0.15fF
C389 a_n644_55# a_n644_553# 0.15fF
C390 a_352_n887# a_352_607# 0.00fF
C391 a_n524_n389# a_644_n389# 0.02fF
C392 a_n524_607# a_466_607# 0.02fF
C393 a_n524_n887# a_n232_n887# 0.07fF
C394 a_n702_n887# a_n118_n887# 0.03fF
C395 a_n644_n943# a_n644_n445# 0.15fF
C396 a_n118_607# a_n994_n887# 0.05fF
C397 a_524_55# a_232_55# 0.04fF
C398 a_n524_n887# a_n524_109# 0.00fF
C399 a_n702_n887# a_644_n887# 0.01fF
C400 a_n994_n887# a_n702_607# 0.33fF
C401 a_60_n389# a_n994_n887# 0.04fF
C402 a_n702_n887# a_n702_109# 0.00fF
C403 a_n410_109# a_466_109# 0.02fF
C404 a_60_n887# a_n994_n887# 0.04fF
C405 a_n232_n887# a_n232_607# 0.00fF
C406 a_n410_607# a_n524_607# 0.25fF
C407 a_466_109# a_466_n389# 0.01fF
C408 a_n644_55# a_758_n887# 0.01fF
C409 a_466_n887# a_466_109# 0.00fF
C410 a_n702_109# a_n410_109# 0.07fF
C411 a_232_n943# a_n994_n887# 0.01fF
C412 a_n232_109# a_n994_n887# 0.06fF
C413 a_466_n389# a_644_n389# 0.13fF
C414 a_n644_553# a_n994_n887# 0.05fF
C415 a_n118_109# a_n994_n887# 0.05fF
C416 a_n118_n887# a_466_n887# 0.03fF
C417 a_n232_n389# a_644_n389# 0.02fF
C418 a_n118_607# a_n524_607# 0.05fF
C419 a_n410_n887# a_n118_n887# 0.07fF
C420 a_n702_n389# a_174_n389# 0.02fF
C421 a_466_n887# a_644_n887# 0.13fF
C422 a_644_607# a_758_n887# 0.33fF
C423 a_n702_n389# a_758_n887# 0.02fF
C424 a_n524_607# a_n702_607# 0.13fF
C425 a_174_607# a_352_607# 0.13fF
C426 a_n410_n887# a_644_n887# 0.02fF
C427 a_n232_109# a_174_109# 0.05fF
C428 a_n118_109# a_174_109# 0.07fF
C429 a_n524_109# a_60_109# 0.03fF
C430 a_644_607# a_60_607# 0.03fF
C431 a_644_n887# VSUBS 0.01fF
C432 a_466_n887# VSUBS 0.01fF
C433 a_352_n887# VSUBS 0.01fF
C434 a_174_n887# VSUBS 0.01fF
C435 a_60_n887# VSUBS 0.01fF
C436 a_n118_n887# VSUBS 0.01fF
C437 a_n232_n887# VSUBS 0.01fF
C438 a_n410_n887# VSUBS 0.01fF
C439 a_n524_n887# VSUBS 0.01fF
C440 a_n702_n887# VSUBS 0.01fF
C441 a_524_n943# VSUBS 0.17fF
C442 a_232_n943# VSUBS 0.19fF
C443 a_n60_n943# VSUBS 0.20fF
C444 a_n352_n943# VSUBS 0.21fF
C445 a_n644_n943# VSUBS 0.22fF
C446 a_644_n389# VSUBS 0.01fF
C447 a_466_n389# VSUBS 0.01fF
C448 a_352_n389# VSUBS 0.01fF
C449 a_174_n389# VSUBS 0.01fF
C450 a_60_n389# VSUBS 0.01fF
C451 a_n118_n389# VSUBS 0.01fF
C452 a_n232_n389# VSUBS 0.01fF
C453 a_n410_n389# VSUBS 0.01fF
C454 a_n524_n389# VSUBS 0.01fF
C455 a_n702_n389# VSUBS 0.01fF
C456 a_524_n445# VSUBS 0.16fF
C457 a_232_n445# VSUBS 0.17fF
C458 a_n60_n445# VSUBS 0.18fF
C459 a_n352_n445# VSUBS 0.19fF
C460 a_n644_n445# VSUBS 0.20fF
C461 a_644_109# VSUBS 0.01fF
C462 a_466_109# VSUBS 0.01fF
C463 a_352_109# VSUBS 0.01fF
C464 a_174_109# VSUBS 0.01fF
C465 a_60_109# VSUBS 0.01fF
C466 a_n118_109# VSUBS 0.01fF
C467 a_n232_109# VSUBS 0.01fF
C468 a_n410_109# VSUBS 0.01fF
C469 a_n524_109# VSUBS 0.01fF
C470 a_n702_109# VSUBS 0.01fF
C471 a_524_55# VSUBS 0.17fF
C472 a_232_55# VSUBS 0.18fF
C473 a_n60_55# VSUBS 0.19fF
C474 a_n352_55# VSUBS 0.20fF
C475 a_n644_55# VSUBS 0.21fF
C476 a_644_607# VSUBS 0.02fF
C477 a_466_607# VSUBS 0.02fF
C478 a_352_607# VSUBS 0.02fF
C479 a_174_607# VSUBS 0.02fF
C480 a_60_607# VSUBS 0.02fF
C481 a_n118_607# VSUBS 0.02fF
C482 a_n232_607# VSUBS 0.02fF
C483 a_n410_607# VSUBS 0.02fF
C484 a_n524_607# VSUBS 0.02fF
C485 a_n702_607# VSUBS 0.02fF
C486 a_758_n887# VSUBS 1.42fF
C487 a_524_553# VSUBS 0.20fF
C488 a_232_553# VSUBS 0.22fF
C489 a_n60_553# VSUBS 0.23fF
C490 a_n352_553# VSUBS 0.24fF
C491 a_n644_553# VSUBS 0.25fF
C492 a_n994_n887# VSUBS 1.66fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EZNTQN a_n830_109# a_n652_n887# a_n652_109# a_n772_55#
+ a_118_553# a_594_n389# a_n772_n445# a_60_607# a_772_n887# a_n474_109# a_772_109#
+ a_n296_109# a_n772_553# a_n296_n389# a_594_109# a_n594_55# a_n594_553# a_n474_n887#
+ a_118_n943# a_60_n389# a_n594_n445# a_n60_55# a_n830_607# a_n772_n943# a_416_n389#
+ a_n652_607# a_594_n887# a_652_n445# a_n416_55# a_n474_607# a_772_607# a_n296_607#
+ a_n60_n445# a_594_607# a_n296_n887# a_n118_n389# a_652_553# a_60_n887# a_n238_55#
+ a_474_553# a_n594_n943# a_238_n389# a_n416_n445# a_416_n887# a_474_n445# a_296_553#
+ a_652_n943# a_n830_n389# a_652_55# a_n118_n887# a_n60_n943# a_n118_109# a_n238_n445#
+ a_416_109# a_n416_553# a_296_n445# a_238_109# a_474_55# a_n238_553# a_238_n887#
+ a_n416_n943# a_n1110_n1061# a_474_n943# a_n652_n389# a_n830_n887# a_60_109# a_772_n389#
+ a_n60_553# a_296_55# a_n118_607# a_n238_n943# a_416_607# a_296_n943# a_n474_n389#
+ a_118_n445# a_118_55# a_238_607#
X0 a_n652_109# a_n772_55# a_n830_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_60_n389# a_n60_n445# a_n118_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_594_n389# a_474_n445# a_416_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1110_n1061# a_n1110_n1061# a_772_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n830_n887# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n474_n887# a_n594_n943# a_n652_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_594_607# a_474_553# a_416_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_109# a_n416_55# a_n474_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_416_n887# a_296_n943# a_238_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n474_607# a_n594_553# a_n652_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n296_n887# a_n416_n943# a_n474_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1110_n1061# a_n1110_n1061# a_772_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1110_n1061# a_n1110_n1061# a_772_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_238_607# a_118_553# a_60_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_238_n887# a_118_n943# a_60_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n830_n389# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n474_n389# a_n594_n445# a_n652_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n830_607# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n118_607# a_n238_553# a_n296_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_594_109# a_474_55# a_416_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_416_n389# a_296_n445# a_238_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_772_n887# a_652_n943# a_594_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n474_109# a_n594_55# a_n652_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n296_n389# a_n416_n445# a_n474_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1110_n1061# a_n1110_n1061# a_772_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_238_109# a_118_55# a_60_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_238_n389# a_118_n445# a_60_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_607# a_296_553# a_238_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n830_109# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n118_109# a_n238_55# a_n296_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n118_n887# a_n238_n943# a_n296_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_60_607# a_n60_553# a_n118_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_772_n389# a_652_n445# a_594_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_772_607# a_652_553# a_594_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_n652_n887# a_n772_n943# a_n830_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_594_n887# a_474_n943# a_416_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_n652_607# a_n772_553# a_n830_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_60_n887# a_n60_n943# a_n118_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_416_109# a_296_55# a_238_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n118_n389# a_n238_n445# a_n296_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_60_109# a_n60_55# a_n118_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X41 a_n296_607# a_n416_553# a_n474_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X42 a_772_109# a_652_55# a_594_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_n652_n389# a_n772_n445# a_n830_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_652_55# a_296_55# 0.03fF
C1 a_n416_553# a_n238_553# 0.10fF
C2 a_n60_n445# a_n60_n943# 0.15fF
C3 a_n772_553# a_n772_n943# 0.01fF
C4 a_n474_109# a_n118_109# 0.03fF
C5 a_652_n445# a_652_55# 0.15fF
C6 a_n652_109# a_n830_109# 0.06fF
C7 a_n474_n887# a_594_n887# 0.01fF
C8 a_n474_n887# a_n118_n887# 0.03fF
C9 a_n238_n943# a_474_n943# 0.01fF
C10 a_416_109# a_594_109# 0.06fF
C11 a_n594_n445# a_n594_553# 0.03fF
C12 a_652_n445# a_n594_n445# 0.01fF
C13 a_n296_607# a_772_607# 0.01fF
C14 a_n652_607# a_n296_607# 0.03fF
C15 a_n118_n887# a_n118_607# 0.00fF
C16 a_n118_n389# a_n830_n389# 0.01fF
C17 a_772_109# a_416_109# 0.03fF
C18 a_n830_n887# a_772_n887# 0.01fF
C19 a_n772_n943# a_n594_n943# 0.10fF
C20 a_60_n389# a_60_607# 0.00fF
C21 a_n60_n445# a_652_n445# 0.01fF
C22 a_n652_109# a_60_109# 0.01fF
C23 a_n238_n943# a_n416_n943# 0.10fF
C24 a_n118_607# a_594_607# 0.01fF
C25 a_238_n887# a_238_109# 0.00fF
C26 a_772_109# a_594_109# 0.06fF
C27 a_n60_55# a_n238_55# 0.10fF
C28 a_n830_607# a_594_607# 0.01fF
C29 a_238_n389# a_n474_n389# 0.01fF
C30 a_296_n445# a_118_n445# 0.10fF
C31 a_594_n887# a_594_109# 0.00fF
C32 a_n238_553# a_296_553# 0.02fF
C33 a_238_n389# a_772_n389# 0.02fF
C34 a_118_55# a_474_55# 0.03fF
C35 a_238_n389# a_n296_n389# 0.02fF
C36 a_n238_n445# a_118_n445# 0.03fF
C37 a_n652_607# a_772_607# 0.01fF
C38 a_296_n445# a_n238_n445# 0.02fF
C39 a_n118_n887# a_594_n887# 0.01fF
C40 a_416_n887# a_772_n887# 0.03fF
C41 a_474_n445# a_n772_n445# 0.01fF
C42 a_n416_55# a_n238_55# 0.10fF
C43 a_594_607# a_594_109# 0.00fF
C44 a_n772_n943# a_n60_n943# 0.01fF
C45 a_118_55# a_n594_55# 0.01fF
C46 a_n238_55# a_296_55# 0.02fF
C47 a_652_55# a_474_55# 0.10fF
C48 a_n772_n943# a_118_n943# 0.01fF
C49 a_n118_n389# a_n118_109# 0.00fF
C50 a_n474_607# a_238_607# 0.01fF
C51 a_n474_n887# a_772_n887# 0.01fF
C52 a_n238_n943# a_652_n943# 0.01fF
C53 a_n118_n389# a_238_n389# 0.03fF
C54 a_594_n887# a_594_607# 0.00fF
C55 a_n416_553# a_n60_553# 0.03fF
C56 a_296_n943# a_474_n943# 0.10fF
C57 a_652_55# a_n594_55# 0.01fF
C58 a_n416_553# a_652_553# 0.01fF
C59 a_416_607# a_n474_607# 0.01fF
C60 a_n594_n445# a_n594_55# 0.15fF
C61 a_296_n943# a_n416_n943# 0.01fF
C62 a_118_n943# a_118_n445# 0.15fF
C63 a_416_n887# a_416_n389# 0.00fF
C64 a_772_n887# a_772_109# 0.00fF
C65 a_n652_109# a_n118_109# 0.02fF
C66 a_594_n887# a_772_n887# 0.06fF
C67 a_n118_n887# a_772_n887# 0.01fF
C68 a_238_607# a_n296_607# 0.02fF
C69 a_n60_553# a_296_553# 0.03fF
C70 a_652_n445# a_118_n445# 0.02fF
C71 a_n416_n445# a_n772_n445# 0.03fF
C72 a_n594_n943# a_n60_n943# 0.02fF
C73 a_n772_553# a_n594_553# 0.10fF
C74 a_296_n943# a_296_553# 0.01fF
C75 a_296_n445# a_296_55# 0.15fF
C76 a_n296_109# a_416_109# 0.01fF
C77 a_652_n445# a_296_n445# 0.03fF
C78 a_n594_n943# a_118_n943# 0.01fF
C79 a_238_109# a_416_109# 0.06fF
C80 a_652_553# a_296_553# 0.03fF
C81 a_n238_55# a_474_55# 0.01fF
C82 a_652_n445# a_n238_n445# 0.01fF
C83 a_416_607# a_n296_607# 0.01fF
C84 a_n652_n887# a_60_n887# 0.01fF
C85 a_416_n389# a_416_109# 0.00fF
C86 a_296_n943# a_652_n943# 0.03fF
C87 a_n296_109# a_594_109# 0.01fF
C88 a_n474_109# a_n474_n887# 0.00fF
C89 a_238_109# a_594_109# 0.03fF
C90 a_n772_553# a_474_553# 0.01fF
C91 a_n594_n943# a_n594_553# 0.01fF
C92 a_652_n943# a_652_553# 0.01fF
C93 a_n416_553# a_118_553# 0.02fF
C94 a_n238_55# a_n594_55# 0.03fF
C95 a_772_109# a_n296_109# 0.01fF
C96 a_772_109# a_238_109# 0.02fF
C97 a_60_109# a_n830_109# 0.01fF
C98 a_n60_55# a_n60_n943# 0.03fF
C99 a_238_607# a_772_607# 0.02fF
C100 a_n238_553# a_n238_55# 0.15fF
C101 a_n652_607# a_238_607# 0.01fF
C102 a_n474_607# a_60_607# 0.02fF
C103 a_594_n389# a_594_109# 0.00fF
C104 a_n474_109# a_416_109# 0.01fF
C105 a_n238_n943# a_n238_55# 0.03fF
C106 a_118_n943# a_n60_n943# 0.10fF
C107 a_n60_55# a_n416_55# 0.03fF
C108 a_n772_55# a_118_55# 0.01fF
C109 a_416_607# a_772_607# 0.03fF
C110 a_416_607# a_n652_607# 0.01fF
C111 a_652_553# a_652_55# 0.15fF
C112 a_n60_55# a_296_55# 0.03fF
C113 a_n594_n445# a_n772_n445# 0.10fF
C114 a_594_n389# a_594_n887# 0.00fF
C115 a_n474_109# a_594_109# 0.01fF
C116 a_n772_n943# a_n238_n943# 0.02fF
C117 a_n296_n887# a_60_n887# 0.03fF
C118 a_n474_n887# a_n474_n389# 0.00fF
C119 a_n60_n445# a_n772_n445# 0.01fF
C120 a_n474_109# a_772_109# 0.01fF
C121 a_n60_n445# a_n60_553# 0.03fF
C122 a_n830_n389# a_n830_109# 0.00fF
C123 a_n772_55# a_652_55# 0.01fF
C124 a_594_n389# a_594_607# 0.00fF
C125 a_n416_55# a_296_55# 0.01fF
C126 a_118_553# a_296_553# 0.10fF
C127 a_n652_n887# a_238_n887# 0.01fF
C128 a_60_607# a_n296_607# 0.03fF
C129 a_n772_553# a_n238_553# 0.02fF
C130 a_118_55# a_118_553# 0.15fF
C131 a_n238_553# a_n238_n445# 0.03fF
C132 a_n118_n389# a_n118_607# 0.00fF
C133 a_n830_n887# a_n652_n887# 0.06fF
C134 a_772_109# a_772_n389# 0.00fF
C135 a_n594_n943# a_n594_55# 0.03fF
C136 a_n238_n943# a_n238_n445# 0.15fF
C137 a_474_553# a_n594_553# 0.01fF
C138 a_n652_607# a_60_607# 0.01fF
C139 a_n118_109# a_n830_109# 0.01fF
C140 a_60_607# a_772_607# 0.01fF
C141 a_n594_n943# a_n238_n943# 0.03fF
C142 a_n60_55# a_474_55# 0.02fF
C143 a_n296_n887# a_238_n887# 0.02fF
C144 a_n772_n943# a_n772_n445# 0.15fF
C145 a_n772_n943# a_296_n943# 0.01fF
C146 a_n772_55# a_n238_55# 0.02fF
C147 a_238_109# a_n296_109# 0.02fF
C148 a_n474_607# a_n474_n887# 0.00fF
C149 a_60_109# a_n118_109# 0.06fF
C150 a_n416_55# a_474_55# 0.01fF
C151 a_n60_55# a_n594_55# 0.02fF
C152 a_n652_n887# a_416_n887# 0.01fF
C153 a_n118_n389# a_n118_n887# 0.00fF
C154 a_60_n887# a_60_109# 0.00fF
C155 a_n474_607# a_n118_607# 0.03fF
C156 a_474_55# a_296_55# 0.10fF
C157 a_n772_n943# a_n772_55# 0.03fF
C158 a_n474_607# a_n830_607# 0.03fF
C159 a_n652_n887# a_n474_n887# 0.06fF
C160 a_n830_n887# a_n296_n887# 0.02fF
C161 a_416_607# a_238_607# 0.06fF
C162 a_474_n445# a_474_n943# 0.15fF
C163 a_n652_109# a_416_109# 0.01fF
C164 a_n416_55# a_n594_55# 0.10fF
C165 a_n238_n943# a_n60_n943# 0.10fF
C166 a_118_n445# a_n772_n445# 0.01fF
C167 a_n772_553# a_n772_n445# 0.03fF
C168 a_n238_n943# a_118_n943# 0.03fF
C169 a_n594_55# a_296_55# 0.01fF
C170 a_n772_553# a_n60_553# 0.01fF
C171 a_60_n389# a_416_n389# 0.03fF
C172 a_296_n445# a_n772_n445# 0.01fF
C173 a_594_n389# a_416_n389# 0.06fF
C174 a_n594_553# a_n594_55# 0.15fF
C175 a_594_n389# a_60_n389# 0.02fF
C176 a_n652_109# a_594_109# 0.01fF
C177 a_n474_109# a_n296_109# 0.06fF
C178 a_n652_n389# a_416_n389# 0.01fF
C179 a_296_n445# a_296_n943# 0.15fF
C180 a_n238_553# a_n594_553# 0.03fF
C181 a_n474_109# a_238_109# 0.01fF
C182 a_n238_n445# a_n772_n445# 0.02fF
C183 a_n772_553# a_652_553# 0.01fF
C184 a_474_55# a_474_553# 0.15fF
C185 a_772_n887# a_772_n389# 0.00fF
C186 a_238_n389# a_n830_n389# 0.01fF
C187 a_n652_n389# a_60_n389# 0.01fF
C188 a_n652_n389# a_594_n389# 0.01fF
C189 a_772_109# a_n652_109# 0.01fF
C190 a_60_607# a_60_109# 0.00fF
C191 a_238_n389# a_238_607# 0.00fF
C192 a_n296_n887# a_416_n887# 0.01fF
C193 a_n772_553# a_n772_55# 0.15fF
C194 a_n594_n943# a_296_n943# 0.01fF
C195 a_n416_553# a_n416_n943# 0.01fF
C196 a_n118_607# a_n296_607# 0.06fF
C197 a_474_n943# a_n416_n943# 0.01fF
C198 a_n238_553# a_474_553# 0.01fF
C199 a_n830_607# a_n296_607# 0.02fF
C200 a_n652_n887# a_594_n887# 0.01fF
C201 a_n652_n887# a_n118_n887# 0.02fF
C202 a_n474_n887# a_n296_n887# 0.06fF
C203 a_474_n445# a_n416_n445# 0.01fF
C204 a_n474_607# a_594_607# 0.01fF
C205 a_n416_553# a_296_553# 0.01fF
C206 a_n296_n389# a_n296_109# 0.00fF
C207 a_n830_n887# a_n830_109# 0.00fF
C208 a_n416_553# a_n416_n445# 0.03fF
C209 a_n60_55# a_n60_553# 0.15fF
C210 a_416_n389# a_n474_n389# 0.01fF
C211 a_238_607# a_60_607# 0.06fF
C212 a_n60_553# a_n60_n943# 0.01fF
C213 a_772_n389# a_416_n389# 0.03fF
C214 a_60_n389# a_n474_n389# 0.02fF
C215 a_594_n389# a_n474_n389# 0.01fF
C216 a_296_n943# a_n60_n943# 0.03fF
C217 a_n296_n389# a_416_n389# 0.01fF
C218 a_n118_607# a_772_607# 0.01fF
C219 a_n118_607# a_n652_607# 0.02fF
C220 a_60_n389# a_772_n389# 0.01fF
C221 a_474_55# a_n594_55# 0.01fF
C222 a_594_n389# a_772_n389# 0.06fF
C223 a_n296_n389# a_60_n389# 0.03fF
C224 a_n652_n389# a_n474_n389# 0.06fF
C225 a_474_n943# a_652_n943# 0.10fF
C226 a_118_n943# a_296_n943# 0.10fF
C227 a_594_n389# a_n296_n389# 0.01fF
C228 a_n830_607# a_772_607# 0.01fF
C229 a_n652_607# a_n830_607# 0.06fF
C230 a_n652_n389# a_772_n389# 0.01fF
C231 a_118_553# a_118_n445# 0.03fF
C232 a_n652_n389# a_n296_n389# 0.03fF
C233 a_n772_553# a_118_553# 0.01fF
C234 a_416_607# a_60_607# 0.03fF
C235 a_n416_n943# a_n416_n445# 0.15fF
C236 a_n60_55# a_n772_55# 0.01fF
C237 a_n474_109# a_n474_n389# 0.00fF
C238 a_n296_n887# a_594_n887# 0.01fF
C239 a_652_n445# a_n772_n445# 0.01fF
C240 a_n296_n887# a_n118_n887# 0.06fF
C241 a_238_n887# a_238_607# 0.00fF
C242 a_296_n943# a_296_55# 0.03fF
C243 a_594_607# a_n296_607# 0.01fF
C244 a_n60_553# a_n594_553# 0.02fF
C245 a_n118_n389# a_416_n389# 0.02fF
C246 a_474_n445# a_n594_n445# 0.01fF
C247 a_652_n943# a_n416_n943# 0.01fF
C248 a_n118_n389# a_60_n389# 0.06fF
C249 a_652_n445# a_652_553# 0.03fF
C250 a_652_553# a_n594_553# 0.01fF
C251 a_n118_n389# a_594_n389# 0.01fF
C252 a_n652_n887# a_772_n887# 0.01fF
C253 a_n416_55# a_n772_55# 0.03fF
C254 a_n118_n389# a_n652_n389# 0.02fF
C255 a_772_109# a_772_607# 0.00fF
C256 a_n60_n445# a_474_n445# 0.02fF
C257 a_n238_n943# a_n238_553# 0.01fF
C258 a_n830_n887# a_n830_n389# 0.00fF
C259 a_n772_55# a_296_55# 0.01fF
C260 a_n60_553# a_474_553# 0.02fF
C261 a_60_n887# a_60_607# 0.00fF
C262 a_n830_607# a_n830_109# 0.00fF
C263 a_416_109# a_n830_109# 0.01fF
C264 a_652_553# a_474_553# 0.10fF
C265 a_n652_109# a_n296_109# 0.03fF
C266 a_594_607# a_772_607# 0.06fF
C267 a_n652_109# a_238_109# 0.01fF
C268 a_n652_607# a_594_607# 0.01fF
C269 a_772_n389# a_n474_n389# 0.01fF
C270 a_n296_n389# a_n474_n389# 0.06fF
C271 a_n296_n389# a_772_n389# 0.01fF
C272 a_238_n389# a_238_n887# 0.00fF
C273 a_n830_109# a_594_109# 0.01fF
C274 a_60_109# a_416_109# 0.03fF
C275 a_60_n887# a_238_n887# 0.06fF
C276 a_118_n943# a_118_553# 0.01fF
C277 a_772_109# a_n830_109# 0.01fF
C278 a_n652_n389# a_n652_109# 0.00fF
C279 a_n296_n887# a_772_n887# 0.01fF
C280 a_n118_n389# a_n474_n389# 0.03fF
C281 a_60_109# a_594_109# 0.02fF
C282 a_n118_n389# a_772_n389# 0.01fF
C283 a_n416_n445# a_n594_n445# 0.10fF
C284 a_n474_109# a_n652_109# 0.06fF
C285 a_n118_n389# a_n296_n389# 0.06fF
C286 a_n474_109# a_n474_607# 0.00fF
C287 a_652_n943# a_652_55# 0.03fF
C288 a_772_109# a_60_109# 0.01fF
C289 a_118_553# a_n594_553# 0.01fF
C290 a_n652_n389# a_n652_n887# 0.00fF
C291 a_416_607# a_416_n887# 0.00fF
C292 a_118_55# a_652_55# 0.02fF
C293 a_n830_n887# a_60_n887# 0.01fF
C294 a_n60_n445# a_n416_n445# 0.03fF
C295 a_772_n887# a_772_607# 0.00fF
C296 a_n830_n389# a_n830_607# 0.00fF
C297 a_n296_109# a_n296_607# 0.00fF
C298 a_n118_607# a_238_607# 0.03fF
C299 a_n60_553# a_n238_553# 0.10fF
C300 a_n772_55# a_474_55# 0.01fF
C301 a_238_607# a_n830_607# 0.01fF
C302 a_n772_n943# a_474_n943# 0.01fF
C303 a_652_553# a_n238_553# 0.01fF
C304 a_n238_n943# a_296_n943# 0.02fF
C305 a_474_553# a_118_553# 0.03fF
C306 a_n296_n887# a_n296_109# 0.00fF
C307 a_416_607# a_n118_607# 0.02fF
C308 a_n772_55# a_n594_55# 0.10fF
C309 a_416_607# a_n830_607# 0.01fF
C310 a_416_607# a_416_109# 0.00fF
C311 a_n474_607# a_n474_n389# 0.00fF
C312 a_60_n887# a_416_n887# 0.03fF
C313 a_474_n445# a_118_n445# 0.03fF
C314 a_n772_n943# a_n416_n943# 0.03fF
C315 a_474_n445# a_296_n445# 0.10fF
C316 a_474_n445# a_n238_n445# 0.01fF
C317 a_n474_n887# a_60_n887# 0.02fF
C318 a_n118_607# a_n118_109# 0.00fF
C319 a_n772_553# a_n416_553# 0.03fF
C320 a_n60_n445# a_n594_n445# 0.02fF
C321 a_416_109# a_n118_109# 0.02fF
C322 a_238_607# a_594_607# 0.03fF
C323 a_n830_n887# a_238_n887# 0.01fF
C324 a_n652_n389# a_n652_607# 0.00fF
C325 a_118_55# a_n238_55# 0.03fF
C326 a_n118_109# a_594_109# 0.01fF
C327 a_n594_n943# a_474_n943# 0.01fF
C328 a_n772_n943# a_652_n943# 0.01fF
C329 a_416_607# a_594_607# 0.06fF
C330 a_n238_553# a_118_553# 0.03fF
C331 a_772_109# a_n118_109# 0.01fF
C332 a_n296_109# a_n830_109# 0.02fF
C333 a_238_109# a_n830_109# 0.01fF
C334 a_n296_n389# a_n296_607# 0.00fF
C335 a_n238_55# a_652_55# 0.01fF
C336 a_n118_n887# a_n118_109# 0.00fF
C337 a_n118_607# a_60_607# 0.06fF
C338 a_n60_553# a_652_553# 0.01fF
C339 a_60_n887# a_594_n887# 0.02fF
C340 a_238_n887# a_416_n887# 0.06fF
C341 a_n118_n887# a_60_n887# 0.06fF
C342 a_n772_553# a_296_553# 0.01fF
C343 a_n830_607# a_60_607# 0.01fF
C344 a_n594_n943# a_n416_n943# 0.10fF
C345 a_n416_n445# a_118_n445# 0.02fF
C346 a_n296_n389# a_n296_n887# 0.00fF
C347 a_60_109# a_n296_109# 0.03fF
C348 a_296_n445# a_296_553# 0.03fF
C349 a_60_109# a_238_109# 0.06fF
C350 a_296_n445# a_n416_n445# 0.01fF
C351 a_n772_55# a_n772_n445# 0.15fF
C352 a_n474_n887# a_238_n887# 0.01fF
C353 a_n416_n445# a_n238_n445# 0.10fF
C354 a_474_n943# a_n60_n943# 0.02fF
C355 a_60_n389# a_60_109# 0.00fF
C356 a_n474_109# a_n830_109# 0.03fF
C357 a_772_n389# a_772_607# 0.00fF
C358 a_652_n445# a_474_n445# 0.10fF
C359 a_118_n943# a_474_n943# 0.03fF
C360 a_118_55# a_118_n445# 0.15fF
C361 a_n652_n887# a_n652_109# 0.00fF
C362 a_n830_n887# a_416_n887# 0.01fF
C363 a_n416_553# a_n416_55# 0.15fF
C364 a_n416_n943# a_n60_n943# 0.03fF
C365 a_n474_109# a_60_109# 0.02fF
C366 a_n416_553# a_n594_553# 0.10fF
C367 a_n830_n887# a_n474_n887# 0.03fF
C368 a_n594_n943# a_652_n943# 0.01fF
C369 a_118_n943# a_n416_n943# 0.02fF
C370 a_474_n445# a_474_553# 0.03fF
C371 a_238_607# a_238_109# 0.00fF
C372 a_60_607# a_594_607# 0.02fF
C373 a_n416_n943# a_n416_55# 0.03fF
C374 a_n830_n389# a_416_n389# 0.01fF
C375 a_n594_n445# a_118_n445# 0.01fF
C376 a_n830_n887# a_n830_607# 0.00fF
C377 a_n830_n389# a_60_n389# 0.01fF
C378 a_n474_607# a_n296_607# 0.06fF
C379 a_594_n389# a_n830_n389# 0.01fF
C380 a_60_n887# a_772_n887# 0.01fF
C381 a_238_n887# a_594_n887# 0.03fF
C382 a_n118_n887# a_238_n887# 0.03fF
C383 a_296_n445# a_n594_n445# 0.01fF
C384 a_n60_553# a_118_553# 0.10fF
C385 a_n416_553# a_474_553# 0.01fF
C386 a_n652_n389# a_n830_n389# 0.06fF
C387 a_n60_n445# a_118_n445# 0.10fF
C388 a_474_n943# a_474_553# 0.01fF
C389 a_n594_n445# a_n238_n445# 0.03fF
C390 a_652_553# a_118_553# 0.02fF
C391 a_n60_n445# a_296_n445# 0.03fF
C392 a_n474_n887# a_416_n887# 0.01fF
C393 a_n60_n445# a_n238_n445# 0.10fF
C394 a_n416_55# a_n416_n445# 0.15fF
C395 a_416_607# a_416_n389# 0.00fF
C396 a_652_n943# a_n60_n943# 0.01fF
C397 a_n60_55# a_118_55# 0.10fF
C398 a_n594_n943# a_n594_n445# 0.15fF
C399 a_296_55# a_296_553# 0.15fF
C400 a_118_n943# a_652_n943# 0.02fF
C401 a_n594_553# a_296_553# 0.01fF
C402 a_474_n445# a_474_55# 0.15fF
C403 a_n830_n887# a_594_n887# 0.01fF
C404 a_n652_n887# a_n296_n887# 0.03fF
C405 a_n830_n887# a_n118_n887# 0.01fF
C406 a_652_n445# a_n416_n445# 0.01fF
C407 a_118_n943# a_118_55# 0.03fF
C408 a_416_n887# a_416_109# 0.00fF
C409 a_n652_607# a_n652_109# 0.00fF
C410 a_n296_109# a_n118_109# 0.06fF
C411 a_238_109# a_n118_109# 0.03fF
C412 a_n474_607# a_772_607# 0.01fF
C413 a_n474_607# a_n652_607# 0.06fF
C414 a_238_n389# a_238_109# 0.00fF
C415 a_n416_55# a_118_55# 0.02fF
C416 a_n60_55# a_652_55# 0.01fF
C417 a_652_n445# a_652_n943# 0.15fF
C418 a_474_n943# a_474_55# 0.03fF
C419 a_118_55# a_296_55# 0.10fF
C420 a_238_n389# a_416_n389# 0.06fF
C421 a_474_553# a_296_553# 0.10fF
C422 a_n652_n887# a_n652_607# 0.00fF
C423 a_n118_607# a_n830_607# 0.01fF
C424 a_238_n389# a_60_n389# 0.06fF
C425 a_238_n389# a_594_n389# 0.03fF
C426 a_60_n887# a_60_n389# 0.00fF
C427 a_n830_n389# a_n474_n389# 0.03fF
C428 a_n416_55# a_652_55# 0.01fF
C429 a_n652_n389# a_238_n389# 0.01fF
C430 a_n830_n389# a_772_n389# 0.01fF
C431 a_416_n887# a_594_n887# 0.06fF
C432 a_n296_n389# a_n830_n389# 0.02fF
C433 a_n296_n887# a_n296_607# 0.00fF
C434 a_238_n887# a_772_n887# 0.02fF
C435 a_n60_n445# a_n60_55# 0.15fF
C436 a_n118_n887# a_416_n887# 0.02fF
C437 a_n238_55# a_n238_n445# 0.15fF
C438 a_772_n887# a_n1110_n1061# 0.10fF
C439 a_594_n887# a_n1110_n1061# 0.06fF
C440 a_416_n887# a_n1110_n1061# 0.05fF
C441 a_238_n887# a_n1110_n1061# 0.05fF
C442 a_60_n887# a_n1110_n1061# 0.04fF
C443 a_n118_n887# a_n1110_n1061# 0.04fF
C444 a_n296_n887# a_n1110_n1061# 0.05fF
C445 a_n474_n887# a_n1110_n1061# 0.05fF
C446 a_n652_n887# a_n1110_n1061# 0.06fF
C447 a_n830_n887# a_n1110_n1061# 0.10fF
C448 a_652_n943# a_n1110_n1061# 0.27fF
C449 a_474_n943# a_n1110_n1061# 0.24fF
C450 a_296_n943# a_n1110_n1061# 0.24fF
C451 a_118_n943# a_n1110_n1061# 0.24fF
C452 a_n60_n943# a_n1110_n1061# 0.25fF
C453 a_n238_n943# a_n1110_n1061# 0.26fF
C454 a_n416_n943# a_n1110_n1061# 0.26fF
C455 a_n594_n943# a_n1110_n1061# 0.27fF
C456 a_n772_n943# a_n1110_n1061# 0.32fF
C457 a_772_n389# a_n1110_n1061# 0.10fF
C458 a_594_n389# a_n1110_n1061# 0.06fF
C459 a_416_n389# a_n1110_n1061# 0.05fF
C460 a_238_n389# a_n1110_n1061# 0.04fF
C461 a_60_n389# a_n1110_n1061# 0.04fF
C462 a_n118_n389# a_n1110_n1061# 0.04fF
C463 a_n296_n389# a_n1110_n1061# 0.04fF
C464 a_n474_n389# a_n1110_n1061# 0.05fF
C465 a_n652_n389# a_n1110_n1061# 0.06fF
C466 a_n830_n389# a_n1110_n1061# 0.10fF
C467 a_652_n445# a_n1110_n1061# 0.22fF
C468 a_474_n445# a_n1110_n1061# 0.19fF
C469 a_296_n445# a_n1110_n1061# 0.19fF
C470 a_118_n445# a_n1110_n1061# 0.19fF
C471 a_n60_n445# a_n1110_n1061# 0.20fF
C472 a_n238_n445# a_n1110_n1061# 0.21fF
C473 a_n416_n445# a_n1110_n1061# 0.21fF
C474 a_n594_n445# a_n1110_n1061# 0.22fF
C475 a_n772_n445# a_n1110_n1061# 0.27fF
C476 a_772_109# a_n1110_n1061# 0.10fF
C477 a_594_109# a_n1110_n1061# 0.06fF
C478 a_416_109# a_n1110_n1061# 0.05fF
C479 a_238_109# a_n1110_n1061# 0.05fF
C480 a_60_109# a_n1110_n1061# 0.04fF
C481 a_n118_109# a_n1110_n1061# 0.04fF
C482 a_n296_109# a_n1110_n1061# 0.05fF
C483 a_n474_109# a_n1110_n1061# 0.05fF
C484 a_n652_109# a_n1110_n1061# 0.06fF
C485 a_n830_109# a_n1110_n1061# 0.10fF
C486 a_652_55# a_n1110_n1061# 0.23fF
C487 a_474_55# a_n1110_n1061# 0.20fF
C488 a_296_55# a_n1110_n1061# 0.20fF
C489 a_118_55# a_n1110_n1061# 0.21fF
C490 a_n60_55# a_n1110_n1061# 0.21fF
C491 a_n238_55# a_n1110_n1061# 0.22fF
C492 a_n416_55# a_n1110_n1061# 0.23fF
C493 a_n594_55# a_n1110_n1061# 0.24fF
C494 a_n772_55# a_n1110_n1061# 0.28fF
C495 a_772_607# a_n1110_n1061# 0.10fF
C496 a_594_607# a_n1110_n1061# 0.06fF
C497 a_416_607# a_n1110_n1061# 0.06fF
C498 a_238_607# a_n1110_n1061# 0.05fF
C499 a_60_607# a_n1110_n1061# 0.05fF
C500 a_n118_607# a_n1110_n1061# 0.05fF
C501 a_n296_607# a_n1110_n1061# 0.05fF
C502 a_n474_607# a_n1110_n1061# 0.06fF
C503 a_n652_607# a_n1110_n1061# 0.07fF
C504 a_n830_607# a_n1110_n1061# 0.10fF
C505 a_652_553# a_n1110_n1061# 0.30fF
C506 a_474_553# a_n1110_n1061# 0.27fF
C507 a_296_553# a_n1110_n1061# 0.27fF
C508 a_118_553# a_n1110_n1061# 0.27fF
C509 a_n60_553# a_n1110_n1061# 0.28fF
C510 a_n238_553# a_n1110_n1061# 0.29fF
C511 a_n416_553# a_n1110_n1061# 0.29fF
C512 a_n594_553# a_n1110_n1061# 0.30fF
C513 a_n772_553# a_n1110_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_JJWXCM a_n207_n140# a_29_n205# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n205# a_563_n205# a_n741_n140# a_n327_n205# a_n563_n140# a_385_n205#
+ w_n777_n241# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n327_n205# a_n385_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_563_n205# a_563_n205# a_505_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n29_n140# a_n149_n205# a_n207_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_505_n140# a_385_n205# a_327_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n207_n140# a_n563_n140# 0.06fF
C1 a_n741_n140# a_327_n140# 0.01fF
C2 a_505_n140# a_n563_n140# 0.02fF
C3 w_n777_n241# a_207_n205# 0.15fF
C4 a_n29_n140# a_149_n140# 0.13fF
C5 a_29_n205# a_n741_n140# 0.01fF
C6 a_n29_n140# a_563_n205# 0.01fF
C7 a_327_n140# a_n385_n140# 0.03fF
C8 a_n149_n205# a_385_n205# 0.02fF
C9 a_n327_n205# a_385_n205# 0.01fF
C10 a_n327_n205# a_n149_n205# 0.10fF
C11 w_n777_n241# a_327_n140# 0.02fF
C12 a_n207_n140# a_327_n140# 0.04fF
C13 a_327_n140# a_505_n140# 0.13fF
C14 a_29_n205# w_n777_n241# 0.16fF
C15 a_n29_n140# a_n563_n140# 0.04fF
C16 a_n741_n140# a_385_n205# 0.01fF
C17 a_n741_n140# a_n149_n205# 0.01fF
C18 a_n741_n140# a_n327_n205# 0.02fF
C19 a_563_n205# a_149_n140# 0.02fF
C20 w_n777_n241# a_385_n205# 0.14fF
C21 w_n777_n241# a_n149_n205# 0.17fF
C22 a_n327_n205# w_n777_n241# 0.18fF
C23 a_n29_n140# a_327_n140# 0.06fF
C24 a_n505_n205# a_563_n205# 0.01fF
C25 a_n741_n140# a_n385_n140# 0.03fF
C26 a_n563_n140# a_149_n140# 0.03fF
C27 a_n741_n140# w_n777_n241# 0.33fF
C28 a_563_n205# a_n563_n140# 0.01fF
C29 a_n207_n140# a_n741_n140# 0.02fF
C30 a_n741_n140# a_505_n140# 0.01fF
C31 w_n777_n241# a_n385_n140# 0.02fF
C32 a_207_n205# a_563_n205# 0.02fF
C33 a_n207_n140# a_n385_n140# 0.13fF
C34 a_505_n140# a_n385_n140# 0.02fF
C35 a_327_n140# a_149_n140# 0.13fF
C36 a_n207_n140# w_n777_n241# 0.02fF
C37 w_n777_n241# a_505_n140# 0.02fF
C38 a_327_n140# a_563_n205# 0.03fF
C39 a_n505_n205# a_207_n205# 0.01fF
C40 a_n207_n140# a_505_n140# 0.03fF
C41 a_29_n205# a_563_n205# 0.01fF
C42 a_n741_n140# a_n29_n140# 0.01fF
C43 a_29_n205# a_n505_n205# 0.02fF
C44 a_n29_n140# a_n385_n140# 0.06fF
C45 a_327_n140# a_n563_n140# 0.02fF
C46 w_n777_n241# a_n29_n140# 0.02fF
C47 a_563_n205# a_385_n205# 0.07fF
C48 a_563_n205# a_n149_n205# 0.01fF
C49 a_n207_n140# a_n29_n140# 0.13fF
C50 a_n29_n140# a_505_n140# 0.04fF
C51 a_n327_n205# a_563_n205# 0.01fF
C52 a_29_n205# a_207_n205# 0.10fF
C53 a_n505_n205# a_385_n205# 0.01fF
C54 a_n505_n205# a_n149_n205# 0.03fF
C55 a_n505_n205# a_n327_n205# 0.10fF
C56 a_n741_n140# a_149_n140# 0.01fF
C57 a_n741_n140# a_563_n205# 0.01fF
C58 a_n385_n140# a_149_n140# 0.04fF
C59 a_207_n205# a_385_n205# 0.10fF
C60 a_207_n205# a_n149_n205# 0.03fF
C61 a_563_n205# a_n385_n140# 0.01fF
C62 w_n777_n241# a_149_n140# 0.02fF
C63 a_n327_n205# a_207_n205# 0.02fF
C64 a_n207_n140# a_149_n140# 0.06fF
C65 a_n741_n140# a_n505_n205# 0.07fF
C66 w_n777_n241# a_563_n205# 0.28fF
C67 a_505_n140# a_149_n140# 0.06fF
C68 a_n207_n140# a_563_n205# 0.01fF
C69 a_505_n140# a_563_n205# 0.06fF
C70 a_29_n205# a_385_n205# 0.03fF
C71 a_29_n205# a_n149_n205# 0.10fF
C72 a_n505_n205# w_n777_n241# 0.19fF
C73 a_n741_n140# a_n563_n140# 0.06fF
C74 a_29_n205# a_n327_n205# 0.03fF
C75 a_n741_n140# a_207_n205# 0.01fF
C76 a_n385_n140# a_n563_n140# 0.13fF
C77 w_n777_n241# a_n563_n140# 0.02fF
C78 w_n777_n241# VSUBS 2.25fF
.ends

.subckt sky130_fd_pr__nfet_01v8_LJREPQ a_n149_n195# a_n207_n140# a_207_n195# a_n29_n140#
+ a_149_n140# a_29_n195# a_n385_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_207_n195# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n385_n140# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n149_n195# a_29_n195# 0.10fF
C1 a_207_n195# a_29_n195# 0.06fF
C2 a_n385_n140# a_n207_n140# 0.06fF
C3 a_n149_n195# a_207_n195# 0.02fF
C4 a_n29_n140# a_n385_n140# 0.03fF
C5 a_n385_n140# a_149_n140# 0.02fF
C6 a_207_n195# a_n207_n140# 0.02fF
C7 a_207_n195# a_n29_n140# 0.03fF
C8 a_207_n195# a_149_n140# 0.06fF
C9 a_n29_n140# a_n207_n140# 0.06fF
C10 a_n385_n140# a_29_n195# 0.02fF
C11 a_149_n140# a_n207_n140# 0.03fF
C12 a_n149_n195# a_n385_n140# 0.06fF
C13 a_207_n195# a_n385_n140# 0.03fF
C14 a_n29_n140# a_149_n140# 0.06fF
C15 a_149_n140# VSUBS 0.01fF
C16 a_n29_n140# VSUBS 0.01fF
C17 a_n207_n140# VSUBS 0.02fF
C18 a_207_n195# VSUBS 0.31fF
C19 a_29_n195# VSUBS 0.19fF
C20 a_n149_n195# VSUBS 0.20fF
C21 a_n385_n140# VSUBS 0.33fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SAWXCM a_n207_n140# a_29_n205# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n205# a_563_n205# a_n741_n140# a_n327_n205# a_n563_n140# a_385_n205#
+ w_n777_n241# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# VSUBS
X0 a_505_n140# a_385_n205# a_327_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n385_n140# a_n505_n205# a_n563_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_327_n140# a_207_n205# a_149_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_149_n140# a_29_n205# a_n29_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n205# a_n385_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_563_n205# a_563_n205# a_505_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n29_n140# a_n149_n205# a_n207_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 w_n777_n241# a_n29_n140# 0.02fF
C1 a_149_n140# a_n29_n140# 0.13fF
C2 a_n505_n205# a_563_n205# 0.01fF
C3 a_207_n205# a_n149_n205# 0.03fF
C4 a_n29_n140# a_n563_n140# 0.04fF
C5 a_n207_n140# a_n741_n140# 0.02fF
C6 a_n741_n140# a_385_n205# 0.01fF
C7 a_29_n205# a_n741_n140# 0.01fF
C8 a_149_n140# a_n207_n140# 0.06fF
C9 w_n777_n241# a_n207_n140# 0.02fF
C10 w_n777_n241# a_385_n205# 0.14fF
C11 w_n777_n241# a_29_n205# 0.16fF
C12 a_n327_n205# a_563_n205# 0.01fF
C13 a_n741_n140# a_n149_n205# 0.01fF
C14 a_n207_n140# a_n563_n140# 0.06fF
C15 a_505_n140# a_327_n140# 0.13fF
C16 a_n741_n140# a_n385_n140# 0.03fF
C17 w_n777_n241# a_n149_n205# 0.17fF
C18 a_505_n140# a_563_n205# 0.06fF
C19 a_149_n140# a_n385_n140# 0.04fF
C20 w_n777_n241# a_n385_n140# 0.02fF
C21 a_385_n205# a_n505_n205# 0.01fF
C22 a_207_n205# a_n741_n140# 0.01fF
C23 a_29_n205# a_n505_n205# 0.02fF
C24 w_n777_n241# a_207_n205# 0.15fF
C25 a_n385_n140# a_n563_n140# 0.13fF
C26 a_n505_n205# a_n149_n205# 0.03fF
C27 a_505_n140# a_n29_n140# 0.04fF
C28 a_563_n205# a_327_n140# 0.03fF
C29 a_207_n205# a_n505_n205# 0.01fF
C30 a_n327_n205# a_385_n205# 0.01fF
C31 a_29_n205# a_n327_n205# 0.03fF
C32 w_n777_n241# a_n741_n140# 0.33fF
C33 a_149_n140# a_n741_n140# 0.01fF
C34 a_505_n140# a_n207_n140# 0.03fF
C35 w_n777_n241# a_149_n140# 0.02fF
C36 a_n29_n140# a_327_n140# 0.06fF
C37 a_n327_n205# a_n149_n205# 0.10fF
C38 a_n29_n140# a_563_n205# 0.01fF
C39 a_n741_n140# a_n563_n140# 0.06fF
C40 a_149_n140# a_n563_n140# 0.03fF
C41 w_n777_n241# a_n563_n140# 0.02fF
C42 a_n741_n140# a_n505_n205# 0.07fF
C43 a_n327_n205# a_207_n205# 0.02fF
C44 a_505_n140# a_n385_n140# 0.02fF
C45 w_n777_n241# a_n505_n205# 0.19fF
C46 a_n207_n140# a_327_n140# 0.04fF
C47 a_n207_n140# a_563_n205# 0.01fF
C48 a_385_n205# a_563_n205# 0.07fF
C49 a_29_n205# a_563_n205# 0.01fF
C50 a_n385_n140# a_327_n140# 0.03fF
C51 a_563_n205# a_n149_n205# 0.01fF
C52 a_n327_n205# a_n741_n140# 0.02fF
C53 a_n207_n140# a_n29_n140# 0.13fF
C54 a_563_n205# a_n385_n140# 0.01fF
C55 w_n777_n241# a_n327_n205# 0.18fF
C56 a_505_n140# a_n741_n140# 0.01fF
C57 a_207_n205# a_563_n205# 0.02fF
C58 w_n777_n241# a_505_n140# 0.02fF
C59 a_505_n140# a_149_n140# 0.06fF
C60 a_n29_n140# a_n385_n140# 0.06fF
C61 a_n327_n205# a_n505_n205# 0.10fF
C62 a_505_n140# a_n563_n140# 0.02fF
C63 a_29_n205# a_385_n205# 0.03fF
C64 a_n741_n140# a_327_n140# 0.01fF
C65 a_149_n140# a_327_n140# 0.13fF
C66 w_n777_n241# a_327_n140# 0.02fF
C67 a_n741_n140# a_563_n205# 0.01fF
C68 a_385_n205# a_n149_n205# 0.02fF
C69 a_29_n205# a_n149_n205# 0.10fF
C70 a_n207_n140# a_n385_n140# 0.13fF
C71 w_n777_n241# a_563_n205# 0.28fF
C72 a_149_n140# a_563_n205# 0.02fF
C73 a_327_n140# a_n563_n140# 0.02fF
C74 a_207_n205# a_385_n205# 0.10fF
C75 a_29_n205# a_207_n205# 0.10fF
C76 a_563_n205# a_n563_n140# 0.01fF
C77 a_n741_n140# a_n29_n140# 0.01fF
C78 w_n777_n241# VSUBS 2.25fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_28TRYY a_385_553# a_n1097_109# a_n149_55# a_919_n445#
+ a_29_55# a_n29_n389# a_n207_n887# a_1097_n943# a_n1555_n1061# a_n1097_n389# a_n327_n445#
+ a_149_n389# a_n207_109# a_385_n445# a_563_55# a_n505_n943# a_n1275_n887# a_327_n887#
+ a_505_109# a_563_n943# a_n505_553# a_n741_n389# a_327_109# a_n327_553# a_n1275_607#
+ a_n1217_55# a_861_n389# a_149_109# a_n149_553# a_n1097_607# a_385_55# a_n149_n445#
+ a_n29_109# a_919_n943# a_n29_n887# a_n327_n943# a_n1097_n887# a_149_n887# a_n207_607#
+ a_207_n445# a_385_n943# a_n563_n389# a_1097_553# a_n1039_55# a_1217_n389# a_207_55#
+ a_n1217_n445# a_505_607# a_n741_n887# a_327_607# a_n861_n445# a_683_n389# a_n861_55#
+ a_149_607# a_861_n887# a_n919_n389# a_207_553# a_n741_109# a_n919_109# a_n29_607#
+ a_n149_n943# a_1217_109# a_n563_109# a_919_55# a_n1217_553# a_n385_n389# a_1039_109#
+ a_1039_n389# a_861_109# a_n1039_n445# a_n385_109# a_207_n943# a_n861_553# a_n683_55#
+ a_n563_n887# a_n1039_553# a_29_n445# a_1217_n887# a_683_109# a_n683_n445# a_n1217_n943#
+ a_n683_553# a_29_553# a_505_n389# a_n861_n943# a_683_n887# a_741_n445# a_n505_55#
+ a_n919_n887# a_n741_607# a_n919_607# a_1217_607# a_n563_607# a_1097_55# a_1097_n445#
+ a_n207_n389# a_n385_n887# a_1039_607# a_1039_n887# a_861_607# a_n1039_n943# a_n385_607#
+ a_29_n943# a_n327_55# a_n1275_n389# a_683_607# a_n505_n445# a_327_n389# a_n683_n943#
+ a_919_553# a_741_553# a_563_n445# a_505_n887# a_563_553# a_741_n943# a_741_55# a_n1275_109#
X0 a_n919_607# a_n1039_553# a_n1097_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1039_607# a_919_553# a_861_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_109# a_29_55# a_n29_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1097_n887# a_n1217_n943# a_n1275_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_683_n887# a_563_n943# a_505_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n207_n389# a_n327_n445# a_n385_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_607# a_n327_553# a_n385_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n1275_109# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=3.248e+12p ps=2.704e+07u w=1.4e+06u l=600000u
X8 a_683_109# a_563_55# a_505_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_1217_n389# a_1097_n445# a_1039_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1275_n389# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n563_109# a_n683_55# a_n741_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1555_n1061# a_n1555_n1061# a_1217_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_n741_n389# a_n861_n445# a_n919_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n29_n887# a_n149_n943# a_n207_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n919_109# a_n1039_55# a_n1097_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_327_109# a_207_55# a_149_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1039_109# a_919_55# a_861_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1097_n389# a_n1217_n445# a_n1275_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_683_n389# a_563_n445# a_505_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_1039_n389# a_919_n445# a_861_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_505_607# a_385_553# a_327_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n207_109# a_n327_55# a_n385_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_n563_n887# a_n683_n943# a_n741_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_1217_607# a_1097_553# a_1039_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n919_n887# a_n1039_n943# a_n1097_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_505_n887# a_385_n943# a_327_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_861_607# a_741_553# a_683_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_n29_n389# a_n149_n445# a_n207_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n385_n887# a_n505_n943# a_n563_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n741_607# a_n861_553# a_n919_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_n1555_n1061# a_n1555_n1061# a_1217_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X32 a_n29_607# a_n149_553# a_n207_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_505_109# a_385_55# a_327_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_327_n887# a_207_n943# a_149_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X35 a_n563_n389# a_n683_n445# a_n741_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_149_n887# a_29_n943# a_n29_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_n1097_607# a_n1217_553# a_n1275_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X38 a_1217_109# a_1097_55# a_1039_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n919_n389# a_n1039_n445# a_n1097_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_505_n389# a_385_n445# a_327_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X41 a_n385_607# a_n505_553# a_n563_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X42 a_861_109# a_741_55# a_683_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_861_n887# a_741_n943# a_683_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X44 a_n385_n389# a_n505_n445# a_n563_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X45 a_n741_109# a_n861_55# a_n919_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X46 a_n1555_n1061# a_n1555_n1061# a_1217_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X47 a_n29_109# a_n149_55# a_n207_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X48 a_327_n389# a_207_n445# a_149_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X49 a_149_n389# a_29_n445# a_n29_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X50 a_149_607# a_29_553# a_n29_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X51 a_n1097_109# a_n1217_55# a_n1275_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X52 a_n207_n887# a_n327_n943# a_n385_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X53 a_n1275_607# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X54 a_683_607# a_563_553# a_505_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X55 a_n385_109# a_n505_55# a_n563_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X56 a_861_n389# a_741_n445# a_683_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X57 a_1217_n887# a_1097_n943# a_1039_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X58 a_n1275_n887# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X59 a_n563_607# a_n683_553# a_n741_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X60 a_n1555_n1061# a_n1555_n1061# a_1217_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X61 a_n741_n887# a_n861_n943# a_n919_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X62 a_327_607# a_207_553# a_149_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X63 a_1039_n887# a_919_n943# a_861_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_149_n389# a_683_n389# 0.02fF
C1 a_n683_n445# a_n683_n943# 0.15fF
C2 a_1039_607# a_1217_607# 0.06fF
C3 a_385_55# a_385_n943# 0.03fF
C4 a_n505_553# a_n149_553# 0.03fF
C5 a_741_55# a_741_n445# 0.15fF
C6 a_n29_109# a_n1097_109# 0.01fF
C7 a_n207_n887# a_327_n887# 0.02fF
C8 a_n741_n887# a_861_n887# 0.01fF
C9 a_n29_n887# a_149_n887# 0.06fF
C10 a_n385_n887# a_505_n887# 0.01fF
C11 a_n563_n887# a_683_n887# 0.01fF
C12 a_207_55# a_207_553# 0.15fF
C13 a_n1217_553# a_n149_553# 0.01fF
C14 a_385_55# a_n683_55# 0.01fF
C15 a_149_n389# a_505_n389# 0.03fF
C16 a_n683_553# a_n861_553# 0.10fF
C17 a_385_55# a_1097_55# 0.01fF
C18 a_n29_109# a_n563_109# 0.02fF
C19 a_n563_n887# a_505_n887# 0.01fF
C20 a_n385_n887# a_327_n887# 0.01fF
C21 a_n741_n887# a_683_n887# 0.01fF
C22 a_n207_n887# a_149_n887# 0.03fF
C23 a_n741_n389# a_n741_109# 0.00fF
C24 a_741_n445# a_n683_n445# 0.01fF
C25 a_n327_55# a_29_55# 0.03fF
C26 a_n741_n389# a_n919_n389# 0.06fF
C27 a_n861_n445# a_n149_n445# 0.01fF
C28 a_n207_n389# a_n207_n887# 0.00fF
C29 a_n1097_109# a_n1275_109# 0.06fF
C30 a_n505_553# a_385_553# 0.01fF
C31 a_n385_n887# a_149_n887# 0.02fF
C32 a_n207_n887# a_n29_n887# 0.06fF
C33 a_n919_n887# a_683_n887# 0.01fF
C34 a_327_109# a_327_n389# 0.00fF
C35 a_207_n445# a_n1217_n445# 0.01fF
C36 a_919_n445# a_1097_n445# 0.10fF
C37 a_n563_n887# a_327_n887# 0.01fF
C38 a_n1097_n389# a_149_n389# 0.01fF
C39 a_n741_n887# a_505_n887# 0.01fF
C40 a_n29_109# a_1039_109# 0.01fF
C41 a_n1097_607# a_327_607# 0.01fF
C42 a_n683_n445# a_n327_n445# 0.03fF
C43 a_385_553# a_n1217_553# 0.01fF
C44 a_n683_553# a_29_553# 0.01fF
C45 a_n1039_553# a_n327_553# 0.01fF
C46 a_n505_n445# a_919_n445# 0.01fF
C47 a_29_n445# a_741_n445# 0.01fF
C48 a_n563_109# a_n1275_109# 0.01fF
C49 a_n919_607# a_n385_607# 0.02fF
C50 a_n327_55# a_n1039_55# 0.01fF
C51 a_327_n389# a_1217_n389# 0.01fF
C52 a_563_553# a_563_n943# 0.01fF
C53 a_n385_109# a_683_109# 0.01fF
C54 a_n385_n887# a_n29_n887# 0.03fF
C55 a_n563_n887# a_149_n887# 0.01fF
C56 a_n741_n887# a_327_n887# 0.01fF
C57 a_n919_n887# a_505_n887# 0.01fF
C58 a_741_553# a_207_553# 0.02fF
C59 a_207_55# a_919_55# 0.01fF
C60 a_1039_607# a_1039_n389# 0.00fF
C61 a_683_109# a_1217_109# 0.02fF
C62 a_n1039_n445# a_n1039_n943# 0.15fF
C63 a_149_607# a_n29_607# 0.06fF
C64 a_919_553# a_207_553# 0.01fF
C65 a_29_n445# a_n327_n445# 0.03fF
C66 a_327_n389# a_1039_n389# 0.01fF
C67 a_n861_55# a_n861_n943# 0.03fF
C68 a_327_109# a_683_109# 0.03fF
C69 a_n563_n887# a_n29_n887# 0.02fF
C70 a_n741_n887# a_149_n887# 0.01fF
C71 a_n919_n887# a_327_n887# 0.01fF
C72 a_n1097_n887# a_505_n887# 0.01fF
C73 a_n385_n887# a_n207_n887# 0.06fF
C74 a_919_553# a_741_553# 0.10fF
C75 a_n1039_n445# a_n327_n445# 0.01fF
C76 a_563_553# a_n327_553# 0.01fF
C77 a_327_n389# a_861_n389# 0.02fF
C78 a_n207_109# a_n919_109# 0.01fF
C79 a_n563_n887# a_n207_n887# 0.03fF
C80 a_n919_n887# a_149_n887# 0.01fF
C81 a_n1097_n887# a_327_n887# 0.01fF
C82 a_n741_n887# a_n29_n887# 0.01fF
C83 a_n861_n445# a_n683_n445# 0.10fF
C84 a_n1097_109# a_n563_109# 0.02fF
C85 a_505_109# a_n741_109# 0.01fF
C86 a_149_n389# a_n385_n389# 0.02fF
C87 a_n207_607# a_n29_607# 0.06fF
C88 a_327_n389# a_683_n389# 0.03fF
C89 a_n1275_n887# a_327_n887# 0.01fF
C90 a_n741_n887# a_n207_n887# 0.02fF
C91 a_n1097_n887# a_149_n887# 0.01fF
C92 a_n563_n887# a_n385_n887# 0.06fF
C93 a_n919_n887# a_n29_n887# 0.01fF
C94 a_861_109# a_n741_109# 0.01fF
C95 a_n505_553# a_n1039_553# 0.02fF
C96 a_861_607# a_861_n887# 0.00fF
C97 a_327_607# a_n385_607# 0.01fF
C98 a_n149_55# a_n149_n445# 0.15fF
C99 a_n563_109# a_n563_n887# 0.00fF
C100 a_n29_607# a_505_607# 0.02fF
C101 a_n1039_553# a_n1217_553# 0.10fF
C102 a_n861_n445# a_29_n445# 0.01fF
C103 a_n29_109# a_149_109# 0.06fF
C104 a_327_n389# a_505_n389# 0.06fF
C105 a_327_607# a_1217_607# 0.01fF
C106 a_563_55# a_n505_55# 0.01fF
C107 a_n29_607# a_861_607# 0.01fF
C108 a_919_553# a_919_55# 0.15fF
C109 a_n1275_607# a_n29_607# 0.01fF
C110 a_n919_n887# a_n207_n887# 0.01fF
C111 a_n741_n887# a_n385_n887# 0.03fF
C112 a_n1097_n887# a_n29_n887# 0.01fF
C113 a_n1275_n887# a_149_n887# 0.01fF
C114 a_n149_55# a_563_55# 0.01fF
C115 a_n861_n445# a_n1039_n445# 0.10fF
C116 a_149_607# a_149_n887# 0.00fF
C117 a_n1275_109# a_n1275_n887# 0.00fF
C118 a_207_n445# a_207_n943# 0.15fF
C119 a_1039_109# a_n563_109# 0.01fF
C120 a_29_553# a_29_55# 0.15fF
C121 a_741_n445# a_919_n445# 0.10fF
C122 a_683_109# a_683_n389# 0.00fF
C123 a_505_607# a_505_n887# 0.00fF
C124 a_n1097_n887# a_n207_n887# 0.01fF
C125 a_n741_n887# a_n563_n887# 0.06fF
C126 a_n1275_n887# a_n29_n887# 0.01fF
C127 a_n919_n887# a_n385_n887# 0.02fF
C128 a_149_109# a_149_n887# 0.00fF
C129 a_207_n445# a_1097_n445# 0.01fF
C130 a_n505_553# a_563_553# 0.01fF
C131 a_n1097_n389# a_327_n389# 0.01fF
C132 a_741_55# a_n505_55# 0.01fF
C133 a_149_109# a_n1275_109# 0.01fF
C134 a_n1097_109# a_n1097_n887# 0.00fF
C135 a_n861_n445# a_n861_55# 0.15fF
C136 a_741_55# a_n149_55# 0.01fF
C137 a_327_109# a_327_607# 0.00fF
C138 a_919_n445# a_n327_n445# 0.01fF
C139 a_n919_n887# a_n563_n887# 0.03fF
C140 a_n505_n445# a_207_n445# 0.01fF
C141 a_n1097_n887# a_n385_n887# 0.01fF
C142 a_n1275_n887# a_n207_n887# 0.01fF
C143 a_n563_n389# a_1039_n389# 0.01fF
C144 a_683_607# a_149_607# 0.02fF
C145 a_n1039_553# a_n1039_n943# 0.01fF
C146 a_n683_n445# a_n683_553# 0.03fF
C147 a_n207_n389# a_n207_607# 0.00fF
C148 a_683_109# a_n919_109# 0.01fF
C149 a_n1097_n887# a_n563_n887# 0.02fF
C150 a_n919_n887# a_n741_n887# 0.06fF
C151 a_n1275_n887# a_n385_n887# 0.01fF
C152 a_1039_607# a_n563_607# 0.01fF
C153 a_n563_n389# a_861_n389# 0.01fF
C154 a_n1275_607# a_n1275_109# 0.00fF
C155 a_149_109# a_n1097_109# 0.01fF
C156 a_n207_607# a_n207_n887# 0.00fF
C157 a_n1275_n887# a_n563_n887# 0.01fF
C158 a_n385_109# a_n741_109# 0.03fF
C159 a_n207_n389# a_n741_n389# 0.02fF
C160 a_n919_607# a_n919_109# 0.00fF
C161 a_n1097_n887# a_n741_n887# 0.03fF
C162 a_861_109# a_861_n887# 0.00fF
C163 a_n563_n389# a_683_n389# 0.01fF
C164 a_n1097_607# a_n29_607# 0.01fF
C165 a_683_607# a_n207_607# 0.01fF
C166 a_n683_553# a_n149_553# 0.02fF
C167 a_n149_55# a_n149_553# 0.15fF
C168 a_149_109# a_n563_109# 0.01fF
C169 a_919_553# a_919_n943# 0.01fF
C170 a_207_55# a_n683_55# 0.01fF
C171 a_n29_n389# a_149_n389# 0.06fF
C172 a_327_n389# a_n385_n389# 0.01fF
C173 a_327_109# a_n741_109# 0.01fF
C174 a_n1275_n887# a_n741_n887# 0.02fF
C175 a_n1097_n887# a_n919_n887# 0.06fF
C176 a_563_55# a_29_55# 0.02fF
C177 a_207_55# a_1097_55# 0.01fF
C178 a_207_55# a_207_n943# 0.03fF
C179 a_683_607# a_505_607# 0.06fF
C180 a_741_553# a_741_n943# 0.01fF
C181 a_n1217_55# a_n861_55# 0.03fF
C182 a_n563_n389# a_505_n389# 0.01fF
C183 a_505_109# a_505_n887# 0.00fF
C184 a_683_607# a_861_607# 0.06fF
C185 a_n29_109# a_505_109# 0.02fF
C186 a_n1275_n887# a_n919_n887# 0.03fF
C187 a_1039_109# a_149_109# 0.01fF
C188 a_n505_55# a_n861_55# 0.03fF
C189 a_1217_607# a_1217_n887# 0.00fF
C190 a_n149_55# a_n861_55# 0.01fF
C191 a_563_55# a_n1039_55# 0.01fF
C192 a_n29_109# a_861_109# 0.01fF
C193 a_n683_553# a_385_553# 0.01fF
C194 a_n919_607# a_n563_607# 0.03fF
C195 a_741_55# a_29_55# 0.01fF
C196 a_n1275_n887# a_n1097_n887# 0.06fF
C197 a_741_n445# a_207_n445# 0.02fF
C198 a_919_55# a_919_n943# 0.03fF
C199 a_n1097_n389# a_n563_n389# 0.02fF
C200 a_1217_109# a_1217_n887# 0.00fF
C201 a_n327_553# a_207_553# 0.02fF
C202 a_207_553# a_207_n943# 0.01fF
C203 a_n1217_55# a_385_55# 0.01fF
C204 a_741_553# a_n327_553# 0.01fF
C205 a_207_n445# a_n327_n445# 0.02fF
C206 a_n741_n389# a_n741_n887# 0.00fF
C207 a_n29_607# a_n385_607# 0.03fF
C208 a_n1097_n389# a_n1275_n389# 0.06fF
C209 a_919_553# a_n327_553# 0.01fF
C210 a_29_553# a_n861_553# 0.01fF
C211 a_1217_607# a_n29_607# 0.01fF
C212 a_n505_55# a_385_55# 0.01fF
C213 a_n327_55# a_563_55# 0.01fF
C214 a_1217_n389# a_1217_n887# 0.00fF
C215 a_563_n445# a_385_n445# 0.10fF
C216 a_n149_55# a_385_55# 0.02fF
C217 a_n919_n389# a_683_n389# 0.01fF
C218 a_n563_607# a_n563_n389# 0.00fF
C219 a_29_n445# a_29_55# 0.15fF
C220 a_149_109# a_149_607# 0.00fF
C221 a_149_607# a_n207_607# 0.03fF
C222 a_n1097_109# a_505_109# 0.01fF
C223 a_n919_n389# a_505_n389# 0.01fF
C224 a_n1097_607# a_n1097_109# 0.00fF
C225 a_n563_607# a_327_607# 0.01fF
C226 a_n563_n389# a_n385_n389# 0.06fF
C227 a_741_55# a_n327_55# 0.01fF
C228 a_n683_55# a_919_55# 0.01fF
C229 a_149_607# a_505_607# 0.03fF
C230 a_n683_553# a_n1039_553# 0.03fF
C231 a_n741_109# a_n919_109# 0.06fF
C232 a_1039_n389# a_1039_n887# 0.00fF
C233 a_919_n943# a_1097_n943# 0.10fF
C234 a_n861_n445# a_207_n445# 0.01fF
C235 a_505_109# a_n563_109# 0.01fF
C236 a_1097_55# a_919_55# 0.10fF
C237 a_n1275_607# a_n1275_n887# 0.00fF
C238 a_149_607# a_861_607# 0.01fF
C239 a_n919_109# a_n919_n389# 0.00fF
C240 a_n1275_607# a_149_607# 0.01fF
C241 a_n29_n389# a_327_n389# 0.03fF
C242 a_n505_553# a_207_553# 0.01fF
C243 a_n1039_n445# a_n1039_55# 0.15fF
C244 a_29_55# a_n861_55# 0.01fF
C245 a_n29_109# a_n385_109# 0.03fF
C246 a_861_109# a_n563_109# 0.01fF
C247 a_n505_553# a_741_553# 0.01fF
C248 a_n1217_553# a_207_553# 0.01fF
C249 a_n1275_n389# a_n385_n389# 0.01fF
C250 a_563_n445# a_n149_n445# 0.01fF
C251 a_741_n943# a_1097_n943# 0.03fF
C252 a_n29_109# a_1217_109# 0.01fF
C253 a_n1097_n389# a_n919_n389# 0.06fF
C254 a_1039_109# a_505_109# 0.02fF
C255 a_n505_553# a_919_553# 0.01fF
C256 a_n29_109# a_327_109# 0.03fF
C257 a_563_n445# a_563_55# 0.15fF
C258 a_n207_607# a_505_607# 0.01fF
C259 a_741_n943# a_919_n943# 0.10fF
C260 a_861_n389# a_861_n887# 0.00fF
C261 a_563_n943# a_1097_n943# 0.02fF
C262 a_1039_109# a_861_109# 0.06fF
C263 a_n1039_55# a_n861_55# 0.10fF
C264 a_n207_607# a_861_607# 0.01fF
C265 a_563_553# a_n683_553# 0.01fF
C266 a_327_109# a_327_n887# 0.00fF
C267 a_n1275_607# a_n207_607# 0.01fF
C268 a_n385_109# a_n1275_109# 0.01fF
C269 a_563_n943# a_919_n943# 0.03fF
C270 a_385_n943# a_1097_n943# 0.01fF
C271 a_861_607# a_505_607# 0.03fF
C272 a_n919_607# a_n741_607# 0.06fF
C273 a_385_55# a_29_55# 0.03fF
C274 a_683_607# a_n385_607# 0.01fF
C275 a_327_109# a_n1275_109# 0.01fF
C276 a_683_607# a_1217_607# 0.02fF
C277 a_n1097_607# a_n1097_n887# 0.00fF
C278 a_n385_607# a_n385_n887# 0.00fF
C279 a_741_n445# a_741_553# 0.03fF
C280 a_683_n389# a_683_n887# 0.00fF
C281 a_385_n943# a_919_n943# 0.02fF
C282 a_563_n943# a_741_n943# 0.10fF
C283 a_1097_55# a_1097_n943# 0.03fF
C284 a_207_n943# a_1097_n943# 0.01fF
C285 a_1097_553# a_29_553# 0.01fF
C286 a_n327_55# a_n861_55# 0.02fF
C287 a_n385_n389# a_n919_n389# 0.02fF
C288 a_563_n445# a_n683_n445# 0.01fF
C289 a_n149_n445# a_385_n445# 0.02fF
C290 a_385_55# a_n1039_55# 0.01fF
C291 a_n207_n389# a_1217_n389# 0.01fF
C292 a_n1097_607# a_149_607# 0.01fF
C293 a_n385_109# a_n1097_109# 0.01fF
C294 a_385_n943# a_741_n943# 0.03fF
C295 a_29_n943# a_1097_n943# 0.01fF
C296 a_207_n943# a_919_n943# 0.01fF
C297 a_n385_109# a_n385_n887# 0.00fF
C298 a_1097_n445# a_1097_n943# 0.15fF
C299 a_n505_n445# a_n1217_n445# 0.01fF
C300 a_n207_n389# a_1039_n389# 0.01fF
C301 a_n385_109# a_n563_109# 0.06fF
C302 a_149_109# a_505_109# 0.03fF
C303 a_327_109# a_n1097_109# 0.01fF
C304 a_n29_n389# a_n563_n389# 0.02fF
C305 a_207_n943# a_741_n943# 0.02fF
C306 a_563_n445# a_29_n445# 0.02fF
C307 a_29_n943# a_919_n943# 0.01fF
C308 a_385_n943# a_563_n943# 0.10fF
C309 a_505_n389# a_505_n887# 0.00fF
C310 a_n149_n943# a_1097_n943# 0.01fF
C311 a_861_109# a_149_109# 0.01fF
C312 a_n1039_n445# a_563_n445# 0.01fF
C313 a_327_109# a_n563_109# 0.01fF
C314 a_n1039_553# a_n1039_55# 0.15fF
C315 a_n207_n389# a_861_n389# 0.01fF
C316 a_149_n389# a_327_n389# 0.06fF
C317 a_n1097_607# a_n207_607# 0.01fF
C318 a_327_607# a_n741_607# 0.01fF
C319 a_n149_553# a_n861_553# 0.01fF
C320 a_n327_55# a_385_55# 0.01fF
C321 a_1039_109# a_n385_109# 0.01fF
C322 a_207_n943# a_563_n943# 0.03fF
C323 a_n149_n943# a_919_n943# 0.01fF
C324 a_n327_n943# a_1097_n943# 0.01fF
C325 a_29_n943# a_741_n943# 0.01fF
C326 a_n1275_n389# a_n29_n389# 0.01fF
C327 a_505_109# a_505_607# 0.00fF
C328 a_1039_109# a_1217_109# 0.06fF
C329 a_n29_109# a_n919_109# 0.01fF
C330 a_n1097_607# a_505_607# 0.01fF
C331 a_n207_n389# a_683_n389# 0.01fF
C332 a_n1217_553# a_n1217_n445# 0.03fF
C333 a_385_n445# a_n683_n445# 0.01fF
C334 a_n149_n943# a_741_n943# 0.01fF
C335 a_29_n943# a_563_n943# 0.02fF
C336 a_n505_n943# a_1097_n943# 0.01fF
C337 a_n327_n943# a_919_n943# 0.01fF
C338 a_207_n943# a_385_n943# 0.10fF
C339 a_1039_109# a_327_109# 0.01fF
C340 a_n1275_607# a_n1097_607# 0.06fF
C341 a_861_109# a_861_607# 0.00fF
C342 a_29_n445# a_29_553# 0.03fF
C343 a_n563_607# a_n29_607# 0.02fF
C344 a_207_55# a_n1217_55# 0.01fF
C345 a_n207_n389# a_505_n389# 0.01fF
C346 a_n861_553# a_n861_55# 0.15fF
C347 a_29_553# a_n149_553# 0.10fF
C348 a_149_607# a_n385_607# 0.02fF
C349 a_n327_n943# a_741_n943# 0.01fF
C350 a_n505_n943# a_919_n943# 0.01fF
C351 a_n149_n943# a_563_n943# 0.01fF
C352 a_29_n943# a_385_n943# 0.03fF
C353 a_385_553# a_n861_553# 0.01fF
C354 a_n919_109# a_n1275_109# 0.03fF
C355 a_683_607# a_683_n389# 0.00fF
C356 a_29_n445# a_385_n445# 0.03fF
C357 a_149_607# a_1217_607# 0.01fF
C358 a_207_55# a_n505_55# 0.01fF
C359 a_n149_55# a_207_55# 0.03fF
C360 a_1039_109# a_1039_n389# 0.00fF
C361 a_n1039_n445# a_385_n445# 0.01fF
C362 a_n327_n943# a_563_n943# 0.01fF
C363 a_29_n943# a_207_n943# 0.10fF
C364 a_n505_n943# a_741_n943# 0.01fF
C365 a_n683_n943# a_919_n943# 0.01fF
C366 a_n149_n943# a_385_n943# 0.02fF
C367 a_1097_n445# a_1097_55# 0.15fF
C368 a_n741_109# a_n741_607# 0.00fF
C369 a_n1097_n389# a_n207_n389# 0.01fF
C370 a_741_55# a_563_55# 0.10fF
C371 a_n29_n389# a_n919_n389# 0.01fF
C372 a_n207_607# a_n385_607# 0.06fF
C373 a_n149_n445# a_n683_n445# 0.02fF
C374 a_563_n445# a_919_n445# 0.03fF
C375 a_n683_n943# a_741_n943# 0.01fF
C376 a_n327_n943# a_385_n943# 0.01fF
C377 a_n149_n943# a_207_n943# 0.03fF
C378 a_385_553# a_29_553# 0.03fF
C379 a_n505_n943# a_563_n943# 0.01fF
C380 a_n207_607# a_1217_607# 0.01fF
C381 a_n385_109# a_149_109# 0.02fF
C382 a_n1217_n445# a_n1217_n943# 0.15fF
C383 a_n385_607# a_505_607# 0.01fF
C384 a_n327_n445# a_n1217_n445# 0.01fF
C385 a_n1097_109# a_n919_109# 0.06fF
C386 a_n327_553# a_n327_n943# 0.01fF
C387 a_n505_n445# a_1097_n445# 0.01fF
C388 a_385_n445# a_385_553# 0.03fF
C389 a_n505_n943# a_385_n943# 0.01fF
C390 a_n149_n943# a_29_n943# 0.10fF
C391 a_n861_n943# a_741_n943# 0.01fF
C392 a_n683_n943# a_563_n943# 0.01fF
C393 a_n327_n943# a_207_n943# 0.02fF
C394 a_149_109# a_1217_109# 0.01fF
C395 a_861_607# a_n385_607# 0.01fF
C396 a_n207_109# a_683_109# 0.01fF
C397 a_n1275_607# a_n385_607# 0.01fF
C398 a_1217_607# a_505_607# 0.01fF
C399 a_n683_553# a_207_553# 0.01fF
C400 a_n1097_n389# a_n1097_109# 0.00fF
C401 a_149_n389# a_n563_n389# 0.01fF
C402 a_n505_553# a_n327_553# 0.10fF
C403 a_n149_n445# a_29_n445# 0.10fF
C404 a_149_109# a_327_109# 0.06fF
C405 a_1217_607# a_861_607# 0.03fF
C406 a_n563_109# a_n919_109# 0.03fF
C407 a_741_n445# a_741_n943# 0.15fF
C408 a_n683_553# a_741_553# 0.01fF
C409 a_n1217_553# a_n327_553# 0.01fF
C410 a_n149_n445# a_n149_553# 0.03fF
C411 a_861_109# a_505_109# 0.03fF
C412 a_n1039_n445# a_n149_n445# 0.01fF
C413 a_n505_n943# a_207_n943# 0.01fF
C414 a_n327_n943# a_29_n943# 0.03fF
C415 a_n683_n943# a_385_n943# 0.01fF
C416 a_n861_n943# a_563_n943# 0.01fF
C417 a_919_553# a_n683_553# 0.01fF
C418 a_1097_553# a_n149_553# 0.01fF
C419 a_n1039_553# a_n861_553# 0.10fF
C420 a_n683_55# a_n683_n943# 0.03fF
C421 a_n207_n389# a_n385_n389# 0.06fF
C422 a_n1275_n389# a_149_n389# 0.01fF
C423 a_n1039_n943# a_563_n943# 0.01fF
C424 a_n861_n943# a_385_n943# 0.01fF
C425 a_n327_n943# a_n149_n943# 0.10fF
C426 a_n683_n943# a_207_n943# 0.01fF
C427 a_n505_n943# a_29_n943# 0.02fF
C428 a_385_n445# a_385_55# 0.15fF
C429 a_683_607# a_n563_607# 0.01fF
C430 a_n505_553# a_n505_n445# 0.03fF
C431 a_919_n445# a_385_n445# 0.02fF
C432 a_n861_n445# a_n1217_n445# 0.03fF
C433 a_207_55# a_29_55# 0.10fF
C434 a_n505_n445# a_n505_n943# 0.15fF
C435 a_563_553# a_563_n445# 0.03fF
C436 a_n861_n943# a_207_n943# 0.01fF
C437 a_n505_n943# a_n149_n943# 0.03fF
C438 a_n1039_n943# a_385_n943# 0.01fF
C439 a_n683_n943# a_29_n943# 0.01fF
C440 a_n919_109# a_n919_n887# 0.00fF
C441 a_563_55# a_n861_55# 0.01fF
C442 a_n1039_553# a_29_553# 0.01fF
C443 a_n505_55# a_919_55# 0.01fF
C444 a_n563_607# a_n563_109# 0.00fF
C445 a_1097_553# a_385_553# 0.01fF
C446 a_n149_55# a_919_55# 0.01fF
C447 a_563_553# a_n861_553# 0.01fF
C448 a_n29_607# a_n741_607# 0.01fF
C449 a_29_n445# a_n683_n445# 0.01fF
C450 a_n563_607# a_n563_n887# 0.00fF
C451 a_n505_n943# a_n327_n943# 0.10fF
C452 a_n1039_n943# a_207_n943# 0.01fF
C453 a_n683_n943# a_n149_n943# 0.02fF
C454 a_n861_n943# a_29_n943# 0.01fF
C455 a_n1217_n943# a_385_n943# 0.01fF
C456 a_n385_n389# a_n385_n887# 0.00fF
C457 a_n29_n389# a_n29_607# 0.00fF
C458 a_207_55# a_n1039_55# 0.01fF
C459 a_n1039_n445# a_n683_n445# 0.03fF
C460 a_n505_553# a_n1217_553# 0.01fF
C461 a_n505_553# a_n505_n943# 0.01fF
C462 a_n1097_607# a_n385_607# 0.01fF
C463 a_n1097_n389# a_n1097_n887# 0.00fF
C464 a_n327_n445# a_n327_553# 0.03fF
C465 a_741_n445# a_1097_n445# 0.03fF
C466 a_741_55# a_n861_55# 0.01fF
C467 a_n1039_n943# a_29_n943# 0.01fF
C468 a_n861_n943# a_n149_n943# 0.01fF
C469 a_n683_n943# a_n327_n943# 0.03fF
C470 a_n1217_n943# a_207_n943# 0.01fF
C471 a_n741_n389# a_861_n389# 0.01fF
C472 a_861_607# a_861_n389# 0.00fF
C473 a_149_n389# a_n919_n389# 0.01fF
C474 a_563_n445# a_207_n445# 0.03fF
C475 a_n149_n445# a_919_n445# 0.01fF
C476 a_n505_n445# a_741_n445# 0.01fF
C477 a_563_553# a_29_553# 0.02fF
C478 a_n385_109# a_505_109# 0.01fF
C479 a_563_55# a_385_55# 0.10fF
C480 a_n1039_n445# a_29_n445# 0.01fF
C481 a_n29_109# a_n29_n389# 0.00fF
C482 a_n861_n943# a_n327_n943# 0.02fF
C483 a_n683_n943# a_n505_n943# 0.10fF
C484 a_n1039_n943# a_n149_n943# 0.01fF
C485 a_n1217_n943# a_29_n943# 0.01fF
C486 a_n327_n445# a_1097_n445# 0.01fF
C487 a_n1217_55# a_n1217_n445# 0.15fF
C488 a_505_109# a_1217_109# 0.01fF
C489 a_n741_n389# a_683_n389# 0.01fF
C490 a_149_109# a_n919_109# 0.01fF
C491 a_861_109# a_n385_109# 0.01fF
C492 a_207_55# a_n327_55# 0.02fF
C493 a_n505_n445# a_n327_n445# 0.10fF
C494 a_327_n389# a_n563_n389# 0.01fF
C495 a_327_109# a_505_109# 0.06fF
C496 a_505_607# a_505_n389# 0.00fF
C497 a_861_109# a_1217_109# 0.03fF
C498 a_n1039_n943# a_n327_n943# 0.01fF
C499 a_n861_n943# a_n505_n943# 0.03fF
C500 a_n1217_n943# a_n149_n943# 0.01fF
C501 a_n741_n389# a_505_n389# 0.01fF
C502 a_1039_607# a_327_607# 0.01fF
C503 a_861_109# a_327_109# 0.02fF
C504 a_741_55# a_385_55# 0.03fF
C505 a_n861_n943# a_n683_n943# 0.10fF
C506 a_n327_n445# a_n327_n943# 0.15fF
C507 a_327_n389# a_327_607# 0.00fF
C508 a_n1217_n943# a_n327_n943# 0.01fF
C509 a_n1039_n943# a_n505_n943# 0.02fF
C510 a_149_607# a_n563_607# 0.01fF
C511 a_n1275_n389# a_327_n389# 0.01fF
C512 a_n207_109# a_n741_109# 0.02fF
C513 a_385_553# a_n149_553# 0.02fF
C514 a_n207_n389# a_n29_n389# 0.06fF
C515 a_n29_n389# a_n29_n887# 0.00fF
C516 a_919_55# a_29_55# 0.01fF
C517 a_385_n445# a_207_n445# 0.10fF
C518 a_919_n445# a_n683_n445# 0.01fF
C519 a_n1097_n389# a_n741_n389# 0.03fF
C520 a_n1217_553# a_n1217_n943# 0.01fF
C521 a_n1039_n943# a_n683_n943# 0.03fF
C522 a_n1217_n943# a_n505_n943# 0.01fF
C523 a_1217_607# a_n385_607# 0.01fF
C524 a_n861_n445# a_n505_n445# 0.03fF
C525 a_683_607# a_n741_607# 0.01fF
C526 a_n207_607# a_n563_607# 0.03fF
C527 a_563_553# a_1097_553# 0.02fF
C528 a_n1039_n943# a_n861_n943# 0.10fF
C529 a_n1217_n943# a_n683_n943# 0.02fF
C530 a_n385_109# a_n385_607# 0.00fF
C531 a_563_553# a_563_55# 0.15fF
C532 a_861_109# a_861_n389# 0.00fF
C533 a_29_n445# a_919_n445# 0.01fF
C534 a_n563_607# a_505_607# 0.01fF
C535 a_1217_607# a_1217_109# 0.00fF
C536 a_n1217_n943# a_n861_n943# 0.03fF
C537 a_n919_607# a_327_607# 0.01fF
C538 a_n1217_55# a_n683_55# 0.02fF
C539 a_n563_607# a_861_607# 0.01fF
C540 a_n1275_607# a_n563_607# 0.01fF
C541 a_505_109# a_505_n389# 0.00fF
C542 a_741_n445# a_n327_n445# 0.01fF
C543 a_327_n389# a_n919_n389# 0.01fF
C544 a_n385_109# a_1217_109# 0.01fF
C545 a_n149_n445# a_207_n445# 0.03fF
C546 a_n1217_n943# a_n1039_n943# 0.10fF
C547 a_n505_55# a_n683_55# 0.10fF
C548 a_n683_553# a_n683_55# 0.15fF
C549 a_n149_55# a_n683_55# 0.02fF
C550 a_n683_553# a_n327_553# 0.03fF
C551 a_n505_55# a_1097_55# 0.01fF
C552 a_385_55# a_n861_55# 0.01fF
C553 a_1217_607# a_1217_n389# 0.00fF
C554 a_n741_607# a_n741_n887# 0.00fF
C555 a_n327_55# a_919_55# 0.01fF
C556 a_n385_109# a_327_109# 0.01fF
C557 a_n741_n389# a_n385_n389# 0.03fF
C558 a_n149_55# a_1097_55# 0.01fF
C559 a_n1039_553# a_n149_553# 0.01fF
C560 a_505_109# a_n919_109# 0.01fF
C561 a_n1039_n445# a_n1039_553# 0.03fF
C562 a_385_553# a_385_55# 0.15fF
C563 a_327_109# a_1217_109# 0.01fF
C564 a_683_109# a_n741_109# 0.01fF
C565 a_n1097_607# a_n1097_n389# 0.00fF
C566 a_1217_109# a_1217_n389# 0.00fF
C567 a_n861_553# a_207_553# 0.01fF
C568 a_n861_n445# a_n861_n943# 0.15fF
C569 a_n1275_n389# a_n563_n389# 0.01fF
C570 a_n505_n445# a_n505_55# 0.15fF
C571 a_149_n389# a_149_n887# 0.00fF
C572 a_741_553# a_n861_553# 0.01fF
C573 a_n861_n445# a_741_n445# 0.01fF
C574 a_n149_55# a_n149_n943# 0.03fF
C575 a_385_553# a_n1039_553# 0.01fF
C576 a_n207_n389# a_149_n389# 0.03fF
C577 a_563_553# a_n149_553# 0.01fF
C578 a_n919_607# a_n919_n389# 0.00fF
C579 a_1039_607# a_1039_n887# 0.00fF
C580 a_n683_n445# a_207_n445# 0.01fF
C581 a_n1217_55# a_n1217_553# 0.15fF
C582 a_149_607# a_n741_607# 0.01fF
C583 a_29_553# a_207_553# 0.10fF
C584 a_n1097_607# a_n563_607# 0.02fF
C585 a_n861_n445# a_n327_n445# 0.02fF
C586 a_n505_553# a_n505_55# 0.15fF
C587 a_n29_109# a_n207_109# 0.06fF
C588 a_n505_553# a_n683_553# 0.10fF
C589 a_29_553# a_741_553# 0.01fF
C590 a_1039_n389# a_1217_n389# 0.06fF
C591 a_n505_55# a_n505_n943# 0.03fF
C592 a_n683_553# a_n1217_553# 0.02fF
C593 a_1039_607# a_n29_607# 0.01fF
C594 a_919_553# a_29_553# 0.01fF
C595 a_29_n445# a_207_n445# 0.10fF
C596 a_563_553# a_385_553# 0.10fF
C597 a_861_n389# a_1217_n389# 0.03fF
C598 a_n563_n389# a_n919_n389# 0.03fF
C599 a_n683_55# a_29_55# 0.01fF
C600 a_n1039_n445# a_207_n445# 0.01fF
C601 a_n683_553# a_n683_n943# 0.01fF
C602 a_207_55# a_563_55# 0.03fF
C603 a_n207_607# a_n741_607# 0.02fF
C604 a_1097_55# a_29_55# 0.01fF
C605 a_n207_109# a_n1275_109# 0.01fF
C606 a_683_n389# a_1217_n389# 0.02fF
C607 a_861_n389# a_1039_n389# 0.06fF
C608 a_n207_n389# a_n207_109# 0.00fF
C609 a_n741_607# a_505_607# 0.01fF
C610 a_n385_109# a_n919_109# 0.02fF
C611 a_861_607# a_n741_607# 0.01fF
C612 a_29_55# a_29_n943# 0.03fF
C613 a_n741_n389# a_n741_607# 0.00fF
C614 a_n1275_607# a_n741_607# 0.02fF
C615 a_n1275_n389# a_n919_n389# 0.03fF
C616 a_n29_n389# a_n741_n389# 0.01fF
C617 a_n683_55# a_n1039_55# 0.03fF
C618 a_505_n389# a_1217_n389# 0.01fF
C619 a_683_n389# a_1039_n389# 0.03fF
C620 a_741_55# a_207_55# 0.02fF
C621 a_683_109# a_683_n887# 0.00fF
C622 a_327_109# a_n919_109# 0.01fF
C623 a_n207_109# a_n207_n887# 0.00fF
C624 a_n1217_55# a_n1217_n943# 0.03fF
C625 a_327_n389# a_327_n887# 0.00fF
C626 a_n563_607# a_n385_607# 0.06fF
C627 a_683_n389# a_861_n389# 0.06fF
C628 a_505_n389# a_1039_n389# 0.02fF
C629 a_1097_553# a_207_553# 0.01fF
C630 a_n1097_109# a_n207_109# 0.01fF
C631 a_n919_607# a_n29_607# 0.01fF
C632 a_1097_553# a_741_553# 0.03fF
C633 a_n29_109# a_683_109# 0.01fF
C634 a_n207_109# a_n563_109# 0.03fF
C635 a_1097_553# a_919_553# 0.10fF
C636 a_n385_n389# a_n385_607# 0.00fF
C637 a_505_n389# a_861_n389# 0.03fF
C638 a_n327_55# a_n683_55# 0.03fF
C639 a_n327_55# a_n327_553# 0.15fF
C640 a_563_553# a_n1039_553# 0.01fF
C641 a_n207_n389# a_327_n389# 0.02fF
C642 a_n327_55# a_1097_55# 0.01fF
C643 a_919_n445# a_207_n445# 0.01fF
C644 a_505_n389# a_683_n389# 0.06fF
C645 a_149_n389# a_149_607# 0.00fF
C646 a_1039_109# a_n207_109# 0.01fF
C647 a_741_55# a_741_553# 0.15fF
C648 a_683_607# a_1039_607# 0.03fF
C649 a_n385_109# a_n385_n389# 0.00fF
C650 a_563_n445# a_563_n943# 0.15fF
C651 a_n1097_607# a_n741_607# 0.03fF
C652 a_563_55# a_919_55# 0.03fF
C653 a_149_109# a_149_n389# 0.00fF
C654 a_385_n445# a_n1217_n445# 0.01fF
C655 a_327_607# a_n29_607# 0.03fF
C656 a_207_55# a_n861_55# 0.01fF
C657 a_n385_n389# a_1217_n389# 0.01fF
C658 a_n327_55# a_n327_n943# 0.03fF
C659 a_n1097_n389# a_505_n389# 0.01fF
C660 a_683_607# a_683_109# 0.00fF
C661 a_n149_553# a_207_553# 0.03fF
C662 a_1039_109# a_1039_607# 0.00fF
C663 a_741_55# a_919_55# 0.10fF
C664 a_741_553# a_n149_553# 0.01fF
C665 a_n385_n389# a_1039_n389# 0.01fF
C666 a_149_n389# a_n741_n389# 0.01fF
C667 a_n327_553# a_n861_553# 0.02fF
C668 a_919_553# a_n149_553# 0.01fF
C669 a_683_109# a_n563_109# 0.01fF
C670 a_683_607# a_n919_607# 0.01fF
C671 a_327_607# a_327_n887# 0.00fF
C672 a_n1039_55# a_n1039_n943# 0.03fF
C673 a_n385_n389# a_861_n389# 0.01fF
C674 a_563_n445# a_1097_n445# 0.02fF
C675 a_n149_n445# a_n1217_n445# 0.01fF
C676 a_207_55# a_385_55# 0.10fF
C677 a_149_109# a_n207_109# 0.03fF
C678 a_n1217_55# a_n505_55# 0.01fF
C679 a_n207_n389# a_n563_n389# 0.03fF
C680 a_563_n445# a_n505_n445# 0.01fF
C681 a_n149_55# a_n1217_55# 0.01fF
C682 a_385_553# a_207_553# 0.10fF
C683 a_1097_553# a_1097_n943# 0.01fF
C684 a_n385_n389# a_683_n389# 0.01fF
C685 a_1039_109# a_683_109# 0.03fF
C686 a_n741_607# a_n385_607# 0.03fF
C687 a_385_553# a_741_553# 0.03fF
C688 a_n207_109# a_n207_607# 0.00fF
C689 a_29_553# a_n327_553# 0.03fF
C690 a_385_n445# a_385_n943# 0.15fF
C691 a_n1275_n389# a_n1275_109# 0.00fF
C692 a_n149_55# a_n505_55# 0.03fF
C693 a_919_553# a_385_553# 0.02fF
C694 a_149_607# a_1039_607# 0.01fF
C695 a_n385_n389# a_505_n389# 0.01fF
C696 a_n1275_n389# a_n207_n389# 0.01fF
C697 a_29_553# a_29_n943# 0.01fF
C698 a_1039_n887# a_1217_n887# 0.06fF
C699 a_n29_109# a_n741_109# 0.01fF
C700 a_n505_553# a_n861_553# 0.03fF
C701 a_n327_n445# a_n327_55# 0.15fF
C702 a_n919_607# a_n919_n887# 0.00fF
C703 a_n563_n389# a_n563_109# 0.00fF
C704 a_683_607# a_327_607# 0.03fF
C705 a_861_n887# a_1217_n887# 0.03fF
C706 a_385_n445# a_1097_n445# 0.01fF
C707 a_n683_n445# a_n1217_n445# 0.02fF
C708 a_n1217_553# a_n861_553# 0.03fF
C709 a_n1097_n389# a_n385_n389# 0.01fF
C710 a_1039_607# a_n207_607# 0.01fF
C711 a_n563_n389# a_n563_n887# 0.00fF
C712 a_563_55# a_563_n943# 0.03fF
C713 a_n505_n445# a_385_n445# 0.01fF
C714 a_919_553# a_919_n445# 0.03fF
C715 a_n29_n389# a_1217_n389# 0.01fF
C716 a_683_n887# a_1217_n887# 0.02fF
C717 a_861_n887# a_1039_n887# 0.06fF
C718 a_n741_109# a_n1275_109# 0.02fF
C719 a_1039_607# a_505_607# 0.02fF
C720 a_741_55# a_741_n943# 0.03fF
C721 a_1039_607# a_861_607# 0.06fF
C722 a_n505_553# a_29_553# 0.02fF
C723 a_n1039_553# a_207_553# 0.01fF
C724 a_29_n445# a_n1217_n445# 0.01fF
C725 a_n29_n389# a_1039_n389# 0.01fF
C726 a_n1217_553# a_29_553# 0.01fF
C727 a_149_109# a_683_109# 0.02fF
C728 a_505_n887# a_1217_n887# 0.01fF
C729 a_683_n887# a_1039_n887# 0.03fF
C730 a_n207_n389# a_n919_n389# 0.01fF
C731 a_n919_607# a_149_607# 0.01fF
C732 a_327_n389# a_n741_n389# 0.01fF
C733 a_n861_553# a_n861_n943# 0.01fF
C734 a_563_n445# a_741_n445# 0.10fF
C735 a_n1039_n445# a_n1217_n445# 0.10fF
C736 a_563_55# a_n683_55# 0.01fF
C737 a_n1217_55# a_29_55# 0.01fF
C738 a_1097_553# a_n327_553# 0.01fF
C739 a_1097_553# a_1097_55# 0.15fF
C740 a_563_55# a_1097_55# 0.02fF
C741 a_385_55# a_919_55# 0.02fF
C742 a_919_n445# a_919_55# 0.15fF
C743 a_n29_n389# a_861_n389# 0.01fF
C744 a_327_n887# a_1217_n887# 0.01fF
C745 a_683_n887# a_861_n887# 0.06fF
C746 a_505_n887# a_1039_n887# 0.02fF
C747 a_n149_n445# a_1097_n445# 0.01fF
C748 a_n505_55# a_29_55# 0.02fF
C749 a_n207_109# a_505_109# 0.01fF
C750 a_n149_55# a_29_55# 0.10fF
C751 a_563_n445# a_n327_n445# 0.01fF
C752 a_n1097_109# a_n741_109# 0.03fF
C753 a_207_n445# a_207_55# 0.15fF
C754 a_n149_n445# a_n505_n445# 0.03fF
C755 a_1097_553# a_1097_n445# 0.03fF
C756 a_563_553# a_207_553# 0.03fF
C757 a_n1217_55# a_n1039_55# 0.10fF
C758 a_n919_607# a_n207_607# 0.01fF
C759 a_n29_n389# a_683_n389# 0.01fF
C760 a_n149_n445# a_n149_n943# 0.15fF
C761 a_861_109# a_n207_109# 0.01fF
C762 a_149_n887# a_1217_n887# 0.01fF
C763 a_505_n887# a_861_n887# 0.03fF
C764 a_327_n887# a_1039_n887# 0.01fF
C765 a_741_55# a_n683_55# 0.01fF
C766 a_563_553# a_741_553# 0.10fF
C767 a_741_55# a_1097_55# 0.03fF
C768 a_n741_109# a_n563_109# 0.06fF
C769 a_n505_55# a_n1039_55# 0.02fF
C770 a_n919_607# a_505_607# 0.01fF
C771 a_563_553# a_919_553# 0.03fF
C772 a_n29_n389# a_505_n389# 0.02fF
C773 a_n149_55# a_n1039_55# 0.01fF
C774 a_n29_109# a_n29_607# 0.00fF
C775 a_n29_n887# a_1217_n887# 0.01fF
C776 a_149_n887# a_1039_n887# 0.01fF
C777 a_505_n887# a_683_n887# 0.06fF
C778 a_327_n887# a_861_n887# 0.02fF
C779 a_n1275_607# a_n919_607# 0.03fF
C780 a_n683_n445# a_n683_55# 0.15fF
C781 a_741_n445# a_385_n445# 0.03fF
C782 a_149_607# a_327_607# 0.06fF
C783 a_n1275_n389# a_n1275_n887# 0.00fF
C784 a_n741_109# a_n741_n887# 0.00fF
C785 a_327_n887# a_683_n887# 0.03fF
C786 a_n505_553# a_1097_553# 0.01fF
C787 a_149_n887# a_861_n887# 0.01fF
C788 a_n207_n887# a_1217_n887# 0.01fF
C789 a_n29_n887# a_1039_n887# 0.01fF
C790 a_n1217_55# a_n327_55# 0.01fF
C791 a_207_n445# a_207_553# 0.03fF
C792 a_n861_n445# a_563_n445# 0.01fF
C793 a_n1097_n389# a_n29_n389# 0.01fF
C794 a_n861_n445# a_n861_553# 0.03fF
C795 a_385_n445# a_n327_n445# 0.01fF
C796 a_n327_55# a_n505_55# 0.10fF
C797 a_n29_n887# a_861_n887# 0.01fF
C798 a_149_n887# a_683_n887# 0.02fF
C799 a_n385_n887# a_1217_n887# 0.01fF
C800 a_n207_n887# a_1039_n887# 0.01fF
C801 a_n327_553# a_n149_553# 0.10fF
C802 a_327_n887# a_505_n887# 0.06fF
C803 a_n505_n445# a_n683_n445# 0.10fF
C804 a_n149_55# a_n327_55# 0.10fF
C805 a_n919_n389# a_n919_n887# 0.00fF
C806 a_149_n389# a_1217_n389# 0.01fF
C807 a_n207_607# a_327_607# 0.02fF
C808 a_n741_n389# a_n563_n389# 0.06fF
C809 a_n29_607# a_n29_n887# 0.00fF
C810 a_919_n445# a_919_n943# 0.15fF
C811 a_29_n445# a_29_n943# 0.15fF
C812 a_n207_n887# a_861_n887# 0.01fF
C813 a_149_n887# a_505_n887# 0.03fF
C814 a_n29_n887# a_683_n887# 0.01fF
C815 a_n385_n887# a_1039_n887# 0.01fF
C816 a_29_n445# a_1097_n445# 0.01fF
C817 a_505_109# a_683_109# 0.06fF
C818 a_327_607# a_505_607# 0.06fF
C819 a_149_n389# a_1039_n389# 0.01fF
C820 a_385_553# a_385_n943# 0.01fF
C821 a_n29_109# a_n1275_109# 0.01fF
C822 a_n563_607# a_n741_607# 0.06fF
C823 a_n149_n445# a_741_n445# 0.01fF
C824 a_n505_n445# a_29_n445# 0.02fF
C825 a_327_607# a_861_607# 0.02fF
C826 a_n1275_607# a_327_607# 0.01fF
C827 a_n683_55# a_n861_55# 0.10fF
C828 a_n385_109# a_n207_109# 0.06fF
C829 a_683_607# a_n29_607# 0.01fF
C830 a_861_109# a_683_109# 0.06fF
C831 a_n563_n887# a_1039_n887# 0.01fF
C832 a_149_n887# a_327_n887# 0.06fF
C833 a_n385_n887# a_861_n887# 0.01fF
C834 a_n207_n887# a_683_n887# 0.01fF
C835 a_n1275_n389# a_n741_n389# 0.02fF
C836 a_n29_n887# a_505_n887# 0.02fF
C837 a_n1275_607# a_n1275_n389# 0.00fF
C838 a_n1039_n445# a_n505_n445# 0.02fF
C839 a_n149_553# a_n149_n943# 0.01fF
C840 a_385_553# a_n327_553# 0.01fF
C841 a_149_n389# a_861_n389# 0.01fF
C842 a_n29_109# a_n29_n887# 0.00fF
C843 a_683_607# a_683_n887# 0.00fF
C844 a_n207_109# a_1217_109# 0.01fF
C845 a_n1097_607# a_n919_607# 0.06fF
C846 a_n861_n445# a_385_n445# 0.01fF
C847 a_n149_n445# a_n327_n445# 0.10fF
C848 a_1039_109# a_1039_n887# 0.00fF
C849 a_n29_n389# a_n385_n389# 0.03fF
C850 a_n207_n887# a_505_n887# 0.01fF
C851 a_n385_n887# a_683_n887# 0.01fF
C852 a_n563_n887# a_861_n887# 0.01fF
C853 a_n1039_55# a_29_55# 0.01fF
C854 a_n29_n887# a_327_n887# 0.03fF
C855 a_327_109# a_n207_109# 0.02fF
C856 a_1039_607# a_n385_607# 0.01fF
C857 a_149_109# a_n741_109# 0.01fF
C858 a_1217_n887# a_n1555_n1061# 0.10fF
C859 a_1039_n887# a_n1555_n1061# 0.05fF
C860 a_861_n887# a_n1555_n1061# 0.04fF
C861 a_683_n887# a_n1555_n1061# 0.03fF
C862 a_505_n887# a_n1555_n1061# 0.03fF
C863 a_327_n887# a_n1555_n1061# 0.03fF
C864 a_149_n887# a_n1555_n1061# 0.03fF
C865 a_n29_n887# a_n1555_n1061# 0.03fF
C866 a_n207_n887# a_n1555_n1061# 0.03fF
C867 a_n385_n887# a_n1555_n1061# 0.03fF
C868 a_n563_n887# a_n1555_n1061# 0.03fF
C869 a_n741_n887# a_n1555_n1061# 0.03fF
C870 a_n919_n887# a_n1555_n1061# 0.04fF
C871 a_n1097_n887# a_n1555_n1061# 0.05fF
C872 a_n1275_n887# a_n1555_n1061# 0.10fF
C873 a_1097_n943# a_n1555_n1061# 0.27fF
C874 a_919_n943# a_n1555_n1061# 0.23fF
C875 a_741_n943# a_n1555_n1061# 0.23fF
C876 a_563_n943# a_n1555_n1061# 0.24fF
C877 a_385_n943# a_n1555_n1061# 0.24fF
C878 a_207_n943# a_n1555_n1061# 0.25fF
C879 a_29_n943# a_n1555_n1061# 0.26fF
C880 a_n149_n943# a_n1555_n1061# 0.26fF
C881 a_n327_n943# a_n1555_n1061# 0.26fF
C882 a_n505_n943# a_n1555_n1061# 0.26fF
C883 a_n683_n943# a_n1555_n1061# 0.26fF
C884 a_n861_n943# a_n1555_n1061# 0.26fF
C885 a_n1039_n943# a_n1555_n1061# 0.27fF
C886 a_n1217_n943# a_n1555_n1061# 0.32fF
C887 a_1217_n389# a_n1555_n1061# 0.10fF
C888 a_1039_n389# a_n1555_n1061# 0.05fF
C889 a_861_n389# a_n1555_n1061# 0.04fF
C890 a_683_n389# a_n1555_n1061# 0.03fF
C891 a_505_n389# a_n1555_n1061# 0.03fF
C892 a_327_n389# a_n1555_n1061# 0.02fF
C893 a_149_n389# a_n1555_n1061# 0.03fF
C894 a_n29_n389# a_n1555_n1061# 0.03fF
C895 a_n207_n389# a_n1555_n1061# 0.03fF
C896 a_n385_n389# a_n1555_n1061# 0.02fF
C897 a_n563_n389# a_n1555_n1061# 0.03fF
C898 a_n741_n389# a_n1555_n1061# 0.03fF
C899 a_n919_n389# a_n1555_n1061# 0.04fF
C900 a_n1097_n389# a_n1555_n1061# 0.05fF
C901 a_n1275_n389# a_n1555_n1061# 0.10fF
C902 a_1097_n445# a_n1555_n1061# 0.22fF
C903 a_919_n445# a_n1555_n1061# 0.18fF
C904 a_741_n445# a_n1555_n1061# 0.18fF
C905 a_563_n445# a_n1555_n1061# 0.19fF
C906 a_385_n445# a_n1555_n1061# 0.19fF
C907 a_207_n445# a_n1555_n1061# 0.20fF
C908 a_29_n445# a_n1555_n1061# 0.21fF
C909 a_n149_n445# a_n1555_n1061# 0.21fF
C910 a_n327_n445# a_n1555_n1061# 0.21fF
C911 a_n505_n445# a_n1555_n1061# 0.21fF
C912 a_n683_n445# a_n1555_n1061# 0.21fF
C913 a_n861_n445# a_n1555_n1061# 0.21fF
C914 a_n1039_n445# a_n1555_n1061# 0.22fF
C915 a_n1217_n445# a_n1555_n1061# 0.27fF
C916 a_1217_109# a_n1555_n1061# 0.10fF
C917 a_1039_109# a_n1555_n1061# 0.05fF
C918 a_861_109# a_n1555_n1061# 0.04fF
C919 a_683_109# a_n1555_n1061# 0.03fF
C920 a_505_109# a_n1555_n1061# 0.03fF
C921 a_327_109# a_n1555_n1061# 0.03fF
C922 a_149_109# a_n1555_n1061# 0.03fF
C923 a_n29_109# a_n1555_n1061# 0.03fF
C924 a_n207_109# a_n1555_n1061# 0.03fF
C925 a_n385_109# a_n1555_n1061# 0.03fF
C926 a_n563_109# a_n1555_n1061# 0.03fF
C927 a_n741_109# a_n1555_n1061# 0.03fF
C928 a_n919_109# a_n1555_n1061# 0.04fF
C929 a_n1097_109# a_n1555_n1061# 0.06fF
C930 a_n1275_109# a_n1555_n1061# 0.10fF
C931 a_1097_55# a_n1555_n1061# 0.23fF
C932 a_919_55# a_n1555_n1061# 0.20fF
C933 a_741_55# a_n1555_n1061# 0.20fF
C934 a_563_55# a_n1555_n1061# 0.20fF
C935 a_385_55# a_n1555_n1061# 0.21fF
C936 a_207_55# a_n1555_n1061# 0.21fF
C937 a_29_55# a_n1555_n1061# 0.22fF
C938 a_n149_55# a_n1555_n1061# 0.22fF
C939 a_n327_55# a_n1555_n1061# 0.22fF
C940 a_n505_55# a_n1555_n1061# 0.22fF
C941 a_n683_55# a_n1555_n1061# 0.22fF
C942 a_n861_55# a_n1555_n1061# 0.23fF
C943 a_n1039_55# a_n1555_n1061# 0.23fF
C944 a_n1217_55# a_n1555_n1061# 0.28fF
C945 a_1217_607# a_n1555_n1061# 0.10fF
C946 a_1039_607# a_n1555_n1061# 0.06fF
C947 a_861_607# a_n1555_n1061# 0.05fF
C948 a_683_607# a_n1555_n1061# 0.04fF
C949 a_505_607# a_n1555_n1061# 0.03fF
C950 a_327_607# a_n1555_n1061# 0.03fF
C951 a_149_607# a_n1555_n1061# 0.03fF
C952 a_n29_607# a_n1555_n1061# 0.04fF
C953 a_n207_607# a_n1555_n1061# 0.03fF
C954 a_n385_607# a_n1555_n1061# 0.03fF
C955 a_n563_607# a_n1555_n1061# 0.03fF
C956 a_n741_607# a_n1555_n1061# 0.04fF
C957 a_n919_607# a_n1555_n1061# 0.05fF
C958 a_n1097_607# a_n1555_n1061# 0.06fF
C959 a_n1275_607# a_n1555_n1061# 0.10fF
C960 a_1097_553# a_n1555_n1061# 0.30fF
C961 a_919_553# a_n1555_n1061# 0.26fF
C962 a_741_553# a_n1555_n1061# 0.26fF
C963 a_563_553# a_n1555_n1061# 0.27fF
C964 a_385_553# a_n1555_n1061# 0.27fF
C965 a_207_553# a_n1555_n1061# 0.28fF
C966 a_29_553# a_n1555_n1061# 0.29fF
C967 a_n149_553# a_n1555_n1061# 0.29fF
C968 a_n327_553# a_n1555_n1061# 0.29fF
C969 a_n505_553# a_n1555_n1061# 0.29fF
C970 a_n683_553# a_n1555_n1061# 0.29fF
C971 a_n861_553# a_n1555_n1061# 0.29fF
C972 a_n1039_553# a_n1555_n1061# 0.30fF
C973 a_n1217_553# a_n1555_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EL6FQZ a_n1008_n140# a_1306_n140# a_n652_n140# a_652_n194#
+ a_n1662_n194# a_772_n140# a_n1720_n140# a_n60_n194# a_2076_n194# a_1008_n194# a_2196_n140#
+ a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194# a_594_n140# a_n1542_n140#
+ a_1720_n194# a_1840_n140# a_n238_n194# a_n296_n140# a_n1898_n140# a_296_n194# a_2018_n140#
+ a_60_n140# a_n1306_n194# a_n1364_n140# a_1542_n194# a_416_n140# a_n950_n194# a_n2432_n140#
+ a_1662_n140# a_1898_n194# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194# a_238_n140#
+ a_n1186_n140# a_n2254_n140# a_1364_n194# a_n772_n194# a_1484_n140# a_n830_n140#
+ a_830_n194# a_n1840_n194# a_950_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2254_n194# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2254_n140# a_n2432_n140# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1542_n140# a_n1720_n140# 0.06fF
C1 a_n60_n194# a_474_n194# 0.02fF
C2 a_594_n140# a_1662_n140# 0.01fF
C3 a_1186_n194# a_2254_n194# 0.01fF
C4 a_830_n194# a_296_n194# 0.02fF
C5 a_1364_n194# a_474_n194# 0.01fF
C6 a_830_n194# a_n772_n194# 0.01fF
C7 a_1898_n194# a_1542_n194# 0.03fF
C8 a_n1128_n194# a_118_n194# 0.01fF
C9 a_n1128_n194# a_n1484_n194# 0.03fF
C10 a_n1662_n194# a_n950_n194# 0.01fF
C11 a_n416_n194# a_1186_n194# 0.01fF
C12 a_1484_n140# a_772_n140# 0.01fF
C13 a_594_n140# a_n830_n140# 0.01fF
C14 a_n2018_n194# a_n416_n194# 0.01fF
C15 a_n60_n194# a_652_n194# 0.01fF
C16 a_n238_n194# a_n1662_n194# 0.01fF
C17 a_n1306_n194# a_n2018_n194# 0.01fF
C18 a_416_n140# a_n118_n140# 0.02fF
C19 a_n594_n194# a_n2018_n194# 0.01fF
C20 a_1306_n140# a_1840_n140# 0.02fF
C21 a_1364_n194# a_652_n194# 0.01fF
C22 a_n652_n140# a_n474_n140# 0.06fF
C23 a_1128_n140# a_1840_n140# 0.01fF
C24 a_1128_n140# a_1306_n140# 0.06fF
C25 a_n1720_n140# a_n2254_n140# 0.02fF
C26 a_n1662_n194# a_n2432_n140# 0.01fF
C27 a_1484_n140# a_2254_n194# 0.01fF
C28 a_n296_n140# a_n474_n140# 0.06fF
C29 a_n2196_n194# a_n1484_n194# 0.01fF
C30 a_n60_n194# a_n950_n194# 0.01fF
C31 a_1720_n194# a_118_n194# 0.01fF
C32 a_n830_n140# a_n118_n140# 0.01fF
C33 a_n474_n140# a_n1008_n140# 0.02fF
C34 a_n60_n194# a_n238_n194# 0.10fF
C35 a_1484_n140# a_594_n140# 0.01fF
C36 a_474_n194# a_652_n194# 0.10fF
C37 a_n830_n140# a_n1720_n140# 0.01fF
C38 a_n474_n140# a_n1364_n140# 0.01fF
C39 a_1008_n194# a_2076_n194# 0.01fF
C40 a_772_n140# a_n474_n140# 0.01fF
C41 a_1720_n194# a_1008_n194# 0.01fF
C42 a_n238_n194# a_1364_n194# 0.01fF
C43 a_n1542_n140# a_n1898_n140# 0.03fF
C44 a_296_n194# a_1186_n194# 0.01fF
C45 a_950_n140# a_60_n140# 0.01fF
C46 a_830_n194# a_2076_n194# 0.01fF
C47 a_n2018_n194# a_n772_n194# 0.01fF
C48 a_830_n194# a_1720_n194# 0.01fF
C49 a_n1662_n194# a_n416_n194# 0.01fF
C50 a_n1306_n194# a_n1662_n194# 0.03fF
C51 a_n594_n194# a_n1662_n194# 0.01fF
C52 a_n1186_n140# a_n652_n140# 0.02fF
C53 a_n1542_n140# a_60_n140# 0.01fF
C54 a_474_n194# a_n950_n194# 0.01fF
C55 a_1484_n140# a_n118_n140# 0.01fF
C56 a_n238_n194# a_474_n194# 0.01fF
C57 a_118_n194# a_1542_n194# 0.01fF
C58 a_n296_n140# a_1306_n140# 0.01fF
C59 a_n1186_n140# a_n296_n140# 0.01fF
C60 a_594_n140# a_n474_n140# 0.01fF
C61 a_n1128_n194# a_n2018_n194# 0.01fF
C62 a_1128_n140# a_n296_n140# 0.01fF
C63 a_1364_n194# a_2254_n194# 0.01fF
C64 a_1008_n194# a_1542_n194# 0.02fF
C65 a_772_n140# a_1840_n140# 0.01fF
C66 a_n1186_n140# a_n1008_n140# 0.06fF
C67 a_n1898_n140# a_n2254_n140# 0.03fF
C68 a_772_n140# a_1306_n140# 0.02fF
C69 a_n1186_n140# a_n1364_n140# 0.06fF
C70 a_n1186_n140# a_n2432_n140# 0.01fF
C71 a_n950_n194# a_652_n194# 0.01fF
C72 a_n60_n194# a_n416_n194# 0.03fF
C73 a_n60_n194# a_n1306_n194# 0.01fF
C74 a_772_n140# a_1128_n140# 0.03fF
C75 a_n238_n194# a_652_n194# 0.01fF
C76 a_n60_n194# a_n594_n194# 0.02fF
C77 a_416_n140# a_60_n140# 0.03fF
C78 a_830_n194# a_1542_n194# 0.01fF
C79 a_2254_n194# a_1840_n140# 0.02fF
C80 a_n1662_n194# a_n772_n194# 0.01fF
C81 a_n1898_n140# a_n830_n140# 0.01fF
C82 a_2254_n194# a_1306_n140# 0.01fF
C83 a_60_n140# a_1662_n140# 0.01fF
C84 a_n1542_n140# a_n2076_n140# 0.02fF
C85 a_n474_n140# a_n118_n140# 0.03fF
C86 a_n2196_n194# a_n2018_n194# 0.10fF
C87 a_1128_n140# a_2254_n194# 0.01fF
C88 a_950_n140# a_238_n140# 0.01fF
C89 a_2076_n194# a_1186_n194# 0.01fF
C90 a_n1720_n140# a_n474_n140# 0.01fF
C91 a_1898_n194# a_1008_n194# 0.01fF
C92 a_1720_n194# a_1186_n194# 0.02fF
C93 a_594_n140# a_1840_n140# 0.01fF
C94 a_n238_n194# a_n950_n194# 0.01fF
C95 a_594_n140# a_1306_n140# 0.01fF
C96 a_n652_n140# a_n296_n140# 0.03fF
C97 a_474_n194# a_n416_n194# 0.01fF
C98 a_60_n140# a_n830_n140# 0.01fF
C99 a_1128_n140# a_594_n140# 0.02fF
C100 a_830_n194# a_1898_n194# 0.01fF
C101 a_2254_n194# a_652_n194# 0.00fF
C102 a_n594_n194# a_474_n194# 0.01fF
C103 a_n652_n140# a_n1008_n140# 0.03fF
C104 a_n1128_n194# a_n1662_n194# 0.02fF
C105 a_n652_n140# a_n1364_n140# 0.01fF
C106 a_772_n140# a_n652_n140# 0.01fF
C107 a_n60_n194# a_296_n194# 0.03fF
C108 a_n60_n194# a_n772_n194# 0.01fF
C109 a_n1840_n194# a_n1484_n194# 0.03fF
C110 a_n2432_n140# a_n950_n194# 0.00fF
C111 a_296_n194# a_1364_n194# 0.01fF
C112 a_n416_n194# a_652_n194# 0.01fF
C113 a_n296_n140# a_n1008_n140# 0.01fF
C114 a_n2076_n140# a_n2254_n140# 0.06fF
C115 a_n594_n194# a_652_n194# 0.01fF
C116 a_n296_n140# a_n1364_n140# 0.01fF
C117 a_772_n140# a_n296_n140# 0.01fF
C118 a_n1364_n140# a_n1008_n140# 0.03fF
C119 a_1306_n140# a_n118_n140# 0.01fF
C120 a_n2432_n140# a_n1008_n140# 0.01fF
C121 a_416_n140# a_238_n140# 0.06fF
C122 a_1186_n194# a_1542_n194# 0.03fF
C123 a_n1186_n140# a_n118_n140# 0.01fF
C124 a_n2432_n140# a_n1364_n140# 0.01fF
C125 a_n1186_n140# a_n1720_n140# 0.02fF
C126 a_1128_n140# a_n118_n140# 0.01fF
C127 a_1484_n140# a_60_n140# 0.01fF
C128 a_n2196_n194# a_n1662_n194# 0.02fF
C129 a_950_n140# a_2018_n140# 0.01fF
C130 a_n1128_n194# a_n60_n194# 0.01fF
C131 a_n830_n140# a_n2076_n140# 0.01fF
C132 a_1662_n140# a_238_n140# 0.01fF
C133 a_594_n140# a_n652_n140# 0.01fF
C134 a_296_n194# a_474_n194# 0.10fF
C135 a_474_n194# a_n772_n194# 0.01fF
C136 a_n416_n194# a_n950_n194# 0.02fF
C137 a_n1306_n194# a_n950_n194# 0.03fF
C138 a_n238_n194# a_n416_n194# 0.10fF
C139 a_n1898_n140# a_n474_n140# 0.01fF
C140 a_n594_n194# a_n950_n194# 0.03fF
C141 a_772_n140# a_2254_n194# 0.01fF
C142 a_n238_n194# a_n1306_n194# 0.01fF
C143 a_n594_n194# a_n238_n194# 0.03fF
C144 a_n830_n140# a_238_n140# 0.01fF
C145 a_594_n140# a_n296_n140# 0.01fF
C146 a_1898_n194# a_1186_n194# 0.01fF
C147 a_296_n194# a_652_n194# 0.03fF
C148 a_n1484_n194# a_118_n194# 0.01fF
C149 a_594_n140# a_n1008_n140# 0.01fF
C150 a_n772_n194# a_652_n194# 0.01fF
C151 a_n1306_n194# a_n2432_n140# 0.01fF
C152 a_118_n194# a_1008_n194# 0.01fF
C153 a_772_n140# a_594_n140# 0.06fF
C154 a_n1128_n194# a_474_n194# 0.01fF
C155 a_60_n140# a_n474_n140# 0.02fF
C156 a_2018_n140# a_2196_n140# 0.06fF
C157 a_n652_n140# a_n118_n140# 0.02fF
C158 a_1364_n194# a_2076_n194# 0.01fF
C159 a_n652_n140# a_n1720_n140# 0.01fF
C160 a_416_n140# a_2018_n140# 0.01fF
C161 a_1720_n194# a_1364_n194# 0.03fF
C162 a_830_n194# a_118_n194# 0.01fF
C163 a_830_n194# a_1008_n194# 0.10fF
C164 a_n296_n140# a_n118_n140# 0.06fF
C165 a_n1840_n194# a_n2018_n194# 0.10fF
C166 a_296_n194# a_n950_n194# 0.01fF
C167 a_1662_n140# a_2018_n140# 0.03fF
C168 a_1484_n140# a_238_n140# 0.01fF
C169 a_n296_n140# a_n1720_n140# 0.01fF
C170 a_n950_n194# a_n772_n194# 0.10fF
C171 a_296_n194# a_n238_n194# 0.02fF
C172 a_n118_n140# a_n1008_n140# 0.01fF
C173 a_n1186_n140# a_n1898_n140# 0.01fF
C174 a_n238_n194# a_n772_n194# 0.02fF
C175 a_n1364_n140# a_n118_n140# 0.01fF
C176 a_772_n140# a_n118_n140# 0.01fF
C177 a_n1720_n140# a_n1008_n140# 0.01fF
C178 a_n1306_n194# a_n416_n194# 0.01fF
C179 a_n1720_n140# a_n2432_n140# 0.01fF
C180 a_n1720_n140# a_n1364_n140# 0.03fF
C181 a_n594_n194# a_n416_n194# 0.10fF
C182 a_474_n194# a_2076_n194# 0.01fF
C183 a_n594_n194# a_n1306_n194# 0.01fF
C184 a_1720_n194# a_474_n194# 0.01fF
C185 a_950_n140# a_2196_n140# 0.01fF
C186 a_n474_n140# a_n2076_n140# 0.01fF
C187 a_950_n140# a_416_n140# 0.02fF
C188 a_n60_n194# a_1542_n194# 0.01fF
C189 a_n2432_n140# a_n772_n194# 0.00fF
C190 a_60_n140# a_1306_n140# 0.01fF
C191 a_n1186_n140# a_60_n140# 0.01fF
C192 a_n1128_n194# a_n950_n194# 0.10fF
C193 a_1364_n194# a_1542_n194# 0.10fF
C194 a_1128_n140# a_60_n140# 0.01fF
C195 a_n1128_n194# a_n238_n194# 0.01fF
C196 a_2076_n194# a_652_n194# 0.01fF
C197 a_1720_n194# a_652_n194# 0.01fF
C198 a_950_n140# a_1662_n140# 0.01fF
C199 a_n474_n140# a_238_n140# 0.01fF
C200 a_594_n140# a_n118_n140# 0.01fF
C201 a_n1542_n140# a_n2254_n140# 0.01fF
C202 a_118_n194# a_1186_n194# 0.01fF
C203 a_n1128_n194# a_n2432_n140# 0.00fF
C204 a_n1840_n194# a_n1662_n194# 0.10fF
C205 a_n1484_n194# a_n2018_n194# 0.02fF
C206 a_1484_n140# a_2018_n140# 0.02fF
C207 a_n652_n140# a_n1898_n140# 0.01fF
C208 a_296_n194# a_n416_n194# 0.01fF
C209 a_1008_n194# a_1186_n194# 0.10fF
C210 a_296_n194# a_n1306_n194# 0.01fF
C211 a_474_n194# a_1542_n194# 0.01fF
C212 a_n416_n194# a_n772_n194# 0.03fF
C213 a_n1306_n194# a_n772_n194# 0.02fF
C214 a_n2196_n194# a_n950_n194# 0.01fF
C215 a_n594_n194# a_296_n194# 0.01fF
C216 a_1364_n194# a_1898_n194# 0.02fF
C217 a_n594_n194# a_n772_n194# 0.10fF
C218 a_n1542_n140# a_n830_n140# 0.01fF
C219 a_n296_n140# a_n1898_n140# 0.01fF
C220 a_n1186_n140# a_n2076_n140# 0.01fF
C221 a_830_n194# a_1186_n194# 0.03fF
C222 a_n652_n140# a_60_n140# 0.01fF
C223 a_n1898_n140# a_n1008_n140# 0.01fF
C224 a_1662_n140# a_2196_n140# 0.02fF
C225 a_652_n194# a_1542_n194# 0.01fF
C226 a_n1898_n140# a_n1364_n140# 0.02fF
C227 a_n1898_n140# a_n2432_n140# 0.02fF
C228 a_416_n140# a_1662_n140# 0.01fF
C229 a_n2196_n194# a_n2432_n140# 0.06fF
C230 a_n1720_n140# a_n118_n140# 0.01fF
C231 a_238_n140# a_1840_n140# 0.01fF
C232 a_n1128_n194# a_n416_n194# 0.01fF
C233 a_n1128_n194# a_n1306_n194# 0.10fF
C234 a_1306_n140# a_238_n140# 0.01fF
C235 a_n1186_n140# a_238_n140# 0.01fF
C236 a_n296_n140# a_60_n140# 0.03fF
C237 a_1484_n140# a_950_n140# 0.02fF
C238 a_n1128_n194# a_n594_n194# 0.02fF
C239 a_474_n194# a_1898_n194# 0.01fF
C240 a_1128_n140# a_238_n140# 0.01fF
C241 a_60_n140# a_n1008_n140# 0.01fF
C242 a_416_n140# a_n830_n140# 0.01fF
C243 a_60_n140# a_n1364_n140# 0.01fF
C244 a_772_n140# a_60_n140# 0.01fF
C245 a_n1484_n194# a_n1662_n194# 0.10fF
C246 a_296_n194# a_n772_n194# 0.01fF
C247 a_2076_n194# a_2254_n194# 0.06fF
C248 a_n830_n140# a_n2254_n140# 0.01fF
C249 a_1720_n194# a_2254_n194# 0.01fF
C250 a_1898_n194# a_652_n194# 0.01fF
C251 a_n652_n140# a_n2076_n140# 0.01fF
C252 a_n2196_n194# a_n1306_n194# 0.01fF
C253 a_n594_n194# a_n2196_n194# 0.01fF
C254 a_950_n140# a_n474_n140# 0.01fF
C255 a_1484_n140# a_2196_n140# 0.01fF
C256 a_n1128_n194# a_296_n194# 0.01fF
C257 a_1484_n140# a_416_n140# 0.01fF
C258 a_n1128_n194# a_n772_n194# 0.03fF
C259 a_n652_n140# a_238_n140# 0.01fF
C260 a_2018_n140# a_1840_n140# 0.06fF
C261 a_594_n140# a_60_n140# 0.02fF
C262 a_n60_n194# a_118_n194# 0.10fF
C263 a_n60_n194# a_n1484_n194# 0.01fF
C264 a_2018_n140# a_1306_n140# 0.01fF
C265 a_n2076_n140# a_n1008_n140# 0.01fF
C266 a_n2076_n140# a_n1364_n140# 0.01fF
C267 a_n2432_n140# a_n2076_n140# 0.03fF
C268 a_1128_n140# a_2018_n140# 0.01fF
C269 a_n1542_n140# a_n474_n140# 0.01fF
C270 a_1364_n194# a_118_n194# 0.01fF
C271 a_n60_n194# a_1008_n194# 0.01fF
C272 a_1484_n140# a_1662_n140# 0.06fF
C273 a_2254_n194# a_1542_n194# 0.01fF
C274 a_1364_n194# a_1008_n194# 0.03fF
C275 a_n296_n140# a_238_n140# 0.02fF
C276 a_n1898_n140# a_n1720_n140# 0.06fF
C277 a_238_n140# a_n1008_n140# 0.01fF
C278 a_830_n194# a_n60_n194# 0.01fF
C279 a_n1364_n140# a_238_n140# 0.01fF
C280 a_772_n140# a_238_n140# 0.02fF
C281 a_830_n194# a_1364_n194# 0.02fF
C282 a_n2196_n194# a_n772_n194# 0.01fF
C283 a_60_n140# a_n118_n140# 0.06fF
C284 a_1720_n194# a_296_n194# 0.01fF
C285 a_n1840_n194# a_n950_n194# 0.01fF
C286 a_950_n140# a_1840_n140# 0.01fF
C287 a_474_n194# a_118_n194# 0.03fF
C288 a_416_n140# a_n474_n140# 0.01fF
C289 a_950_n140# a_1306_n140# 0.03fF
C290 a_n238_n194# a_n1840_n194# 0.01fF
C291 a_474_n194# a_1008_n194# 0.02fF
C292 a_950_n140# a_1128_n140# 0.06fF
C293 a_1898_n194# a_2254_n194# 0.02fF
C294 a_n2018_n194# a_n1662_n194# 0.03fF
C295 a_n1186_n140# a_n1542_n140# 0.03fF
C296 a_n1840_n194# a_n2432_n140# 0.01fF
C297 a_n1128_n194# a_n2196_n194# 0.01fF
C298 a_118_n194# a_652_n194# 0.02fF
C299 a_830_n194# a_474_n194# 0.03fF
C300 a_594_n140# a_238_n140# 0.03fF
C301 a_1008_n194# a_652_n194# 0.03fF
C302 a_n830_n140# a_n474_n140# 0.03fF
C303 a_2196_n140# a_1840_n140# 0.03fF
C304 a_296_n194# a_1542_n194# 0.01fF
C305 a_772_n140# a_2018_n140# 0.01fF
C306 a_830_n194# a_652_n194# 0.10fF
C307 a_1306_n140# a_2196_n140# 0.01fF
C308 a_n1720_n140# a_n2076_n140# 0.03fF
C309 a_416_n140# a_1840_n140# 0.01fF
C310 a_n60_n194# a_1186_n194# 0.01fF
C311 a_1128_n140# a_2196_n140# 0.01fF
C312 a_416_n140# a_1306_n140# 0.01fF
C313 a_n1186_n140# a_416_n140# 0.01fF
C314 a_118_n194# a_n950_n194# 0.01fF
C315 a_950_n140# a_n652_n140# 0.01fF
C316 a_1128_n140# a_416_n140# 0.01fF
C317 a_n1484_n194# a_n950_n194# 0.02fF
C318 a_1364_n194# a_1186_n194# 0.10fF
C319 a_n1840_n194# a_n416_n194# 0.01fF
C320 a_n238_n194# a_118_n194# 0.03fF
C321 a_n1840_n194# a_n1306_n194# 0.02fF
C322 a_n238_n194# a_n1484_n194# 0.01fF
C323 a_1662_n140# a_1840_n140# 0.06fF
C324 a_n1186_n140# a_n2254_n140# 0.01fF
C325 a_238_n140# a_n118_n140# 0.03fF
C326 a_1662_n140# a_1306_n140# 0.03fF
C327 a_2018_n140# a_2254_n194# 0.03fF
C328 a_n594_n194# a_n1840_n194# 0.01fF
C329 a_n238_n194# a_1008_n194# 0.01fF
C330 a_1720_n194# a_2076_n194# 0.03fF
C331 a_1128_n140# a_1662_n140# 0.02fF
C332 a_n652_n140# a_n1542_n140# 0.01fF
C333 a_950_n140# a_n296_n140# 0.01fF
C334 a_296_n194# a_1898_n194# 0.01fF
C335 a_n1484_n194# a_n2432_n140# 0.01fF
C336 a_830_n194# a_n238_n194# 0.01fF
C337 a_772_n140# a_950_n140# 0.06fF
C338 a_594_n140# a_2018_n140# 0.01fF
C339 a_n1186_n140# a_n830_n140# 0.03fF
C340 a_474_n194# a_1186_n194# 0.01fF
C341 a_n1542_n140# a_n296_n140# 0.01fF
C342 a_n1542_n140# a_n1008_n140# 0.02fF
C343 a_n1542_n140# a_n1364_n140# 0.06fF
C344 a_n1542_n140# a_n2432_n140# 0.01fF
C345 a_416_n140# a_n652_n140# 0.01fF
C346 a_950_n140# a_2254_n194# 0.01fF
C347 a_1008_n194# a_2254_n194# 0.00fF
C348 a_n60_n194# a_n1662_n194# 0.01fF
C349 a_1186_n194# a_652_n194# 0.02fF
C350 a_n1840_n194# a_n772_n194# 0.01fF
C351 a_n652_n140# a_n2254_n140# 0.01fF
C352 a_2076_n194# a_1542_n194# 0.02fF
C353 a_118_n194# a_n416_n194# 0.02fF
C354 a_1720_n194# a_1542_n194# 0.10fF
C355 a_n1484_n194# a_n416_n194# 0.01fF
C356 a_n1306_n194# a_118_n194# 0.01fF
C357 a_n1484_n194# a_n1306_n194# 0.10fF
C358 a_1484_n140# a_1840_n140# 0.03fF
C359 a_416_n140# a_n296_n140# 0.01fF
C360 a_n1898_n140# a_n2076_n140# 0.06fF
C361 a_n594_n194# a_118_n194# 0.01fF
C362 a_830_n194# a_2254_n194# 0.00fF
C363 a_n416_n194# a_1008_n194# 0.01fF
C364 a_1484_n140# a_1306_n140# 0.06fF
C365 a_n594_n194# a_n1484_n194# 0.01fF
C366 a_950_n140# a_594_n140# 0.03fF
C367 a_772_n140# a_2196_n140# 0.01fF
C368 a_1484_n140# a_1128_n140# 0.03fF
C369 a_416_n140# a_n1008_n140# 0.01fF
C370 a_n594_n194# a_1008_n194# 0.01fF
C371 a_772_n140# a_416_n140# 0.03fF
C372 a_n652_n140# a_n830_n140# 0.06fF
C373 a_830_n194# a_n416_n194# 0.01fF
C374 a_n1008_n140# a_n2254_n140# 0.01fF
C375 a_n1128_n194# a_n1840_n194# 0.01fF
C376 a_n1364_n140# a_n2254_n140# 0.01fF
C377 a_n2432_n140# a_n2254_n140# 0.06fF
C378 a_830_n194# a_n594_n194# 0.01fF
C379 a_n2018_n194# a_n950_n194# 0.01fF
C380 a_772_n140# a_1662_n140# 0.01fF
C381 a_n238_n194# a_1186_n194# 0.01fF
C382 a_1898_n194# a_2076_n194# 0.10fF
C383 a_2254_n194# a_2196_n140# 0.06fF
C384 a_1720_n194# a_1898_n194# 0.10fF
C385 a_n60_n194# a_1364_n194# 0.01fF
C386 a_n296_n140# a_n830_n140# 0.02fF
C387 a_950_n140# a_n118_n140# 0.01fF
C388 a_n830_n140# a_n1008_n140# 0.06fF
C389 a_60_n140# a_238_n140# 0.06fF
C390 a_n830_n140# a_n1364_n140# 0.02fF
C391 a_772_n140# a_n830_n140# 0.01fF
C392 a_n830_n140# a_n2432_n140# 0.01fF
C393 a_n1186_n140# a_n474_n140# 0.01fF
C394 a_296_n194# a_118_n194# 0.10fF
C395 a_594_n140# a_2196_n140# 0.01fF
C396 a_1662_n140# a_2254_n194# 0.01fF
C397 a_n2018_n194# a_n2432_n140# 0.02fF
C398 a_118_n194# a_n772_n194# 0.01fF
C399 a_1128_n140# a_n474_n140# 0.01fF
C400 a_594_n140# a_416_n140# 0.06fF
C401 a_n1484_n194# a_n772_n194# 0.01fF
C402 a_296_n194# a_1008_n194# 0.01fF
C403 a_n1542_n140# a_n118_n140# 0.01fF
C404 a_n2196_n194# a_n1840_n194# 0.03fF
C405 a_2196_n140# VSUBS 0.01fF
C406 a_2018_n140# VSUBS 0.01fF
C407 a_1840_n140# VSUBS 0.02fF
C408 a_1662_n140# VSUBS 0.02fF
C409 a_1484_n140# VSUBS 0.02fF
C410 a_1306_n140# VSUBS 0.02fF
C411 a_1128_n140# VSUBS 0.02fF
C412 a_950_n140# VSUBS 0.02fF
C413 a_772_n140# VSUBS 0.02fF
C414 a_594_n140# VSUBS 0.02fF
C415 a_416_n140# VSUBS 0.02fF
C416 a_238_n140# VSUBS 0.02fF
C417 a_60_n140# VSUBS 0.02fF
C418 a_n118_n140# VSUBS 0.02fF
C419 a_n296_n140# VSUBS 0.02fF
C420 a_n474_n140# VSUBS 0.02fF
C421 a_n652_n140# VSUBS 0.02fF
C422 a_n830_n140# VSUBS 0.02fF
C423 a_n1008_n140# VSUBS 0.02fF
C424 a_n1186_n140# VSUBS 0.02fF
C425 a_n1364_n140# VSUBS 0.02fF
C426 a_n1542_n140# VSUBS 0.02fF
C427 a_n1720_n140# VSUBS 0.02fF
C428 a_n1898_n140# VSUBS 0.02fF
C429 a_n2076_n140# VSUBS 0.02fF
C430 a_n2254_n140# VSUBS 0.02fF
C431 a_2254_n194# VSUBS 0.31fF
C432 a_2076_n194# VSUBS 0.19fF
C433 a_1898_n194# VSUBS 0.20fF
C434 a_1720_n194# VSUBS 0.21fF
C435 a_1542_n194# VSUBS 0.22fF
C436 a_1364_n194# VSUBS 0.23fF
C437 a_1186_n194# VSUBS 0.23fF
C438 a_1008_n194# VSUBS 0.24fF
C439 a_830_n194# VSUBS 0.24fF
C440 a_652_n194# VSUBS 0.24fF
C441 a_474_n194# VSUBS 0.24fF
C442 a_296_n194# VSUBS 0.24fF
C443 a_118_n194# VSUBS 0.24fF
C444 a_n60_n194# VSUBS 0.24fF
C445 a_n238_n194# VSUBS 0.24fF
C446 a_n416_n194# VSUBS 0.24fF
C447 a_n594_n194# VSUBS 0.24fF
C448 a_n772_n194# VSUBS 0.24fF
C449 a_n950_n194# VSUBS 0.24fF
C450 a_n1128_n194# VSUBS 0.24fF
C451 a_n1306_n194# VSUBS 0.24fF
C452 a_n1484_n194# VSUBS 0.24fF
C453 a_n1662_n194# VSUBS 0.24fF
C454 a_n1840_n194# VSUBS 0.24fF
C455 a_n2018_n194# VSUBS 0.24fF
C456 a_n2196_n194# VSUBS 0.24fF
C457 a_n2432_n140# VSUBS 0.36fF
.ends

.subckt bias_circuit bias_c bias_e i_bias VDD m1_7347_1428# m1_7639_1420# li_3433_399#
+ bias_a m1_7169_923# m1_7461_921# m1_7347_423# m1_7639_427# bias_b VSS m1_1243_5997#
+ m1_3443_5997# m1_3551_3596# m1_5643_5997# bias_d
Xsky130_fd_pr__nfet_01v8_6RUDQZ_0 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_1 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_2 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_SD55Q9_0 m1_7347_1428# m1_7639_1420# bias_e m1_7055_1417#
+ bias_e m1_6763_422# bias_e m1_6471_422# bias_e VSS VSS VSS m1_7639_427# m1_7347_423#
+ m1_7055_433# bias_e bias_e bias_e m1_6763_422# m1_6471_422# m1_7169_923# bias_e
+ m1_7461_921# bias_e bias_e m1_7639_427# m1_7347_423# m1_6877_922# m1_7055_433# VSS
+ bias_e VSS VSS bias_e bias_e bias_e m1_6877_922# m1_6585_923# VSS bias_e m1_6763_1422#
+ m1_6293_922# bias_e m1_6471_1426# m1_7347_1428# bias_e bias_e m1_7639_1420# m1_7169_923#
+ m1_7055_1417# bias_e bias_e m1_7461_921# bias_e bias_e bias_e m1_6585_923# bias_e
+ m1_6293_922# m1_6763_1422# bias_e m1_6471_1426# VSS sky130_fd_pr__nfet_01v8_SD55Q9
Xsky130_fd_pr__nfet_01v8_6RUDQZ_3 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_EZNTQN_0 bias_c VSS VSS i_bias i_bias i_bias i_bias VSS VSS
+ bias_c VSS VSS i_bias VSS bias_c i_bias i_bias i_bias i_bias VSS i_bias i_bias bias_c
+ i_bias VSS VSS i_bias i_bias i_bias bias_c VSS VSS i_bias bias_c VSS i_bias i_bias
+ VSS i_bias i_bias i_bias i_bias i_bias VSS i_bias i_bias i_bias i_bias i_bias i_bias
+ i_bias bias_c i_bias VSS i_bias i_bias bias_c i_bias i_bias i_bias i_bias VSS i_bias
+ VSS i_bias VSS VSS i_bias i_bias bias_c i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ sky130_fd_pr__nfet_01v8_EZNTQN
Xsky130_fd_pr__pfet_01v8_JJWXCM_0 bias_b bias_c m1_1243_5997# m1_1243_5997# bias_b
+ bias_c VDD VDD bias_c bias_b bias_c VDD bias_c m1_1243_5997# bias_c bias_b VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_1 m1_3551_3596# bias_c m1_3443_5997# m1_3443_5997#
+ m1_3551_3596# bias_c VDD VDD bias_c m1_3551_3596# bias_c VDD bias_c m1_3443_5997#
+ bias_c m1_3551_3596# VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_2 bias_e bias_c m1_5643_5997# m1_5643_5997# bias_e
+ bias_c VDD VDD bias_c bias_e bias_c VDD bias_c m1_5643_5997# bias_c bias_e VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__nfet_01v8_LJREPQ_0 m1_3551_3596# bias_d VSS bias_a bias_d m1_3551_3596#
+ VSS VSS sky130_fd_pr__nfet_01v8_LJREPQ
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_0 m1_1243_5997# bias_b VDD VDD m1_1243_5997# bias_b
+ VDD VDD bias_b m1_1243_5997# bias_b VDD bias_b VDD bias_b m1_1243_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_2 m1_5643_5997# bias_b VDD VDD m1_5643_5997# bias_b
+ VDD VDD bias_b m1_5643_5997# bias_b VDD bias_b VDD bias_b m1_5643_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_1 m1_3443_5997# bias_b VDD VDD m1_3443_5997# bias_b
+ VDD VDD bias_b m1_3443_5997# bias_b VDD bias_b VDD bias_b m1_3443_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__nfet_01v8_lvt_28TRYY_0 bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b VSS bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_c bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_c bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_b bias_c bias_b bias_b bias_b
+ bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_c
+ bias_c bias_b bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c
+ bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_c bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b sky130_fd_pr__nfet_01v8_lvt_28TRYY
Xsky130_fd_pr__nfet_01v8_EL6FQZ_0 bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d VSS m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
Xsky130_fd_pr__nfet_01v8_EL6FQZ_1 bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d VSS m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
C0 bias_e VDD 0.26fF
C1 bias_e m1_7347_423# 0.26fF
C2 m1_6763_1422# m1_7639_1420# 0.01fF
C3 bias_a m1_7461_921# 0.00fF
C4 bias_d bias_e 0.26fF
C5 m1_6763_422# m1_7055_433# 0.03fF
C6 bias_c m1_5643_5997# 0.44fF
C7 m1_7055_1417# bias_e 0.33fF
C8 bias_e m1_6763_1422# 0.33fF
C9 bias_a m1_7055_433# 0.01fF
C10 bias_d li_3433_399# 5.36fF
C11 m1_7461_921# m1_6585_923# 0.01fF
C12 m1_7169_923# m1_6877_922# 0.03fF
C13 bias_a i_bias 0.02fF
C14 m1_6471_1426# m1_7347_1428# 0.01fF
C15 bias_a m1_7639_1420# 0.00fF
C16 bias_c bias_b 22.44fF
C17 m1_7055_433# m1_7639_427# 0.01fF
C18 VDD m1_3443_5997# 0.84fF
C19 bias_c i_bias 5.62fF
C20 m1_7639_427# m1_7639_1420# -0.00fF
C21 m1_1243_5997# m1_3551_3596# 0.03fF
C22 bias_d m1_6293_922# 0.00fF
C23 bias_e m1_6763_422# 0.26fF
C24 m1_7347_423# m1_6471_422# 0.01fF
C25 bias_d m1_3443_5997# 0.03fF
C26 bias_e bias_a 0.24fF
C27 bias_e bias_c 0.65fF
C28 bias_e m1_7639_427# 0.18fF
C29 bias_a li_3433_399# 7.53fF
C30 bias_e m1_6585_923# 0.22fF
C31 bias_a m1_6293_922# 0.01fF
C32 li_3433_399# m1_6585_923# 0.01fF
C33 VDD m1_3551_3596# 0.64fF
C34 m1_6763_422# m1_6471_422# 0.03fF
C35 bias_c m1_3443_5997# 0.44fF
C36 m1_5643_5997# bias_b 0.63fF
C37 m1_6293_922# m1_6585_923# 0.03fF
C38 m1_7347_423# m1_7347_1428# -0.00fF
C39 bias_a m1_6471_422# 0.01fF
C40 bias_d m1_3551_3596# 18.83fF
C41 m1_7639_427# m1_6471_422# 0.01fF
C42 bias_d m1_6471_1426# 0.01fF
C43 bias_d m1_7347_1428# 0.00fF
C44 VDD m1_1243_5997# 1.50fF
C45 i_bias bias_b 0.60fF
C46 m1_7055_1417# m1_6471_1426# 0.01fF
C47 m1_7055_1417# m1_7347_1428# 0.03fF
C48 m1_6763_1422# m1_6471_1426# 0.03fF
C49 m1_6763_1422# m1_7347_1428# 0.01fF
C50 bias_e m1_5643_5997# 0.71fF
C51 bias_e m1_7461_921# 0.21fF
C52 bias_a m1_7169_923# 0.00fF
C53 bias_e bias_b 0.07fF
C54 bias_e m1_7055_433# 0.26fF
C55 bias_a m1_3551_3596# 0.26fF
C56 bias_e m1_7639_1420# 0.18fF
C57 bias_c m1_3551_3596# 2.13fF
C58 bias_a m1_6471_1426# 0.01fF
C59 m1_7461_921# m1_6293_922# 0.01fF
C60 m1_7169_923# m1_6585_923# 0.01fF
C61 bias_a m1_7347_1428# 0.00fF
C62 li_3433_399# i_bias 0.03fF
C63 m1_3443_5997# m1_5643_5997# 0.11fF
C64 bias_a m1_6877_922# 0.00fF
C65 bias_c m1_1243_5997# 0.52fF
C66 m1_3443_5997# bias_b 0.65fF
C67 bias_d VDD 0.07fF
C68 bias_e li_3433_399# 0.02fF
C69 m1_6585_923# m1_6877_922# 0.03fF
C70 m1_7055_433# m1_6471_422# 0.01fF
C71 bias_e m1_6293_922# 0.18fF
C72 bias_d m1_7055_1417# 0.00fF
C73 m1_7169_923# m1_7461_921# 0.03fF
C74 bias_e m1_3443_5997# 0.02fF
C75 bias_d m1_6763_1422# 0.00fF
C76 li_3433_399# m1_6293_922# 0.02fF
C77 m1_6763_422# m1_7347_423# 0.01fF
C78 m1_7055_1417# m1_6763_1422# 0.03fF
C79 m1_5643_5997# m1_3551_3596# 0.08fF
C80 bias_e m1_6471_422# 0.25fF
C81 bias_a m1_7347_423# 0.01fF
C82 bias_c VDD 4.90fF
C83 m1_7347_423# m1_7639_427# 0.03fF
C84 li_3433_399# m1_6471_422# 0.01fF
C85 bias_b m1_3551_3596# 0.71fF
C86 m1_6763_1422# m1_6763_422# -0.00fF
C87 bias_d bias_a 7.33fF
C88 m1_7055_1417# bias_a 0.00fF
C89 m1_7461_921# m1_6877_922# 0.01fF
C90 bias_d bias_c 0.90fF
C91 m1_6471_1426# m1_7639_1420# 0.01fF
C92 m1_7347_1428# m1_7639_1420# 0.03fF
C93 m1_6763_1422# bias_a 0.00fF
C94 bias_e m1_7169_923# 0.22fF
C95 bias_d m1_6585_923# 0.00fF
C96 m1_1243_5997# bias_b 0.77fF
C97 bias_e m1_3551_3596# 0.76fF
C98 bias_a m1_6763_422# 0.01fF
C99 bias_e m1_6471_1426# 0.34fF
C100 bias_e m1_7347_1428# 0.32fF
C101 li_3433_399# m1_3551_3596# 0.03fF
C102 m1_6763_422# m1_7639_427# 0.01fF
C103 m1_7169_923# m1_6293_922# 0.01fF
C104 li_3433_399# m1_6471_1426# 0.01fF
C105 bias_a bias_c 0.02fF
C106 bias_a m1_7639_427# 0.01fF
C107 bias_e m1_6877_922# 0.22fF
C108 VDD m1_5643_5997# 1.16fF
C109 bias_a m1_6585_923# 0.00fF
C110 m1_3443_5997# m1_3551_3596# 0.98fF
C111 VDD bias_b 8.29fF
C112 bias_d m1_5643_5997# 0.03fF
C113 m1_7055_433# m1_7347_423# 0.03fF
C114 m1_6293_922# m1_6877_922# 0.01fF
C115 m1_6471_1426# m1_6471_422# -0.00fF
C116 m1_1243_5997# m1_3443_5997# 0.07fF
C117 bias_d bias_b 0.26fF
C118 bias_d i_bias 0.00fF
C119 bias_d m1_7639_1420# 0.00fF
C120 m1_7055_1417# m1_7055_433# -0.00fF
C121 m1_7055_1417# m1_7639_1420# 0.01fF
C122 m1_3551_3596# VSS -340.53fF
C123 bias_b VSS -284.38fF
C124 m1_5643_5997# VSS 38.06fF
C125 m1_3443_5997# VSS 35.86fF
C126 m1_1243_5997# VSS 25.05fF
C127 VDD VSS 131.75fF
C128 i_bias VSS -59.70fF
C129 bias_c VSS -50.79fF
C130 m1_7639_427# VSS 0.32fF
C131 m1_7347_423# VSS 0.27fF
C132 m1_7461_921# VSS 0.22fF
C133 m1_7169_923# VSS 0.20fF
C134 m1_7055_433# VSS 0.28fF
C135 m1_6763_422# VSS 0.35fF
C136 m1_6471_422# VSS 0.38fF
C137 m1_7639_1420# VSS 0.31fF
C138 m1_7347_1428# VSS 0.20fF
C139 m1_6877_922# VSS 0.21fF
C140 m1_6585_923# VSS 0.29fF
C141 m1_6293_922# VSS 0.32fF
C142 m1_7055_1417# VSS 0.20fF
C143 m1_6763_1422# VSS 0.29fF
C144 m1_6471_1426# VSS 0.30fF
C145 bias_e VSS 7.90fF
C146 bias_d VSS -76.91fF
C147 li_3433_399# VSS 5.57fF
C148 bias_a VSS -48.09fF
.ends

.subckt sky130_fd_pr__pfet_01v8_YVTMSC a_n207_n140# a_29_n205# a_327_n140# a_n683_n205#
+ a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_n505_n205# a_n741_n140# a_563_n205#
+ a_861_n140# a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_683_n140# w_n1133_n241#
+ a_n919_n140# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_861_n140# a_741_n205# a_683_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n205# a_n385_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n741_n140# a_n861_n205# a_n919_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_683_n140# a_563_n205# a_505_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_919_n205# a_919_n205# a_861_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_n29_n140# a_n149_n205# a_n207_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n563_n140# a_n683_n205# a_n741_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_n919_n140# a_n1097_n140# a_n1097_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_505_n140# a_385_n205# a_327_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_861_n140# a_n741_n140# 0.01fF
C1 w_n1133_n241# a_919_n205# 0.28fF
C2 a_n1097_n140# a_n505_n205# 0.01fF
C3 a_n385_n140# a_327_n140# 0.01fF
C4 a_n385_n140# a_505_n140# 0.01fF
C5 a_149_n140# a_n385_n140# 0.02fF
C6 a_919_n205# a_29_n205# 0.01fF
C7 w_n1133_n241# a_n385_n140# 0.02fF
C8 a_n861_n205# a_207_n205# 0.01fF
C9 a_n1097_n140# a_n327_n205# 0.01fF
C10 a_n1097_n140# a_n683_n205# 0.02fF
C11 a_n1097_n140# a_327_n140# 0.01fF
C12 a_n1097_n140# a_505_n140# 0.01fF
C13 a_207_n205# a_385_n205# 0.10fF
C14 a_n1097_n140# a_149_n140# 0.01fF
C15 a_n861_n205# a_385_n205# 0.01fF
C16 a_207_n205# a_563_n205# 0.03fF
C17 a_n861_n205# a_563_n205# 0.01fF
C18 a_683_n140# a_n919_n140# 0.01fF
C19 w_n1133_n241# a_n1097_n140# 0.33fF
C20 a_385_n205# a_563_n205# 0.10fF
C21 a_n207_n140# a_n919_n140# 0.01fF
C22 a_n1097_n140# a_29_n205# 0.01fF
C23 a_683_n140# a_n563_n140# 0.01fF
C24 a_207_n205# a_n505_n205# 0.01fF
C25 a_n861_n205# a_n505_n205# 0.03fF
C26 a_861_n140# a_327_n140# 0.02fF
C27 a_861_n140# a_505_n140# 0.03fF
C28 a_683_n140# a_n29_n140# 0.01fF
C29 a_741_n205# a_207_n205# 0.02fF
C30 a_861_n140# a_149_n140# 0.01fF
C31 a_741_n205# a_n861_n205# 0.01fF
C32 a_n207_n140# a_n563_n140# 0.03fF
C33 a_n505_n205# a_385_n205# 0.01fF
C34 a_n505_n205# a_563_n205# 0.01fF
C35 w_n1133_n241# a_861_n140# 0.01fF
C36 a_741_n205# a_385_n205# 0.03fF
C37 a_207_n205# a_n327_n205# 0.02fF
C38 a_207_n205# a_n683_n205# 0.01fF
C39 a_n207_n140# a_n29_n140# 0.06fF
C40 a_n861_n205# a_n327_n205# 0.02fF
C41 a_n861_n205# a_n683_n205# 0.10fF
C42 a_741_n205# a_563_n205# 0.10fF
C43 a_327_n140# a_n741_n140# 0.01fF
C44 a_n741_n140# a_505_n140# 0.01fF
C45 a_149_n140# a_n741_n140# 0.01fF
C46 a_919_n205# a_n563_n140# 0.01fF
C47 a_n919_n140# a_n385_n140# 0.02fF
C48 a_n327_n205# a_385_n205# 0.01fF
C49 a_385_n205# a_n683_n205# 0.01fF
C50 a_n327_n205# a_563_n205# 0.01fF
C51 a_n683_n205# a_563_n205# 0.01fF
C52 w_n1133_n241# a_n741_n140# 0.02fF
C53 a_919_n205# a_n29_n140# 0.01fF
C54 w_n1133_n241# a_207_n205# 0.17fF
C55 w_n1133_n241# a_n861_n205# 0.20fF
C56 a_741_n205# a_n505_n205# 0.01fF
C57 a_n385_n140# a_n563_n140# 0.06fF
C58 a_919_n205# a_n149_n205# 0.01fF
C59 a_207_n205# a_29_n205# 0.10fF
C60 w_n1133_n241# a_385_n205# 0.16fF
C61 a_n861_n205# a_29_n205# 0.01fF
C62 a_n1097_n140# a_n919_n140# 0.06fF
C63 w_n1133_n241# a_563_n205# 0.15fF
C64 a_n385_n140# a_n29_n140# 0.03fF
C65 a_n505_n205# a_n327_n205# 0.10fF
C66 a_n505_n205# a_n683_n205# 0.10fF
C67 a_385_n205# a_29_n205# 0.03fF
C68 a_741_n205# a_n327_n205# 0.01fF
C69 a_741_n205# a_n683_n205# 0.01fF
C70 a_29_n205# a_563_n205# 0.02fF
C71 a_n1097_n140# a_n563_n140# 0.02fF
C72 a_n327_n205# a_n683_n205# 0.03fF
C73 w_n1133_n241# a_n505_n205# 0.20fF
C74 a_n1097_n140# a_n29_n140# 0.01fF
C75 a_n207_n140# a_683_n140# 0.01fF
C76 w_n1133_n241# a_741_n205# 0.14fF
C77 a_n505_n205# a_29_n205# 0.02fF
C78 a_n1097_n140# a_n149_n205# 0.01fF
C79 a_327_n140# a_505_n140# 0.06fF
C80 a_149_n140# a_327_n140# 0.06fF
C81 a_149_n140# a_505_n140# 0.03fF
C82 a_741_n205# a_29_n205# 0.01fF
C83 w_n1133_n241# a_n327_n205# 0.19fF
C84 w_n1133_n241# a_n683_n205# 0.20fF
C85 a_919_n205# a_683_n140# 0.03fF
C86 w_n1133_n241# a_327_n140# 0.02fF
C87 w_n1133_n241# a_505_n140# 0.02fF
C88 a_n919_n140# a_n741_n140# 0.06fF
C89 a_861_n140# a_n563_n140# 0.01fF
C90 w_n1133_n241# a_149_n140# 0.02fF
C91 a_n327_n205# a_29_n205# 0.03fF
C92 a_n683_n205# a_29_n205# 0.01fF
C93 a_861_n140# a_n29_n140# 0.01fF
C94 a_n207_n140# a_919_n205# 0.01fF
C95 a_683_n140# a_n385_n140# 0.01fF
C96 a_n563_n140# a_n741_n140# 0.06fF
C97 w_n1133_n241# a_29_n205# 0.18fF
C98 a_n29_n140# a_n741_n140# 0.01fF
C99 a_n207_n140# a_n385_n140# 0.06fF
C100 a_207_n205# a_n149_n205# 0.03fF
C101 a_n861_n205# a_n149_n205# 0.01fF
C102 a_919_n205# a_n385_n140# 0.01fF
C103 a_n207_n140# a_n1097_n140# 0.01fF
C104 a_n149_n205# a_385_n205# 0.02fF
C105 a_n149_n205# a_563_n205# 0.01fF
C106 a_n919_n140# a_327_n140# 0.01fF
C107 a_n919_n140# a_505_n140# 0.01fF
C108 a_149_n140# a_n919_n140# 0.01fF
C109 a_861_n140# a_683_n140# 0.06fF
C110 a_n505_n205# a_n149_n205# 0.03fF
C111 w_n1133_n241# a_n919_n140# 0.02fF
C112 a_n207_n140# a_861_n140# 0.01fF
C113 a_741_n205# a_n149_n205# 0.01fF
C114 a_327_n140# a_n563_n140# 0.01fF
C115 a_n563_n140# a_505_n140# 0.01fF
C116 a_n1097_n140# a_n385_n140# 0.01fF
C117 a_149_n140# a_n563_n140# 0.01fF
C118 a_683_n140# a_n741_n140# 0.01fF
C119 a_n29_n140# a_327_n140# 0.03fF
C120 a_n29_n140# a_505_n140# 0.02fF
C121 a_149_n140# a_n29_n140# 0.06fF
C122 w_n1133_n241# a_n563_n140# 0.02fF
C123 a_n149_n205# a_n327_n205# 0.10fF
C124 a_n149_n205# a_n683_n205# 0.02fF
C125 a_861_n140# a_919_n205# 0.06fF
C126 a_n207_n140# a_n741_n140# 0.02fF
C127 w_n1133_n241# a_n29_n140# 0.02fF
C128 w_n1133_n241# a_n149_n205# 0.19fF
C129 a_861_n140# a_n385_n140# 0.01fF
C130 a_919_n205# a_207_n205# 0.01fF
C131 a_n149_n205# a_29_n205# 0.10fF
C132 a_919_n205# a_385_n205# 0.01fF
C133 a_919_n205# a_563_n205# 0.02fF
C134 a_n385_n140# a_n741_n140# 0.03fF
C135 a_683_n140# a_327_n140# 0.03fF
C136 a_683_n140# a_505_n140# 0.06fF
C137 a_149_n140# a_683_n140# 0.02fF
C138 a_n1097_n140# a_n741_n140# 0.03fF
C139 a_919_n205# a_n505_n205# 0.00fF
C140 a_n1097_n140# a_207_n205# 0.00fF
C141 a_n1097_n140# a_n861_n205# 0.07fF
C142 a_n919_n140# a_n563_n140# 0.03fF
C143 a_741_n205# a_919_n205# 0.07fF
C144 w_n1133_n241# a_683_n140# 0.01fF
C145 a_n207_n140# a_327_n140# 0.02fF
C146 a_n207_n140# a_505_n140# 0.01fF
C147 a_n207_n140# a_149_n140# 0.03fF
C148 a_n919_n140# a_n29_n140# 0.01fF
C149 a_n1097_n140# a_385_n205# 0.00fF
C150 a_n1097_n140# a_563_n205# 0.00fF
C151 a_919_n205# a_n327_n205# 0.00fF
C152 a_919_n205# a_n683_n205# 0.00fF
C153 w_n1133_n241# a_n207_n140# 0.02fF
C154 a_919_n205# a_327_n140# 0.01fF
C155 a_919_n205# a_505_n140# 0.02fF
C156 a_149_n140# a_919_n205# 0.01fF
C157 a_n29_n140# a_n563_n140# 0.02fF
C158 w_n1133_n241# VSUBS 3.28fF
.ends

.subckt ota_v2_without_cmfb in bias_c bias_e op on i_bias VDD bias_d m1_18877_3928#
+ m1_15613_3568# bias_circuit_0/li_3433_399# li_11121_570# cmc li_8434_570# li_8436_5651#
+ li_11122_5650# bias_circuit_0/m1_1243_5997# li_14138_570# bias_circuit_0/m1_3443_5997#
+ bias_a ip VSS bias_circuit_0/m1_5643_5997# VSUBS bias_b bias_circuit_0/m1_3551_3596#
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_0 VDD bias_b bias_b li_8436_5651# bias_b VDD bias_b
+ li_8436_5651# VDD li_8436_5651# VDD bias_b li_8436_5651# bias_b VDD VDD bias_b bias_b
+ VDD bias_b li_8436_5651# VDD bias_b li_8436_5651# li_8436_5651# bias_b VDD bias_b
+ VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_8 bias_d li_8434_570# bias_d on VSS bias_d on li_8434_570#
+ on bias_d bias_d bias_d on bias_d li_8434_570# VSS li_8434_570# bias_d bias_d on
+ li_8434_570# bias_d on on bias_d bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_1 VDD bias_b bias_b li_11122_5650# bias_b VDD
+ bias_b li_11122_5650# VDD li_11122_5650# VDD bias_b li_11122_5650# bias_b VDD VDD
+ bias_b bias_b VDD bias_b li_11122_5650# VDD bias_b li_11122_5650# li_11122_5650#
+ bias_b VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_9 bias_d li_11121_570# bias_d op VSS bias_d op li_11121_570#
+ op bias_d bias_d bias_d op bias_d li_11121_570# VSS li_11121_570# bias_d bias_d
+ op li_11121_570# bias_d op op bias_d bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_2 VDD bias_b bias_b li_8436_5651# bias_b VDD bias_b
+ li_8436_5651# VDD li_8436_5651# VDD bias_b li_8436_5651# bias_b VDD VDD bias_b bias_b
+ VDD bias_b li_8436_5651# VDD bias_b li_8436_5651# li_8436_5651# bias_b VDD bias_b
+ VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_3 VDD bias_b bias_b li_11122_5650# bias_b VDD
+ bias_b li_11122_5650# VDD li_11122_5650# VDD bias_b li_11122_5650# bias_b VDD VDD
+ bias_b bias_b VDD bias_b li_11122_5650# VDD bias_b li_11122_5650# li_11122_5650#
+ bias_b VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_0 VSS li_8436_5651# li_14138_570# ip li_8436_5651#
+ li_8436_5651# ip li_14138_570# li_8436_5651# li_14138_570# li_14138_570# li_8436_5651#
+ li_8436_5651# ip ip li_14138_570# ip li_14138_570# ip VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_1 VSS li_11122_5650# li_14138_570# in li_11122_5650#
+ li_11122_5650# in li_14138_570# li_11122_5650# li_14138_570# li_14138_570# li_11122_5650#
+ li_11122_5650# in in li_14138_570# in li_14138_570# in VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_AKSJZW_10 bias_d li_11121_570# bias_d op VSS bias_d op li_11121_570#
+ op bias_d bias_d bias_d op bias_d li_11121_570# VSS li_11121_570# bias_d bias_d
+ op li_11121_570# bias_d op op bias_d bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_0 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_AKSJZW_11 bias_d li_11121_570# bias_d op VSS bias_d op li_11121_570#
+ op bias_d bias_d bias_d op bias_d li_11121_570# VSS li_11121_570# bias_d bias_d
+ op li_11121_570# bias_d op op bias_d bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_1 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_2 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_3 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_4 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_5 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_6 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_7 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_8 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_9 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_10 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_11 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xbias_circuit_0 bias_c bias_e i_bias VDD bias_circuit_0/m1_7347_1428# bias_circuit_0/m1_7639_1420#
+ bias_circuit_0/li_3433_399# bias_a bias_circuit_0/m1_7169_923# bias_circuit_0/m1_7461_921#
+ bias_circuit_0/m1_7347_423# bias_circuit_0/m1_7639_427# bias_b VSS bias_circuit_0/m1_1243_5997#
+ bias_circuit_0/m1_3443_5997# bias_circuit_0/m1_3551_3596# bias_circuit_0/m1_5643_5997#
+ bias_d bias_circuit
Xsky130_fd_pr__pfet_01v8_YVTMSC_0 on bias_c li_8436_5651# bias_c bias_c li_8436_5651#
+ on VDD bias_c li_8436_5651# bias_c on VDD bias_c on bias_c li_8436_5651# VDD on
+ bias_c li_8436_5651# bias_c on bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_1 on bias_c li_8436_5651# bias_c bias_c li_8436_5651#
+ on VDD bias_c li_8436_5651# bias_c on VDD bias_c on bias_c li_8436_5651# VDD on
+ bias_c li_8436_5651# bias_c on bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_0 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_YVTMSC_2 op bias_c li_11122_5650# bias_c bias_c li_11122_5650#
+ op VDD bias_c li_11122_5650# bias_c op VDD bias_c op bias_c li_11122_5650# VDD op
+ bias_c li_11122_5650# bias_c op bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_3 op bias_c li_11122_5650# bias_c bias_c li_11122_5650#
+ op VDD bias_c li_11122_5650# bias_c op VDD bias_c op bias_c li_11122_5650# VDD op
+ bias_c li_11122_5650# bias_c op bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_2 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_1 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_3 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_4 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_5 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_6 bias_d li_8434_570# bias_d on VSS bias_d on li_8434_570#
+ on bias_d bias_d bias_d on bias_d li_8434_570# VSS li_8434_570# bias_d bias_d on
+ li_8434_570# bias_d on on bias_d bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_7 bias_d li_8434_570# bias_d on VSS bias_d on li_8434_570#
+ on bias_d bias_d bias_d on bias_d li_8434_570# VSS li_8434_570# bias_d bias_d on
+ li_8434_570# bias_d on on bias_d bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
C0 bias_d li_8436_5651# 0.66fF
C1 on bias_b 0.27fF
C2 bias_a li_8436_5651# 0.14fF
C3 li_14138_570# bias_d 0.02fF
C4 li_14138_570# bias_a 27.43fF
C5 cmc li_11122_5650# 0.13fF
C6 ip m1_15613_3568# 0.01fF
C7 on li_8436_5651# 2.52fF
C8 li_14138_570# m1_15613_3568# 0.01fF
C9 bias_c li_11122_5650# 3.17fF
C10 VDD bias_circuit_0/m1_3551_3596# 0.15fF
C11 op bias_b 0.27fF
C12 li_8434_570# bias_c 0.12fF
C13 in ip 0.03fF
C14 li_8434_570# bias_circuit_0/m1_7639_427# 0.01fF
C15 bias_d VDD 1.89fF
C16 bias_c li_11121_570# 0.12fF
C17 op li_8436_5651# 0.12fF
C18 li_11122_5650# li_11121_570# 0.16fF
C19 li_8434_570# bias_circuit_0/m1_7639_1420# 0.01fF
C20 in li_8436_5651# 0.01fF
C21 op li_14138_570# 0.08fF
C22 in li_14138_570# 1.51fF
C23 li_8436_5651# bias_b 4.47fF
C24 ip li_8436_5651# 1.22fF
C25 on VDD 0.63fF
C26 li_8434_570# li_11121_570# 0.52fF
C27 ip li_14138_570# 1.47fF
C28 li_14138_570# li_8436_5651# 0.80fF
C29 cmc bias_a 0.78fF
C30 op VDD 0.65fF
C31 bias_c bias_circuit_0/m1_3551_3596# 0.00fF
C32 m1_17393_3568# li_11122_5650# 0.00fF
C33 VDD bias_b 12.46fF
C34 bias_d bias_c 2.13fF
C35 bias_d li_11122_5650# 0.28fF
C36 bias_a bias_circuit_0/m1_7639_427# 0.01fF
C37 VDD li_8436_5651# 4.66fF
C38 bias_e li_8434_570# 0.00fF
C39 bias_d li_8434_570# 6.56fF
C40 in m1_18877_3928# 0.01fF
C41 bias_a li_8434_570# 10.56fF
C42 bias_d bias_circuit_0/m1_7639_1420# 0.00fF
C43 bias_a bias_circuit_0/m1_7639_1420# 0.00fF
C44 bias_c on 4.65fF
C45 on li_11122_5650# 0.12fF
C46 bias_d li_11121_570# 6.30fF
C47 bias_a li_11121_570# 10.56fF
C48 VDD bias_circuit_0/m1_5643_5997# -0.00fF
C49 li_8434_570# on 4.15fF
C50 in cmc 0.31fF
C51 bias_circuit_0/m1_7639_1420# on 0.00fF
C52 li_14138_570# m1_18877_3928# 0.00fF
C53 on li_11121_570# 0.17fF
C54 li_8434_570# bias_circuit_0/m1_7461_921# 0.01fF
C55 cmc li_14138_570# 26.78fF
C56 op bias_c 4.25fF
C57 op li_11122_5650# 2.52fF
C58 in li_11122_5650# 1.14fF
C59 bias_c bias_b 1.94fF
C60 bias_b li_11122_5650# 4.74fF
C61 ip li_11122_5650# 0.01fF
C62 op li_8434_570# 0.17fF
C63 bias_d bias_circuit_0/m1_3551_3596# 0.03fF
C64 op li_11121_570# 4.14fF
C65 bias_c li_8436_5651# 4.18fF
C66 li_8436_5651# li_11122_5650# 1.47fF
C67 li_14138_570# li_11122_5650# 0.78fF
C68 bias_a bias_e 0.00fF
C69 bias_a bias_d 2.86fF
C70 li_8434_570# li_8436_5651# 0.16fF
C71 on bias_circuit_0/m1_3551_3596# 0.00fF
C72 bias_e on 0.01fF
C73 bias_d on 10.13fF
C74 li_14138_570# li_11121_570# 0.23fF
C75 bias_a on 0.48fF
C76 bias_a m1_15613_3568# 0.01fF
C77 cmc m1_18877_3928# 0.01fF
C78 in m1_17097_3928# 0.00fF
C79 bias_c VDD 6.20fF
C80 VDD li_11122_5650# 4.01fF
C81 ip m1_17097_3928# 0.01fF
C82 in m1_17393_3568# 0.01fF
C83 li_8434_570# VDD 0.03fF
C84 ip m1_17393_3568# 0.00fF
C85 op bias_d 9.36fF
C86 op bias_a 0.52fF
C87 bias_d bias_b 0.02fF
C88 li_14138_570# m1_17097_3928# 0.00fF
C89 VDD li_11121_570# 0.02fF
C90 ip bias_a 0.31fF
C91 li_14138_570# m1_17393_3568# 0.01fF
C92 op on 0.59fF
C93 m1_17393_3568# VSS 0.09fF $ **FLOATING
C94 m1_15613_3568# VSS 0.12fF
C95 m1_18877_3928# VSS 0.10fF
C96 m1_17097_3928# VSS 0.06fF $ **FLOATING
C97 on VSS 5.53fF
C98 li_11121_570# VSS 11.01fF
C99 li_11122_5650# VSS -32.46fF
C100 li_8434_570# VSS 10.89fF
C101 li_8436_5651# VSS 5.93fF
C102 bias_circuit_0/m1_3551_3596# VSS -342.21fF
C103 bias_b VSS -361.08fF
C104 bias_circuit_0/m1_5643_5997# VSS 38.05fF
C105 bias_circuit_0/m1_3443_5997# VSS 35.85fF
C106 bias_circuit_0/m1_1243_5997# VSS 25.03fF
C107 VDD VSS 288.14fF
C108 i_bias VSS -60.67fF
C109 bias_c VSS -128.39fF
C110 bias_circuit_0/m1_7639_427# VSS 0.13fF
C111 bias_circuit_0/m1_7347_423# VSS 0.13fF
C112 bias_circuit_0/m1_7461_921# VSS 0.14fF
C113 bias_circuit_0/m1_7169_923# VSS 0.14fF
C114 bias_circuit_0/m1_7055_433# VSS 0.14fF
C115 bias_circuit_0/m1_6763_422# VSS 0.20fF
C116 bias_circuit_0/m1_6471_422# VSS 0.20fF
C117 bias_circuit_0/m1_7639_1420# VSS 0.13fF
C118 bias_circuit_0/m1_7347_1428# VSS 0.14fF
C119 bias_circuit_0/m1_6877_922# VSS 0.14fF
C120 bias_circuit_0/m1_6585_923# VSS 0.22fF
C121 bias_circuit_0/m1_6293_922# VSS 0.16fF
C122 bias_circuit_0/m1_7055_1417# VSS 0.14fF
C123 bias_circuit_0/m1_6763_1422# VSS 0.22fF
C124 bias_circuit_0/m1_6471_1426# VSS 0.22fF
C125 bias_e VSS 3.21fF
C126 bias_d VSS -235.00fF
C127 bias_circuit_0/li_3433_399# VSS 4.65fF
C128 bias_a VSS -295.16fF
C129 li_14138_570# VSS 42.14fF
C130 cmc VSS -107.95fF
C131 op VSS 5.33fF
C132 in VSS -27.58fF
C133 ip VSS -28.74fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 c1_n530_n480# m3_n630_n580# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_20/m3_n630_n580#
+ unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_24/c1_n530_n480#
+ unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480# transmission_gate_6/in
+ bias_a unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_27/m3_n630_n580# transmission_gate_8/in
+ unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# p2 on transmission_gate_4/out
+ transmission_gate_3/out p1 VDD unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480#
+ unit_cap_mim_m3m4_18/m3_n630_n580# cmc unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_7/in transmission_gate_9/in
+ cm unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# p1_b VSS
+ op p2_b
Xtransmission_gate_10 p1 VDD VSS transmission_gate_3/out on p1_b VSS transmission_gate
Xtransmission_gate_11 p1 VDD VSS transmission_gate_4/out op p1_b VSS transmission_gate
Xtransmission_gate_0 p1 VDD transmission_gate_0/nmos_tgate_0/w_n646_n262# cm transmission_gate_7/in
+ p1_b VSS transmission_gate
Xtransmission_gate_1 p1 VDD transmission_gate_1/nmos_tgate_0/w_n646_n262# cm transmission_gate_6/in
+ p1_b VSS transmission_gate
Xtransmission_gate_2 p1 VDD VSS bias_a transmission_gate_8/in p1_b VSS transmission_gate
Xtransmission_gate_3 p2 VDD VSS cm transmission_gate_3/out p2_b VSS transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 VDD transmission_gate_4/nmos_tgate_0/w_n646_n262# cm transmission_gate_4/out
+ p2_b VSS transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 VDD transmission_gate_5/nmos_tgate_0/w_n646_n262# bias_a transmission_gate_9/in
+ p2_b VSS transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 VDD VSS transmission_gate_6/in op p2_b VSS transmission_gate
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 VDD VSS transmission_gate_7/in on p2_b VSS transmission_gate
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 VDD VSS transmission_gate_8/in cmc p2_b VSS transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 VDD VSS transmission_gate_9/in cmc p1_b VSS transmission_gate
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.10fF
C1 p1 unit_cap_mim_m3m4_27/c1_n530_n480# 0.11fF
C2 op unit_cap_mim_m3m4_27/m3_n630_n580# 0.48fF
C3 p2 unit_cap_mim_m3m4_16/m3_n630_n580# 0.05fF
C4 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C5 op unit_cap_mim_m3m4_31/c1_n530_n480# 0.05fF
C6 transmission_gate_8/in transmission_gate_9/in 3.35fF
C7 bias_a transmission_gate_7/in 0.11fF
C8 cm transmission_gate_3/out 0.17fF
C9 p2 p1_b 5.94fF
C10 transmission_gate_4/out unit_cap_mim_m3m4_31/m3_n630_n580# 0.32fF
C11 cmc p1_b 0.53fF
C12 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_3/out -0.30fF
C13 transmission_gate_6/in transmission_gate_9/in 0.09fF
C14 unit_cap_mim_m3m4_34/c1_n530_n480# transmission_gate_7/in 0.06fF
C15 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_24/c1_n530_n480# -0.30fF
C16 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C17 unit_cap_mim_m3m4_18/m3_n630_n580# p1_b 0.06fF
C18 transmission_gate_6/in transmission_gate_8/in -0.31fF
C19 p2_b transmission_gate_9/in 0.01fF
C20 unit_cap_mim_m3m4_32/m3_n630_n580# cmc 0.12fF
C21 transmission_gate_4/out cm 0.07fF
C22 op on 2.00fF
C23 p2_b transmission_gate_8/in 0.40fF
C24 transmission_gate_7/in transmission_gate_9/in 0.02fF
C25 op VDD 0.89fF
C26 p1 unit_cap_mim_m3m4_29/m3_n630_n580# 0.06fF
C27 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.17fF
C28 p1 op 0.52fF
C29 cm p2 1.33fF
C30 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C31 transmission_gate_6/in p2_b 0.42fF
C32 transmission_gate_8/in transmission_gate_7/in 0.81fF
C33 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C34 unit_cap_mim_m3m4_21/m3_n630_n580# cmc 0.69fF
C35 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_16/c1_n530_n480# -0.21fF
C36 transmission_gate_8/in unit_cap_mim_m3m4_35/m3_n630_n580# -0.15fF
C37 transmission_gate_6/in transmission_gate_7/in 0.45fF
C38 bias_a p1_b 0.52fF
C39 on unit_cap_mim_m3m4_23/c1_n530_n480# 0.19fF
C40 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580# -0.21fF
C41 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C42 p2 unit_cap_mim_m3m4_27/c1_n530_n480# 0.04fF
C43 unit_cap_mim_m3m4_30/c1_n530_n480# transmission_gate_4/out -0.37fF
C44 p1 unit_cap_mim_m3m4_24/c1_n530_n480# 0.11fF
C45 p1_b unit_cap_mim_m3m4_17/m3_n630_n580# 0.06fF
C46 op transmission_gate_3/out 0.56fF
C47 p1 unit_cap_mim_m3m4_22/m3_n630_n580# 0.06fF
C48 p2_b transmission_gate_7/in 0.41fF
C49 unit_cap_mim_m3m4_29/c1_n530_n480# p1_b 0.06fF
C50 on unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C51 on unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C52 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580# -0.14fF
C53 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C54 op unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C55 unit_cap_mim_m3m4_16/m3_n630_n580# transmission_gate_9/in 0.17fF
C56 transmission_gate_6/in unit_cap_mim_m3m4_28/c1_n530_n480# 0.05fF
C57 p1_b transmission_gate_9/in 0.59fF
C58 p1 unit_cap_mim_m3m4_30/m3_n630_n580# 0.06fF
C59 unit_cap_mim_m3m4_23/c1_n530_n480# transmission_gate_3/out -0.24fF
C60 op transmission_gate_4/out 1.08fF
C61 cm bias_a 1.15fF
C62 unit_cap_mim_m3m4_25/c1_n530_n480# p1_b 0.06fF
C63 unit_cap_mim_m3m4_25/m3_n630_n580# transmission_gate_9/in 0.38fF
C64 transmission_gate_8/in p1_b 0.17fF
C65 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_25/c1_n530_n480# -0.32fF
C66 op p2 0.16fF
C67 unit_cap_mim_m3m4_31/m3_n630_n580# transmission_gate_9/in 0.12fF
C68 op cmc 4.24fF
C69 transmission_gate_6/in p1_b 0.41fF
C70 unit_cap_mim_m3m4_34/m3_n630_n580# transmission_gate_8/in 0.57fF
C71 transmission_gate_7/in unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C72 transmission_gate_4/out unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C73 p1 unit_cap_mim_m3m4_24/m3_n630_n580# 0.08fF
C74 on unit_cap_mim_m3m4_20/m3_n630_n580# 0.61fF
C75 p1 unit_cap_mim_m3m4_19/m3_n630_n580# 0.08fF
C76 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_31/c1_n530_n480# 0.06fF
C77 transmission_gate_8/in unit_cap_mim_m3m4_28/m3_n630_n580# 0.10fF
C78 p2_b p1_b 2.92fF
C79 p1 unit_cap_mim_m3m4_20/m3_n630_n580# 0.06fF
C80 cm transmission_gate_9/in 0.04fF
C81 p2 unit_cap_mim_m3m4_24/c1_n530_n480# 0.04fF
C82 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_9/in 0.17fF
C83 transmission_gate_6/in unit_cap_mim_m3m4_28/m3_n630_n580# -0.13fF
C84 transmission_gate_7/in p1_b 0.40fF
C85 cm transmission_gate_8/in 0.03fF
C86 unit_cap_mim_m3m4_22/m3_n630_n580# cmc 0.71fF
C87 transmission_gate_4/out unit_cap_mim_m3m4_30/m3_n630_n580# -0.80fF
C88 p1_b unit_cap_mim_m3m4_35/m3_n630_n580# 0.01fF
C89 transmission_gate_8/in unit_cap_mim_m3m4_21/m3_n630_n580# -1.15fF
C90 transmission_gate_6/in cm 0.17fF
C91 unit_cap_mim_m3m4_21/c1_n530_n480# cmc 0.13fF
C92 unit_cap_mim_m3m4_22/c1_n530_n480# cmc 0.13fF
C93 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# 0.17fF
C94 unit_cap_mim_m3m4_32/c1_n530_n480# on 0.06fF
C95 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480# -0.20fF
C96 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580# -0.13fF
C97 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580# -0.18fF
C98 on VDD 0.88fF
C99 cm p2_b 1.01fF
C100 p1 on 0.49fF
C101 transmission_gate_6/in unit_cap_mim_m3m4_27/c1_n530_n480# -0.13fF
C102 unit_cap_mim_m3m4_28/c1_n530_n480# p1_b 0.06fF
C103 p1 VDD 1.10fF
C104 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C105 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580# -0.29fF
C106 cm transmission_gate_7/in 0.10fF
C107 op unit_cap_mim_m3m4_29/c1_n530_n480# 0.03fF
C108 unit_cap_mim_m3m4_16/m3_n630_n580# p1_b 0.06fF
C109 transmission_gate_4/out unit_cap_mim_m3m4_31/c1_n530_n480# 0.05fF
C110 unit_cap_mim_m3m4_24/m3_n630_n580# p2 0.05fF
C111 unit_cap_mim_m3m4_33/m3_n630_n580# cmc 0.12fF
C112 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C113 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580# -0.33fF
C114 op transmission_gate_9/in 0.67fF
C115 on transmission_gate_3/out 0.40fF
C116 VDD transmission_gate_3/out -0.05fF
C117 unit_cap_mim_m3m4_27/m3_n630_n580# cmc 0.10fF
C118 p1 transmission_gate_3/out 0.72fF
C119 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C120 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C121 op transmission_gate_8/in 0.86fF
C122 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C123 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580# -0.20fF
C124 transmission_gate_6/in unit_cap_mim_m3m4_29/m3_n630_n580# -0.80fF
C125 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580# -0.19fF
C126 transmission_gate_6/in op 0.60fF
C127 on unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C128 transmission_gate_4/out on 3.24fF
C129 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C130 transmission_gate_4/out VDD -0.06fF
C131 unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_9/in -0.80fF
C132 p1 unit_cap_mim_m3m4_26/c1_n530_n480# 0.11fF
C133 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C134 p1 transmission_gate_4/out 0.80fF
C135 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C136 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.12fF
C137 op p2_b 0.40fF
C138 cm p1_b 1.15fF
C139 on p2 0.24fF
C140 unit_cap_mim_m3m4_23/m3_n630_n580# p1_b 0.05fF
C141 on cmc 1.91fF
C142 VDD p2 4.16fF
C143 unit_cap_mim_m3m4_21/m3_n630_n580# p1_b 0.05fF
C144 unit_cap_mim_m3m4_22/c1_n530_n480# transmission_gate_9/in -0.37fF
C145 VDD cmc 1.23fF
C146 p1 p2 2.82fF
C147 op transmission_gate_7/in 2.63fF
C148 p1 cmc 0.49fF
C149 unit_cap_mim_m3m4_21/c1_n530_n480# transmission_gate_8/in -0.41fF
C150 p1_b unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C151 p1 unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C152 on unit_cap_mim_m3m4_20/c1_n530_n480# 0.15fF
C153 transmission_gate_4/out transmission_gate_3/out 0.37fF
C154 p2 transmission_gate_3/out 0.15fF
C155 transmission_gate_3/out cmc 0.97fF
C156 op unit_cap_mim_m3m4_28/c1_n530_n480# 0.17fF
C157 unit_cap_mim_m3m4_24/m3_n630_n580# transmission_gate_9/in 0.17fF
C158 transmission_gate_8/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C159 VDD bias_a 0.99fF
C160 p2 unit_cap_mim_m3m4_26/c1_n530_n480# 0.04fF
C161 p1 bias_a 0.81fF
C162 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_8/in 0.17fF
C163 transmission_gate_4/out p2 0.15fF
C164 p1_b unit_cap_mim_m3m4_29/m3_n630_n580# 0.05fF
C165 transmission_gate_4/out cmc 0.10fF
C166 op p1_b 0.28fF
C167 transmission_gate_6/in unit_cap_mim_m3m4_27/m3_n630_n580# 0.13fF
C168 p1 unit_cap_mim_m3m4_17/m3_n630_n580# 0.08fF
C169 p1 unit_cap_mim_m3m4_29/c1_n530_n480# 0.11fF
C170 unit_cap_mim_m3m4_19/c1_n530_n480# transmission_gate_7/in 0.06fF
C171 p2 cmc 0.25fF
C172 op unit_cap_mim_m3m4_31/m3_n630_n580# 0.03fF
C173 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.17fF
C174 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_26/c1_n530_n480# -0.35fF
C175 op unit_cap_mim_m3m4_28/m3_n630_n580# 0.66fF
C176 bias_a transmission_gate_3/out 0.07fF
C177 on transmission_gate_9/in 1.05fF
C178 unit_cap_mim_m3m4_18/m3_n630_n580# cmc 0.17fF
C179 unit_cap_mim_m3m4_24/c1_n530_n480# p1_b 0.06fF
C180 transmission_gate_7/in unit_cap_mim_m3m4_19/m3_n630_n580# -0.28fF
C181 VDD transmission_gate_9/in -0.11fF
C182 unit_cap_mim_m3m4_22/m3_n630_n580# p1_b 0.05fF
C183 p1 transmission_gate_9/in 0.70fF
C184 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_7/in -0.56fF
C185 transmission_gate_3/out unit_cap_mim_m3m4_17/m3_n630_n580# -0.23fF
C186 on transmission_gate_8/in 0.88fF
C187 p1 unit_cap_mim_m3m4_25/c1_n530_n480# 0.11fF
C188 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# 0.12fF
C189 VDD transmission_gate_8/in -0.07fF
C190 cmc unit_cap_mim_m3m4_26/m3_n630_n580# 0.10fF
C191 p1 transmission_gate_8/in 0.39fF
C192 transmission_gate_6/in on 0.40fF
C193 transmission_gate_6/in VDD 0.03fF
C194 transmission_gate_4/out bias_a 0.10fF
C195 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C196 transmission_gate_6/in p1 0.38fF
C197 unit_cap_mim_m3m4_30/m3_n630_n580# p1_b 0.01fF
C198 transmission_gate_4/out unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C199 op unit_cap_mim_m3m4_27/c1_n530_n480# 0.01fF
C200 transmission_gate_3/out transmission_gate_9/in 1.40fF
C201 on p2_b 0.34fF
C202 p2 bias_a 0.60fF
C203 VDD p2_b 1.67fF
C204 p1 p2_b 2.16fF
C205 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_23/c1_n530_n480# -0.19fF
C206 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.17fF
C207 transmission_gate_8/in transmission_gate_3/out 0.24fF
C208 unit_cap_mim_m3m4_30/c1_n530_n480# op 0.18fF
C209 on transmission_gate_7/in 3.12fF
C210 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.10fF
C211 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.12fF
C212 p2 unit_cap_mim_m3m4_17/m3_n630_n580# 0.04fF
C213 VDD transmission_gate_7/in -0.16fF
C214 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C215 cmc unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C216 p1 transmission_gate_7/in 0.39fF
C217 p2 unit_cap_mim_m3m4_29/c1_n530_n480# 0.04fF
C218 transmission_gate_6/in transmission_gate_3/out 0.76fF
C219 unit_cap_mim_m3m4_24/m3_n630_n580# p1_b 0.06fF
C220 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C221 unit_cap_mim_m3m4_19/m3_n630_n580# p1_b 0.06fF
C222 transmission_gate_4/out transmission_gate_9/in 3.02fF
C223 p1 unit_cap_mim_m3m4_35/m3_n630_n580# 0.07fF
C224 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C225 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C226 unit_cap_mim_m3m4_20/m3_n630_n580# p1_b 0.05fF
C227 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C228 transmission_gate_4/out unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C229 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580# -0.19fF
C230 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.17fF
C231 transmission_gate_4/out transmission_gate_8/in 0.26fF
C232 p2_b transmission_gate_3/out 0.10fF
C233 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580# 0.12fF
C234 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C235 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C236 p2 transmission_gate_9/in 0.14fF
C237 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C238 op unit_cap_mim_m3m4_29/m3_n630_n580# 0.39fF
C239 cmc transmission_gate_9/in 6.62fF
C240 unit_cap_mim_m3m4_25/c1_n530_n480# p2 0.04fF
C241 transmission_gate_6/in transmission_gate_4/out 0.46fF
C242 transmission_gate_3/out transmission_gate_7/in 0.29fF
C243 p2 transmission_gate_8/in 0.63fF
C244 p1 unit_cap_mim_m3m4_28/c1_n530_n480# 0.11fF
C245 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# -0.25fF
C246 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.12fF
C247 transmission_gate_8/in cmc 8.44fF
C248 transmission_gate_6/in p2 0.61fF
C249 transmission_gate_4/out p2_b 0.05fF
C250 transmission_gate_6/in cmc 1.15fF
C251 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580# -0.12fF
C252 p1 unit_cap_mim_m3m4_16/m3_n630_n580# 0.08fF
C253 on p1_b 0.45fF
C254 op unit_cap_mim_m3m4_23/c1_n530_n480# 0.13fF
C255 VDD p1_b 1.01fF
C256 transmission_gate_4/out transmission_gate_7/in 0.61fF
C257 transmission_gate_6/in unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C258 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C259 p1 p1_b 8.88fF
C260 p2 p2_b 6.58fF
C261 p2_b cmc 0.12fF
C262 op unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C263 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_27/c1_n530_n480# -0.37fF
C264 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_32/c1_n530_n480# -0.20fF
C265 p2 transmission_gate_7/in 0.60fF
C266 cmc transmission_gate_7/in 0.07fF
C267 op unit_cap_mim_m3m4_22/c1_n530_n480# 0.07fF
C268 bias_a transmission_gate_9/in 0.02fF
C269 op unit_cap_mim_m3m4_30/m3_n630_n580# 0.56fF
C270 bias_a transmission_gate_8/in 0.04fF
C271 transmission_gate_3/out p1_b 0.59fF
C272 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_31/c1_n530_n480# 0.06fF
C273 unit_cap_mim_m3m4_20/c1_n530_n480# transmission_gate_7/in -0.18fF
C274 VDD cm 1.83fF
C275 unit_cap_mim_m3m4_23/m3_n630_n580# on 0.47fF
C276 p1 cm 1.50fF
C277 transmission_gate_6/in bias_a 0.07fF
C278 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C279 unit_cap_mim_m3m4_23/m3_n630_n580# p1 0.06fF
C280 p2 unit_cap_mim_m3m4_28/c1_n530_n480# 0.04fF
C281 p1 unit_cap_mim_m3m4_21/m3_n630_n580# 0.06fF
C282 transmission_gate_4/out unit_cap_mim_m3m4_16/m3_n630_n580# -0.28fF
C283 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480# -0.19fF
C284 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C285 p1_b unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C286 transmission_gate_4/out p1_b 0.55fF
C287 p2_b bias_a 0.48fF
C288 transmission_gate_6/in unit_cap_mim_m3m4_29/c1_n530_n480# -0.37fF
C289 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C290 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C291 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.39fF
C292 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C293 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.51fF
C294 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C295 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.74fF
C296 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.51fF
C297 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.51fF
C298 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.82fF
C299 cmc VSS -31.94fF
C300 transmission_gate_9/in VSS 3.96fF
C301 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.60fF
C302 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.61fF
C303 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.61fF
C304 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C305 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C306 p2 VSS 148.24fF
C307 p2_b VSS 41.62fF
C308 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.84fF
C309 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C310 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.39fF
C311 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C312 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.04fF
C313 transmission_gate_3/out VSS 2.28fF
C314 transmission_gate_8/in VSS 2.29fF
C315 bias_a VSS 11.61fF
C316 transmission_gate_6/in VSS -13.31fF
C317 transmission_gate_7/in VSS 9.28fF
C318 cm VSS 13.12fF
C319 p1 VSS 112.15fF
C320 op VSS -1.36fF
C321 transmission_gate_4/out VSS -3.74fF
C322 p1_b VSS 173.84fF
C323 VDD VSS 71.01fF
C324 on VSS -23.21fF
.ends

.subckt ota_v2 ip in op i_bias ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580#
+ ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# ota_v2_without_cmfb_0/li_11122_5650#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_8/in ota_v2_without_cmfb_0/li_11121_570# sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480#
+ ota_v2_without_cmfb_0/li_8434_570# sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580#
+ on sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# ota_v2_without_cmfb_0/li_8436_5651#
+ sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# sc_cmfb_0/transmission_gate_6/in ota_v2_without_cmfb_0/bias_c
+ sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/bias_a
+ VDD sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ ota_v2_without_cmfb_0/bias_b p1_b sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480#
+ ota_v2_without_cmfb_0/li_14138_570# sc_cmfb_0/transmission_gate_9/in sc_cmfb_0/cmc
+ ota_v2_without_cmfb_0/m1_18877_3928# sc_cmfb_0/transmission_gate_4/out cm p2_b p2
+ ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# p1 ota_v2_without_cmfb_0/bias_d
+ ota_v2_without_cmfb_0/m1_15613_3568# VSS
Xota_v2_without_cmfb_0 in ota_v2_without_cmfb_0/bias_c cm op on i_bias VDD ota_v2_without_cmfb_0/bias_d
+ ota_v2_without_cmfb_0/m1_18877_3928# ota_v2_without_cmfb_0/m1_15613_3568# ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399#
+ ota_v2_without_cmfb_0/li_11121_570# sc_cmfb_0/cmc ota_v2_without_cmfb_0/li_8434_570#
+ ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997#
+ ota_v2_without_cmfb_0/li_14138_570# ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997#
+ sc_cmfb_0/bias_a ip VSS ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS ota_v2_without_cmfb_0/bias_b
+ ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# ota_v2_without_cmfb
Xsc_cmfb_0 sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# sc_cmfb_0/transmission_gate_6/in sc_cmfb_0/bias_a
+ sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580#
+ p2 on sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_3/out p1 VDD
+ sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# sc_cmfb_0/cmc sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/transmission_gate_9/in cm sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# p1_b VSS op p2_b sc_cmfb
C0 ip op 0.01fF
C1 sc_cmfb_0/bias_a VDD 0.02fF
C2 sc_cmfb_0/cmc on 0.31fF
C3 VDD p1_b -0.00fF
C4 sc_cmfb_0/bias_a p1_b 0.00fF
C5 ota_v2_without_cmfb_0/bias_c cm 2.51fF
C6 VDD cm -0.07fF
C7 sc_cmfb_0/bias_a cm 3.22fF
C8 sc_cmfb_0/transmission_gate_4/out p1 0.05fF
C9 cm p1_b 0.01fF
C10 ota_v2_without_cmfb_0/li_14138_570# in -0.00fF
C11 cm ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# 0.23fF
C12 VDD sc_cmfb_0/transmission_gate_8/in 0.02fF
C13 sc_cmfb_0/bias_a sc_cmfb_0/transmission_gate_8/in 0.00fF
C14 VDD sc_cmfb_0/transmission_gate_7/in 0.01fF
C15 op ota_v2_without_cmfb_0/li_8436_5651# 0.40fF
C16 op sc_cmfb_0/transmission_gate_4/out -0.00fF
C17 cm ota_v2_without_cmfb_0/li_8434_570# 0.38fF
C18 sc_cmfb_0/bias_a p1 0.00fF
C19 p1_b p1 0.00fF
C20 op ota_v2_without_cmfb_0/li_14138_570# 0.00fF
C21 ota_v2_without_cmfb_0/bias_c ota_v2_without_cmfb_0/bias_b 0.26fF
C22 ota_v2_without_cmfb_0/li_8436_5651# on 0.37fF
C23 ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/bias_b -0.00fF
C24 VDD ota_v2_without_cmfb_0/bias_b 0.16fF
C25 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_b 0.15fF
C26 ota_v2_without_cmfb_0/li_14138_570# on 0.01fF
C27 op ota_v2_without_cmfb_0/bias_c 1.56fF
C28 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_d -0.00fF
C29 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_4/out -0.02fF
C30 op ota_v2_without_cmfb_0/li_11122_5650# 0.36fF
C31 p1 sc_cmfb_0/transmission_gate_8/in 0.00fF
C32 sc_cmfb_0/cmc ota_v2_without_cmfb_0/li_14138_570# 0.03fF
C33 ota_v2_without_cmfb_0/bias_c i_bias 0.00fF
C34 cm ota_v2_without_cmfb_0/bias_b 3.45fF
C35 op VDD 3.19fF
C36 op p1_b 0.00fF
C37 ip ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C38 ota_v2_without_cmfb_0/bias_d cm 4.24fF
C39 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.00fF
C40 ota_v2_without_cmfb_0/bias_c on -0.00fF
C41 op cm 1.43fF
C42 ota_v2_without_cmfb_0/li_11121_570# cm 0.39fF
C43 p2_b p1 0.00fF
C44 ip ota_v2_without_cmfb_0/li_14138_570# 0.00fF
C45 ota_v2_without_cmfb_0/li_11122_5650# on 0.22fF
C46 VDD on 0.45fF
C47 p1_b on 0.01fF
C48 sc_cmfb_0/cmc VDD -0.08fF
C49 ota_v2_without_cmfb_0/bias_d ota_v2_without_cmfb_0/li_8434_570# -0.00fF
C50 cm on 3.11fF
C51 sc_cmfb_0/cmc cm -2.78fF
C52 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# 0.00fF
C53 op p1 0.01fF
C54 ota_v2_without_cmfb_0/li_8434_570# on 0.00fF
C55 ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/li_14138_570# 0.00fF
C56 on p1 0.01fF
C57 ota_v2_without_cmfb_0/li_11121_570# ota_v2_without_cmfb_0/bias_d -0.00fF
C58 op ota_v2_without_cmfb_0/bias_d -0.00fF
C59 ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/bias_c -0.00fF
C60 ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/li_11122_5650# -0.00fF
C61 op ota_v2_without_cmfb_0/li_11121_570# 0.00fF
C62 ota_v2_without_cmfb_0/li_8436_5651# VDD -0.00fF
C63 VDD sc_cmfb_0/transmission_gate_4/out 0.04fF
C64 p1_b sc_cmfb_0/transmission_gate_4/out 0.00fF
C65 ota_v2_without_cmfb_0/bias_d on 7.34fF
C66 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# 0.00fF
C67 ota_v2_without_cmfb_0/li_11121_570# on 0.01fF
C68 op on 3.51fF
C69 op sc_cmfb_0/cmc 0.37fF
C70 ota_v2_without_cmfb_0/li_14138_570# cm 1.29fF
C71 ota_v2_without_cmfb_0/bias_c ota_v2_without_cmfb_0/li_11122_5650# 0.00fF
C72 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_c 2.52fF
C73 VDD ota_v2_without_cmfb_0/li_11122_5650# 0.23fF
C74 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C75 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C76 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C77 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C78 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C79 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C80 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C81 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C82 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C83 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.37fF
C84 sc_cmfb_0/transmission_gate_9/in VSS 2.58fF
C85 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C86 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C87 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C88 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C89 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C90 p2 VSS 147.84fF
C91 p2_b VSS 39.93fF
C92 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C93 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C94 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C95 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C96 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.86fF
C97 sc_cmfb_0/transmission_gate_3/out VSS 1.19fF
C98 sc_cmfb_0/transmission_gate_8/in VSS 1.29fF
C99 sc_cmfb_0/transmission_gate_6/in VSS -14.72fF
C100 sc_cmfb_0/transmission_gate_7/in VSS 7.87fF
C101 cm VSS 36.42fF
C102 p1 VSS 111.00fF
C103 op VSS 4.21fF
C104 sc_cmfb_0/transmission_gate_4/out VSS -4.84fF
C105 p1_b VSS 172.94fF
C106 on VSS -20.78fF
C107 ota_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C108 ota_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF
C109 ota_v2_without_cmfb_0/m1_18877_3928# VSS 0.05fF
C110 ota_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C111 ota_v2_without_cmfb_0/li_11121_570# VSS 9.29fF
C112 ota_v2_without_cmfb_0/li_11122_5650# VSS -32.55fF
C113 ota_v2_without_cmfb_0/li_8434_570# VSS 9.00fF
C114 ota_v2_without_cmfb_0/li_8436_5651# VSS 5.90fF
C115 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -342.20fF
C116 ota_v2_without_cmfb_0/bias_b VSS -361.14fF
C117 ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C118 ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.85fF
C119 ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C120 VDD VSS 358.85fF
C121 i_bias VSS -61.81fF
C122 ota_v2_without_cmfb_0/bias_c VSS -128.70fF
C123 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C124 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C125 ota_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C126 ota_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C127 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C128 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C129 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C130 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C131 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.13fF
C132 ota_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C133 ota_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C134 ota_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C135 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.14fF
C136 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C137 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C138 ota_v2_without_cmfb_0/bias_d VSS -236.30fF
C139 ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 4.65fF
C140 sc_cmfb_0/bias_a VSS -319.09fF
C141 ota_v2_without_cmfb_0/li_14138_570# VSS 33.89fF
C142 sc_cmfb_0/cmc VSS -143.12fF
C143 in VSS -28.56fF
C144 ip VSS -29.73fF
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y w_82_21# VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 A Y 0.88fF
C1 VPB A 0.21fF
C2 VPB Y 0.05fF
C3 VPWR A 0.13fF
C4 VPWR Y 1.13fF
C5 VPWR VPB 0.34fF
C6 VGND A 0.13fF
C7 VGND Y 0.56fF
C8 VGND VPWR 0.10fF
C9 VGND VNB 0.40fF
C10 Y VNB 0.10fF
C11 VPWR VNB 0.14fF
C12 A VNB 0.47fF
C13 VPB VNB 0.69fF
.ends

.subckt onebit_dac v VDD v_hi v_b v_lo out VSS
Xtransmission_gate_0 v VDD transmission_gate_0/nmos_tgate_0/w_n646_n262# v_hi out
+ v_b VSS transmission_gate
Xtransmission_gate_1 v_b VDD transmission_gate_1/nmos_tgate_0/w_n646_n262# v_lo out
+ v VSS transmission_gate
C0 v v_hi 0.49fF
C1 out v_hi 0.20fF
C2 v_b v_lo 0.40fF
C3 out v 0.29fF
C4 VDD v_lo -0.13fF
C5 v_b VDD 0.62fF
C6 v_hi v_lo 0.47fF
C7 v_b v_hi 0.45fF
C8 VDD v_hi 0.20fF
C9 v v_lo 0.46fF
C10 out v_lo 0.30fF
C11 v_b v 0.53fF
C12 v_b out 1.55fF
C13 VDD v 0.33fF
C14 out VDD -0.09fF
C15 v_b VSS 0.47fF
C16 v_lo VSS 1.40fF
C17 v VSS 1.66fF
C18 VDD VSS 7.83fF
C19 out VSS 1.99fF
C20 v_hi VSS 1.57fF
.ends

.subckt nmos_PDN_mux2 a_n33_32# a_15_n90# a_n73_n90# VSUBS
X0 a_15_n90# a_n33_32# a_n73_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
C0 a_n73_n90# a_n33_32# 0.01fF
C1 a_15_n90# a_n33_32# 0.01fF
C2 a_n73_n90# a_15_n90# 0.14fF
C3 a_15_n90# VSUBS 0.02fF
C4 a_n73_n90# VSUBS 0.02fF
C5 a_n33_32# VSUBS 0.15fF
.ends

.subckt switch_5t_mux2 in out en_b VDD transmission_gate_0/nmos_tgate_0/w_n646_n262#
+ en VSS transmission_gate_1/in
Xnmos_PDN_mux2_0 en_b transmission_gate_1/in VSS VSS nmos_PDN_mux2
Xtransmission_gate_0 en VDD transmission_gate_0/nmos_tgate_0/w_n646_n262# in transmission_gate_1/in
+ en_b VSS transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/nmos_tgate_0/w_n646_n262# transmission_gate_1/in
+ out en_b VSS transmission_gate
C0 transmission_gate_1/in en_b 0.67fF
C1 in transmission_gate_1/in 0.68fF
C2 VDD en_b 0.59fF
C3 in VDD 0.10fF
C4 en transmission_gate_1/in 0.51fF
C5 in en_b 0.50fF
C6 en en_b 0.19fF
C7 en in 0.51fF
C8 out transmission_gate_1/in 0.72fF
C9 out VDD -0.13fF
C10 out en_b 0.11fF
C11 out in 0.43fF
C12 out en 0.10fF
C13 transmission_gate_1/in VDD 0.19fF
C14 en VSS 4.27fF
C15 out VSS 0.81fF
C16 en_b VSS 0.43fF
C17 VDD VSS 10.97fF
C18 transmission_gate_1/in VSS 1.85fF
C19 in VSS 0.97fF
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
C0 VPB A 0.08fF
C1 VPWR Y 0.22fF
C2 VGND Y 0.17fF
C3 VGND VPWR 0.05fF
C4 VPB Y 0.06fF
C5 VPWR VPB 0.21fF
C6 A Y 0.05fF
C7 VPWR A 0.05fF
C8 VGND A 0.05fF
C9 VGND VNB 0.25fF
C10 Y VNB 0.06fF
C11 VPWR VNB 0.06fF
C12 A VNB 0.13fF
C13 VPB VNB 0.34fF
.ends

.subckt a_mux2_en en in0 in1 out transmission_gate_1/en_b switch_5t_mux2_0/transmission_gate_1/in
+ switch_5t_mux2_1/en VDD switch_5t_mux2_1/transmission_gate_1/in switch_5t_mux2_1/in
+ VSS s0 switch_5t_mux2_0/in
Xswitch_5t_mux2_0 switch_5t_mux2_0/in out switch_5t_mux2_1/en VDD switch_5t_mux2_0/transmission_gate_0/nmos_tgate_0/w_n646_n262#
+ s0 VSS switch_5t_mux2_0/transmission_gate_1/in switch_5t_mux2
Xswitch_5t_mux2_1 switch_5t_mux2_1/in out s0 VDD switch_5t_mux2_1/transmission_gate_0/nmos_tgate_0/w_n646_n262#
+ switch_5t_mux2_1/en VSS switch_5t_mux2_1/transmission_gate_1/in switch_5t_mux2
Xtransmission_gate_0 en VDD transmission_gate_0/nmos_tgate_0/w_n646_n262# in0 switch_5t_mux2_1/in
+ transmission_gate_1/en_b VSS transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/nmos_tgate_0/w_n646_n262# in1 switch_5t_mux2_0/in
+ transmission_gate_1/en_b VSS transmission_gate
Xsky130_fd_sc_hd__inv_1_1 switch_5t_mux2_1/en s0 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 transmission_gate_1/en_b en VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
C0 VDD s0 0.92fF
C1 transmission_gate_1/en_b switch_5t_mux2_1/en 0.05fF
C2 switch_5t_mux2_1/in switch_5t_mux2_0/transmission_gate_1/in 0.07fF
C3 en switch_5t_mux2_1/transmission_gate_0/nmos_tgate_0/w_n646_n262# 0.00fF
C4 in1 switch_5t_mux2_0/in 0.01fF
C5 transmission_gate_1/en_b s0 0.03fF
C6 switch_5t_mux2_1/en switch_5t_mux2_0/transmission_gate_1/in 0.02fF
C7 switch_5t_mux2_0/transmission_gate_0/nmos_tgate_0/w_n646_n262# switch_5t_mux2_0/in 0.00fF
C8 switch_5t_mux2_0/transmission_gate_1/in s0 0.04fF
C9 switch_5t_mux2_1/transmission_gate_1/in switch_5t_mux2_0/in 0.06fF
C10 out switch_5t_mux2_1/transmission_gate_1/in 0.21fF
C11 en in1 0.09fF
C12 en switch_5t_mux2_0/in 0.40fF
C13 switch_5t_mux2_1/in switch_5t_mux2_1/en 0.21fF
C14 in1 in0 0.49fF
C15 in1 VDD -0.10fF
C16 in0 switch_5t_mux2_0/in 0.08fF
C17 VDD switch_5t_mux2_0/in 0.22fF
C18 out VDD 0.28fF
C19 switch_5t_mux2_1/in s0 0.19fF
C20 transmission_gate_1/en_b in1 0.14fF
C21 switch_5t_mux2_1/transmission_gate_1/in VDD 0.39fF
C22 switch_5t_mux2_1/en s0 0.78fF
C23 transmission_gate_1/en_b switch_5t_mux2_0/in 0.16fF
C24 switch_5t_mux2_1/transmission_gate_0/nmos_tgate_0/w_n646_n262# switch_5t_mux2_1/in 0.00fF
C25 en in0 0.07fF
C26 en VDD 0.65fF
C27 switch_5t_mux2_0/transmission_gate_1/in switch_5t_mux2_0/in 0.06fF
C28 out switch_5t_mux2_0/transmission_gate_1/in 0.15fF
C29 in0 VDD 0.18fF
C30 en transmission_gate_1/en_b 0.43fF
C31 switch_5t_mux2_1/transmission_gate_1/in switch_5t_mux2_0/transmission_gate_1/in 0.32fF
C32 switch_5t_mux2_1/in in1 0.08fF
C33 transmission_gate_1/en_b in0 0.13fF
C34 transmission_gate_1/en_b VDD 0.62fF
C35 en switch_5t_mux2_0/transmission_gate_1/in 0.01fF
C36 switch_5t_mux2_1/in switch_5t_mux2_0/in 0.35fF
C37 switch_5t_mux2_0/transmission_gate_1/in VDD 0.22fF
C38 switch_5t_mux2_1/in switch_5t_mux2_1/transmission_gate_1/in 0.03fF
C39 switch_5t_mux2_1/en switch_5t_mux2_0/in 0.06fF
C40 out switch_5t_mux2_1/en 0.01fF
C41 en switch_5t_mux2_1/in 0.13fF
C42 switch_5t_mux2_1/en switch_5t_mux2_1/transmission_gate_1/in 0.10fF
C43 transmission_gate_1/en_b switch_5t_mux2_0/transmission_gate_1/in 0.01fF
C44 switch_5t_mux2_0/in s0 -0.00fF
C45 out s0 0.08fF
C46 switch_5t_mux2_1/in in0 0.00fF
C47 switch_5t_mux2_1/in VDD 0.53fF
C48 en switch_5t_mux2_1/en 0.22fF
C49 switch_5t_mux2_1/transmission_gate_1/in s0 0.12fF
C50 switch_5t_mux2_1/en in0 0.03fF
C51 en s0 0.15fF
C52 switch_5t_mux2_1/en VDD 1.15fF
C53 switch_5t_mux2_1/in transmission_gate_1/en_b 0.11fF
C54 in0 s0 0.02fF
C55 VDD VSS 5.36fF
C56 en VSS 12.78fF
C57 switch_5t_mux2_0/in VSS 1.12fF
C58 in1 VSS 1.31fF
C59 transmission_gate_1/en_b VSS -0.92fF
C60 switch_5t_mux2_1/in VSS -1.08fF
C61 in0 VSS 1.93fF
C62 switch_5t_mux2_1/en VSS 12.04fF
C63 s0 VSS 10.75fF
C64 switch_5t_mux2_1/transmission_gate_1/in VSS 1.71fF
C65 out VSS 1.48fF
C66 switch_5t_mux2_0/transmission_gate_1/in VSS 1.47fF
.ends

.subckt ota_w_test_v2 ip in op sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/li_11122_5650# sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997#
+ sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997#
+ sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_v2_without_cmfb_0/li_8434_570#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_v2_without_cmfb_0/bias_b on sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580#
+ sc_cmfb_0/bias_a sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_6/in sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# sc_cmfb_0/transmission_gate_7/in VDD
+ sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# sc_cmfb_0/cmc sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580#
+ ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ p1_b sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480#
+ i_bias sc_cmfb_0/transmission_gate_9/in ota_v2_without_cmfb_0/m1_18877_3928# sc_cmfb_0/transmission_gate_4/out
+ VSS cm p2_b ota_v2_without_cmfb_0/li_14138_570# p2 ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399#
+ ota_v2_without_cmfb_0/bias_c p1 ota_v2_without_cmfb_0/bias_d ota_v2_without_cmfb_0/m1_15613_3568#
Xota_v2_without_cmfb_0 in ota_v2_without_cmfb_0/bias_c cm op on i_bias VDD ota_v2_without_cmfb_0/bias_d
+ ota_v2_without_cmfb_0/m1_18877_3928# ota_v2_without_cmfb_0/m1_15613_3568# ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399#
+ ota_v2_without_cmfb_0/li_11121_570# sc_cmfb_0/cmc ota_v2_without_cmfb_0/li_8434_570#
+ ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997#
+ ota_v2_without_cmfb_0/li_14138_570# ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997#
+ sc_cmfb_0/bias_a ip VSS ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# ota_v2_without_cmfb_0/VSUBS
+ ota_v2_without_cmfb_0/bias_b ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596#
+ ota_v2_without_cmfb
Xsc_cmfb_0 sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# sc_cmfb_0/transmission_gate_6/in sc_cmfb_0/bias_a
+ sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580#
+ p2 on sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_3/out p1 VDD
+ sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# sc_cmfb_0/cmc sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/transmission_gate_9/in cm sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# p1_b VSS op p2_b sc_cmfb
C0 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.00fF
C1 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_4/out -0.00fF
C2 ota_v2_without_cmfb_0/bias_c i_bias 0.00fF
C3 ota_v2_without_cmfb_0/bias_c ota_v2_without_cmfb_0/bias_b 0.29fF
C4 p1_b cm 0.01fF
C5 on ota_v2_without_cmfb_0/li_11121_570# 0.01fF
C6 ota_v2_without_cmfb_0/li_14138_570# cm 1.02fF
C7 sc_cmfb_0/transmission_gate_8/in p1 0.00fF
C8 VDD ota_v2_without_cmfb_0/bias_b 0.16fF
C9 in ota_v2_without_cmfb_0/li_14138_570# -0.00fF
C10 on ota_v2_without_cmfb_0/li_8436_5651# 0.44fF
C11 VDD p1_b 0.00fF
C12 p1_b op 0.00fF
C13 sc_cmfb_0/cmc ota_v2_without_cmfb_0/li_14138_570# 0.03fF
C14 ota_v2_without_cmfb_0/li_14138_570# op 0.01fF
C15 ota_v2_without_cmfb_0/bias_d cm 4.20fF
C16 ota_v2_without_cmfb_0/li_8434_570# cm 0.38fF
C17 sc_cmfb_0/transmission_gate_8/in VDD 0.07fF
C18 ota_v2_without_cmfb_0/bias_d op -0.00fF
C19 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# 0.00fF
C20 on p1_b 0.23fF
C21 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_b 0.15fF
C22 ota_v2_without_cmfb_0/li_14138_570# on 0.02fF
C23 sc_cmfb_0/bias_a p1_b 0.00fF
C24 p1 sc_cmfb_0/transmission_gate_4/out 0.05fF
C25 ip op 0.01fF
C26 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# cm 0.23fF
C27 ota_v2_without_cmfb_0/li_14138_570# ota_v2_without_cmfb_0/li_8436_5651# 0.00fF
C28 ota_v2_without_cmfb_0/bias_d on 4.96fF
C29 on sc_cmfb_0/transmission_gate_3/out 0.00fF
C30 ota_v2_without_cmfb_0/li_8434_570# on 0.00fF
C31 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/bias_a 0.00fF
C32 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_d -0.00fF
C33 ota_v2_without_cmfb_0/bias_d ota_v2_without_cmfb_0/li_11121_570# -0.00fF
C34 VDD sc_cmfb_0/transmission_gate_4/out 0.03fF
C35 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# 0.00fF
C36 sc_cmfb_0/transmission_gate_4/out op -0.00fF
C37 p1 op 0.00fF
C38 ota_v2_without_cmfb_0/bias_c cm 1.19fF
C39 ota_v2_without_cmfb_0/bias_c ota_v2_without_cmfb_0/li_11122_5650# 0.00fF
C40 VDD cm -0.07fF
C41 sc_cmfb_0/cmc cm -1.06fF
C42 ota_v2_without_cmfb_0/li_11122_5650# VDD 0.23fF
C43 ip ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C44 op cm 1.43fF
C45 ota_v2_without_cmfb_0/li_11122_5650# op 0.34fF
C46 ota_v2_without_cmfb_0/bias_c op -0.51fF
C47 sc_cmfb_0/cmc VDD 0.14fF
C48 sc_cmfb_0/transmission_gate_7/in cm -0.03fF
C49 VDD op 3.66fF
C50 sc_cmfb_0/cmc op 0.38fF
C51 on p1 0.01fF
C52 sc_cmfb_0/bias_a p1 0.00fF
C53 VDD sc_cmfb_0/transmission_gate_7/in 0.01fF
C54 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# -0.01fF
C55 on cm 2.94fF
C56 ota_v2_without_cmfb_0/li_11122_5650# on 1.38fF
C57 ota_v2_without_cmfb_0/bias_c on -0.00fF
C58 sc_cmfb_0/bias_a cm 3.29fF
C59 ota_v2_without_cmfb_0/li_11121_570# cm 0.39fF
C60 ip ota_v2_without_cmfb_0/li_14138_570# -0.01fF
C61 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_c 0.74fF
C62 VDD on 0.32fF
C63 sc_cmfb_0/cmc on 0.49fF
C64 ota_v2_without_cmfb_0/bias_d ota_v2_without_cmfb_0/li_8434_570# -0.00fF
C65 on op 1.99fF
C66 sc_cmfb_0/bias_a VDD 0.00fF
C67 ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C68 ota_v2_without_cmfb_0/bias_c ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C69 op ota_v2_without_cmfb_0/li_11121_570# 0.00fF
C70 VDD ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C71 op ota_v2_without_cmfb_0/li_8436_5651# 0.39fF
C72 p1_b sc_cmfb_0/transmission_gate_4/out 0.00fF
C73 p1 p1_b 0.00fF
C74 p2_b p1 0.00fF
C75 ota_v2_without_cmfb_0/bias_b cm 2.71fF
C76 ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/bias_b -0.00fF
C77 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C78 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C79 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C80 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C81 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C82 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C83 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C84 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C85 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C86 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.50fF
C87 sc_cmfb_0/transmission_gate_9/in VSS 2.58fF
C88 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C89 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C90 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C91 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C92 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C93 p2 VSS 147.84fF
C94 p2_b VSS 39.88fF
C95 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C96 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C97 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C98 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C99 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.77fF
C100 sc_cmfb_0/transmission_gate_3/out VSS 1.19fF
C101 sc_cmfb_0/transmission_gate_8/in VSS 1.33fF
C102 sc_cmfb_0/transmission_gate_6/in VSS -14.72fF
C103 sc_cmfb_0/transmission_gate_7/in VSS 7.87fF
C104 cm VSS 24.75fF
C105 p1 VSS 110.99fF
C106 op VSS 2.48fF
C107 sc_cmfb_0/transmission_gate_4/out VSS -4.84fF
C108 p1_b VSS 172.45fF
C109 on VSS -19.61fF
C110 ota_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C111 ota_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF
C112 ota_v2_without_cmfb_0/m1_18877_3928# VSS 0.05fF
C113 ota_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C114 ota_v2_without_cmfb_0/li_11121_570# VSS 9.29fF
C115 ota_v2_without_cmfb_0/li_11122_5650# VSS -32.55fF
C116 ota_v2_without_cmfb_0/li_8434_570# VSS 9.00fF
C117 ota_v2_without_cmfb_0/li_8436_5651# VSS 5.90fF
C118 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -342.20fF
C119 ota_v2_without_cmfb_0/bias_b VSS -361.14fF
C120 ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C121 ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.85fF
C122 ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C123 VDD VSS 361.99fF
C124 i_bias VSS -62.81fF
C125 ota_v2_without_cmfb_0/bias_c VSS -128.72fF
C126 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C127 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C128 ota_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C129 ota_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C130 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C131 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C132 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C133 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C134 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.13fF
C135 ota_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C136 ota_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C137 ota_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C138 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.14fF
C139 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C140 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C141 ota_v2_without_cmfb_0/bias_d VSS -236.30fF
C142 ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 4.65fF
C143 sc_cmfb_0/bias_a VSS -313.39fF
C144 ota_v2_without_cmfb_0/li_14138_570# VSS 33.90fF
C145 sc_cmfb_0/cmc VSS -141.20fF
C146 in VSS -28.57fF
C147 ip VSS -29.73fF
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VPWR X a_1290_413# a_757_363#
+ a_1478_413# a_277_47# VNB VPB a_750_97# a_27_413# a_923_363# a_193_47# a_834_97#
+ a_247_21# a_668_97# a_193_413# a_27_47#
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=6.142e+11p pd=7.3e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=7.039e+11p ps=8e+06u w=420000u l=150000u
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=2.7965e+11p ps=3.21e+06u w=420000u l=150000u
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.8025e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=150000u
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_750_97# a_668_97# 0.11fF
C1 VPB S1 0.17fF
C2 S1 a_1478_413# 0.02fF
C3 S1 a_277_47# 0.06fF
C4 a_1290_413# S0 0.02fF
C5 a_247_21# X 0.01fF
C6 a_1290_413# a_668_97# 0.01fF
C7 a_247_21# a_750_97# 0.24fF
C8 VGND a_1478_413# 0.31fF
C9 VGND a_277_47# 0.54fF
C10 VPB VPWR 0.82fF
C11 VPWR a_1478_413# 0.34fF
C12 VPWR a_277_47# 0.26fF
C13 a_193_413# VPB 0.05fF
C14 a_193_413# a_1478_413# 0.00fF
C15 a_193_413# a_277_47# 0.12fF
C16 X a_834_97# 0.01fF
C17 A0 A1 0.17fF
C18 a_757_363# VPB 0.04fF
C19 a_834_97# a_750_97# 0.08fF
C20 a_757_363# a_1478_413# 0.01fF
C21 a_27_47# a_1478_413# 0.01fF
C22 a_757_363# a_277_47# 0.03fF
C23 a_1290_413# a_247_21# 0.04fF
C24 a_27_47# a_277_47# 0.14fF
C25 A0 A3 0.01fF
C26 S1 X 0.01fF
C27 S1 a_750_97# 0.06fF
C28 A3 A1 0.01fF
C29 a_1290_413# a_834_97# 0.02fF
C30 X VGND 0.08fF
C31 X VPWR 0.09fF
C32 VGND a_750_97# 0.22fF
C33 a_193_413# X 0.00fF
C34 VPWR a_750_97# 0.32fF
C35 a_1290_413# S1 0.22fF
C36 a_193_413# a_750_97# 0.01fF
C37 VPB a_1478_413# 0.11fF
C38 a_757_363# X 0.01fF
C39 a_27_47# X 0.00fF
C40 VPB a_277_47# 0.05fF
C41 A0 a_27_413# 0.08fF
C42 A0 A2 0.01fF
C43 a_277_47# a_1478_413# 0.18fF
C44 a_757_363# a_750_97# 0.21fF
C45 a_27_47# a_750_97# 0.01fF
C46 a_1290_413# VGND 0.17fF
C47 A2 A1 0.01fF
C48 a_27_413# A1 0.06fF
C49 a_1290_413# VPWR 0.17fF
C50 a_1290_413# a_193_413# 0.01fF
C51 a_923_363# VPWR 0.01fF
C52 a_1290_413# a_757_363# 0.03fF
C53 A2 A3 0.20fF
C54 A0 S0 0.03fF
C55 a_27_47# a_1290_413# 0.01fF
C56 a_923_363# a_757_363# 0.02fF
C57 S0 A1 0.02fF
C58 VPB X 0.05fF
C59 X a_1478_413# 0.22fF
C60 X a_277_47# 0.04fF
C61 VPB a_750_97# 0.08fF
C62 a_750_97# a_1478_413# 0.24fF
C63 a_750_97# a_277_47# 0.44fF
C64 A3 S0 0.04fF
C65 A3 a_668_97# 0.02fF
C66 A0 a_247_21# 0.12fF
C67 a_247_21# A1 0.05fF
C68 a_1290_413# VPB 0.13fF
C69 a_1290_413# a_1478_413# 0.15fF
C70 a_1290_413# a_277_47# 0.60fF
C71 a_247_21# A3 0.09fF
C72 a_27_413# S0 0.00fF
C73 A2 S0 0.03fF
C74 X a_750_97# 0.04fF
C75 A0 S1 0.01fF
C76 a_834_97# A3 0.05fF
C77 S1 A1 0.01fF
C78 A0 VGND 0.04fF
C79 A0 VPWR 0.04fF
C80 a_1290_413# X 0.03fF
C81 A0 a_193_413# 0.01fF
C82 S1 A3 0.05fF
C83 A1 VGND 0.03fF
C84 S0 a_668_97# 0.03fF
C85 a_27_413# a_247_21# 0.02fF
C86 a_1290_413# a_750_97# 0.23fF
C87 a_247_21# A2 0.04fF
C88 VPWR A1 0.04fF
C89 a_923_363# a_750_97# 0.00fF
C90 A0 a_27_47# 0.07fF
C91 A3 VGND 0.02fF
C92 A3 VPWR 0.02fF
C93 A2 a_834_97# 0.07fF
C94 a_27_47# A1 0.06fF
C95 a_247_21# S0 0.45fF
C96 a_247_21# a_668_97# 0.04fF
C97 a_757_363# A3 0.04fF
C98 S1 A2 0.09fF
C99 a_834_97# a_668_97# 0.11fF
C100 A0 VPB 0.10fF
C101 A0 a_1478_413# 0.00fF
C102 A2 VGND 0.02fF
C103 a_27_413# VGND 0.03fF
C104 A0 a_277_47# 0.11fF
C105 A2 VPWR 0.04fF
C106 a_27_413# VPWR 0.15fF
C107 a_27_413# a_193_413# 0.12fF
C108 VPB A1 0.14fF
C109 S1 S0 0.03fF
C110 A1 a_277_47# 0.02fF
C111 a_757_363# A2 0.05fF
C112 a_27_413# a_757_363# 0.01fF
C113 a_27_47# a_27_413# 0.04fF
C114 a_247_21# a_834_97# 0.05fF
C115 VPB A3 0.07fF
C116 A3 a_1478_413# 0.01fF
C117 S0 VGND 0.06fF
C118 A3 a_277_47# 0.02fF
C119 VGND a_668_97# 0.37fF
C120 VPWR S0 0.07fF
C121 VPWR a_668_97# 0.02fF
C122 a_193_413# S0 0.02fF
C123 S1 a_247_21# 0.04fF
C124 a_757_363# S0 0.04fF
C125 a_27_47# S0 0.02fF
C126 a_757_363# a_668_97# 0.02fF
C127 a_27_47# a_668_97# 0.02fF
C128 A0 a_750_97# 0.01fF
C129 a_247_21# VGND 0.23fF
C130 a_193_47# VGND 0.00fF
C131 a_247_21# VPWR 0.21fF
C132 A1 a_750_97# 0.01fF
C133 a_27_413# VPB 0.04fF
C134 a_27_413# a_1478_413# 0.00fF
C135 VPB A2 0.07fF
C136 A2 a_1478_413# 0.01fF
C137 a_27_413# a_277_47# 0.11fF
C138 A2 a_277_47# 0.02fF
C139 a_193_413# a_247_21# 0.17fF
C140 X A3 0.00fF
C141 A0 a_1290_413# 0.01fF
C142 A3 a_750_97# 0.05fF
C143 a_757_363# a_247_21# 0.06fF
C144 a_834_97# VGND 0.18fF
C145 a_27_47# a_247_21# 0.07fF
C146 a_834_97# VPWR 0.03fF
C147 a_27_47# a_193_47# 0.02fF
C148 a_1290_413# A1 0.01fF
C149 VPB S0 0.30fF
C150 S0 a_1478_413# 0.01fF
C151 S0 a_277_47# 0.07fF
C152 a_668_97# a_1478_413# 0.01fF
C153 S1 VGND 0.04fF
C154 a_757_363# a_834_97# 0.04fF
C155 a_668_97# a_277_47# 0.01fF
C156 a_27_47# a_834_97# 0.01fF
C157 S1 VPWR 0.05fF
C158 a_1290_413# A3 0.02fF
C159 A2 X 0.00fF
C160 a_27_413# X 0.00fF
C161 VPWR VGND 0.27fF
C162 a_27_413# a_750_97# 0.01fF
C163 A2 a_750_97# 0.03fF
C164 a_193_413# VGND 0.02fF
C165 VPB a_247_21# 0.23fF
C166 a_247_21# a_1478_413# 0.02fF
C167 a_193_413# VPWR 0.31fF
C168 a_247_21# a_277_47# 0.60fF
C169 a_757_363# VGND 0.03fF
C170 a_27_47# VGND 0.39fF
C171 a_757_363# VPWR 0.40fF
C172 a_27_47# VPWR 0.03fF
C173 X S0 0.00fF
C174 a_1290_413# A2 0.03fF
C175 a_1290_413# a_27_413# 0.00fF
C176 a_193_413# a_757_363# 0.03fF
C177 X a_668_97# 0.00fF
C178 a_27_47# a_193_413# 0.02fF
C179 a_834_97# a_1478_413# 0.01fF
C180 S0 a_750_97# 0.16fF
C181 a_834_97# a_277_47# 0.05fF
C182 VGND VNB 1.06fF
C183 X VNB 0.05fF
C184 S1 VNB 0.21fF
C185 A2 VNB 0.08fF
C186 A3 VNB 0.09fF
C187 S0 VNB 0.34fF
C188 VPWR VNB 0.41fF
C189 A0 VNB 0.10fF
C190 A1 VNB 0.15fF
C191 VPB VNB 1.93fF
C192 a_834_97# VNB 0.02fF
C193 a_668_97# VNB 0.03fF
C194 a_27_47# VNB 0.03fF
C195 a_1478_413# VNB 0.11fF
C196 a_1290_413# VNB 0.15fF
C197 a_750_97# VNB 0.03fF
C198 a_277_47# VNB 0.07fF
C199 a_247_21# VNB 0.27fF
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_XAYTAL a_n129_n203# a_n173_n100# w_n311_n319#
+ VSUBS
X0 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=1.28e+12p pd=1.056e+07u as=0p ps=0u w=1e+06u l=150000u
X1 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n173_n100# a_n129_n203# 0.30fF
C1 a_n129_n203# w_n311_n319# 0.51fF
C2 a_n173_n100# w_n311_n319# 0.42fF
C3 w_n311_n319# VSUBS 1.19fF
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X a_110_47# VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 A a_110_47# 0.51fF
C1 a_110_47# X 2.36fF
C2 VGND VPWR 0.28fF
C3 VPB VPWR 0.78fF
C4 A VPWR 0.07fF
C5 VPWR X 2.96fF
C6 A VGND 0.10fF
C7 VGND X 1.95fF
C8 A VPB 0.23fF
C9 VPB X 0.03fF
C10 A X 0.00fF
C11 a_110_47# VPWR 0.98fF
C12 VGND a_110_47# 0.78fF
C13 a_110_47# VPB 0.81fF
C14 VGND VNB 1.05fF
C15 X VNB 0.10fF
C16 VPWR VNB 0.39fF
C17 A VNB 0.43fF
C18 VPB VNB 1.85fF
C19 a_110_47# VNB 1.28fF
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
C0 VPB VGND 0.25fF
C1 VPWR VGND 0.82fF
C2 VPWR VPB 0.27fF
C3 VPWR VNB 0.41fF
C4 VGND VNB 0.37fF
C5 VPB VNB 0.43fF
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
C0 VPWR VPB 0.37fF
C1 VGND VPWR 1.92fF
C2 VGND VPB 0.55fF
C3 VPWR VNB 0.86fF
C4 VGND VNB 0.56fF
C5 VPB VNB 0.78fF
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VPWR X VNB VPB a_283_47# a_390_47#
+ a_27_47#
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=6.517e+11p ps=5.37e+06u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=4.027e+11p pd=3.97e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
C0 A a_283_47# 0.02fF
C1 VPWR A 0.02fF
C2 VGND X 0.14fF
C3 A X 0.00fF
C4 a_27_47# a_390_47# 0.05fF
C5 A VGND 0.02fF
C6 a_27_47# a_283_47# 0.18fF
C7 a_27_47# VPWR 0.31fF
C8 a_27_47# X 0.02fF
C9 a_27_47# VGND 0.24fF
C10 a_390_47# VPB 0.06fF
C11 a_27_47# A 0.29fF
C12 a_283_47# VPB 0.12fF
C13 VPWR VPB 0.32fF
C14 X VPB 0.05fF
C15 A VPB 0.06fF
C16 a_27_47# VPB 0.16fF
C17 a_283_47# a_390_47# 0.44fF
C18 VPWR a_390_47# 0.16fF
C19 VPWR a_283_47# 0.17fF
C20 a_390_47# X 0.12fF
C21 a_390_47# VGND 0.14fF
C22 a_283_47# X 0.04fF
C23 a_283_47# VGND 0.14fF
C24 VPWR X 0.19fF
C25 A a_390_47# 0.01fF
C26 VPWR VGND 0.11fF
C27 VGND VNB 0.43fF
C28 X VNB 0.05fF
C29 VPWR VNB 0.16fF
C30 A VNB 0.13fF
C31 VPB VNB 0.78fF
C32 a_390_47# VNB 0.10fF
C33 a_283_47# VNB 0.18fF
C34 a_27_47# VNB 0.18fF
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB a_27_47#
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 Y VGND 0.13fF
C1 A VPWR 0.09fF
C2 VPWR B 0.12fF
C3 Y A 0.35fF
C4 Y B 0.30fF
C5 VGND a_27_47# 0.77fF
C6 A a_27_47# 0.10fF
C7 a_27_47# B 0.33fF
C8 Y VPWR 1.44fF
C9 A VPB 0.18fF
C10 VPB B 0.21fF
C11 VGND A 0.08fF
C12 VGND B 0.10fF
C13 VPWR a_27_47# 0.07fF
C14 Y a_27_47# 0.41fF
C15 A B 0.16fF
C16 VPB VPWR 0.43fF
C17 Y VPB 0.02fF
C18 VGND VPWR 0.12fF
C19 VGND VNB 0.48fF
C20 Y VNB 0.01fF
C21 VPWR VNB 0.18fF
C22 A VNB 0.26fF
C23 B VNB 0.30fF
C24 VPB VNB 0.87fF
C25 a_27_47# VNB 0.06fF
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
C0 VGND VPWR 0.54fF
C1 VPB VPWR 0.24fF
C2 VPB VGND 0.16fF
C3 VPWR VNB 0.28fF
C4 VGND VNB 0.31fF
C5 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__dfxbp_1 CLK D VGND VPWR Q Q_N a_975_413# a_891_413# VNB VPB
+ a_466_413# a_592_47# a_1059_315# a_193_47# a_561_413# a_634_159# a_381_47# a_1017_47#
+ a_1490_369# a_27_47#
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=9.432e+11p ps=1.006e+07u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.32905e+12p pd=1.228e+07u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X6 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1059_315# a_1490_369# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X17 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23 Q_N a_1490_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q_N a_1490_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 VPWR a_1059_315# a_1490_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
C0 a_1059_315# a_1490_369# 0.18fF
C1 a_381_47# D 0.21fF
C2 VGND a_381_47# 0.09fF
C3 VPB D 0.13fF
C4 VGND a_592_47# 0.00fF
C5 a_634_159# a_466_413# 0.36fF
C6 a_466_413# a_1490_369# 0.02fF
C7 VPWR D 0.03fF
C8 VGND VPWR 0.26fF
C9 a_634_159# CLK 0.01fF
C10 a_1490_369# CLK 0.00fF
C11 a_193_47# a_634_159# 0.21fF
C12 a_193_47# a_1490_369# 0.03fF
C13 a_634_159# a_27_47# 0.29fF
C14 Q_N a_1059_315# 0.03fF
C15 a_1490_369# a_27_47# 0.03fF
C16 a_891_413# a_634_159# 0.10fF
C17 a_891_413# a_1490_369# 0.04fF
C18 Q_N a_466_413# 0.01fF
C19 a_1059_315# a_466_413# 0.05fF
C20 Q a_634_159# 0.02fF
C21 VPB a_381_47# 0.03fF
C22 Q a_1490_369# 0.31fF
C23 a_561_413# VPWR 0.01fF
C24 Q_N CLK 0.00fF
C25 a_1059_315# CLK 0.01fF
C26 a_193_47# Q_N 0.02fF
C27 VPWR a_381_47# 0.13fF
C28 a_891_413# a_1017_47# 0.01fF
C29 VPB VPWR 0.73fF
C30 a_193_47# a_1059_315# 0.13fF
C31 Q_N a_27_47# 0.02fF
C32 a_634_159# D 0.04fF
C33 a_1059_315# a_27_47# 0.14fF
C34 VGND a_634_159# 0.18fF
C35 a_1490_369# D 0.01fF
C36 a_975_413# VPWR 0.01fF
C37 VGND a_1490_369# 0.12fF
C38 a_466_413# CLK 0.01fF
C39 a_891_413# Q_N 0.02fF
C40 a_193_47# a_466_413# 0.20fF
C41 a_891_413# a_1059_315# 0.44fF
C42 a_466_413# a_27_47# 0.51fF
C43 Q Q_N 0.05fF
C44 Q a_1059_315# 0.19fF
C45 a_891_413# a_466_413# 0.04fF
C46 VGND a_1017_47# 0.00fF
C47 a_193_47# CLK 0.06fF
C48 a_27_47# CLK 0.33fF
C49 a_193_47# a_27_47# 1.69fF
C50 Q a_466_413# 0.02fF
C51 Q_N D 0.00fF
C52 VGND Q_N 0.11fF
C53 a_891_413# CLK 0.01fF
C54 a_1059_315# D 0.02fF
C55 VGND a_1059_315# 0.22fF
C56 a_193_47# a_891_413# 0.38fF
C57 a_891_413# a_27_47# 0.09fF
C58 Q CLK 0.00fF
C59 a_634_159# a_381_47# 0.03fF
C60 a_466_413# D 0.03fF
C61 a_1490_369# a_381_47# 0.01fF
C62 a_634_159# VPB 0.08fF
C63 VGND a_466_413# 0.15fF
C64 Q a_193_47# 0.03fF
C65 a_1490_369# VPB 0.06fF
C66 Q a_27_47# 0.03fF
C67 a_634_159# VPWR 0.21fF
C68 a_1490_369# VPWR 0.29fF
C69 CLK D 0.04fF
C70 Q a_891_413# 0.04fF
C71 VGND CLK 0.04fF
C72 a_193_47# D 0.30fF
C73 a_193_47# VGND 0.24fF
C74 a_27_47# D 0.17fF
C75 VGND a_27_47# 0.30fF
C76 a_891_413# D 0.01fF
C77 Q_N a_381_47# 0.01fF
C78 VGND a_891_413# 0.18fF
C79 Q_N VPB 0.05fF
C80 a_1059_315# a_381_47# 0.01fF
C81 a_1059_315# VPB 0.24fF
C82 a_466_413# a_561_413# 0.01fF
C83 Q D 0.00fF
C84 Q VGND 0.14fF
C85 Q_N VPWR 0.25fF
C86 a_466_413# a_381_47# 0.09fF
C87 a_1059_315# VPWR 0.37fF
C88 a_466_413# VPB 0.08fF
C89 a_466_413# a_592_47# 0.01fF
C90 a_466_413# VPWR 0.31fF
C91 VGND D 0.05fF
C92 CLK a_381_47# 0.01fF
C93 CLK VPB 0.14fF
C94 a_634_159# a_1490_369# 0.02fF
C95 a_193_47# a_381_47# 0.22fF
C96 a_193_47# VPB 0.21fF
C97 a_27_47# a_381_47# 0.16fF
C98 a_27_47# VPB 0.30fF
C99 CLK VPWR 0.03fF
C100 a_193_47# VPWR 0.37fF
C101 a_891_413# a_381_47# 0.02fF
C102 a_891_413# VPB 0.08fF
C103 a_27_47# VPWR 0.60fF
C104 a_891_413# a_975_413# 0.02fF
C105 Q a_381_47# 0.01fF
C106 Q VPB 0.02fF
C107 a_891_413# VPWR 0.20fF
C108 Q_N a_634_159# 0.01fF
C109 Q_N a_1490_369# 0.14fF
C110 a_1059_315# a_634_159# 0.06fF
C111 Q VPWR 0.24fF
C112 Q_N VNB 0.05fF
C113 Q VNB 0.01fF
C114 VGND VNB 0.95fF
C115 VPWR VNB 0.37fF
C116 D VNB 0.12fF
C117 CLK VNB 0.18fF
C118 VPB VNB 1.76fF
C119 a_381_47# VNB 0.03fF
C120 a_1490_369# VNB 0.09fF
C121 a_891_413# VNB 0.12fF
C122 a_1059_315# VNB 0.24fF
C123 a_466_413# VNB 0.11fF
C124 a_634_159# VNB 0.12fF
C125 a_193_47# VNB 0.21fF
C126 a_27_47# VNB 0.31fF
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 B VGND 0.06fF
C1 Y VGND 0.21fF
C2 VGND A 0.02fF
C3 B VPWR 0.06fF
C4 Y VPWR 0.40fF
C5 A VPWR 0.05fF
C6 B VPB 0.06fF
C7 VGND VPWR 0.05fF
C8 VPB Y 0.02fF
C9 VPB A 0.06fF
C10 Y a_113_47# 0.01fF
C11 B Y 0.05fF
C12 a_113_47# VGND 0.01fF
C13 B A 0.07fF
C14 Y A 0.11fF
C15 VPB VPWR 0.24fF
C16 VGND VNB 0.23fF
C17 Y VNB 0.05fF
C18 VPWR VNB 0.06fF
C19 A VNB 0.10fF
C20 B VNB 0.10fF
C21 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 VGND A 0.05fF
C1 Y VPWR 0.35fF
C2 Y VPB 0.00fF
C3 Y A 0.26fF
C4 VPWR VPB 0.23fF
C5 VPWR A 0.04fF
C6 Y VGND 0.17fF
C7 VPB A 0.14fF
C8 VPWR VGND 0.04fF
C9 VGND VNB 0.23fF
C10 Y VNB 0.04fF
C11 VPWR VNB 0.06fF
C12 A VNB 0.24fF
C13 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB a_505_21# a_535_374# a_439_47#
+ a_218_47# a_76_199# a_218_374#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 X a_505_21# 0.02fF
C1 a_76_199# VPB 0.08fF
C2 S VPB 0.24fF
C3 A1 A0 0.41fF
C4 VGND A1 0.12fF
C5 a_76_199# A0 0.14fF
C6 A1 a_439_47# 0.00fF
C7 A1 VPWR 0.04fF
C8 A0 S 0.09fF
C9 VGND a_76_199# 0.24fF
C10 a_76_199# VPWR 0.15fF
C11 VGND S 0.07fF
C12 A0 VPB 0.08fF
C13 S VPWR 0.64fF
C14 A1 X 0.04fF
C15 VPWR VPB 0.44fF
C16 a_76_199# X 0.18fF
C17 S X 0.08fF
C18 X VPB 0.06fF
C19 A1 a_505_21# 0.16fF
C20 VGND A0 0.08fF
C21 A0 VPWR 0.01fF
C22 A0 a_439_47# 0.01fF
C23 a_218_47# a_76_199# 0.01fF
C24 a_76_199# a_505_21# 0.04fF
C25 S a_505_21# 0.26fF
C26 VGND a_439_47# 0.01fF
C27 VGND VPWR 0.12fF
C28 VPB a_505_21# 0.09fF
C29 A0 X 0.02fF
C30 VGND X 0.09fF
C31 VPWR X 0.23fF
C32 A0 a_505_21# 0.08fF
C33 S a_535_374# 0.01fF
C34 a_76_199# a_218_374# 0.00fF
C35 a_218_374# S 0.01fF
C36 A1 a_76_199# 0.41fF
C37 VGND a_218_47# 0.01fF
C38 VGND a_505_21# 0.16fF
C39 A1 S 0.25fF
C40 VPWR a_505_21# 0.12fF
C41 a_76_199# S 0.54fF
C42 A1 VPB 0.06fF
C43 VGND VNB 0.48fF
C44 A1 VNB 0.09fF
C45 A0 VNB 0.08fF
C46 S VNB 0.17fF
C47 VPWR VNB 0.18fF
C48 X VNB 0.06fF
C49 VPB VNB 0.87fF
C50 a_505_21# VNB 0.15fF
C51 a_76_199# VNB 0.11fF
.ends

.subckt clock_v2 clk p2d_b p2d p2_b p2 p1d_b p1d p1_b p1 Ad_b Ad A_b A Bd_b Bd B_b
+ B sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__mux2_1_0/a_439_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47#
+ sky130_fd_sc_hd__mux2_1_0/a_218_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47#
+ sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__mux2_1_0/a_218_374#
+ sky130_fd_sc_hd__clkinv_1_2/Y sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__dfxbp_1_1/a_27_47#
+ sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A
+ sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47#
+ sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__nand2_4_2/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__nand2_4_0/B
+ sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47#
+ sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkinv_1_1/Y
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_1_3/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__dfxbp_1_1/D
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxbp_1_1/a_592_47# sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
+ sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__mux2_1_0/a_505_21#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__mux2_1_0/a_535_374# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47#
+ sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47#
+ sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_131/A
+ sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47#
+ sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A
+ sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_20/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__nand2_4_0/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkinv_4_7/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_3/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A
+ sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
+ sky130_fd_sc_hd__nand2_1_2/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_2/Y
Xsky130_fd_sc_hd__clkbuf_16_11 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD p1d_b sky130_fd_sc_hd__clkbuf_16_11/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_226 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_204 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_12 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD p2d_b sky130_fd_sc_hd__clkbuf_16_12/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_13 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD p2d sky130_fd_sc_hd__clkbuf_16_13/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_217 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_0 sky130_fd_sc_hd__clkinv_1_0/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_14 sky130_fd_sc_hd__clkinv_4_10/Y VSS VDD p2_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_10 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_4_10/Y
+ sky130_fd_sc_hd__clkinv_4_10/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_1 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_140 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_162 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_15 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD p2 sky130_fd_sc_hd__clkbuf_16_15/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_11 sky130_fd_sc_hd__nand2_4_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/A
+ sky130_fd_sc_hd__clkinv_4_11/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_2 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_3 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS VDD sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/A
+ sky130_fd_sc_hd__clkinv_4_0/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_165 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_2 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__nand2_4_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__nand2_4_2/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_190 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_5 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__clkinv_4_1/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_111 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_166 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_180 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_4_3 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__nand2_4_3/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_6 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__clkinv_4_2/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__clkinv_4_3/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_168 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_157 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_193 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_8 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__clkinv_4_4/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_158 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_172 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_183 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_5/Y
+ sky130_fd_sc_hd__clkinv_4_5/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_159 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_195 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_140 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_162 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_6 sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/A
+ sky130_fd_sc_hd__clkinv_4_6/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_190 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_196 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_90 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_7 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__clkinv_4_7/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_191 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_180 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_186 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_80 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_8 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__clkinv_4_8/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_165 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_198 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_92 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_9 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__clkinv_4_9/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_193 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_182 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_111 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_166 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_188 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_71 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_82 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_93 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_0 p2 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__mux2_1_0/S
+ sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__dfxbp_1_0/a_975_413# sky130_fd_sc_hd__dfxbp_1_0/a_891_413#
+ VSS VDD sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_592_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__dfxbp_1_0/a_1017_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_172 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_150 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_178 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_189 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_50 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_61 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_1 clk sky130_fd_sc_hd__dfxbp_1_1/D VSS VDD sky130_fd_sc_hd__nand2_1_1/A
+ sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__dfxbp_1_1/a_975_413# sky130_fd_sc_hd__dfxbp_1_1/a_891_413#
+ VSS VDD sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_592_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# sky130_fd_sc_hd__dfxbp_1_1/a_1017_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_195 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_184 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_173 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_140 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_162 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_157 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_168 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_179 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_73 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_84 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_95 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_141 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_196 sky130_fd_sc_hd__clkinv_1_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_174 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_152 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_163 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_158 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_52 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_63 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_96 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_197 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_186 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_164 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_131 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_142 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD B sky130_fd_sc_hd__clkbuf_16_0/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_159 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_42 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_20 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_31 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_75 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_86 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_97 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_1/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_198 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_187 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_121 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_132 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_154 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD Bd sky130_fd_sc_hd__clkbuf_16_1/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_10 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_54 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_32 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_65 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_87 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_199 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_3/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_177 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_100 sky130_fd_sc_hd__clkinv_1_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_122 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD
+ sky130_fd_sc_hd__nand2_1_4/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD B_b sky130_fd_sc_hd__clkbuf_16_2/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_22 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_44 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_11 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_77 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_99 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_178 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_167 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_112 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_101 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_123 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_134 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD Bd_b sky130_fd_sc_hd__clkbuf_16_3/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_56 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_34 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_67 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_78 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_89 sky130_fd_sc_hd__clkinv_1_1/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_157 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_102 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_113 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_146 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_168 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_4 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD Ad_b sky130_fd_sc_hd__clkbuf_16_4/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_24 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_13 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_68 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_0/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_169 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_2/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_103 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_2/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_125 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_136 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_147 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_158 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_5 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD Ad sky130_fd_sc_hd__clkbuf_16_5/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_25 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_47 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_58 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_36 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_69 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_104 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_159 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_6 sky130_fd_sc_hd__clkinv_4_4/Y VSS VDD A_b sky130_fd_sc_hd__clkbuf_16_6/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_15 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_48 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_59 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_116 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_127 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_138 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_149 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_7 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD A sky130_fd_sc_hd__clkbuf_16_7/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_49 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_1/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_27 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_38 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_250 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_117 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_8 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD p1 sky130_fd_sc_hd__clkbuf_16_8/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_17 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_39 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_107 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_118 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_129 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_9 sky130_fd_sc_hd__clkinv_4_7/Y VSS VDD p1_b sky130_fd_sc_hd__clkbuf_16_9/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_1_0/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_18 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_29 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_108 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__nand2_1_2/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_1_1/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_109 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_1_3/A clk VSS VDD sky130_fd_sc_hd__nand2_4_3/A
+ VSS VDD sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_254 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_232 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_210 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/B
+ VSS VDD sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1_4/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_211 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_200 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux2_1_0 Ad_b Bd_b sky130_fd_sc_hd__mux2_1_0/S VSS VDD sky130_fd_sc_hd__mux2_1_0/X
+ VSS VDD sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/a_535_374#
+ sky130_fd_sc_hd__mux2_1_0/a_439_47# sky130_fd_sc_hd__mux2_1_0/a_218_47# sky130_fd_sc_hd__mux2_1_0/a_76_199#
+ sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_234 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_246 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_224 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_10 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD p1d sky130_fd_sc_hd__clkbuf_16_10/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_6 clk VSS VDD sky130_fd_sc_hd__nand2_1_2/A VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_247 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_225 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
C0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C1 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C2 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C3 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C4 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.05fF
C5 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C6 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.02fF
C7 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C8 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C9 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C10 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C11 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.13fF
C12 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C13 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.14fF
C14 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C15 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C16 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C17 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C18 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C19 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VDD 0.12fF
C20 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_4/B 0.23fF
C21 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C22 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C23 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C24 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C25 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C26 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.05fF
C27 VDD sky130_fd_sc_hd__nand2_1_0/B 1.07fF
C28 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C29 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C30 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C31 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C32 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C33 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C34 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C35 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C36 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C37 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C38 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.02fF
C39 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.04fF
C40 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.04fF
C41 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.04fF
C42 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.04fF
C43 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C44 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C45 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C46 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clk 0.01fF
C47 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C48 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C49 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C50 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C51 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C52 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C53 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C54 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C55 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.02fF
C56 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.04fF
C57 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.03fF
C58 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C59 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.03fF
C60 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C61 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C62 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.09fF
C63 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0.00fF
C64 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.02fF
C65 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.04fF
C66 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.02fF
C67 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C68 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C69 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.01fF
C70 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.01fF
C71 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VDD 5.72fF
C72 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.02fF
C73 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0.08fF
C74 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C75 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C76 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C77 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C78 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C79 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.11fF
C80 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.31fF
C81 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C82 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C83 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C84 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.02fF
C85 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.04fF
C86 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.09fF
C87 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C88 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C89 p2 sky130_fd_sc_hd__nand2_4_1/Y 0.00fF
C90 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C91 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# Ad_b 0.01fF
C92 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C93 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C94 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C95 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.04fF
C96 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.04fF
C97 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C98 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C99 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C100 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C101 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C102 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VDD 0.23fF
C103 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C104 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C105 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.01fF
C106 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# Bd -0.04fF
C107 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# VDD 0.15fF
C108 B sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.06fF
C109 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# Bd 0.06fF
C110 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# B -0.04fF
C111 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C112 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.05fF
C113 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C114 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C115 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# VDD 0.35fF
C116 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C117 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C118 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C119 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C120 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.00fF
C121 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C122 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C123 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C124 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/A 1.18fF
C125 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C126 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.04fF
C127 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C128 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.06fF
C129 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C130 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C131 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.04fF
C132 p2 VDD 4.22fF
C133 p2d p2 0.20fF
C134 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C135 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.04fF
C136 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.04fF
C137 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C138 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C139 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C140 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.04fF
C141 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C142 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C143 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C144 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C145 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C146 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkinv_4_1/A 0.11fF
C147 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C148 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.04fF
C149 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C150 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C151 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C152 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C153 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__dfxbp_1_0/a_1017_47# -0.00fF
C154 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/A 0.70fF
C155 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C156 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C157 sky130_fd_sc_hd__clkinv_1_3/Y VDD -1.28fF
C158 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C159 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C160 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C161 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.04fF
C162 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.04fF
C163 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.04fF
C164 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Bd_b 0.07fF
C165 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.03fF
C166 sky130_fd_sc_hd__nand2_1_1/A Bd_b 1.60fF
C167 sky130_fd_sc_hd__clkinv_4_5/Y A 0.00fF
C168 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C169 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.12fF
C170 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C171 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.15fF
C172 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.30fF
C173 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C174 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C175 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.05fF
C176 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C177 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.19fF
C178 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C179 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C180 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 1.10fF
C181 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C182 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.02fF
C183 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C184 p2 sky130_fd_sc_hd__nand2_4_3/B 0.06fF
C185 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# VDD 0.15fF
C186 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C187 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C188 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# VDD 0.17fF
C189 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.04fF
C190 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.04fF
C191 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C192 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C193 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C194 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.04fF
C195 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.04fF
C196 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C197 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C198 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VDD 0.36fF
C199 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.04fF
C200 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.03fF
C201 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C202 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C203 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.00fF
C204 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.09fF
C205 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C206 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C207 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C208 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C209 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C210 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C211 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C212 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C213 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C214 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.05fF
C215 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C216 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C217 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.02fF
C218 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C219 p1d_b sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.12fF
C220 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VDD 0.30fF
C221 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.04fF
C222 A_b sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.12fF
C223 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# A 0.12fF
C224 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.06fF
C225 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.02fF
C226 p2 sky130_fd_sc_hd__nand2_4_3/A 0.34fF
C227 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VDD 0.15fF
C228 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.04fF
C229 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C230 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C231 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C232 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C233 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C234 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C235 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.01fF
C236 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C237 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# VDD 0.11fF
C238 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C239 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.04fF
C240 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# VDD 0.30fF
C241 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.06fF
C242 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C243 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C244 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C245 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C246 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C247 sky130_fd_sc_hd__clkinv_4_8/Y VDD 0.77fF
C248 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.08fF
C249 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.01fF
C250 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C251 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C252 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# VDD 0.16fF
C253 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C254 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_4_3/A 0.73fF
C255 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C256 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C257 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C258 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X -0.00fF
C259 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VDD 0.12fF
C260 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C261 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0.01fF
C262 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 1.56fF
C263 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C264 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.02fF
C265 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.14fF
C266 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 2.25fF
C267 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_1/A 0.37fF
C268 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C269 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.16fF
C270 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C271 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.02fF
C272 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C273 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C274 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.10fF
C275 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 2.22fF
C276 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# VDD 0.21fF
C277 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.03fF
C278 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C279 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C280 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C281 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.02fF
C282 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.02fF
C283 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# -0.00fF
C284 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# VDD 0.21fF
C285 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C286 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C287 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C288 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.01fF
C289 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C290 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C291 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C292 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C293 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C294 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.09fF
C295 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.15fF
C296 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C297 VDD sky130_fd_sc_hd__nand2_1_1/B 1.41fF
C298 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.16fF
C299 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.30fF
C300 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.11fF
C301 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# p1_b 0.07fF
C302 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C303 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.15fF
C304 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.10fF
C305 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.35fF
C306 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C307 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C308 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.18fF
C309 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C310 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.12fF
C311 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C312 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.07fF
C313 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.02fF
C314 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C315 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C316 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C317 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C318 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.09fF
C319 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C320 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.02fF
C321 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C322 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.06fF
C323 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.11fF
C324 Bd_b sky130_fd_sc_hd__clkinv_4_2/Y 0.10fF
C325 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C326 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.05fF
C327 VDD sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.43fF
C328 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C329 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C330 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.12fF
C331 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C332 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X -0.00fF
C333 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C334 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VDD 0.22fF
C335 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_1_0/A 0.06fF
C336 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.02fF
C337 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.02fF
C338 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.01fF
C339 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.02fF
C340 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C341 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C342 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C343 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C344 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C345 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.05fF
C346 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VDD 1.46fF
C347 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C348 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C349 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C350 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.08fF
C351 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Ad_b 0.12fF
C352 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__nand2_4_2/A 2.12fF
C353 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# VDD 0.15fF
C354 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.31fF
C355 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.04fF
C356 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# VDD 0.19fF
C357 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# VDD 0.15fF
C358 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C359 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C360 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.08fF
C361 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C362 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C363 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C364 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# -0.00fF
C365 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C366 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C367 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C368 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C369 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.01fF
C370 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.05fF
C371 p2d sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C372 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__nand2_4_0/Y 0.16fF
C373 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.05fF
C374 sky130_fd_sc_hd__nand2_4_3/Y VDD 9.78fF
C375 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.02fF
C376 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.02fF
C377 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.15fF
C378 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C379 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C380 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C381 sky130_fd_sc_hd__clkinv_4_1/w_82_21# sky130_fd_sc_hd__clkinv_4_1/A 0.03fF
C382 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C383 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C384 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# VDD 0.16fF
C385 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.01fF
C386 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C387 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C388 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C389 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.00fF
C390 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# VDD 0.34fF
C391 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C392 sky130_fd_sc_hd__nand2_4_2/Y VDD 9.42fF
C393 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C394 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_1_3/A 0.04fF
C395 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.05fF
C396 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C397 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C398 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C399 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.00fF
C400 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C401 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.02fF
C402 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C403 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C404 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C405 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C406 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.13fF
C407 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.04fF
C408 p2 Ad_b 1.13fF
C409 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.05fF
C410 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.15fF
C411 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C412 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C413 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C414 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C415 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.00fF
C416 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.00fF
C417 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C418 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C419 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C420 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C421 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.05fF
C422 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C423 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.03fF
C424 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C425 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C426 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B 0.16fF
C427 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.09fF
C428 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.21fF
C429 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0.06fF
C430 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C431 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C432 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C433 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C434 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C435 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# VDD 0.15fF
C436 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.02fF
C437 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# VDD 0.15fF
C438 p1d_b p2d_b 0.11fF
C439 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.12fF
C440 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C441 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C442 sky130_fd_sc_hd__clkinv_4_10/Y VDD -0.41fF
C443 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# p2 0.02fF
C444 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C445 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C446 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C447 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C448 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C449 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C450 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C451 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C452 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.03fF
C453 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.03fF
C454 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C455 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C456 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C457 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C458 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C459 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.08fF
C460 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C461 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C462 Bd VDD 1.51fF
C463 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.02fF
C464 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C465 B VDD 1.52fF
C466 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.02fF
C467 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.15fF
C468 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.02fF
C469 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.02fF
C470 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.02fF
C471 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C472 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C473 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.29fF
C474 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A 0.62fF
C475 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C476 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.03fF
C477 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# -0.01fF
C478 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C479 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C480 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C481 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C482 sky130_fd_sc_hd__mux2_1_0/a_439_47# Ad_b 0.02fF
C483 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C484 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C485 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C486 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C487 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X -0.00fF
C488 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C489 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C490 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C491 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C492 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C493 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.07fF
C494 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C495 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C496 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C497 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C498 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C499 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C500 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.04fF
C501 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C502 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C503 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C504 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C505 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C506 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C507 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.02fF
C508 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C509 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 1.41fF
C510 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C511 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C512 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A -0.00fF
C513 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# -0.00fF
C514 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.03fF
C515 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C516 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C517 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.08fF
C518 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.00fF
C519 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C520 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C521 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C522 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.02fF
C523 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C524 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C525 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VDD 1.38fF
C526 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.08fF
C527 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C528 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C529 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.05fF
C530 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.05fF
C531 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.08fF
C532 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.02fF
C533 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A -0.00fF
C534 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.01fF
C535 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C536 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C537 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C538 p2 sky130_fd_sc_hd__nand2_4_1/B 0.04fF
C539 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_1_1/A 0.05fF
C540 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.18fF
C541 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C542 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C543 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C544 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# -0.00fF
C545 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.34fF
C546 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.19fF
C547 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C548 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C549 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C550 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# Bd_b 0.02fF
C551 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# Ad_b 0.00fF
C552 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/S 0.06fF
C553 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.08fF
C554 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C555 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.01fF
C556 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C557 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C558 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C559 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C560 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C561 p2d sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.06fF
C562 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# VDD 0.15fF
C563 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.02fF
C564 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.02fF
C565 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C566 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.03fF
C567 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VDD 0.51fF
C568 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C569 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C570 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C571 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.18fF
C572 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.03fF
C573 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C574 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# VDD 0.23fF
C575 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C576 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C577 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C578 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C579 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# VDD 0.31fF
C580 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C581 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.19fF
C582 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.07fF
C583 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C584 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C585 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C586 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.03fF
C587 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C588 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C589 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C590 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_2/Y 0.68fF
C591 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A -0.00fF
C592 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C593 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.15fF
C594 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C595 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C596 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C597 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C598 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C599 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C600 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C601 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.08fF
C602 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C603 sky130_fd_sc_hd__clkinv_1_3/A clk 0.00fF
C604 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.02fF
C605 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C606 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C607 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.04fF
C608 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.04fF
C609 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.01fF
C610 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C611 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C612 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C613 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C614 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C615 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y 0.32fF
C616 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C617 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# p2 0.06fF
C618 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C619 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.03fF
C620 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.03fF
C621 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C622 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C623 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C624 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C625 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.06fF
C626 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C627 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C628 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C629 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C630 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.11fF
C631 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C632 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.08fF
C633 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.15fF
C634 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C635 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C636 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C637 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C638 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.01fF
C639 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.02fF
C640 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.12fF
C641 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C642 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C643 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C644 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.40fF
C645 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.09fF
C646 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C647 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.02fF
C648 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C649 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.97fF
C650 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Ad -0.01fF
C651 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD 1.41fF
C652 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.07fF
C653 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.00fF
C654 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.00fF
C655 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A -0.00fF
C656 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C657 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C658 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# VDD 0.15fF
C659 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C660 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C661 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.02fF
C662 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C663 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C664 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# p2 0.12fF
C665 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C666 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.00fF
C667 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.00fF
C668 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# VDD 0.21fF
C669 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C670 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C671 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.22fF
C672 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# 0.01fF
C673 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.07fF
C674 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_4/B 0.40fF
C675 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD 1.01fF
C676 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.11fF
C677 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.02fF
C678 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.04fF
C679 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.04fF
C680 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C681 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C682 sky130_fd_sc_hd__nand2_4_3/Y Ad_b 0.00fF
C683 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C684 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VDD 0.15fF
C685 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VDD 0.36fF
C686 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C687 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# 0.05fF
C688 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# -0.01fF
C689 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C690 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C691 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.03fF
C692 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C693 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C694 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A -0.00fF
C695 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.07fF
C696 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C697 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VDD 0.29fF
C698 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# VDD 0.15fF
C699 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.04fF
C700 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.04fF
C701 sky130_fd_sc_hd__nand2_4_1/Y Ad 0.00fF
C702 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C703 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C704 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# VDD 0.35fF
C705 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.04fF
C706 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_3/Y 0.01fF
C707 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C708 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C709 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C710 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.12fF
C711 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C712 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C713 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C714 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.62fF
C715 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VDD 0.10fF
C716 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.02fF
C717 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.07fF
C718 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C719 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 1.14fF
C720 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/B 0.07fF
C721 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C722 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C723 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C724 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__nand2_1_1/A 0.05fF
C725 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C726 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VDD 0.38fF
C727 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.07fF
C728 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# -0.01fF
C729 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C730 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VDD 0.16fF
C731 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.14fF
C732 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C733 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C734 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C735 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.08fF
C736 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C737 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# VDD 0.15fF
C738 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2d 0.12fF
C739 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A -0.00fF
C740 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VDD 0.40fF
C741 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_1_4/B 0.07fF
C742 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C743 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# VDD 0.09fF
C744 VDD Ad 1.63fF
C745 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# VDD 0.26fF
C746 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C747 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C748 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C749 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C750 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C751 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C752 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C753 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C754 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C755 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.05fF
C756 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C757 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.15fF
C758 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_1_2/B 0.00fF
C759 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C760 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/A 0.46fF
C761 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C762 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C763 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C764 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C765 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.15fF
C766 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.07fF
C767 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C768 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__nand2_1_4/B 0.03fF
C769 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.15fF
C770 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C771 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.22fF
C772 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C773 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C774 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C775 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.06fF
C776 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.39fF
C777 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C778 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C779 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.03fF
C780 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C781 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C782 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.07fF
C783 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C784 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C785 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.06fF
C786 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 1.21fF
C787 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A -0.00fF
C788 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C789 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C790 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_1/B 0.00fF
C791 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.05fF
C792 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C793 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.18fF
C794 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.19fF
C795 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C796 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C797 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C798 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C799 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C800 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C801 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C802 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.04fF
C803 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C804 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C805 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Bd_b 0.14fF
C806 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.18fF
C807 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# VDD 0.15fF
C808 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.33fF
C809 VDD sky130_fd_sc_hd__nand2_1_4/B 2.33fF
C810 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C811 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.04fF
C812 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.04fF
C813 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.08fF
C814 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C815 sky130_fd_sc_hd__nand2_4_0/Y Bd 0.00fF
C816 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C817 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C818 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C819 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X -0.00fF
C820 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.02fF
C821 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.02fF
C822 sky130_fd_sc_hd__clkinv_4_10/w_82_21# sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C823 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.00fF
C824 sky130_fd_sc_hd__clkinv_4_9/w_82_21# sky130_fd_sc_hd__nand2_4_3/Y 0.03fF
C825 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A -0.00fF
C826 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C827 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C828 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.04fF
C829 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C830 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C831 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.03fF
C832 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# VDD 0.22fF
C833 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C834 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C835 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.07fF
C836 VDD sky130_fd_sc_hd__clkinv_4_4/Y -0.31fF
C837 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C838 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C839 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.00fF
C840 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C841 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C842 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__nand2_4_2/Y 0.04fF
C843 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A -0.00fF
C844 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.00fF
C845 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C846 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C847 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C848 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C849 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_3/A 0.13fF
C850 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.31fF
C851 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C852 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C853 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# VDD 0.15fF
C854 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.01fF
C855 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C856 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.01fF
C857 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C858 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.02fF
C859 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C860 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.05fF
C861 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.04fF
C862 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.04fF
C863 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# 0.09fF
C864 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C865 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C866 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.07fF
C867 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C868 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.03fF
C869 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C870 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 2.38fF
C871 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.10fF
C872 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.09fF
C873 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C874 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.05fF
C875 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.67fF
C876 p2 Bd_b 0.56fF
C877 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C878 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 2.38fF
C879 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.05fF
C880 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# -0.01fF
C881 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C882 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.10fF
C883 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VDD 0.06fF
C884 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C885 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.08fF
C886 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.00fF
C887 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.00fF
C888 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.01fF
C889 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.02fF
C890 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_1_2/B 0.03fF
C891 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.11fF
C892 sky130_fd_sc_hd__nand2_4_2/a_27_47# VDD 0.04fF
C893 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.08fF
C894 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C895 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C896 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C897 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C898 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C899 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.08fF
C900 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0.05fF
C901 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.04fF
C902 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.04fF
C903 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.02fF
C904 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.19fF
C905 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.79fF
C906 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C907 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C908 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C909 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C910 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C911 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C912 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C913 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 2.27fF
C914 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C915 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# VDD 0.15fF
C916 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.16fF
C917 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_3/A 0.16fF
C918 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C919 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.12fF
C920 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.13fF
C921 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C922 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C923 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C924 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C925 sky130_fd_sc_hd__clkinv_4_3/Y VDD 1.02fF
C926 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_1_4/B 0.25fF
C927 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C928 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.02fF
C929 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C930 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.03fF
C931 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.45fF
C932 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C933 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C934 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.10fF
C935 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C936 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Ad_b 0.05fF
C937 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.04fF
C938 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.04fF
C939 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C940 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.25fF
C941 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 1.21fF
C942 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C943 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C944 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.01fF
C945 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C946 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.03fF
C947 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C948 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C949 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C950 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C951 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C952 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.34fF
C953 sky130_fd_sc_hd__mux2_1_0/a_439_47# Bd_b 0.00fF
C954 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.05fF
C955 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C956 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C957 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C958 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.11fF
C959 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.02fF
C960 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.04fF
C961 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.04fF
C962 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.02fF
C963 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C964 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C965 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C966 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C967 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C968 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C969 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C970 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C971 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 1.12fF
C972 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Ad_b 0.05fF
C973 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C974 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C975 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C976 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# VDD 0.22fF
C977 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkinv_4_1/A 0.05fF
C978 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.02fF
C979 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.02fF
C980 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C981 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C982 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.03fF
C983 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C984 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.00fF
C985 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.02fF
C986 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C987 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C988 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C989 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkinv_4_10/Y 0.08fF
C990 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C991 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.08fF
C992 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.34fF
C993 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.02fF
C994 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C995 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C996 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C997 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/A 0.45fF
C998 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C999 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# 0.07fF
C1000 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.14fF
C1001 p2 sky130_fd_sc_hd__clkinv_4_5/Y 0.16fF
C1002 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C1003 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C1004 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C1005 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VDD 0.41fF
C1006 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0.04fF
C1007 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.04fF
C1008 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.10fF
C1009 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.15fF
C1010 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.04fF
C1011 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.04fF
C1012 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD 1.95fF
C1013 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C1014 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.03fF
C1015 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# 0.00fF
C1016 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.15fF
C1017 p1 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.06fF
C1018 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1d 0.06fF
C1019 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C1020 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.05fF
C1021 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.04fF
C1022 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.30fF
C1023 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# Bd_b 0.01fF
C1024 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# Ad_b 0.01fF
C1025 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C1026 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.02fF
C1027 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C1028 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C1029 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C1030 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.05fF
C1031 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.03fF
C1032 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.05fF
C1033 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.05fF
C1034 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C1035 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C1036 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.03fF
C1037 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.05fF
C1038 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.05fF
C1039 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.10fF
C1040 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# VDD 0.16fF
C1041 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.01fF
C1042 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C1043 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C1044 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C1045 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# VDD 0.18fF
C1046 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkinv_4_1/A 0.06fF
C1047 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.05fF
C1048 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C1049 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# -0.05fF
C1050 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# VDD 0.29fF
C1051 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.08fF
C1052 Ad Ad_b 0.60fF
C1053 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.07fF
C1054 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_1_0/B 0.00fF
C1055 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.02fF
C1056 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C1057 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C1058 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C1059 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.08fF
C1060 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 1.58fF
C1061 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C1062 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C1063 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C1064 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C1065 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C1066 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C1067 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.19fF
C1068 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C1069 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.05fF
C1070 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C1071 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C1072 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C1073 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C1074 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C1075 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.00fF
C1076 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.00fF
C1077 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# -0.05fF
C1078 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C1079 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C1080 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.41fF
C1081 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.02fF
C1082 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C1083 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C1084 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.31fF
C1085 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.01fF
C1086 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C1087 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C1088 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VDD 5.36fF
C1089 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C1090 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.04fF
C1091 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.18fF
C1092 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C1093 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C1094 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C1095 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.31fF
C1096 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C1097 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C1098 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C1099 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C1100 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.14fF
C1101 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.04fF
C1102 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.04fF
C1103 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C1104 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C1105 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.16fF
C1106 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C1107 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C1108 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C1109 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C1110 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.00fF
C1111 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 2.22fF
C1112 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C1113 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.03fF
C1114 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.18fF
C1115 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C1116 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C1117 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C1118 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C1119 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1120 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C1121 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.03fF
C1122 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C1123 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VDD 1.38fF
C1124 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkinv_4_1/A 0.11fF
C1125 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C1126 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C1127 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C1128 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A -0.00fF
C1129 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.11fF
C1130 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.04fF
C1131 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.02fF
C1132 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.04fF
C1133 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C1134 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C1135 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C1136 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.02fF
C1137 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.02fF
C1138 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C1139 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.00fF
C1140 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.01fF
C1141 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C1142 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C1143 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# VDD 0.16fF
C1144 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C1145 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C1146 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C1147 sky130_fd_sc_hd__nand2_1_4/B Ad_b 0.02fF
C1148 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.08fF
C1149 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.05fF
C1150 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VDD 1.46fF
C1151 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.03fF
C1152 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.02fF
C1153 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C1154 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.01fF
C1155 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.41fF
C1156 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.01fF
C1157 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C1158 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.02fF
C1159 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C1160 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C1161 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.08fF
C1162 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C1163 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C1164 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C1165 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C1166 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C1167 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1168 sky130_fd_sc_hd__nand2_4_3/Y Bd_b 0.00fF
C1169 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C1170 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C1171 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C1172 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VDD 0.16fF
C1173 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C1174 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.00fF
C1175 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VDD 0.18fF
C1176 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C1177 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Ad 0.12fF
C1178 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# VDD 0.29fF
C1179 sky130_fd_sc_hd__clkinv_4_7/A p1 0.00fF
C1180 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.07fF
C1181 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_1_1/Y 0.12fF
C1182 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.04fF
C1183 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C1184 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C1185 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C1186 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C1187 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C1188 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkinv_4_2/Y 0.03fF
C1189 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C1190 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.08fF
C1191 sky130_fd_sc_hd__nand2_1_3/A clk 0.02fF
C1192 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C1193 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C1194 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C1195 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__mux2_1_0/S 0.02fF
C1196 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.02fF
C1197 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C1198 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C1199 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# VDD 0.16fF
C1200 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.01fF
C1201 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.01fF
C1202 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.01fF
C1203 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C1204 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# VDD 0.18fF
C1205 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.02fF
C1206 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C1207 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C1208 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C1209 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C1210 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VDD 0.47fF
C1211 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_3/A 2.16fF
C1212 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C1213 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C1214 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VDD 0.06fF
C1215 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A -0.00fF
C1216 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.04fF
C1217 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.04fF
C1218 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1219 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C1220 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C1221 sky130_fd_sc_hd__nand2_1_2/B clk 0.04fF
C1222 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.08fF
C1223 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C1224 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C1225 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C1226 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C1227 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_4/Y 0.23fF
C1228 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C1229 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 1.38fF
C1230 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C1231 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C1232 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VDD 0.24fF
C1233 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.03fF
C1234 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C1235 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_12/a_110_47# 0.04fF
C1236 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.08fF
C1237 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.02fF
C1238 VDD sky130_fd_sc_hd__nand2_4_2/B 0.40fF
C1239 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.02fF
C1240 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C1241 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C1242 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C1243 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C1244 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.07fF
C1245 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C1246 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C1247 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C1248 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C1249 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C1250 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# VDD 0.11fF
C1251 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.02fF
C1252 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.02fF
C1253 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C1254 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# VDD 0.13fF
C1255 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C1256 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C1257 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.14fF
C1258 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C1259 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.05fF
C1260 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C1261 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# VDD 0.30fF
C1262 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.02fF
C1263 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VDD 0.37fF
C1264 sky130_fd_sc_hd__clkinv_4_3/Y Ad_b 0.07fF
C1265 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C1266 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_1_2/A 0.01fF
C1267 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C1268 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X -0.00fF
C1269 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.16fF
C1270 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.07fF
C1271 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C1272 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.31fF
C1273 Bd Bd_b 0.47fF
C1274 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C1275 B Bd_b 0.08fF
C1276 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.04fF
C1277 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C1278 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.16fF
C1279 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.02fF
C1280 VDD sky130_fd_sc_hd__clkinv_1_1/Y -1.16fF
C1281 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.04fF
C1282 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C1283 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.06fF
C1284 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# VDD 0.31fF
C1285 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VDD 0.40fF
C1286 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C1287 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C1288 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C1289 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C1290 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.17fF
C1291 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.03fF
C1292 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.10fF
C1293 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.04fF
C1294 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.02fF
C1295 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C1296 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 1.12fF
C1297 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C1298 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1299 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C1300 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C1301 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.03fF
C1302 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C1303 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.09fF
C1304 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 1.14fF
C1305 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C1306 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.03fF
C1307 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C1308 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.19fF
C1309 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C1310 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C1311 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.09fF
C1312 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C1313 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.07fF
C1314 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C1315 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.07fF
C1316 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C1317 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.02fF
C1318 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C1319 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C1320 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A -0.00fF
C1321 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C1322 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_3/A 0.04fF
C1323 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.95fF
C1324 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.05fF
C1325 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C1326 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C1327 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Ad_b 0.04fF
C1328 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__nand2_4_2/A 0.42fF
C1329 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C1330 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.31fF
C1331 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.09fF
C1332 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.08fF
C1333 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.31fF
C1334 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C1335 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C1336 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C1337 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.08fF
C1338 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.19fF
C1339 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.34fF
C1340 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C1341 sky130_fd_sc_hd__nand2_4_0/a_27_47# VDD 0.04fF
C1342 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.02fF
C1343 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.03fF
C1344 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C1345 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C1346 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.01fF
C1347 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A -0.00fF
C1348 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.07fF
C1349 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# VDD 0.10fF
C1350 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.08fF
C1351 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C1352 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C1353 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__nand2_1_0/A 0.10fF
C1354 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C1355 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C1356 sky130_fd_sc_hd__clkinv_4_9/Y VDD 0.74fF
C1357 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C1358 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.08fF
C1359 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# VDD 0.31fF
C1360 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C1361 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C1362 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C1363 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.02fF
C1364 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C1365 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.11fF
C1366 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# 0.35fF
C1367 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.30fF
C1368 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A -0.00fF
C1369 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C1370 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C1371 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X -0.00fF
C1372 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VDD 0.15fF
C1373 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C1374 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# VDD 0.32fF
C1375 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C1376 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C1377 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.01fF
C1378 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.07fF
C1379 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C1380 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C1381 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1382 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C1383 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.03fF
C1384 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD 1.51fF
C1385 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C1386 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.04fF
C1387 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 2.27fF
C1388 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C1389 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C1390 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C1391 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C1392 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C1393 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C1394 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C1395 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C1396 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C1397 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C1398 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.19fF
C1399 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_3/w_82_21# 0.03fF
C1400 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.11fF
C1401 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C1402 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C1403 p2 A 0.02fF
C1404 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C1405 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C1406 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C1407 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C1408 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1409 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C1410 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_0/B 0.12fF
C1411 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.01fF
C1412 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.00fF
C1413 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C1414 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkinv_4_1/A 0.01fF
C1415 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C1416 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.12fF
C1417 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.05fF
C1418 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.02fF
C1419 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.12fF
C1420 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# VDD 0.34fF
C1421 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.08fF
C1422 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C1423 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C1424 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C1425 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1426 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C1427 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.44fF
C1428 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C1429 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.00fF
C1430 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C1431 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C1432 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C1433 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C1434 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VDD 0.35fF
C1435 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.11fF
C1436 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C1437 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C1438 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Ad_b 0.09fF
C1439 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.09fF
C1440 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C1441 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C1442 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C1443 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C1444 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C1445 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.03fF
C1446 p2_b p2d 0.53fF
C1447 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.06fF
C1448 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.04fF
C1449 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.04fF
C1450 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# p2 0.00fF
C1451 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C1452 p2_b VDD 0.90fF
C1453 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.05fF
C1454 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C1455 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C1456 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C1457 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.16fF
C1458 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.19fF
C1459 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C1460 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C1461 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C1462 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.11fF
C1463 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.07fF
C1464 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_1/A 0.37fF
C1465 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VDD 0.19fF
C1466 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__nand2_1_0/A 0.02fF
C1467 p1_b sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.15fF
C1468 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# p1d 0.15fF
C1469 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_1_4/B 0.11fF
C1470 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.26fF
C1471 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Bd_b 0.05fF
C1472 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C1473 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C1474 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C1475 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C1476 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C1477 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C1478 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.13fF
C1479 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C1480 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.19fF
C1481 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A -0.00fF
C1482 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C1483 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C1484 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.17fF
C1485 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C1486 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.35fF
C1487 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C1488 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C1489 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.03fF
C1490 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.22fF
C1491 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.04fF
C1492 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.04fF
C1493 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.63fF
C1494 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.09fF
C1495 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.02fF
C1496 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C1497 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.01fF
C1498 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.11fF
C1499 VDD sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.08fF
C1500 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A -0.00fF
C1501 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C1502 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.05fF
C1503 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C1504 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C1505 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.01fF
C1506 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.03fF
C1507 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Bd_b 0.05fF
C1508 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# VDD 0.10fF
C1509 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C1510 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.03fF
C1511 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.09fF
C1512 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C1513 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# VDD 0.19fF
C1514 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C1515 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C1516 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.03fF
C1517 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__nand2_1_4/B 0.12fF
C1518 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_4/Y 0.04fF
C1519 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C1520 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C1521 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C1522 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD 1.08fF
C1523 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1524 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.30fF
C1525 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C1526 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.03fF
C1527 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C1528 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C1529 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.00fF
C1530 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.00fF
C1531 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.23fF
C1532 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.03fF
C1533 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C1534 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C1535 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.04fF
C1536 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.04fF
C1537 p2 sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C1538 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C1539 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C1540 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# VDD 0.20fF
C1541 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C1542 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.05fF
C1543 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.05fF
C1544 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VDD 1.52fF
C1545 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C1546 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C1547 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C1548 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C1549 sky130_fd_sc_hd__nand2_4_2/Y p1d 0.00fF
C1550 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VDD 0.33fF
C1551 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.01fF
C1552 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.15fF
C1553 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.17fF
C1554 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# Bd_b 0.01fF
C1555 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.00fF
C1556 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.00fF
C1557 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.07fF
C1558 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C1559 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C1560 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C1561 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_1_3/Y 0.04fF
C1562 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C1563 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C1564 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# VDD 0.34fF
C1565 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.00fF
C1566 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C1567 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.02fF
C1568 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C1569 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.04fF
C1570 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C1571 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C1572 sky130_fd_sc_hd__clkinv_4_1/A B 0.00fF
C1573 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X -0.00fF
C1574 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C1575 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C1576 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C1577 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C1578 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.05fF
C1579 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C1580 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C1581 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# VDD 0.16fF
C1582 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C1583 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.01fF
C1584 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C1585 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# VDD 0.11fF
C1586 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C1587 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C1588 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.05fF
C1589 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C1590 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.01fF
C1591 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# -0.05fF
C1592 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C1593 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C1594 p1d_b p1 0.08fF
C1595 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C1596 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.03fF
C1597 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C1598 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 1.08fF
C1599 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__mux2_1_0/S 0.05fF
C1600 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C1601 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C1602 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.10fF
C1603 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C1604 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C1605 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C1606 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.07fF
C1607 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.04fF
C1608 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.04fF
C1609 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.04fF
C1610 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C1611 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1612 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C1613 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# -0.04fF
C1614 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# Ad_b 0.02fF
C1615 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C1616 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C1617 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.00fF
C1618 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C1619 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.05fF
C1620 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.05fF
C1621 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C1622 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C1623 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C1624 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C1625 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C1626 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C1627 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.03fF
C1628 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C1629 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.33fF
C1630 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.13fF
C1631 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.02fF
C1632 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C1633 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C1634 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C1635 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C1636 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C1637 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.02fF
C1638 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.27fF
C1639 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.07fF
C1640 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/a_27_47# 0.00fF
C1641 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.04fF
C1642 sky130_fd_sc_hd__clkinv_4_7/A VDD 3.56fF
C1643 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.02fF
C1644 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C1645 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C1646 Bd B_b 0.53fF
C1647 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.08fF
C1648 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C1649 B B_b 0.47fF
C1650 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C1651 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C1652 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C1653 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.03fF
C1654 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C1655 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C1656 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C1657 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C1658 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.04fF
C1659 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.04fF
C1660 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C1661 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.03fF
C1662 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VDD 0.35fF
C1663 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C1664 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C1665 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C1666 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C1667 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.00fF
C1668 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C1669 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.02fF
C1670 VDD sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.27fF
C1671 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C1672 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C1673 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 2.24fF
C1674 sky130_fd_sc_hd__nand2_1_4/B Bd_b 0.02fF
C1675 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.06fF
C1676 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.04fF
C1677 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.04fF
C1678 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/D -0.28fF
C1679 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.05fF
C1680 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C1681 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C1682 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C1683 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C1684 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C1685 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.05fF
C1686 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C1687 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C1688 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.04fF
C1689 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C1690 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1691 sky130_fd_sc_hd__clkinv_4_9/Y Ad_b 0.03fF
C1692 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C1693 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C1694 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C1695 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C1696 sky130_fd_sc_hd__clkinv_4_4/Y Bd_b 0.08fF
C1697 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C1698 sky130_fd_sc_hd__nand2_4_3/a_27_47# VDD 0.05fF
C1699 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C1700 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.03fF
C1701 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VDD 0.15fF
C1702 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C1703 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# VDD 0.16fF
C1704 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.07fF
C1705 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# VDD 0.23fF
C1706 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 1.83fF
C1707 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.12fF
C1708 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.08fF
C1709 sky130_fd_sc_hd__dfxbp_1_1/a_592_47# sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C1710 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# sky130_fd_sc_hd__clkinv_4_1/Y 0.08fF
C1711 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C1712 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C1713 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B 0.69fF
C1714 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Ad_b 0.02fF
C1715 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C1716 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.01fF
C1717 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.02fF
C1718 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.02fF
C1719 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# VDD 0.16fF
C1720 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C1721 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# VDD 0.30fF
C1722 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C1723 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C1724 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.07fF
C1725 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.04fF
C1726 sky130_fd_sc_hd__dfxbp_1_0/a_561_413# VDD 0.00fF
C1727 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.02fF
C1728 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/A 0.62fF
C1729 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C1730 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C1731 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C1732 sky130_fd_sc_hd__nand2_1_2/A clk 0.07fF
C1733 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C1734 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C1735 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C1736 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# -0.17fF
C1737 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.04fF
C1738 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C1739 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C1740 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C1741 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C1742 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C1743 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C1744 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C1745 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C1746 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# VDD -0.10fF
C1747 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C1748 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C1749 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.11fF
C1750 p2d_b p2d 0.52fF
C1751 p2d_b VDD 0.91fF
C1752 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.08fF
C1753 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.05fF
C1754 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C1755 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C1756 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C1757 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C1758 Ad sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.15fF
C1759 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# A_b 0.15fF
C1760 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C1761 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C1762 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C1763 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# VDD 0.12fF
C1764 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C1765 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C1766 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# VDD 0.15fF
C1767 sky130_fd_sc_hd__clkinv_4_3/Y Bd_b 0.18fF
C1768 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C1769 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C1770 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1771 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C1772 VDD sky130_fd_sc_hd__nand2_4_1/A 12.32fF
C1773 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.10fF
C1774 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.01fF
C1775 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C1776 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_4/B 0.14fF
C1777 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C1778 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C1779 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C1780 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C1781 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C1782 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.08fF
C1783 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# VDD 0.18fF
C1784 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.07fF
C1785 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.26fF
C1786 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C1787 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C1788 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C1789 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C1790 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C1791 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.04fF
C1792 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C1793 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C1794 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C1795 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.31fF
C1796 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1797 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# VDD 0.30fF
C1798 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C1799 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C1800 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# -0.00fF
C1801 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkinv_4_4/Y 0.02fF
C1802 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.08fF
C1803 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C1804 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.06fF
C1805 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkinv_4_8/Y 0.03fF
C1806 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD 1.59fF
C1807 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Ad_b 0.07fF
C1808 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C1809 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C1810 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C1811 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C1812 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C1813 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1814 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C1815 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C1816 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 1.47fF
C1817 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.08fF
C1818 sky130_fd_sc_hd__clkinv_1_3/A VDD 4.21fF
C1819 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Bd_b 0.05fF
C1820 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.04fF
C1821 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.04fF
C1822 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.07fF
C1823 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.08fF
C1824 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.14fF
C1825 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.03fF
C1826 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C1827 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.02fF
C1828 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.17fF
C1829 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.01fF
C1830 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C1831 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.05fF
C1832 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.01fF
C1833 sky130_fd_sc_hd__clkinv_4_9/w_82_21# sky130_fd_sc_hd__clkinv_4_9/Y 0.05fF
C1834 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.19fF
C1835 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.07fF
C1836 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C1837 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.03fF
C1838 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# VDD 0.11fF
C1839 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.06fF
C1840 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.02fF
C1841 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.15fF
C1842 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C1843 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C1844 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.00fF
C1845 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C1846 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C1847 VDD A_b 0.94fF
C1848 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VDD 0.34fF
C1849 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# VDD 0.15fF
C1850 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C1851 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C1852 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C1853 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C1854 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_1_2/Y 0.36fF
C1855 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# 0.10fF
C1856 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.17fF
C1857 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# VDD 0.26fF
C1858 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__nand2_4_2/A 0.59fF
C1859 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.36fF
C1860 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C1861 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_3/A 0.32fF
C1862 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C1863 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# VDD 0.19fF
C1864 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C1865 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.04fF
C1866 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.64fF
C1867 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.05fF
C1868 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.05fF
C1869 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C1870 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# VDD 0.31fF
C1871 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C1872 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C1873 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VDD 0.35fF
C1874 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/B 0.11fF
C1875 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A -0.00fF
C1876 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C1877 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C1878 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.05fF
C1879 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# 0.05fF
C1880 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C1881 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C1882 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C1883 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkinv_4_3/Y 0.04fF
C1884 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.07fF
C1885 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.07fF
C1886 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C1887 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.03fF
C1888 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X -0.00fF
C1889 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C1890 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C1891 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.11fF
C1892 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C1893 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C1894 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C1895 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C1896 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.03fF
C1897 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.11fF
C1898 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C1899 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.00fF
C1900 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C1901 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.04fF
C1902 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.01fF
C1903 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C1904 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C1905 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C1906 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C1907 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C1908 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.04fF
C1909 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.04fF
C1910 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C1911 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.04fF
C1912 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C1913 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C1914 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.10fF
C1915 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C1916 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# VDD 0.19fF
C1917 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C1918 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.02fF
C1919 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C1920 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C1921 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.01fF
C1922 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C1923 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C1924 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VDD 0.19fF
C1925 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A -0.00fF
C1926 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C1927 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C1928 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C1929 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C1930 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.10fF
C1931 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# VDD 0.23fF
C1932 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C1933 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Bd_b 0.07fF
C1934 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.08fF
C1935 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.19fF
C1936 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C1937 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C1938 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C1939 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C1940 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.03fF
C1941 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.19fF
C1942 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.00fF
C1943 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.05fF
C1944 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C1945 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C1946 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C1947 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C1948 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C1949 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# p2 0.00fF
C1950 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A 1.17fF
C1951 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.41fF
C1952 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C1953 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.08fF
C1954 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.06fF
C1955 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C1956 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C1957 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C1958 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.01fF
C1959 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C1960 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.07fF
C1961 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__nand2_4_1/B 0.07fF
C1962 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.08fF
C1963 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C1964 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C1965 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD 1.66fF
C1966 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.05fF
C1967 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C1968 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.08fF
C1969 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.07fF
C1970 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C1971 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C1972 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C1973 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C1974 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C1975 p2_b sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.15fF
C1976 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C1977 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C1978 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.81fF
C1979 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C1980 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C1981 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C1982 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C1983 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.15fF
C1984 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C1985 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.31fF
C1986 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# Ad_b 0.12fF
C1987 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C1988 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C1989 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.03fF
C1990 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.10fF
C1991 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C1992 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C1993 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C1994 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.01fF
C1995 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C1996 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.02fF
C1997 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C1998 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.03fF
C1999 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C2000 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.30fF
C2001 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C2002 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.02fF
C2003 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C2004 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.04fF
C2005 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.04fF
C2006 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C2007 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.03fF
C2008 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C2009 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# VDD 0.11fF
C2010 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C2011 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C2012 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C2013 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C2014 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C2015 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C2016 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C2017 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C2018 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.03fF
C2019 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.04fF
C2020 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.04fF
C2021 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# VDD 0.06fF
C2022 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C2023 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.04fF
C2024 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.04fF
C2025 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.18fF
C2026 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C2027 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 1.35fF
C2028 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# VDD 0.33fF
C2029 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C2030 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__nand2_1_4/B -0.30fF
C2031 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C2032 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C2033 p1d_b p1_b 0.19fF
C2034 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C2035 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C2036 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# -0.00fF
C2037 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C2038 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkinv_4_1/A 0.08fF
C2039 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# p2_b 0.09fF
C2040 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.14fF
C2041 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.04fF
C2042 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C2043 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.04fF
C2044 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.04fF
C2045 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C2046 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.12fF
C2047 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/A 0.48fF
C2048 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_8/Y 0.04fF
C2049 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.00fF
C2050 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C2051 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C2052 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C2053 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C2054 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C2055 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C2056 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.04fF
C2057 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.15fF
C2058 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C2059 sky130_fd_sc_hd__dfxbp_1_1/D clk 0.04fF
C2060 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C2061 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C2062 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C2063 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.01fF
C2064 p1d_b VDD 0.92fF
C2065 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C2066 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C2067 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C2068 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.04fF
C2069 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C2070 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C2071 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C2072 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C2073 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C2074 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.15fF
C2075 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.04fF
C2076 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.04fF
C2077 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C2078 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C2079 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C2080 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.02fF
C2081 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.02fF
C2082 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C2083 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2084 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C2085 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.02fF
C2086 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# VDD 0.15fF
C2087 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/B 0.02fF
C2088 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.02fF
C2089 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.02fF
C2090 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C2091 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# VDD 0.31fF
C2092 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C2093 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C2094 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.03fF
C2095 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C2096 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C2097 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C2098 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.03fF
C2099 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C2100 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C2101 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C2102 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.15fF
C2103 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.08fF
C2104 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# 0.04fF
C2105 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# VDD 0.14fF
C2106 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C2107 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C2108 Ad A 0.19fF
C2109 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C2110 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.09fF
C2111 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C2112 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C2113 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C2114 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.14fF
C2115 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C2116 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C2117 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C2118 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.09fF
C2119 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X -0.00fF
C2120 sky130_fd_sc_hd__nand2_4_1/A Ad_b 0.48fF
C2121 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C2122 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2123 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2124 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.01fF
C2125 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.09fF
C2126 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.04fF
C2127 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C2128 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C2129 VDD clk 2.29fF
C2130 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_2/A 0.26fF
C2131 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C2132 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C2133 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.01fF
C2134 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C2135 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.01fF
C2136 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.04fF
C2137 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 1.83fF
C2138 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C2139 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# Bd_b 0.46fF
C2140 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C2141 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C2142 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C2143 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C2144 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C2145 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C2146 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C2147 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C2148 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.08fF
C2149 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C2150 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C2151 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.00fF
C2152 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VDD 0.32fF
C2153 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.06fF
C2154 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.07fF
C2155 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.07fF
C2156 sky130_fd_sc_hd__clkinv_4_2/w_82_21# sky130_fd_sc_hd__nand2_4_0/Y 0.03fF
C2157 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.13fF
C2158 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C2159 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.03fF
C2160 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C2161 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.01fF
C2162 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C2163 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C2164 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.00fF
C2165 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# -0.01fF
C2166 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.15fF
C2167 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C2168 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.30fF
C2169 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C2170 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C2171 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C2172 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Ad_b 0.02fF
C2173 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.05fF
C2174 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.11fF
C2175 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C2176 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C2177 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VDD 0.00fF
C2178 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.04fF
C2179 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 1.10fF
C2180 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.08fF
C2181 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C2182 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C2183 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C2184 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C2185 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C2186 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C2187 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C2188 sky130_fd_sc_hd__clkinv_1_3/A Ad_b 0.25fF
C2189 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C2190 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.02fF
C2191 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C2192 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.01fF
C2193 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.05fF
C2194 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C2195 VDD sky130_fd_sc_hd__mux2_1_0/X 0.62fF
C2196 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C2197 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C2198 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C2199 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C2200 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C2201 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C2202 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C2203 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_4/Y 0.04fF
C2204 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.04fF
C2205 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C2206 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C2207 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.01fF
C2208 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.01fF
C2209 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.01fF
C2210 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C2211 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD 1.17fF
C2212 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__nand2_1_1/A 0.08fF
C2213 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/D 0.02fF
C2214 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.01fF
C2215 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C2216 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.04fF
C2217 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.04fF
C2218 sky130_fd_sc_hd__clkinv_4_4/w_82_21# sky130_fd_sc_hd__clkinv_4_5/Y 0.03fF
C2219 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C2220 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.06fF
C2221 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C2222 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.10fF
C2223 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C2224 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C2225 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C2226 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.06fF
C2227 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD -0.61fF
C2228 sky130_fd_sc_hd__clkinv_4_9/Y Bd_b 0.00fF
C2229 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C2230 A_b Ad_b 0.33fF
C2231 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C2232 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.09fF
C2233 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.15fF
C2234 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C2235 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# VDD 0.13fF
C2236 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C2237 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.05fF
C2238 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.08fF
C2239 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C2240 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.04fF
C2241 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.02fF
C2242 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# VDD 0.12fF
C2243 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C2244 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C2245 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C2246 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.16fF
C2247 sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C2248 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.05fF
C2249 sky130_fd_sc_hd__nand2_4_3/A clk 0.03fF
C2250 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C2251 sky130_fd_sc_hd__clkinv_4_5/w_82_21# sky130_fd_sc_hd__clkinv_4_5/Y -0.00fF
C2252 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Bd_b 0.02fF
C2253 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# VDD 0.34fF
C2254 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.04fF
C2255 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.04fF
C2256 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.04fF
C2257 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C2258 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C2259 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C2260 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_1/A 0.66fF
C2261 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C2262 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C2263 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C2264 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# VDD 0.17fF
C2265 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkinv_1_1/Y 0.37fF
C2266 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.18fF
C2267 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# VDD 0.33fF
C2268 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C2269 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.08fF
C2270 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.97fF
C2271 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C2272 sky130_fd_sc_hd__dfxbp_1_0/a_975_413# VDD 0.00fF
C2273 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VDD 0.10fF
C2274 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C2275 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C2276 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C2277 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C2278 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.00fF
C2279 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.10fF
C2280 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C2281 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p2d_b 0.02fF
C2282 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C2283 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C2284 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.03fF
C2285 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.02fF
C2286 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C2287 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# VDD 0.09fF
C2288 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C2289 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C2290 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C2291 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.05fF
C2292 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C2293 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C2294 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C2295 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C2296 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.03fF
C2297 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VDD 1.12fF
C2298 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.01fF
C2299 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C2300 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.01fF
C2301 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C2302 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.19fF
C2303 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C2304 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__mux2_1_0/X 0.07fF
C2305 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C2306 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C2307 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.01fF
C2308 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C2309 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C2310 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C2311 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# VDD 0.31fF
C2312 p2d_b sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.14fF
C2313 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C2314 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C2315 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A 1.05fF
C2316 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.10fF
C2317 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_4/B 0.92fF
C2318 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X -0.00fF
C2319 sky130_fd_sc_hd__clkinv_4_7/Y p1_b 0.03fF
C2320 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.03fF
C2321 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C2322 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.09fF
C2323 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# VDD 0.31fF
C2324 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C2325 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.05fF
C2326 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C2327 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# A_b 0.06fF
C2328 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_2/B 0.07fF
C2329 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.03fF
C2330 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C2331 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.62fF
C2332 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.19fF
C2333 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.98fF
C2334 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.09fF
C2335 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.05fF
C2336 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.04fF
C2337 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.04fF
C2338 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# VDD 0.17fF
C2339 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C2340 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C2341 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C2342 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C2343 VDD sky130_fd_sc_hd__clkinv_4_7/Y -0.33fF
C2344 p2d_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.07fF
C2345 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.08fF
C2346 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.05fF
C2347 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.08fF
C2348 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C2349 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C2350 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C2351 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C2352 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C2353 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.03fF
C2354 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C2355 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.31fF
C2356 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.02fF
C2357 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C2358 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.00fF
C2359 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Bd_b 0.07fF
C2360 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VDD 1.15fF
C2361 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C2362 VDD sky130_fd_sc_hd__nand2_1_0/A 1.26fF
C2363 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C2364 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C2365 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.11fF
C2366 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 1.12fF
C2367 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C2368 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.06fF
C2369 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C2370 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2371 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VDD 0.11fF
C2372 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.19fF
C2373 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# Bd_b 0.06fF
C2374 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.07fF
C2375 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C2376 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C2377 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.01fF
C2378 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.00fF
C2379 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.02fF
C2380 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.01fF
C2381 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C2382 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.08fF
C2383 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.15fF
C2384 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD 1.55fF
C2385 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C2386 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C2387 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C2388 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C2389 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C2390 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C2391 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C2392 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkinv_4_1/A 0.01fF
C2393 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C2394 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C2395 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C2396 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VDD 0.17fF
C2397 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.08fF
C2398 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C2399 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C2400 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C2401 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C2402 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C2403 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# VDD 0.15fF
C2404 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.12fF
C2405 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.25fF
C2406 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.31fF
C2407 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C2408 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C2409 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# VDD 0.13fF
C2410 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.17fF
C2411 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C2412 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C2413 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C2414 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C2415 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# VDD 0.15fF
C2416 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# VDD 0.36fF
C2417 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C2418 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.03fF
C2419 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_1_0/B 0.06fF
C2420 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C2421 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.26fF
C2422 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.10fF
C2423 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C2424 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# VDD 0.18fF
C2425 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.01fF
C2426 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.02fF
C2427 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.01fF
C2428 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C2429 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C2430 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.05fF
C2431 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C2432 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C2433 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.04fF
C2434 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.04fF
C2435 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# VDD 0.31fF
C2436 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C2437 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C2438 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C2439 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.04fF
C2440 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# -0.05fF
C2441 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.02fF
C2442 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C2443 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X -0.00fF
C2444 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.11fF
C2445 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C2446 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C2447 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.01fF
C2448 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.07fF
C2449 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__nand2_1_2/B 0.03fF
C2450 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C2451 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.02fF
C2452 sky130_fd_sc_hd__clkinv_1_0/Y VDD -1.31fF
C2453 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X -0.00fF
C2454 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C2455 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.05fF
C2456 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C2457 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.05fF
C2458 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C2459 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C2460 sky130_fd_sc_hd__clkinv_4_6/w_82_21# sky130_fd_sc_hd__clkinv_4_7/A -0.00fF
C2461 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C2462 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.08fF
C2463 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.19fF
C2464 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C2465 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C2466 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C2467 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C2468 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C2469 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C2470 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.07fF
C2471 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C2472 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# VDD 0.14fF
C2473 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C2474 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C2475 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C2476 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C2477 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C2478 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C2479 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C2480 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C2481 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C2482 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VDD 0.15fF
C2483 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# VDD 0.12fF
C2484 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C2485 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C2486 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C2487 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.10fF
C2488 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C2489 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# VDD 0.41fF
C2490 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C2491 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C2492 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C2493 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C2494 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.04fF
C2495 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.04fF
C2496 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C2497 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C2498 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# p2 -0.00fF
C2499 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C2500 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C2501 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C2502 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C2503 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 2.23fF
C2504 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C2505 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.07fF
C2506 VDD sky130_fd_sc_hd__nand2_1_3/A 4.50fF
C2507 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.05fF
C2508 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C2509 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.08fF
C2510 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C2511 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.00fF
C2512 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.08fF
C2513 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C2514 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.07fF
C2515 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C2516 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.01fF
C2517 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C2518 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.03fF
C2519 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C2520 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.11fF
C2521 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.14fF
C2522 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C2523 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C2524 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C2525 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C2526 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VDD 0.50fF
C2527 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C2528 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C2529 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C2530 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C2531 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C2532 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C2533 VDD sky130_fd_sc_hd__nand2_1_2/B 1.60fF
C2534 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.01fF
C2535 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C2536 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C2537 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C2538 B_b sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.06fF
C2539 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.03fF
C2540 sky130_fd_sc_hd__mux2_1_0/X Ad_b 0.00fF
C2541 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# Bd_b 0.10fF
C2542 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C2543 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.11fF
C2544 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C2545 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C2546 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.08fF
C2547 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C2548 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C2549 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C2550 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C2551 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.15fF
C2552 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.11fF
C2553 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C2554 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C2555 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C2556 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C2557 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C2558 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.00fF
C2559 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.30fF
C2560 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C2561 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/B 0.05fF
C2562 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C2563 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# -0.00fF
C2564 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.04fF
C2565 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C2566 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# VDD 0.11fF
C2567 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C2568 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.02fF
C2569 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.02fF
C2570 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C2571 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C2572 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.03fF
C2573 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# VDD 0.17fF
C2574 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C2575 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.03fF
C2576 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C2577 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.09fF
C2578 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_1_4/B 0.04fF
C2579 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C2580 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# VDD 0.30fF
C2581 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C2582 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C2583 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C2584 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C2585 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C2586 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.01fF
C2587 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C2588 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C2589 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C2590 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C2591 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C2592 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.11fF
C2593 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.08fF
C2594 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C2595 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C2596 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.07fF
C2597 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD 1.55fF
C2598 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C2599 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C2600 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1d_b 0.07fF
C2601 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.05fF
C2602 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C2603 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C2604 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C2605 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C2606 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.04fF
C2607 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.04fF
C2608 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C2609 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.01fF
C2610 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C2611 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C2612 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.00fF
C2613 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C2614 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C2615 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C2616 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/Y -0.11fF
C2617 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C2618 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.13fF
C2619 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_4_3/A 0.69fF
C2620 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# VDD 0.16fF
C2621 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C2622 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C2623 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C2624 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# VDD 0.18fF
C2625 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C2626 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C2627 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C2628 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C2629 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C2630 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkinv_1_2/Y 0.05fF
C2631 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 1.36fF
C2632 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# VDD 0.32fF
C2633 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.00fF
C2634 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C2635 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.06fF
C2636 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C2637 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C2638 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C2639 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C2640 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C2641 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C2642 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# 0.04fF
C2643 p2 sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C2644 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C2645 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C2646 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.00fF
C2647 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C2648 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.08fF
C2649 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X -0.00fF
C2650 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C2651 sky130_fd_sc_hd__nand2_4_1/A Bd_b 0.66fF
C2652 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.14fF
C2653 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2654 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C2655 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.01fF
C2656 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C2657 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C2658 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C2659 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C2660 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C2661 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.04fF
C2662 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C2663 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A -0.00fF
C2664 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C2665 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.02fF
C2666 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C2667 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C2668 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C2669 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 1.49fF
C2670 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C2671 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.36fF
C2672 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C2673 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.05fF
C2674 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C2675 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C2676 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.02fF
C2677 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.02fF
C2678 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.19fF
C2679 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.00fF
C2680 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C2681 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.04fF
C2682 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C2683 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VDD 0.17fF
C2684 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C2685 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C2686 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C2687 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C2688 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C2689 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.08fF
C2690 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.03fF
C2691 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C2692 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C2693 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C2694 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.08fF
C2695 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C2696 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.03fF
C2697 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.15fF
C2698 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.02fF
C2699 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.04fF
C2700 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.04fF
C2701 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C2702 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C2703 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C2704 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# p1d -0.01fF
C2705 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.09fF
C2706 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C2707 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.17fF
C2708 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C2709 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.05fF
C2710 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Bd_b 0.02fF
C2711 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.32fF
C2712 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C2713 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.05fF
C2714 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C2715 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C2716 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C2717 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C2718 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C2719 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C2720 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C2721 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C2722 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C2723 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C2724 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.31fF
C2725 sky130_fd_sc_hd__clkinv_1_3/A Bd_b 0.22fF
C2726 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C2727 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.03fF
C2728 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C2729 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C2730 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C2731 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Ad_b 0.04fF
C2732 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C2733 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__nand2_1_1/A 0.07fF
C2734 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C2735 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C2736 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.02fF
C2737 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.02fF
C2738 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C2739 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C2740 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.07fF
C2741 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C2742 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C2743 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.02fF
C2744 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/D 0.10fF
C2745 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__nand2_1_1/A 0.13fF
C2746 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.06fF
C2747 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C2748 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C2749 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C2750 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C2751 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C2752 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C2753 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C2754 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VDD 1.35fF
C2755 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C2756 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C2757 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C2758 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C2759 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C2760 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.04fF
C2761 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.04fF
C2762 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# -0.00fF
C2763 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C2764 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C2765 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C2766 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C2767 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C2768 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/w_82_21# 0.03fF
C2769 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# VDD 0.11fF
C2770 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C2771 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.06fF
C2772 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.01fF
C2773 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C2774 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.06fF
C2775 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# B_b 0.09fF
C2776 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_4_1/A 1.17fF
C2777 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.02fF
C2778 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# VDD 0.31fF
C2779 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C2780 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.02fF
C2781 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C2782 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.02fF
C2783 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C2784 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C2785 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C2786 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C2787 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C2788 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_1_1/Y 0.12fF
C2789 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# VDD 0.15fF
C2790 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C2791 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.15fF
C2792 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# VDD 0.29fF
C2793 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C2794 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.65fF
C2795 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C2796 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C2797 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C2798 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C2799 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C2800 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.10fF
C2801 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.00fF
C2802 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C2803 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C2804 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# VDD 0.19fF
C2805 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C2806 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C2807 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.08fF
C2808 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C2809 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X -0.00fF
C2810 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C2811 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.04fF
C2812 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C2813 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C2814 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.09fF
C2815 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.04fF
C2816 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.04fF
C2817 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.00fF
C2818 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.01fF
C2819 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C2820 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.08fF
C2821 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C2822 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C2823 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 2.39fF
C2824 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.04fF
C2825 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C2826 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.14fF
C2827 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C2828 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.03fF
C2829 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VDD 1.35fF
C2830 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C2831 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C2832 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.12fF
C2833 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# p2 -0.04fF
C2834 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C2835 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C2836 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.08fF
C2837 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.08fF
C2838 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X -0.00fF
C2839 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD 1.38fF
C2840 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.04fF
C2841 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C2842 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C2843 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/A 0.41fF
C2844 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/B 0.02fF
C2845 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.05fF
C2846 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C2847 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_1_1/Y 0.05fF
C2848 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0.09fF
C2849 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C2850 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2851 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_2/A 0.00fF
C2852 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C2853 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 1.10fF
C2854 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# 0.15fF
C2855 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C2856 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C2857 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C2858 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C2859 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# VDD 0.15fF
C2860 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.03fF
C2861 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.08fF
C2862 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C2863 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.19fF
C2864 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C2865 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C2866 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.08fF
C2867 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.03fF
C2868 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.02fF
C2869 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C2870 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C2871 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# VDD 0.34fF
C2872 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C2873 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C2874 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# VDD 0.37fF
C2875 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2876 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C2877 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C2878 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C2879 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.99fF
C2880 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.04fF
C2881 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C2882 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C2883 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.05fF
C2884 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2885 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C2886 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2887 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A -0.00fF
C2888 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.05fF
C2889 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C2890 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C2891 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.08fF
C2892 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VDD 1.17fF
C2893 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C2894 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.04fF
C2895 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.03fF
C2896 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.01fF
C2897 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C2898 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C2899 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C2900 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C2901 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C2902 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.02fF
C2903 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C2904 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.15fF
C2905 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.05fF
C2906 p1 p1_b 0.47fF
C2907 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# A_b 0.06fF
C2908 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.02fF
C2909 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C2910 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C2911 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C2912 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C2913 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VDD 0.15fF
C2914 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C2915 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C2916 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# VDD 0.12fF
C2917 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.32fF
C2918 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C2919 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C2920 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C2921 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_3/Y 0.03fF
C2922 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.15fF
C2923 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C2924 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# VDD 0.21fF
C2925 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C2926 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.08fF
C2927 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.04fF
C2928 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.04fF
C2929 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.13fF
C2930 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.04fF
C2931 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C2932 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C2933 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C2934 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.02fF
C2935 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.02fF
C2936 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# VDD 0.15fF
C2937 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.07fF
C2938 VDD p1 1.43fF
C2939 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.00fF
C2940 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C2941 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.01fF
C2942 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.01fF
C2943 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.02fF
C2944 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C2945 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C2946 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C2947 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C2948 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# VDD 0.11fF
C2949 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C2950 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C2951 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.03fF
C2952 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C2953 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C2954 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C2955 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.08fF
C2956 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.05fF
C2957 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X -0.00fF
C2958 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/S 0.05fF
C2959 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C2960 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.08fF
C2961 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.08fF
C2962 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C2963 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.08fF
C2964 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C2965 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C2966 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.11fF
C2967 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C2968 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C2969 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C2970 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C2971 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C2972 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.00fF
C2973 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.00fF
C2974 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C2975 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.07fF
C2976 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.02fF
C2977 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.11fF
C2978 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# VDD 0.33fF
C2979 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# VDD 0.51fF
C2980 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C2981 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C2982 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.02fF
C2983 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.07fF
C2984 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# -0.00fF
C2985 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# VDD 0.11fF
C2986 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.02fF
C2987 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__nand2_4_3/Y 0.19fF
C2988 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.04fF
C2989 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VDD 0.25fF
C2990 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C2991 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C2992 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C2993 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C2994 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C2995 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C2996 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C2997 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C2998 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/S 0.02fF
C2999 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C3000 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/X -0.19fF
C3001 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.04fF
C3002 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C3003 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.00fF
C3004 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C3005 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.05fF
C3006 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C3007 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C3008 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__nand2_1_1/A 0.03fF
C3009 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.18fF
C3010 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.14fF
C3011 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C3012 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C3013 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.04fF
C3014 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.02fF
C3015 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C3016 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.03fF
C3017 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C3018 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C3019 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C3020 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C3021 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C3022 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3023 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2 0.02fF
C3024 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.09fF
C3025 VDD sky130_fd_sc_hd__nand2_1_2/A 1.62fF
C3026 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_11/w_82_21# 0.05fF
C3027 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C3028 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C3029 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C3030 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.05fF
C3031 sky130_fd_sc_hd__mux2_1_0/X Bd_b 0.01fF
C3032 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C3033 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C3034 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C3035 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C3036 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C3037 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.02fF
C3038 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C3039 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# A -0.03fF
C3040 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.31fF
C3041 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C3042 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.07fF
C3043 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C3044 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C3045 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C3046 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C3047 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C3048 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.15fF
C3049 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C3050 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C3051 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C3052 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C3053 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C3054 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C3055 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C3056 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C3057 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.01fF
C3058 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.02fF
C3059 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.02fF
C3060 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C3061 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C3062 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C3063 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C3064 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.03fF
C3065 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# VDD 0.15fF
C3066 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C3067 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C3068 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C3069 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.98fF
C3070 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# VDD 0.15fF
C3071 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C3072 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C3073 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C3074 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C3075 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# VDD 0.31fF
C3076 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C3077 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C3078 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C3079 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.04fF
C3080 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VDD 1.56fF
C3081 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.02fF
C3082 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.02fF
C3083 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.04fF
C3084 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.04fF
C3085 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.05fF
C3086 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C3087 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C3088 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.00fF
C3089 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C3090 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C3091 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C3092 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C3093 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C3094 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C3095 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.04fF
C3096 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.04fF
C3097 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.02fF
C3098 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.11fF
C3099 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C3100 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.09fF
C3101 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.01fF
C3102 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C3103 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C3104 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.02fF
C3105 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.02fF
C3106 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C3107 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C3108 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C3109 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C3110 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C3111 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C3112 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.14fF
C3113 B Bd 0.20fF
C3114 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C3115 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.05fF
C3116 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.05fF
C3117 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C3118 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C3119 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C3120 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.07fF
C3121 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# VDD 0.16fF
C3122 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C3123 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.00fF
C3124 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C3125 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C3126 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C3127 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# VDD 0.14fF
C3128 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.00fF
C3129 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C3130 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C3131 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.01fF
C3132 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.08fF
C3133 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C3134 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VDD 0.08fF
C3135 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C3136 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_561_413# 0.01fF
C3137 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.07fF
C3138 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C3139 sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD 0.20fF
C3140 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C3141 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_1_2/B 0.05fF
C3142 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C3143 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C3144 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.07fF
C3145 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/X -0.32fF
C3146 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X sky130_fd_sc_hd__clkinv_4_2/Y 0.04fF
C3147 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.03fF
C3148 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.01fF
C3149 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C3150 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C3151 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C3152 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C3153 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 1.12fF
C3154 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.00fF
C3155 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.00fF
C3156 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C3157 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C3158 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C3159 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A -0.00fF
C3160 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C3161 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.07fF
C3162 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.19fF
C3163 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.17fF
C3164 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C3165 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.01fF
C3166 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.01fF
C3167 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.04fF
C3168 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.04fF
C3169 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.04fF
C3170 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VDD 0.14fF
C3171 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C3172 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C3173 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C3174 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.00fF
C3175 VDD sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.16fF
C3176 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.08fF
C3177 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.01fF
C3178 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C3179 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.04fF
C3180 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.04fF
C3181 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.33fF
C3182 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C3183 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X -0.00fF
C3184 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.01fF
C3185 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.01fF
C3186 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.01fF
C3187 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C3188 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C3189 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.02fF
C3190 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.00fF
C3191 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.15fF
C3192 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.06fF
C3193 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C3194 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C3195 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.04fF
C3196 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/Y 0.13fF
C3197 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C3198 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.10fF
C3199 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.16fF
C3200 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.03fF
C3201 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3202 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C3203 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C3204 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.04fF
C3205 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C3206 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.08fF
C3207 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 2.27fF
C3208 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C3209 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C3210 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C3211 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C3212 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.02fF
C3213 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.00fF
C3214 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C3215 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C3216 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.02fF
C3217 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.00fF
C3218 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C3219 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Bd_b 0.05fF
C3220 VDD sky130_fd_sc_hd__mux2_1_0/S 0.97fF
C3221 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C3222 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C3223 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C3224 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.08fF
C3225 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C3226 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.07fF
C3227 p2 sky130_fd_sc_hd__clkinv_4_3/Y 0.03fF
C3228 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.26fF
C3229 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C3230 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C3231 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD 0.75fF
C3232 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.14fF
C3233 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C3234 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__nand2_1_1/A 0.08fF
C3235 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/D 0.07fF
C3236 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.11fF
C3237 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.10fF
C3238 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C3239 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C3240 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# -0.01fF
C3241 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C3242 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C3243 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C3244 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C3245 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.03fF
C3246 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.05fF
C3247 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C3248 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/A 0.46fF
C3249 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.05fF
C3250 p1d_b p1d 0.47fF
C3251 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C3252 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C3253 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C3254 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C3255 A_b A 0.47fF
C3256 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# 0.11fF
C3257 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.05fF
C3258 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# 0.10fF
C3259 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.04fF
C3260 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VDD 0.53fF
C3261 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3262 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.02fF
C3263 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C3264 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C3265 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C3266 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.02fF
C3267 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C3268 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C3269 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C3270 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.05fF
C3271 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.05fF
C3272 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C3273 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_4_1/A 1.35fF
C3274 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C3275 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.02fF
C3276 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.02fF
C3277 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# VDD 0.14fF
C3278 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C3279 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C3280 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.03fF
C3281 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C3282 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.00fF
C3283 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C3284 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.02fF
C3285 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C3286 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C3287 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C3288 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C3289 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.05fF
C3290 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__nand2_1_2/B 0.02fF
C3291 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# VDD 0.14fF
C3292 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C3293 VDD sky130_fd_sc_hd__clkbuf_16_5/a_110_47# -0.09fF
C3294 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C3295 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.03fF
C3296 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C3297 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__nand2_4_2/A 0.13fF
C3298 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C3299 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.03fF
C3300 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C3301 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C3302 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C3303 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.09fF
C3304 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.02fF
C3305 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# VDD 0.11fF
C3306 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C3307 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C3308 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__nand2_4_3/Y 0.04fF
C3309 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.02fF
C3310 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD -0.23fF
C3311 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.15fF
C3312 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C3313 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C3314 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C3315 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C3316 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C3317 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C3318 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C3319 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C3320 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C3321 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_1/A 0.08fF
C3322 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C3323 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__mux2_1_0/S 0.11fF
C3324 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C3325 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C3326 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C3327 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C3328 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C3329 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.04fF
C3330 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.02fF
C3331 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C3332 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.15fF
C3333 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3334 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_1/A 0.18fF
C3335 sky130_fd_sc_hd__dfxbp_1_1/D VDD 0.62fF
C3336 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.08fF
C3337 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C3338 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# -0.17fF
C3339 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.02fF
C3340 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C3341 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C3342 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.41fF
C3343 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.02fF
C3344 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.02fF
C3345 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.07fF
C3346 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C3347 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C3348 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.08fF
C3349 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C3350 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.05fF
C3351 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/B 0.03fF
C3352 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# VDD 0.35fF
C3353 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.01fF
C3354 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD 1.66fF
C3355 sky130_fd_sc_hd__nand2_4_1/Y VDD 9.94fF
C3356 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.02fF
C3357 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.11fF
C3358 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.19fF
C3359 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# 0.07fF
C3360 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.00fF
C3361 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C3362 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C3363 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C3364 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.07fF
C3365 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C3366 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C3367 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.02fF
C3368 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.05fF
C3369 VDD p1_b 1.39fF
C3370 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3371 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C3372 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.30fF
C3373 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# VDD 0.15fF
C3374 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.04fF
C3375 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.03fF
C3376 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.02fF
C3377 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C3378 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkinv_1_2/Y 0.12fF
C3379 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# VDD 0.24fF
C3380 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C3381 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# VDD 0.25fF
C3382 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C3383 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C3384 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C3385 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# VDD 0.33fF
C3386 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C3387 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C3388 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C3389 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C3390 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VDD 0.35fF
C3391 p2d VDD 1.51fF
C3392 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C3393 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.03fF
C3394 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C3395 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C3396 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C3397 sky130_fd_sc_hd__clkinv_4_2/w_82_21# sky130_fd_sc_hd__clkinv_4_2/Y 0.05fF
C3398 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C3399 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C3400 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C3401 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C3402 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C3403 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C3404 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.04fF
C3405 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.08fF
C3406 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 1.39fF
C3407 sky130_fd_sc_hd__clkinv_4_7/w_82_21# sky130_fd_sc_hd__clkinv_4_7/Y -0.00fF
C3408 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3409 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C3410 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C3411 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C3412 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.04fF
C3413 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X -0.00fF
C3414 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C3415 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C3416 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.14fF
C3417 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C3418 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C3419 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C3420 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C3421 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.11fF
C3422 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C3423 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C3424 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C3425 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_3/A 0.07fF
C3426 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1 0.02fF
C3427 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.03fF
C3428 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# VDD 0.16fF
C3429 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3430 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C3431 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C3432 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C3433 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.12fF
C3434 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.02fF
C3435 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C3436 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# VDD 0.37fF
C3437 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C3438 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# VDD 0.14fF
C3439 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.02fF
C3440 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.02fF
C3441 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C3442 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C3443 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.04fF
C3444 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Ad_b 0.03fF
C3445 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C3446 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD -1.31fF
C3447 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C3448 sky130_fd_sc_hd__nand2_4_3/B VDD 0.47fF
C3449 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C3450 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C3451 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C3452 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.33fF
C3453 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.07fF
C3454 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C3455 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C3456 sky130_fd_sc_hd__dfxbp_1_0/Q_N Ad_b 0.01fF
C3457 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C3458 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.00fF
C3459 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C3460 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C3461 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C3462 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C3463 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C3464 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C3465 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C3466 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# -0.05fF
C3467 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_1_0/A 0.01fF
C3468 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C3469 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3470 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.01fF
C3471 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_0/A 0.22fF
C3472 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C3473 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# VDD 0.33fF
C3474 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.05fF
C3475 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.05fF
C3476 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/Y 0.05fF
C3477 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VDD 0.18fF
C3478 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.02fF
C3479 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C3480 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.02fF
C3481 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C3482 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C3483 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.18fF
C3484 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C3485 sky130_fd_sc_hd__mux2_1_0/a_76_199# Ad_b 0.02fF
C3486 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C3487 VDD sky130_fd_sc_hd__nand2_4_3/A 12.82fF
C3488 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C3489 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_3/A 0.47fF
C3490 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.03fF
C3491 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C3492 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 1.38fF
C3493 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C3494 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.04fF
C3495 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.04fF
C3496 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A -0.00fF
C3497 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.03fF
C3498 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C3499 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.13fF
C3500 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VDD 0.10fF
C3501 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.03fF
C3502 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.01fF
C3503 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3504 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.04fF
C3505 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C3506 sky130_fd_sc_hd__mux2_1_0/S Ad_b 0.17fF
C3507 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C3508 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C3509 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C3510 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C3511 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C3512 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C3513 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.45fF
C3514 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.04fF
C3515 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C3516 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C3517 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# -0.00fF
C3518 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C3519 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C3520 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.07fF
C3521 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C3522 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C3523 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C3524 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C3525 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C3526 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.15fF
C3527 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C3528 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C3529 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C3530 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.08fF
C3531 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.02fF
C3532 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.11fF
C3533 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C3534 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.01fF
C3535 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C3536 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C3537 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkinv_4_1/A 0.37fF
C3538 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C3539 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.18fF
C3540 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C3541 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/A 0.65fF
C3542 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.07fF
C3543 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.05fF
C3544 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__nand2_4_0/A 0.75fF
C3545 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# VDD 0.31fF
C3546 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C3547 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C3548 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.07fF
C3549 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# Ad_b 0.06fF
C3550 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C3551 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.03fF
C3552 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# VDD 0.15fF
C3553 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C3554 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.01fF
C3555 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.03fF
C3556 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C3557 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C3558 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C3559 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.03fF
C3560 sky130_fd_sc_hd__clkinv_4_1/Y VDD -0.41fF
C3561 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C3562 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.09fF
C3563 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C3564 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.04fF
C3565 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.04fF
C3566 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C3567 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.00fF
C3568 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.00fF
C3569 sky130_fd_sc_hd__nand2_1_1/A clk 0.06fF
C3570 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C3571 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C3572 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C3573 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C3574 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.05fF
C3575 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C3576 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C3577 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C3578 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C3579 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C3580 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C3581 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C3582 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.14fF
C3583 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C3584 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.02fF
C3585 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.02fF
C3586 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.01fF
C3587 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.00fF
C3588 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Ad_b 0.22fF
C3589 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C3590 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.06fF
C3591 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C3592 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C3593 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C3594 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C3595 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C3596 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.19fF
C3597 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C3598 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C3599 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C3600 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C3601 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C3602 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.08fF
C3603 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C3604 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.11fF
C3605 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.03fF
C3606 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.19fF
C3607 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.02fF
C3608 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# VDD 0.14fF
C3609 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.00fF
C3610 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# -0.04fF
C3611 VDD sky130_fd_sc_hd__clkinv_1_2/Y -1.35fF
C3612 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.08fF
C3613 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C3614 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C3615 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C3616 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C3617 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.00fF
C3618 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.02fF
C3619 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C3620 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.01fF
C3621 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.00fF
C3622 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C3623 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C3624 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.03fF
C3625 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C3626 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.01fF
C3627 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.07fF
C3628 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.05fF
C3629 p2 sky130_fd_sc_hd__clkinv_4_9/Y 0.04fF
C3630 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C3631 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C3632 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C3633 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C3634 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C3635 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__mux2_1_0/X 0.05fF
C3636 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C3637 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C3638 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C3639 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C3640 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.03fF
C3641 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C3642 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C3643 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.08fF
C3644 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_4_2/A 0.15fF
C3645 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A -0.00fF
C3646 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C3647 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.15fF
C3648 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C3649 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.00fF
C3650 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C3651 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VDD 0.31fF
C3652 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C3653 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.01fF
C3654 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C3655 sky130_fd_sc_hd__nand2_4_1/Y Ad_b 0.00fF
C3656 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C3657 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C3658 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.01fF
C3659 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# -0.00fF
C3660 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.03fF
C3661 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.01fF
C3662 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.01fF
C3663 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.01fF
C3664 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C3665 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C3666 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VDD 1.47fF
C3667 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.02fF
C3668 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.19fF
C3669 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C3670 VDD sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.34fF
C3671 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.11fF
C3672 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X -0.00fF
C3673 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A -0.00fF
C3674 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.31fF
C3675 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C3676 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C3677 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.02fF
C3678 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C3679 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C3680 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.02fF
C3681 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.02fF
C3682 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X -0.00fF
C3683 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_561_413# 0.01fF
C3684 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C3685 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C3686 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C3687 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A -0.00fF
C3688 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.15fF
C3689 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C3690 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C3691 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C3692 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.02fF
C3693 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C3694 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.04fF
C3695 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C3696 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.01fF
C3697 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C3698 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C3699 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.03fF
C3700 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Ad_b 0.03fF
C3701 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C3702 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.02fF
C3703 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C3704 VDD Ad_b 5.02fF
C3705 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C3706 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.38fF
C3707 p2_b p2 0.47fF
C3708 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.01fF
C3709 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C3710 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C3711 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C3712 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.62fF
C3713 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# VDD 0.36fF
C3714 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.04fF
C3715 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.03fF
C3716 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C3717 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.03fF
C3718 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C3719 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VDD 0.34fF
C3720 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__dfxbp_1_1/D 0.07fF
C3721 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__nand2_1_1/A 0.06fF
C3722 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C3723 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.06fF
C3724 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# -0.00fF
C3725 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.03fF
C3726 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.03fF
C3727 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C3728 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C3729 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C3730 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C3731 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_0/Y 0.03fF
C3732 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C3733 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C3734 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C3735 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.10fF
C3736 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.05fF
C3737 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VDD 0.36fF
C3738 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.02fF
C3739 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C3740 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C3741 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C3742 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.08fF
C3743 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C3744 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C3745 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C3746 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.06fF
C3747 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.04fF
C3748 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.04fF
C3749 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C3750 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C3751 sky130_fd_sc_hd__nand2_4_3/B Ad_b 0.04fF
C3752 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# 0.00fF
C3753 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C3754 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__nand2_4_2/A 0.13fF
C3755 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C3756 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.05fF
C3757 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C3758 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C3759 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.04fF
C3760 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C3761 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.03fF
C3762 sky130_fd_sc_hd__nand2_4_0/Y VDD 9.78fF
C3763 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.03fF
C3764 VDD sky130_fd_sc_hd__nand2_1_4/Y 0.44fF
C3765 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C3766 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.22fF
C3767 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_1_1/B 0.05fF
C3768 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C3769 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C3770 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C3771 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C3772 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.03fF
C3773 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/B 0.16fF
C3774 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# VDD 0.12fF
C3775 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# -0.05fF
C3776 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C3777 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C3778 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# Bd_b 0.12fF
C3779 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.05fF
C3780 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 1.84fF
C3781 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C3782 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# Bd_b 0.02fF
C3783 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C3784 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C3785 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C3786 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C3787 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C3788 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.11fF
C3789 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_1_3/A 0.09fF
C3790 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/B 0.14fF
C3791 sky130_fd_sc_hd__nand2_4_3/A Ad_b 0.32fF
C3792 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__nand2_1_4/B 0.16fF
C3793 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C3794 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_0/A 0.21fF
C3795 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C3796 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C3797 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C3798 VDD sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.65fF
C3799 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C3800 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.10fF
C3801 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C3802 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C3803 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C3804 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.02fF
C3805 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C3806 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.08fF
C3807 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.11fF
C3808 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.02fF
C3809 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.08fF
C3810 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.03fF
C3811 sky130_fd_sc_hd__nand2_4_1/B VDD 0.58fF
C3812 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.08fF
C3813 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# -0.16fF
C3814 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.06fF
C3815 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C3816 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C3817 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.10fF
C3818 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# VDD 0.31fF
C3819 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/Y 0.07fF
C3820 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.19fF
C3821 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C3822 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD 1.23fF
C3823 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.00fF
C3824 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# VDD 0.31fF
C3825 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# 0.05fF
C3826 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.02fF
C3827 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C3828 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C3829 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.03fF
C3830 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C3831 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1_b 0.06fF
C3832 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# -0.00fF
C3833 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# 0.07fF
C3834 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.03fF
C3835 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.00fF
C3836 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.01fF
C3837 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.01fF
C3838 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.10fF
C3839 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.03fF
C3840 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD 0.06fF
C3841 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C3842 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.15fF
C3843 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C3844 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C3845 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# VDD 0.15fF
C3846 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C3847 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C3848 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD 0.95fF
C3849 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VDD 5.27fF
C3850 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# VDD 0.17fF
C3851 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C3852 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C3853 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C3854 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C3855 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.01fF
C3856 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C3857 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C3858 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VDD 0.74fF
C3859 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.08fF
C3860 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# VDD 0.15fF
C3861 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C3862 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C3863 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C3864 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.03fF
C3865 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C3866 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# VDD 0.30fF
C3867 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# VDD 0.17fF
C3868 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.06fF
C3869 sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.05fF
C3870 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.07fF
C3871 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C3872 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X -0.00fF
C3873 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C3874 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkinv_1_1/Y 0.03fF
C3875 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C3876 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C3877 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C3878 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C3879 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.03fF
C3880 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C3881 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C3882 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C3883 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.01fF
C3884 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.15fF
C3885 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# VDD 0.32fF
C3886 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C3887 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.02fF
C3888 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.66fF
C3889 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# VDD 0.33fF
C3890 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C3891 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# p2d -0.04fF
C3892 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.02fF
C3893 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VDD 0.33fF
C3894 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.19fF
C3895 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.08fF
C3896 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C3897 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C3898 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C3899 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C3900 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.15fF
C3901 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.04fF
C3902 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.04fF
C3903 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.07fF
C3904 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.02fF
C3905 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_3/A 0.21fF
C3906 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C3907 Bd sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.12fF
C3908 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C3909 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C3910 B sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.02fF
C3911 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.05fF
C3912 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.05fF
C3913 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# VDD 0.21fF
C3914 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C3915 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C3916 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# VDD 0.31fF
C3917 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.08fF
C3918 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Bd_b 0.03fF
C3919 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3920 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.10fF
C3921 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C3922 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.07fF
C3923 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C3924 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C3925 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C3926 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.14fF
C3927 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.14fF
C3928 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C3929 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.08fF
C3930 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.08fF
C3931 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.07fF
C3932 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# -0.03fF
C3933 sky130_fd_sc_hd__dfxbp_1_0/Q_N Bd_b 0.01fF
C3934 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C3935 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3936 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# p2d 0.15fF
C3937 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C3938 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VDD 0.20fF
C3939 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374# 0.01fF
C3940 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C3941 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C3942 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.03fF
C3943 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C3944 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C3945 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_1/Y 0.20fF
C3946 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C3947 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C3948 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C3949 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C3950 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C3951 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.00fF
C3952 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C3953 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C3954 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C3955 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_1/A 2.16fF
C3956 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.34fF
C3957 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C3958 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C3959 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C3960 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C3961 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C3962 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C3963 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C3964 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C3965 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C3966 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.14fF
C3967 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# VDD 0.29fF
C3968 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C3969 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C3970 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C3971 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.04fF
C3972 sky130_fd_sc_hd__mux2_1_0/a_76_199# Bd_b 0.02fF
C3973 sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C3974 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.01fF
C3975 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C3976 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C3977 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.14fF
C3978 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.14fF
C3979 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__nand2_1_2/B 0.02fF
C3980 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C3981 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C3982 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# 0.10fF
C3983 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C3984 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C3985 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C3986 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C3987 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C3988 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C3989 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.04fF
C3990 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.04fF
C3991 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.02fF
C3992 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C3993 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A -0.00fF
C3994 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD 0.88fF
C3995 p2d_b p2 0.09fF
C3996 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.08fF
C3997 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.01fF
C3998 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C3999 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C4000 VDD sky130_fd_sc_hd__nand2_4_2/A 6.98fF
C4001 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VDD 1.12fF
C4002 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.02fF
C4003 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.18fF
C4004 sky130_fd_sc_hd__mux2_1_0/S Bd_b 0.12fF
C4005 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C4006 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C4007 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C4008 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C4009 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C4010 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C4011 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C4012 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C4013 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_8/Y 0.68fF
C4014 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.02fF
C4015 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C4016 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C4017 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C4018 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.03fF
C4019 p2 sky130_fd_sc_hd__nand2_4_1/A 0.17fF
C4020 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__nand2_4_2/A 0.13fF
C4021 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# VDD 0.27fF
C4022 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C4023 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.10fF
C4024 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C4025 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.00fF
C4026 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.00fF
C4027 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# VDD 0.38fF
C4028 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.03fF
C4029 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C4030 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C4031 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.09fF
C4032 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# Bd_b 0.05fF
C4033 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# Ad_b 0.07fF
C4034 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4035 sky130_fd_sc_hd__clkinv_4_10/Y p2_b 0.03fF
C4036 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# VDD 0.15fF
C4037 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.00fF
C4038 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C4039 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C4040 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C4041 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C4042 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.03fF
C4043 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C4044 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.04fF
C4045 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.04fF
C4046 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.08fF
C4047 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0.02fF
C4048 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C4049 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C4050 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.01fF
C4051 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.05fF
C4052 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C4053 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C4054 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C4055 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.00fF
C4056 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# -0.04fF
C4057 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C4058 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C4059 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C4060 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C4061 p1 p1d 0.20fF
C4062 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# -0.00fF
C4063 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__nand2_1_1/B 0.03fF
C4064 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.07fF
C4065 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C4066 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkinv_1_2/Y 0.03fF
C4067 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Bd_b 0.10fF
C4068 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.02fF
C4069 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.10fF
C4070 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C4071 Ad_b sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C4072 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.02fF
C4073 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.02fF
C4074 sky130_fd_sc_hd__clkinv_1_3/A p2 0.24fF
C4075 p1d_b sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.02fF
C4076 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.04fF
C4077 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.08fF
C4078 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C4079 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C4080 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.00fF
C4081 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.03fF
C4082 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.15fF
C4083 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.00fF
C4084 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.02fF
C4085 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C4086 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C4087 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.00fF
C4088 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.05fF
C4089 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C4090 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C4091 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C4092 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_592_47# -0.00fF
C4093 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C4094 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.04fF
C4095 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.05fF
C4096 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.37fF
C4097 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C4098 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C4099 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Ad_b 0.13fF
C4100 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__mux2_1_0/S 0.03fF
C4101 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.05fF
C4102 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_4/B 0.04fF
C4103 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.51fF
C4104 sky130_fd_sc_hd__nand2_4_1/B Ad_b 0.06fF
C4105 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 1.84fF
C4106 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.04fF
C4107 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C4108 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C4109 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VDD 0.18fF
C4110 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# VDD 0.30fF
C4111 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C4112 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C4113 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C4114 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C4115 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C4116 Bd sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.15fF
C4117 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# B_b 0.15fF
C4118 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C4119 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C4120 sky130_fd_sc_hd__nand2_4_1/Y Bd_b 0.22fF
C4121 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C4122 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_7/Y 0.02fF
C4123 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# B_b 0.12fF
C4124 B sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.12fF
C4125 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.08fF
C4126 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.02fF
C4127 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.02fF
C4128 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C4129 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C4130 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C4131 p2_b sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.12fF
C4132 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.01fF
C4133 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C4134 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C4135 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VDD 1.41fF
C4136 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C4137 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.02fF
C4138 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.14fF
C4139 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VDD 0.16fF
C4140 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C4141 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.03fF
C4142 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C4143 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A -0.00fF
C4144 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.10fF
C4145 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C4146 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C4147 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C4148 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C4149 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C4150 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C4151 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C4152 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4153 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C4154 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C4155 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C4156 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C4157 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C4158 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.01fF
C4159 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_7/A 0.72fF
C4160 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C4161 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Bd_b 0.03fF
C4162 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.02fF
C4163 VDD Bd_b 8.03fF
C4164 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C4165 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C4166 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C4167 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C4168 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C4169 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# VDD 0.17fF
C4170 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C4171 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C4172 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.04fF
C4173 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.15fF
C4174 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# VDD 0.31fF
C4175 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C4176 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C4177 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C4178 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4179 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__nand2_1_1/A 0.06fF
C4180 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.03fF
C4181 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.05fF
C4182 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VDD 0.35fF
C4183 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C4184 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C4185 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C4186 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.08fF
C4187 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C4188 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C4189 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 2.28fF
C4190 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.10fF
C4191 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# VDD 0.25fF
C4192 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.10fF
C4193 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C4194 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C4195 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VDD 0.08fF
C4196 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 1.55fF
C4197 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_1_4/B 0.04fF
C4198 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_1_2/Y 0.69fF
C4199 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C4200 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.08fF
C4201 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C4202 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C4203 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C4204 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C4205 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.03fF
C4206 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C4207 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C4208 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C4209 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# -0.03fF
C4210 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VDD 0.23fF
C4211 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C4212 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C4213 sky130_fd_sc_hd__clkinv_4_0/w_82_21# sky130_fd_sc_hd__clkinv_4_1/A 0.05fF
C4214 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C4215 sky130_fd_sc_hd__nand2_4_3/B Bd_b 0.03fF
C4216 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.04fF
C4217 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.04fF
C4218 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C4219 sky130_fd_sc_hd__clkinv_4_0/w_82_21# sky130_fd_sc_hd__nand2_4_0/A -0.43fF
C4220 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.34fF
C4221 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.03fF
C4222 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# 0.10fF
C4223 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C4224 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C4225 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.73fF
C4226 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C4227 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C4228 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.10fF
C4229 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C4230 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C4231 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__nand2_4_1/B 0.02fF
C4232 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.07fF
C4233 sky130_fd_sc_hd__clkinv_4_4/w_82_21# sky130_fd_sc_hd__clkinv_4_4/Y -0.00fF
C4234 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.32fF
C4235 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# VDD 0.07fF
C4236 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.15fF
C4237 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0.04fF
C4238 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.04fF
C4239 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.08fF
C4240 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C4241 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C4242 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VDD 0.53fF
C4243 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C4244 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C4245 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C4246 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C4247 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C4248 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C4249 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C4250 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C4251 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C4252 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_1_4/B 0.08fF
C4253 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD 1.53fF
C4254 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.08fF
C4255 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.00fF
C4256 sky130_fd_sc_hd__nand2_4_3/A Bd_b 0.27fF
C4257 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C4258 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C4259 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.07fF
C4260 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C4261 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C4262 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C4263 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.00fF
C4264 sky130_fd_sc_hd__clkinv_4_5/Y VDD 3.93fF
C4265 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C4266 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C4267 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C4268 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C4269 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/A -0.18fF
C4270 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.00fF
C4271 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.05fF
C4272 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C4273 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C4274 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.10fF
C4275 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VDD 0.32fF
C4276 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C4277 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VDD 0.38fF
C4278 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C4279 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.07fF
C4280 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# VDD 0.16fF
C4281 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.04fF
C4282 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.04fF
C4283 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.19fF
C4284 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# VDD 0.18fF
C4285 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.02fF
C4286 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C4287 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.02fF
C4288 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.29fF
C4289 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.02fF
C4290 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.19fF
C4291 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# VDD 0.33fF
C4292 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C4293 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.05fF
C4294 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# -0.01fF
C4295 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.03fF
C4296 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C4297 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.30fF
C4298 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.01fF
C4299 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C4300 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# -0.05fF
C4301 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C4302 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2_b 0.06fF
C4303 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C4304 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C4305 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# VDD 0.11fF
C4306 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C4307 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C4308 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C4309 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.08fF
C4310 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/Y 0.73fF
C4311 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C4312 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# VDD 0.15fF
C4313 VDD sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.42fF
C4314 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# VDD 0.11fF
C4315 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C4316 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.03fF
C4317 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C4318 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# VDD 0.26fF
C4319 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C4320 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.03fF
C4321 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C4322 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.04fF
C4323 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.04fF
C4324 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.02fF
C4325 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C4326 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C4327 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__nand2_1_1/B 0.03fF
C4328 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C4329 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C4330 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A -0.00fF
C4331 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.04fF
C4332 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# VDD 0.28fF
C4333 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C4334 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C4335 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 1.10fF
C4336 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C4337 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# VDD 0.15fF
C4338 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.08fF
C4339 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.08fF
C4340 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.19fF
C4341 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C4342 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C4343 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C4344 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__nand2_1_1/B 0.07fF
C4345 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.01fF
C4346 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.12fF
C4347 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4348 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C4349 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C4350 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.08fF
C4351 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C4352 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C4353 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C4354 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C4355 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C4356 p1d_b sky130_fd_sc_hd__clkinv_4_8/Y 0.03fF
C4357 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C4358 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C4359 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C4360 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.01fF
C4361 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.02fF
C4362 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# VDD 0.15fF
C4363 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.15fF
C4364 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.07fF
C4365 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# VDD 0.18fF
C4366 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C4367 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4368 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# VDD 0.27fF
C4369 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C4370 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.08fF
C4371 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.14fF
C4372 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C4373 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C4374 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.05fF
C4375 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A -0.00fF
C4376 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A 0.32fF
C4377 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C4378 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C4379 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C4380 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C4381 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C4382 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C4383 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C4384 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C4385 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C4386 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C4387 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C4388 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.03fF
C4389 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.01fF
C4390 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.00fF
C4391 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4392 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X -0.00fF
C4393 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C4394 p2d_b sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.03fF
C4395 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.11fF
C4396 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.03fF
C4397 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C4398 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C4399 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C4400 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C4401 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C4402 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C4403 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# -0.00fF
C4404 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.34fF
C4405 sky130_fd_sc_hd__clkinv_4_1/A VDD 4.19fF
C4406 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# VDD 0.14fF
C4407 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C4408 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C4409 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C4410 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.18fF
C4411 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C4412 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C4413 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C4414 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C4415 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C4416 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C4417 VDD sky130_fd_sc_hd__nand2_4_0/A 18.48fF
C4418 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B 0.12fF
C4419 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.19fF
C4420 sky130_fd_sc_hd__mux2_1_0/a_505_21# Bd_b 0.04fF
C4421 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C4422 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C4423 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C4424 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C4425 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.03fF
C4426 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C4427 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C4428 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.02fF
C4429 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C4430 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C4431 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C4432 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C4433 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C4434 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C4435 p1_b p1d 0.52fF
C4436 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C4437 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.02fF
C4438 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.07fF
C4439 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C4440 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C4441 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C4442 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C4443 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.08fF
C4444 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C4445 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C4446 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.05fF
C4447 p1d_b sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.06fF
C4448 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C4449 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C4450 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4451 Ad_b Bd_b 4.81fF
C4452 sky130_fd_sc_hd__nand2_4_0/B VDD 0.44fF
C4453 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C4454 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.08fF
C4455 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C4456 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C4457 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C4458 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C4459 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C4460 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.03fF
C4461 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C4462 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C4463 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.08fF
C4464 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.04fF
C4465 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C4466 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C4467 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C4468 VDD p1d 1.50fF
C4469 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C4470 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C4471 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C4472 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.02fF
C4473 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C4474 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# VDD 0.16fF
C4475 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C4476 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C4477 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C4478 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C4479 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C4480 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C4481 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.02fF
C4482 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# VDD 0.14fF
C4483 sky130_fd_sc_hd__nand2_1_1/B clk 0.00fF
C4484 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C4485 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A -0.00fF
C4486 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C4487 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C4488 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.08fF
C4489 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C4490 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C4491 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C4492 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# Bd_b 0.06fF
C4493 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4494 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C4495 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.02fF
C4496 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.13fF
C4497 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.03fF
C4498 B_b VDD 0.90fF
C4499 sky130_fd_sc_hd__clkinv_4_3/w_82_21# sky130_fd_sc_hd__clkinv_4_3/Y -0.00fF
C4500 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.07fF
C4501 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C4502 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C4503 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C4504 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.05fF
C4505 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.02fF
C4506 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.02fF
C4507 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C4508 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C4509 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C4510 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.00fF
C4511 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C4512 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C4513 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C4514 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.06fF
C4515 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C4516 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C4517 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.08fF
C4518 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.04fF
C4519 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C4520 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.01fF
C4521 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C4522 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C4523 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4524 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.03fF
C4525 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.01fF
C4526 sky130_fd_sc_hd__nand2_4_0/Y Bd_b 0.00fF
C4527 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# A 0.06fF
C4528 Ad sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.06fF
C4529 Bd_b sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C4530 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C4531 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C4532 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.02fF
C4533 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C4534 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.03fF
C4535 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.12fF
C4536 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.05fF
C4537 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VDD 1.41fF
C4538 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.05fF
C4539 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C4540 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C4541 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C4542 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C4543 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C4544 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C4545 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C4546 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C4547 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD 0.82fF
C4548 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C4549 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.00fF
C4550 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.09fF
C4551 sky130_fd_sc_hd__clkinv_4_11/w_82_21# sky130_fd_sc_hd__nand2_4_3/A -0.43fF
C4552 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C4553 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C4554 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__dfxbp_1_0/a_975_413# 0.01fF
C4555 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4556 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C4557 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C4558 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C4559 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C4560 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C4561 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Bd_b 0.14fF
C4562 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C4563 sky130_fd_sc_hd__clkinv_4_5/Y Ad_b 0.31fF
C4564 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C4565 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C4566 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.08fF
C4567 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C4568 sky130_fd_sc_hd__nand2_4_1/B Bd_b 0.07fF
C4569 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.01fF
C4570 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C4571 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C4572 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C4573 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VDD 0.16fF
C4574 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C4575 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# VDD 0.15fF
C4576 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.00fF
C4577 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.02fF
C4578 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C4579 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.04fF
C4580 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C4581 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C4582 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 2.24fF
C4583 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C4584 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.07fF
C4585 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C4586 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# VDD 0.34fF
C4587 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.02fF
C4588 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VDD 1.01fF
C4589 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C4590 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C4591 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.13fF
C4592 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.00fF
C4593 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_1/Y 0.33fF
C4594 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C4595 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C4596 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C4597 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C4598 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.04fF
C4599 p2d_b sky130_fd_sc_hd__clkbuf_16_12/a_110_47# 0.09fF
C4600 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_1_1/A 0.06fF
C4601 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.01fF
C4602 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C4603 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C4604 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.02fF
C4605 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4606 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_1_2/A 0.00fF
C4607 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.15fF
C4608 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.18fF
C4609 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C4610 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C4611 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_592_47# 0.00fF
C4612 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C4613 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C4614 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.04fF
C4615 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C4616 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 2.22fF
C4617 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C4618 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C4619 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C4620 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.07fF
C4621 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C4622 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A -0.00fF
C4623 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4624 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD 1.06fF
C4625 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.07fF
C4626 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.01fF
C4627 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# Ad_b 0.16fF
C4628 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_7/Y 0.14fF
C4629 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C4630 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C4631 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# -0.06fF
C4632 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.12fF
C4633 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X -0.00fF
C4634 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C4635 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VDD 0.34fF
C4636 VDD A 1.52fF
C4637 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# VDD 0.15fF
C4638 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C4639 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.14fF
C4640 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C4641 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.05fF
C4642 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 1.21fF
C4643 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C4644 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C4645 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# VDD 0.16fF
C4646 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C4647 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__nand2_1_1/A 0.07fF
C4648 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VDD 0.17fF
C4649 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# VDD 0.23fF
C4650 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.03fF
C4651 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C4652 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C4653 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C4654 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.03fF
C4655 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.03fF
C4656 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C4657 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C4658 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C4659 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.12fF
C4660 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.08fF
C4661 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# VDD 0.15fF
C4662 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C4663 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C4664 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# VDD 0.36fF
C4665 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_1_3/A 0.12fF
C4666 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VDD 0.11fF
C4667 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.05fF
C4668 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X -0.00fF
C4669 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.04fF
C4670 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__nand2_1_4/Y -0.05fF
C4671 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.03fF
C4672 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.01fF
C4673 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.33fF
C4674 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_1/A 0.91fF
C4675 sky130_fd_sc_hd__clkinv_4_1/Y B_b 0.03fF
C4676 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.18fF
C4677 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.02fF
C4678 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.02fF
C4679 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.15fF
C4680 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C4681 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C4682 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C4683 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C4684 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C4685 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C4686 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_4_1/B 0.11fF
C4687 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C4688 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C4689 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C4690 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C4691 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C4692 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.05fF
C4693 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.05fF
C4694 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C4695 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C4696 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C4697 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C4698 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.07fF
C4699 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.13fF
C4700 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C4701 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C4702 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.11fF
C4703 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_1/B 0.95fF
C4704 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C4705 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C4706 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C4707 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.14fF
C4708 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C4709 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C4710 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.08fF
C4711 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.08fF
C4712 sky130_fd_sc_hd__dfxbp_1_1/a_561_413# VDD 0.01fF
C4713 sky130_fd_sc_hd__clkinv_4_6/w_82_21# sky130_fd_sc_hd__nand2_4_2/A -0.43fF
C4714 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.00fF
C4715 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.31fF
C4716 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# 0.05fF
C4717 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.01fF
C4718 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C4719 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0.01fF
C4720 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.01fF
C4721 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_4/B 0.31fF
C4722 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.07fF
C4723 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C4724 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C4725 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C4726 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.03fF
C4727 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C4728 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C4729 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C4730 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C4731 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C4732 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C4733 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C4734 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C4735 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C4736 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VDD 1.12fF
C4737 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.02fF
C4738 Ad A_b 0.53fF
C4739 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C4740 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.14fF
C4741 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C4742 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C4743 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.03fF
C4744 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C4745 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.02fF
C4746 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD 1.38fF
C4747 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.10fF
C4748 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkinv_4_1/A 0.08fF
C4749 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.07fF
C4750 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C4751 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C4752 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.00fF
C4753 sky130_fd_sc_hd__nand2_1_1/A VDD 14.92fF
C4754 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD 1.48fF
C4755 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/A 0.48fF
C4756 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.04fF
C4757 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C4758 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C4759 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.09fF
C4760 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C4761 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A -0.00fF
C4762 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C4763 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C4764 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C4765 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C4766 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C4767 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.04fF
C4768 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C4769 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C4770 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C4771 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X -0.00fF
C4772 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.07fF
C4773 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.05fF
C4774 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.05fF
C4775 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C4776 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C4777 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.02fF
C4778 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C4779 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C4780 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C4781 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# -0.01fF
C4782 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# VDD 0.15fF
C4783 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C4784 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.01fF
C4785 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.03fF
C4786 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.13fF
C4787 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.16fF
C4788 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# VDD 0.17fF
C4789 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C4790 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# VDD 0.34fF
C4791 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_4/B 0.12fF
C4792 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# VDD 0.34fF
C4793 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C4794 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VDD 0.42fF
C4795 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C4796 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C4797 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C4798 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.10fF
C4799 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.01fF
C4800 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C4801 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C4802 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.18fF
C4803 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_7/Y 0.19fF
C4804 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C4805 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/Y 0.73fF
C4806 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C4807 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.04fF
C4808 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.09fF
C4809 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A 0.73fF
C4810 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.01fF
C4811 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.04fF
C4812 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.04fF
C4813 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# VDD 0.15fF
C4814 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C4815 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.02fF
C4816 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C4817 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# VDD 0.13fF
C4818 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.01fF
C4819 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.01fF
C4820 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.01fF
C4821 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# VDD 0.30fF
C4822 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C4823 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C4824 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.03fF
C4825 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VDD 1.17fF
C4826 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C4827 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C4828 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C4829 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C4830 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# VDD 0.14fF
C4831 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4832 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C4833 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VDD 1.36fF
C4834 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C4835 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C4836 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C4837 sky130_fd_sc_hd__clkinv_4_4/Y A_b 0.03fF
C4838 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.04fF
C4839 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.04fF
C4840 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# VDD 0.15fF
C4841 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C4842 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C4843 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y 0.16fF
C4844 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# -0.17fF
C4845 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.05fF
C4846 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# -0.04fF
C4847 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C4848 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C4849 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C4850 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_4_3/A 0.30fF
C4851 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.00fF
C4852 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C4853 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C4854 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C4855 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.09fF
C4856 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.05fF
C4857 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.05fF
C4858 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.03fF
C4859 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.13fF
C4860 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# VDD 0.31fF
C4861 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C4862 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.04fF
C4863 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.03fF
C4864 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.02fF
C4865 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# VDD 0.16fF
C4866 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C4867 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# VDD 0.36fF
C4868 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C4869 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C4870 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C4871 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C4872 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.05fF
C4873 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C4874 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1 -0.09fF
C4875 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.02fF
C4876 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.05fF
C4877 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.05fF
C4878 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_47# -0.00fF
C4879 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C4880 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C4881 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C4882 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C4883 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C4884 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C4885 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C4886 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C4887 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.02fF
C4888 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C4889 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4890 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C4891 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C4892 p1d_b sky130_fd_sc_hd__clkbuf_16_12/a_110_47# 0.02fF
C4893 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkinv_4_1/A 0.45fF
C4894 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_1/A 0.47fF
C4895 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.08fF
C4896 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_4_10/w_82_21# 0.04fF
C4897 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__nand2_4_0/A 2.18fF
C4898 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.05fF
C4899 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C4900 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C4901 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.02fF
C4902 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.02fF
C4903 sky130_fd_sc_hd__clkinv_4_1/w_82_21# sky130_fd_sc_hd__clkinv_4_1/Y 0.04fF
C4904 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.10fF
C4905 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C4906 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.04fF
C4907 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.04fF
C4908 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4909 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A -0.00fF
C4910 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.03fF
C4911 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C4912 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C4913 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C4914 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.07fF
C4915 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.01fF
C4916 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VDD 0.17fF
C4917 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X -0.00fF
C4918 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C4919 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C4920 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.02fF
C4921 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C4922 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VDD 0.32fF
C4923 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C4924 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C4925 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C4926 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C4927 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C4928 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C4929 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C4930 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C4931 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C4932 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C4933 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C4934 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# -0.00fF
C4935 VDD sky130_fd_sc_hd__clkinv_4_2/Y 0.80fF
C4936 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C4937 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.03fF
C4938 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.11fF
C4939 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C4940 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C4941 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C4942 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C4943 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C4944 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.02fF
C4945 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C4946 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clk 0.05fF
C4947 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C4948 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C4949 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C4950 sky130_fd_sc_hd__clkinv_4_8/w_82_21# sky130_fd_sc_hd__clkinv_4_8/Y -0.00fF
C4951 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C4952 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C4953 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C4954 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C4955 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C4956 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4957 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C4958 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.01fF
C4959 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.02fF
C4960 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C4961 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C4962 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C4963 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1d 0.12fF
C4964 A Ad_b 0.26fF
C4965 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C4966 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C4967 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C4968 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C4969 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C4970 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.08fF
C4971 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.00fF
C4972 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.00fF
C4973 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.02fF
C4974 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C4975 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# VDD 0.12fF
C4976 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C4977 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C4978 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C4979 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C4980 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# VDD 0.26fF
C4981 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C4982 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C4983 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# 0.11fF
C4984 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C4985 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C4986 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C4987 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.05fF
C4988 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__nand2_4_0/Y 0.26fF
C4989 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C4990 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C4991 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C4992 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C4993 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/B 0.11fF
C4994 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C4995 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C4996 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C4997 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.04fF
C4998 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.04fF
C4999 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_1/A 0.10fF
C5000 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# VDD 0.30fF
C5001 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VDD 0.25fF
C5002 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.01fF
C5003 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C5004 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C5005 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C5006 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.03fF
C5007 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.05fF
C5008 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C5009 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C5010 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C5011 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C5012 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C5013 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C5014 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C5015 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C5016 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C5017 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C5018 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C5019 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.05fF
C5020 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.01fF
C5021 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.01fF
C5022 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C5023 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.05fF
C5024 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.06fF
C5025 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.36fF
C5026 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C5027 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.02fF
C5028 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.18fF
C5029 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.15fF
C5030 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.04fF
C5031 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C5032 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.04fF
C5033 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C5034 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C5035 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.11fF
C5036 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VDD 1.58fF
C5037 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.02fF
C5038 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C5039 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C5040 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkinv_4_3/Y -0.00fF
C5041 sky130_fd_sc_hd__nand2_1_4/B clk 0.07fF
C5042 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C5043 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C5044 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C5045 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C5046 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C5047 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C5048 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C5049 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C5050 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C5051 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD 1.14fF
C5052 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.45fF
C5053 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C5054 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.04fF
C5055 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C5056 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Ad_b 0.07fF
C5057 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C5058 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C5059 sky130_fd_sc_hd__nand2_1_1/A Ad_b 0.55fF
C5060 sky130_fd_sc_hd__clkinv_4_5/Y Bd_b 0.46fF
C5061 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C5062 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# A 0.02fF
C5063 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C5064 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.23fF
C5065 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VDD 0.41fF
C5066 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C5067 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C5068 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C5069 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C5070 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C5071 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.01fF
C5072 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.02fF
C5073 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X Bd_b 0.00fF
C5074 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.02fF
C5075 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C5076 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C5077 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.11fF
C5078 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C5079 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C5080 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# VDD 0.16fF
C5081 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C5082 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.02fF
C5083 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C5084 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C5085 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# VDD 0.17fF
C5086 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.04fF
C5087 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C5088 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C5089 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C5090 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C5091 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# VDD 0.34fF
C5092 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.08fF
C5093 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.07fF
C5094 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C5095 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C5096 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_1_1/A 0.10fF
C5097 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VDD 1.12fF
C5098 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C5099 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C5100 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# -0.00fF
C5101 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C5102 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.11fF
C5103 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/a_975_413# 0.00fF
C5104 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_8/w_82_21# 0.03fF
C5105 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.19fF
C5106 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.14fF
C5107 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C5108 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.09fF
C5109 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C5110 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C5111 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C5112 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C5113 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C5114 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C5115 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C5116 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C5117 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.01fF
C5118 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VDD 0.33fF
C5119 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C5120 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.07fF
C5121 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.04fF
C5122 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C5123 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.03fF
C5124 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.07fF
C5125 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C5126 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C5127 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.11fF
C5128 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C5129 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# Bd_b 0.10fF
C5130 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C5131 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C5132 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.06fF
C5133 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C5134 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C5135 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VDD 0.17fF
C5136 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C5137 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# -0.03fF
C5138 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.01fF
C5139 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_4/Y 0.06fF
C5140 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C5141 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C5142 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C5143 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C5144 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# VDD 0.15fF
C5145 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 1.53fF
C5146 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C5147 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C5148 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C5149 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C5150 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VDD 0.15fF
C5151 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# VDD 0.12fF
C5152 sky130_fd_sc_hd__clkinv_4_5/w_82_21# sky130_fd_sc_hd__nand2_4_1/A -0.43fF
C5153 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VDD 5.11fF
C5154 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C5155 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C5156 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C5157 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C5158 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C5159 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C5160 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.06fF
C5161 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.04fF
C5162 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.04fF
C5163 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.02fF
C5164 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C5165 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# VDD 0.11fF
C5166 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C5167 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_1/Y 0.73fF
C5168 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C5169 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.02fF
C5170 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.04fF
C5171 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.04fF
C5172 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C5173 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# VDD 0.34fF
C5174 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VDD 0.31fF
C5175 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C5176 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C5177 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.07fF
C5178 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# 0.01fF
C5179 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.03fF
C5180 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.02fF
C5181 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.31fF
C5182 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 1.58fF
C5183 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.01fF
C5184 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.15fF
C5185 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.02fF
C5186 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.05fF
C5187 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.33fF
C5188 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C5189 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C5190 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C5191 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C5192 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C5193 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C5194 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.02fF
C5195 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.02fF
C5196 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# VDD 0.33fF
C5197 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.04fF
C5198 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.03fF
C5199 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C5200 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.02fF
C5201 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C5202 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C5203 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C5204 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.03fF
C5205 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C5206 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.00fF
C5207 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C5208 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C5209 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C5210 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 2.24fF
C5211 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C5212 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C5213 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C5214 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C5215 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C5216 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C5217 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C5218 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C5219 p2d_b sky130_fd_sc_hd__clkinv_4_9/Y 0.03fF
C5220 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C5221 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.05fF
C5222 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C5223 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.14fF
C5224 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C5225 sky130_fd_sc_hd__dfxbp_1_1/a_975_413# VDD 0.01fF
C5226 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.31fF
C5227 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C5228 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.18fF
C5229 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C5230 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.02fF
C5231 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.02fF
C5232 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C5233 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.32fF
C5234 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C5235 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.03fF
C5236 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C5237 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A -0.00fF
C5238 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.14fF
C5239 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C5240 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C5241 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C5242 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 1.46fF
C5243 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C5244 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.04fF
C5245 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C5246 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.12fF
C5247 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C5248 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C5249 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C5250 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD 1.51fF
C5251 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C5252 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C5253 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C5254 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C5255 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.14fF
C5256 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C5257 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C5258 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.18fF
C5259 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C5260 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C5261 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.03fF
C5262 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C5263 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C5264 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C5265 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C5266 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C5267 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C5268 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C5269 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C5270 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C5271 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C5272 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C5273 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.15fF
C5274 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C5275 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# VDD 0.14fF
C5276 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C5277 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C5278 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C5279 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# VDD 0.15fF
C5280 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C5281 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VDD 1.05fF
C5282 p2d_b p2_b 0.22fF
C5283 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# VDD 0.35fF
C5284 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# VDD 0.15fF
C5285 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C5286 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# -0.00fF
C5287 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C5288 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C5289 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.07fF
C5290 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C5291 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.04fF
C5292 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C5293 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.03fF
C5294 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.04fF
C5295 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.04fF
C5296 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C5297 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C5298 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.19fF
C5299 p1 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.12fF
C5300 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1_b 0.12fF
C5301 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.08fF
C5302 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_9/Y 0.68fF
C5303 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C5304 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C5305 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C5306 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C5307 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C5308 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C5309 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# VDD 0.12fF
C5310 B_b Bd_b 0.20fF
C5311 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.02fF
C5312 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.02fF
C5313 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C5314 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.11fF
C5315 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# VDD 0.15fF
C5316 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.66fF
C5317 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C5318 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.26fF
C5319 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.00fF
C5320 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C5321 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C5322 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# VDD 0.35fF
C5323 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C5324 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.15fF
C5325 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VDD 0.32fF
C5326 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C5327 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 2.38fF
C5328 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.04fF
C5329 VDD sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.22fF
C5330 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C5331 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C5332 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C5333 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C5334 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.07fF
C5335 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C5336 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C5337 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C5338 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VDD 0.11fF
C5339 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VDD 0.72fF
C5340 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.09fF
C5341 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C5342 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.00fF
C5343 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.00fF
C5344 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C5345 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C5346 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C5347 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.10fF
C5348 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C5349 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.10fF
C5350 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# -0.03fF
C5351 p2 sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C5352 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C5353 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.01fF
C5354 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C5355 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C5356 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.00fF
C5357 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C5358 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C5359 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C5360 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.02fF
C5361 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C5362 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.04fF
C5363 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C5364 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C5365 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.03fF
C5366 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C5367 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C5368 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# VDD 0.12fF
C5369 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C5370 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# 0.16fF
C5371 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C5372 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C5373 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.08fF
C5374 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# VDD 0.17fF
C5375 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C5376 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C5377 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# -0.00fF
C5378 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C5379 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__mux2_1_0/X 0.05fF
C5380 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkinv_1_2/Y 0.00fF
C5381 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.05fF
C5382 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# VDD 0.33fF
C5383 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C5384 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C5385 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C5386 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# p2 0.02fF
C5387 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C5388 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.00fF
C5389 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C5390 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C5391 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C5392 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C5393 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_1_4/B 0.49fF
C5394 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C5395 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.05fF
C5396 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.05fF
C5397 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C5398 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C5399 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C5400 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.00fF
C5401 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C5402 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.08fF
C5403 sky130_fd_sc_hd__clkinv_4_2/Y VSS 30.37fF
C5404 clk VSS 14.35fF
C5405 p1d VSS 14.33fF
C5406 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# VSS 1.44fF
C5407 sky130_fd_sc_hd__nand2_1_0/B VSS 19.83fF
C5408 sky130_fd_sc_hd__nand2_1_4/Y VSS 22.59fF
C5409 Bd_b VSS 34.14fF
C5410 Ad_b VSS 21.84fF
C5411 sky130_fd_sc_hd__mux2_1_0/S VSS -1.88fF
C5412 sky130_fd_sc_hd__mux2_1_0/X VSS 22.73fF
C5413 sky130_fd_sc_hd__mux2_1_0/a_439_47# VSS 0.18fF
C5414 sky130_fd_sc_hd__mux2_1_0/a_218_47# VSS 0.01fF
C5415 sky130_fd_sc_hd__mux2_1_0/a_505_21# VSS 0.30fF
C5416 sky130_fd_sc_hd__mux2_1_0/a_76_199# VSS 0.29fF
C5417 sky130_fd_sc_hd__nand2_1_4/B VSS 44.30fF
C5418 sky130_fd_sc_hd__nand2_1_4/a_113_47# VSS 0.01fF
C5419 sky130_fd_sc_hd__clkinv_1_2/Y VSS 21.34fF
C5420 sky130_fd_sc_hd__nand2_4_3/A VSS 35.15fF
C5421 sky130_fd_sc_hd__nand2_1_3/A VSS 29.65fF
C5422 sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS -0.00fF
C5423 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS 9.04fF
C5424 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# VSS 0.20fF
C5425 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# VSS 0.27fF
C5426 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# VSS 0.38fF
C5427 sky130_fd_sc_hd__clkinv_1_1/Y VSS 27.91fF
C5428 sky130_fd_sc_hd__nand2_4_2/A VSS 23.60fF
C5429 sky130_fd_sc_hd__nand2_1_2/A VSS 19.96fF
C5430 sky130_fd_sc_hd__nand2_1_2/B VSS 11.62fF
C5431 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS 9.08fF
C5432 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# VSS 0.20fF
C5433 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# VSS 0.27fF
C5434 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# VSS 0.38fF
C5435 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS 26.72fF
C5436 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# VSS 0.21fF
C5437 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# VSS 0.27fF
C5438 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# VSS 0.41fF
C5439 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS 23.14fF
C5440 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# VSS 0.20fF
C5441 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# VSS 0.27fF
C5442 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# VSS 0.41fF
C5443 p1_b VSS 14.95fF
C5444 sky130_fd_sc_hd__clkinv_4_7/Y VSS 20.23fF
C5445 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# VSS 1.58fF
C5446 sky130_fd_sc_hd__nand2_4_1/A VSS 35.42fF
C5447 sky130_fd_sc_hd__nand2_1_1/B VSS 13.67fF
C5448 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.01fF
C5449 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS 21.12fF
C5450 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# VSS 0.21fF
C5451 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# VSS 0.28fF
C5452 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# VSS 0.39fF
C5453 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS 24.98fF
C5454 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# VSS 0.22fF
C5455 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# VSS 0.29fF
C5456 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# VSS 0.42fF
C5457 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS 11.12fF
C5458 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# VSS 0.20fF
C5459 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# VSS 0.28fF
C5460 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# VSS 0.37fF
C5461 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS 20.04fF
C5462 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS 25.47fF
C5463 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# VSS 0.22fF
C5464 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# VSS 0.48fF
C5465 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# VSS 0.40fF
C5466 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS 14.40fF
C5467 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# VSS 0.22fF
C5468 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# VSS 0.28fF
C5469 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# VSS 0.36fF
C5470 p1 VSS 6.91fF
C5471 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# VSS 1.39fF
C5472 sky130_fd_sc_hd__nand2_4_0/A VSS 31.98fF
C5473 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS -0.00fF
C5474 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS 21.32fF
C5475 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# VSS 0.21fF
C5476 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# VSS 0.29fF
C5477 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# VSS 0.42fF
C5478 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS 23.36fF
C5479 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# VSS 0.22fF
C5480 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# VSS 0.28fF
C5481 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# VSS 0.36fF
C5482 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS 21.25fF
C5483 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# VSS 0.20fF
C5484 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# VSS 0.27fF
C5485 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# VSS 0.41fF
C5486 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# VSS 0.37fF
C5487 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# VSS 0.35fF
C5488 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# VSS 0.44fF
C5489 A VSS 27.07fF
C5490 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# VSS 1.44fF
C5491 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS 10.33fF
C5492 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# VSS 0.22fF
C5493 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# VSS 0.30fF
C5494 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# VSS 0.40fF
C5495 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS 26.70fF
C5496 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# VSS 0.22fF
C5497 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# VSS 0.29fF
C5498 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# VSS 0.42fF
C5499 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS 21.20fF
C5500 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# VSS 0.21fF
C5501 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# VSS 0.28fF
C5502 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# VSS 0.39fF
C5503 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS 14.63fF
C5504 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# VSS 0.21fF
C5505 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# VSS 0.29fF
C5506 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# VSS 0.42fF
C5507 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS 15.73fF
C5508 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# VSS 0.39fF
C5509 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# VSS 0.29fF
C5510 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# VSS 0.41fF
C5511 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS 14.89fF
C5512 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# VSS 0.21fF
C5513 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# VSS 0.47fF
C5514 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# VSS 0.39fF
C5515 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS 20.98fF
C5516 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# VSS 0.23fF
C5517 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# VSS 0.31fF
C5518 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# VSS 0.40fF
C5519 A_b VSS 15.02fF
C5520 sky130_fd_sc_hd__clkinv_4_4/Y VSS 20.23fF
C5521 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# VSS 1.58fF
C5522 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS 32.19fF
C5523 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS 23.70fF
C5524 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# VSS 0.38fF
C5525 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# VSS 0.27fF
C5526 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# VSS 0.41fF
C5527 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS 11.05fF
C5528 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS 5.11fF
C5529 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# VSS 0.21fF
C5530 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# VSS 0.47fF
C5531 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# VSS 0.37fF
C5532 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS 14.27fF
C5533 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS 16.07fF
C5534 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# VSS 0.20fF
C5535 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# VSS 0.46fF
C5536 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# VSS 0.38fF
C5537 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS 41.68fF
C5538 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# VSS 0.23fF
C5539 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# VSS 0.31fF
C5540 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# VSS 0.40fF
C5541 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# VSS 0.21fF
C5542 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# VSS 0.26fF
C5543 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# VSS 0.35fF
C5544 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS 17.03fF
C5545 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS 14.28fF
C5546 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# VSS 0.38fF
C5547 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# VSS 0.27fF
C5548 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# VSS 0.41fF
C5549 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS 21.61fF
C5550 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# VSS 0.20fF
C5551 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# VSS 0.27fF
C5552 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# VSS 0.41fF
C5553 Ad VSS 11.70fF
C5554 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# VSS 1.45fF
C5555 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# VSS 0.21fF
C5556 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# VSS 0.26fF
C5557 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# VSS 0.35fF
C5558 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS 41.81fF
C5559 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# VSS 0.21fF
C5560 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# VSS 0.28fF
C5561 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# VSS 0.39fF
C5562 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS 21.23fF
C5563 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# VSS 0.21fF
C5564 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# VSS 0.29fF
C5565 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# VSS 0.42fF
C5566 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS 10.76fF
C5567 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# VSS 0.21fF
C5568 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# VSS 0.28fF
C5569 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# VSS 0.39fF
C5570 sky130_fd_sc_hd__nand2_4_2/B VSS 38.23fF
C5571 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# VSS 0.19fF
C5572 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# VSS 0.27fF
C5573 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# VSS 0.39fF
C5574 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# VSS 0.37fF
C5575 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# VSS 0.35fF
C5576 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# VSS 0.44fF
C5577 sky130_fd_sc_hd__nand2_1_0/A VSS 18.50fF
C5578 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS 14.93fF
C5579 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# VSS 0.37fF
C5580 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# VSS 0.35fF
C5581 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# VSS 0.45fF
C5582 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS 21.04fF
C5583 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# VSS 0.22fF
C5584 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# VSS 0.30fF
C5585 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# VSS 0.40fF
C5586 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# VSS 0.18fF
C5587 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# VSS 0.26fF
C5588 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# VSS 0.41fF
C5589 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# VSS 1.64fF
C5590 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS 14.89fF
C5591 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# VSS 0.21fF
C5592 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# VSS 0.47fF
C5593 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# VSS 0.39fF
C5594 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS 24.99fF
C5595 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# VSS 0.22fF
C5596 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# VSS 0.30fF
C5597 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# VSS 0.40fF
C5598 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS 15.73fF
C5599 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# VSS 0.39fF
C5600 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# VSS 0.29fF
C5601 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# VSS 0.41fF
C5602 VDD VSS -37522.19fF
C5603 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS 11.40fF
C5604 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# VSS 0.19fF
C5605 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# VSS 0.26fF
C5606 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# VSS 0.37fF
C5607 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS 19.93fF
C5608 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# VSS 0.22fF
C5609 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# VSS 0.28fF
C5610 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# VSS 0.36fF
C5611 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# VSS 0.23fF
C5612 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# VSS 0.35fF
C5613 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# VSS 0.47fF
C5614 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS 15.73fF
C5615 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# VSS 0.39fF
C5616 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# VSS 0.29fF
C5617 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# VSS 0.42fF
C5618 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS 14.37fF
C5619 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# VSS 0.20fF
C5620 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# VSS 0.28fF
C5621 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# VSS 0.42fF
C5622 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS 19.55fF
C5623 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# VSS 0.22fF
C5624 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# VSS 0.30fF
C5625 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# VSS 0.40fF
C5626 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS 21.38fF
C5627 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# VSS 0.21fF
C5628 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# VSS 0.29fF
C5629 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# VSS 0.40fF
C5630 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VSS 1.55fF
C5631 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS 21.59fF
C5632 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# VSS 0.21fF
C5633 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# VSS 0.29fF
C5634 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# VSS 0.42fF
C5635 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS 14.27fF
C5636 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS 16.07fF
C5637 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# VSS 0.20fF
C5638 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# VSS 0.46fF
C5639 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# VSS 0.38fF
C5640 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS 11.06fF
C5641 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS 9.57fF
C5642 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# VSS 0.20fF
C5643 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# VSS 0.27fF
C5644 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# VSS 0.38fF
C5645 sky130_fd_sc_hd__clkinv_4_8/Y VSS 2.45fF
C5646 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# VSS 0.20fF
C5647 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# VSS 0.25fF
C5648 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# VSS 0.33fF
C5649 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# VSS 0.18fF
C5650 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# VSS 0.26fF
C5651 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# VSS 0.42fF
C5652 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS 16.79fF
C5653 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS 20.13fF
C5654 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# VSS 0.38fF
C5655 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# VSS 0.28fF
C5656 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# VSS 0.41fF
C5657 sky130_fd_sc_hd__clkinv_4_3/Y VSS 35.69fF
C5658 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# VSS 0.21fF
C5659 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# VSS 0.25fF
C5660 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# VSS 0.34fF
C5661 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# VSS 0.21fF
C5662 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# VSS 0.26fF
C5663 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# VSS 0.35fF
C5664 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS 10.65fF
C5665 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# VSS 0.22fF
C5666 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# VSS 0.30fF
C5667 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# VSS 0.40fF
C5668 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS 27.14fF
C5669 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS 20.30fF
C5670 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# VSS 0.38fF
C5671 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# VSS 0.27fF
C5672 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# VSS 0.41fF
C5673 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS 39.94fF
C5674 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# VSS 0.21fF
C5675 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# VSS 0.27fF
C5676 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# VSS 0.41fF
C5677 B_b VSS 20.35fF
C5678 sky130_fd_sc_hd__clkinv_4_1/Y VSS 38.67fF
C5679 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# VSS 1.51fF
C5680 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS 14.93fF
C5681 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# VSS 0.36fF
C5682 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# VSS 0.33fF
C5683 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# VSS 0.43fF
C5684 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# VSS 0.20fF
C5685 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# VSS 0.28fF
C5686 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# VSS 0.39fF
C5687 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS 14.39fF
C5688 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# VSS 0.22fF
C5689 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# VSS 0.28fF
C5690 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# VSS 0.36fF
C5691 sky130_fd_sc_hd__nand2_4_3/B VSS 50.93fF
C5692 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VSS 0.20fF
C5693 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VSS 0.28fF
C5694 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# VSS 0.41fF
C5695 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS 19.82fF
C5696 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS 16.63fF
C5697 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# VSS 0.22fF
C5698 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# VSS 0.47fF
C5699 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# VSS 0.39fF
C5700 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS 26.70fF
C5701 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# VSS 0.22fF
C5702 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# VSS 0.29fF
C5703 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# VSS 0.42fF
C5704 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS 48.73fF
C5705 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# VSS 0.22fF
C5706 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# VSS 0.30fF
C5707 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# VSS 0.40fF
C5708 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS 10.31fF
C5709 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# VSS 0.21fF
C5710 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# VSS 0.28fF
C5711 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# VSS 0.40fF
C5712 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS 24.89fF
C5713 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# VSS 0.22fF
C5714 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# VSS 0.31fF
C5715 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# VSS 0.40fF
C5716 Bd VSS 14.43fF
C5717 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# VSS 1.51fF
C5718 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS 35.95fF
C5719 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# VSS 0.21fF
C5720 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# VSS 0.29fF
C5721 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# VSS 0.40fF
C5722 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS 15.73fF
C5723 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# VSS 0.39fF
C5724 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# VSS 0.29fF
C5725 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# VSS 0.41fF
C5726 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS 14.44fF
C5727 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# VSS 0.20fF
C5728 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# VSS 0.28fF
C5729 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# VSS 0.42fF
C5730 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS 12.08fF
C5731 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# VSS 0.23fF
C5732 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# VSS 0.49fF
C5733 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# VSS 0.41fF
C5734 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS 15.06fF
C5735 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VSS 0.22fF
C5736 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VSS 0.31fF
C5737 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VSS 0.45fF
C5738 sky130_fd_sc_hd__nand2_4_1/B VSS 50.87fF
C5739 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# VSS 0.21fF
C5740 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# VSS 0.29fF
C5741 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# VSS 0.42fF
C5742 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS 14.41fF
C5743 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# VSS 0.20fF
C5744 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# VSS 0.28fF
C5745 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# VSS 0.42fF
C5746 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS 21.12fF
C5747 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# VSS 0.21fF
C5748 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# VSS 0.28fF
C5749 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# VSS 0.39fF
C5750 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# VSS 0.18fF
C5751 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# VSS 0.26fF
C5752 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# VSS 0.42fF
C5753 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS 36.15fF
C5754 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# VSS 0.20fF
C5755 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# VSS 0.27fF
C5756 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# VSS 0.41fF
C5757 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS 8.03fF
C5758 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# VSS 0.22fF
C5759 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# VSS 0.49fF
C5760 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# VSS 0.39fF
C5761 B VSS 14.35fF
C5762 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# VSS 1.48fF
C5763 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS 23.60fF
C5764 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# VSS 0.21fF
C5765 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# VSS 0.46fF
C5766 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# VSS 0.39fF
C5767 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# VSS 0.21fF
C5768 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# VSS 0.26fF
C5769 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# VSS 0.35fF
C5770 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS 52.63fF
C5771 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# VSS 0.21fF
C5772 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# VSS 0.27fF
C5773 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# VSS 0.41fF
C5774 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# VSS 0.18fF
C5775 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# VSS 0.26fF
C5776 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# VSS 0.41fF
C5777 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS 14.75fF
C5778 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# VSS 0.21fF
C5779 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# VSS 0.28fF
C5780 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# VSS 0.40fF
C5781 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS 41.52fF
C5782 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# VSS 0.21fF
C5783 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# VSS 0.29fF
C5784 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# VSS 0.40fF
C5785 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS 21.23fF
C5786 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# VSS 0.21fF
C5787 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# VSS 0.29fF
C5788 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# VSS 0.42fF
C5789 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS 24.97fF
C5790 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# VSS 0.21fF
C5791 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# VSS 0.28fF
C5792 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# VSS 0.39fF
C5793 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS 42.90fF
C5794 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# VSS 0.20fF
C5795 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# VSS 0.27fF
C5796 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# VSS 0.41fF
C5797 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS 21.16fF
C5798 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# VSS 0.23fF
C5799 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# VSS 0.31fF
C5800 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# VSS 0.40fF
C5801 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS 20.98fF
C5802 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# VSS 0.23fF
C5803 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# VSS 0.31fF
C5804 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# VSS 0.40fF
C5805 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS 13.86fF
C5806 sky130_fd_sc_hd__clkinv_1_3/Y VSS 27.99fF
C5807 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# VSS 0.21fF
C5808 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# VSS 0.29fF
C5809 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VSS 0.43fF
C5810 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS 14.67fF
C5811 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS 12.74fF
C5812 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# VSS 0.22fF
C5813 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# VSS 0.48fF
C5814 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# VSS 0.40fF
C5815 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS 15.00fF
C5816 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# VSS 0.23fF
C5817 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# VSS 0.33fF
C5818 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# VSS 0.46fF
C5819 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS 24.98fF
C5820 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# VSS 0.22fF
C5821 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# VSS 0.30fF
C5822 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# VSS 0.43fF
C5823 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS 21.20fF
C5824 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# VSS 0.21fF
C5825 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# VSS 0.28fF
C5826 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# VSS 0.39fF
C5827 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS 42.77fF
C5828 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# VSS 0.20fF
C5829 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# VSS 0.27fF
C5830 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# VSS 0.41fF
C5831 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS 20.42fF
C5832 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# VSS 0.20fF
C5833 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# VSS 0.28fF
C5834 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# VSS 0.42fF
C5835 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS 21.04fF
C5836 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# VSS 0.22fF
C5837 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# VSS 0.30fF
C5838 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# VSS 0.40fF
C5839 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS 24.95fF
C5840 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# VSS 0.21fF
C5841 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# VSS 0.28fF
C5842 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# VSS 0.42fF
C5843 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# VSS 0.22fF
C5844 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# VSS 0.28fF
C5845 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# VSS 0.36fF
C5846 sky130_fd_sc_hd__nand2_1_1/A VSS 54.21fF
C5847 sky130_fd_sc_hd__dfxbp_1_1/D VSS 7.77fF
C5848 sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# VSS -0.00fF
C5849 sky130_fd_sc_hd__dfxbp_1_1/a_592_47# VSS -0.08fF
C5850 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# VSS 0.05fF
C5851 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# VSS 0.16fF
C5852 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# VSS 0.19fF
C5853 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# VSS 0.35fF
C5854 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# VSS 0.16fF
C5855 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# VSS 0.16fF
C5856 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VSS 0.33fF
C5857 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VSS 0.53fF
C5858 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS 21.59fF
C5859 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# VSS 0.21fF
C5860 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# VSS 0.29fF
C5861 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# VSS 0.42fF
C5862 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS 14.84fF
C5863 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# VSS 0.21fF
C5864 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# VSS 0.46fF
C5865 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# VSS 0.39fF
C5866 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS 14.58fF
C5867 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# VSS 0.21fF
C5868 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# VSS 0.28fF
C5869 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# VSS 0.40fF
C5870 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS 10.65fF
C5871 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# VSS 0.22fF
C5872 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# VSS 0.30fF
C5873 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# VSS 0.40fF
C5874 sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS 0.21fF
C5875 sky130_fd_sc_hd__dfxbp_1_0/a_1017_47# VSS 0.01fF
C5876 sky130_fd_sc_hd__dfxbp_1_0/a_592_47# VSS 0.01fF
C5877 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VSS 0.08fF
C5878 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VSS 0.15fF
C5879 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VSS 0.21fF
C5880 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VSS 0.54fF
C5881 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VSS 0.19fF
C5882 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VSS 0.20fF
C5883 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VSS 0.39fF
C5884 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VSS 0.57fF
C5885 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS 14.69fF
C5886 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS 13.48fF
C5887 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# VSS 0.24fF
C5888 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# VSS 0.34fF
C5889 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# VSS 0.46fF
C5890 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS 21.33fF
C5891 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# VSS 0.22fF
C5892 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# VSS 0.29fF
C5893 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# VSS 0.42fF
C5894 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS 10.76fF
C5895 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# VSS 0.21fF
C5896 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# VSS 0.28fF
C5897 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# VSS 0.39fF
C5898 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS 21.28fF
C5899 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# VSS 0.20fF
C5900 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# VSS 0.27fF
C5901 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# VSS 0.41fF
C5902 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS 35.40fF
C5903 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# VSS 0.23fF
C5904 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# VSS 0.31fF
C5905 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# VSS 0.41fF
C5906 sky130_fd_sc_hd__clkinv_4_9/Y VSS 56.73fF
C5907 sky130_fd_sc_hd__nand2_4_3/Y VSS 101.42fF
C5908 sky130_fd_sc_hd__clkinv_4_9/w_82_21# VSS 0.00fF
C5909 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS 41.96fF
C5910 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# VSS 0.21fF
C5911 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# VSS 0.28fF
C5912 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# VSS 0.39fF
C5913 sky130_fd_sc_hd__clkinv_4_8/w_82_21# VSS 0.01fF
C5914 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS 14.64fF
C5915 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VSS 0.22fF
C5916 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VSS 0.29fF
C5917 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VSS 0.42fF
C5918 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS 14.65fF
C5919 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VSS 0.20fF
C5920 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VSS 0.27fF
C5921 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VSS 0.41fF
C5922 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS 35.74fF
C5923 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VSS 0.23fF
C5924 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VSS 0.31fF
C5925 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VSS 0.41fF
C5926 sky130_fd_sc_hd__clkinv_4_7/w_82_21# VSS 0.01fF
C5927 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS 48.87fF
C5928 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VSS 0.21fF
C5929 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VSS 0.29fF
C5930 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VSS 0.40fF
C5931 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS 41.21fF
C5932 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VSS 0.22fF
C5933 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VSS 0.31fF
C5934 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VSS 0.41fF
C5935 sky130_fd_sc_hd__clkinv_4_7/A VSS 65.30fF
C5936 sky130_fd_sc_hd__clkinv_4_6/w_82_21# VSS 0.00fF
C5937 sky130_fd_sc_hd__clkinv_4_5/Y VSS 85.79fF
C5938 sky130_fd_sc_hd__clkinv_4_5/w_82_21# VSS 0.01fF
C5939 sky130_fd_sc_hd__clkinv_4_4/w_82_21# VSS 0.01fF
C5940 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS 21.09fF
C5941 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VSS 0.22fF
C5942 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VSS 0.30fF
C5943 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VSS 0.40fF
C5944 sky130_fd_sc_hd__clkinv_4_3/w_82_21# VSS 0.01fF
C5945 sky130_fd_sc_hd__nand2_4_0/Y VSS 55.37fF
C5946 sky130_fd_sc_hd__clkinv_4_2/w_82_21# VSS 0.00fF
C5947 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS 20.81fF
C5948 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VSS 0.22fF
C5949 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VSS 0.30fF
C5950 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VSS 0.40fF
C5951 sky130_fd_sc_hd__nand2_4_3/a_27_47# VSS 0.33fF
C5952 sky130_fd_sc_hd__clkinv_4_1/A VSS 103.48fF
C5953 sky130_fd_sc_hd__clkinv_4_1/w_82_21# VSS -0.03fF
C5954 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VSS 0.22fF
C5955 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VSS 0.28fF
C5956 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VSS 0.35fF
C5957 sky130_fd_sc_hd__nand2_4_2/Y VSS 53.92fF
C5958 sky130_fd_sc_hd__nand2_4_2/a_27_47# VSS 0.30fF
C5959 sky130_fd_sc_hd__clkinv_4_0/w_82_21# VSS -0.00fF
C5960 sky130_fd_sc_hd__nand2_4_1/Y VSS 54.07fF
C5961 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.40fF
C5962 sky130_fd_sc_hd__nand2_4_0/B VSS 50.88fF
C5963 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VSS 0.19fF
C5964 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VSS 0.27fF
C5965 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VSS 0.39fF
C5966 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.31fF
C5967 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS 15.02fF
C5968 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VSS 0.19fF
C5969 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VSS 0.26fF
C5970 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VSS 0.38fF
C5971 sky130_fd_sc_hd__clkinv_4_11/w_82_21# VSS -0.00fF
C5972 p2 VSS 78.75fF
C5973 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VSS 1.51fF
C5974 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS 14.69fF
C5975 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS 13.72fF
C5976 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VSS 0.20fF
C5977 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VSS 0.27fF
C5978 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VSS 0.39fF
C5979 sky130_fd_sc_hd__clkinv_1_3/A VSS 78.59fF
C5980 sky130_fd_sc_hd__clkinv_4_10/w_82_21# VSS 0.00fF
C5981 p2_b VSS 14.93fF
C5982 sky130_fd_sc_hd__clkinv_4_10/Y VSS 20.31fF
C5983 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VSS 1.51fF
C5984 sky130_fd_sc_hd__clkinv_1_0/Y VSS 27.91fF
C5985 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VSS 0.19fF
C5986 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VSS 0.28fF
C5987 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VSS 0.40fF
C5988 p2d VSS 14.43fF
C5989 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VSS 1.51fF
C5990 p2d_b VSS 22.31fF
C5991 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VSS 1.56fF
C5992 p1d_b VSS 12.16fF
C5993 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VSS 1.63fF
.ends

.subckt switch_5t_mux4_flat in out en en_b a_300_216# VDD VSS
X0 out en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=1.0088e+12p pd=1.012e+07u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X1 a_300_216# en in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X2 in en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3 a_300_216# en in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 in en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X5 a_300_216# en_b in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_300_216# en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X7 a_300_216# en_b in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X8 in en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X9 in en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X10 a_300_216# en_b in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X11 a_300_216# en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.6384e+12p ps=2.02e+07u w=1.36e+06u l=150000u
X12 out en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X13 out en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X14 a_300_216# en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X15 out en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X16 in en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X17 a_300_216# en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X18 a_300_216# en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X19 out en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X20 out en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X21 in en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X22 a_300_216# en_b in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X23 a_300_216# en_b in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X24 a_300_216# en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X25 out en_b a_300_216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X26 a_300_216# en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
X27 in en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X28 in en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X29 a_300_216# en in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X30 a_300_216# en in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X31 out en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X32 a_300_216# en in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X33 in en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X34 in en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X35 a_300_216# en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X36 a_300_216# en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X37 out en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X38 a_300_216# en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X39 out en a_300_216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X40 a_300_216# en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 out in 0.43fF
C1 a_300_216# en_b 1.13fF
C2 out en_b 0.28fF
C3 VDD a_300_216# 2.14fF
C4 out VDD 0.86fF
C5 in en_b 0.78fF
C6 VDD in 1.13fF
C7 VDD en_b 3.32fF
C8 en a_300_216# 0.95fF
C9 out en 0.28fF
C10 en in 0.77fF
C11 en en_b 0.34fF
C12 out a_300_216# 7.40fF
C13 en VDD 0.24fF
C14 a_300_216# in 7.36fF
C15 en VSS 3.84fF
C16 out VSS 0.68fF
C17 in VSS 1.30fF
C18 en_b VSS 0.41fF
C19 VDD VSS 6.77fF
C20 a_300_216# VSS 2.12fF
.ends

.subckt a_mux4_en en in0 in1 in2 in3 sky130_fd_sc_hd__inv_1_0/Y switch_5t_mux4_1/en
+ sky130_fd_sc_hd__nand2_1_2/a_113_47# switch_5t_mux4_1/in switch_5t_mux4_1/en_b switch_5t_mux4_0/a_300_216#
+ switch_5t_mux4_3/en switch_5t_mux4_0/en sky130_fd_sc_hd__nand2_1_3/a_113_47# switch_5t_mux4_1/a_300_216#
+ switch_5t_mux4_2/a_300_216# sky130_fd_sc_hd__inv_1_1/Y switch_5t_mux4_3/a_300_216#
+ transmission_gate_3/en_b sky130_fd_sc_hd__nand2_1_0/a_113_47# switch_5t_mux4_2/en_b
+ switch_5t_mux4_3/in switch_5t_mux4_2/en out switch_5t_mux4_0/en_b s1 switch_5t_mux4_0/in
+ VDD s0 switch_5t_mux4_2/in switch_5t_mux4_3/en_b VSS sky130_fd_sc_hd__nand2_1_1/a_113_47#
Xswitch_5t_mux4_3 switch_5t_mux4_3/in out switch_5t_mux4_3/en switch_5t_mux4_3/en_b
+ switch_5t_mux4_3/a_300_216# VDD VSS switch_5t_mux4_flat
Xsky130_fd_sc_hd__inv_1_4 switch_5t_mux4_0/en switch_5t_mux4_0/en_b VSS VDD VSS VDD
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_5 switch_5t_mux4_2/en switch_5t_mux4_2/en_b VSS VDD VSS VDD
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_6 switch_5t_mux4_3/en switch_5t_mux4_3/en_b VSS VDD VSS VDD
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_8 transmission_gate_3/en_b en VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xtransmission_gate_0 en VDD transmission_gate_0/nmos_tgate_0/w_n646_n262# in0 switch_5t_mux4_0/in
+ transmission_gate_3/en_b VSS transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/nmos_tgate_0/w_n646_n262# in1 switch_5t_mux4_1/in
+ transmission_gate_3/en_b VSS transmission_gate
Xtransmission_gate_2 en VDD transmission_gate_2/nmos_tgate_0/w_n646_n262# in2 switch_5t_mux4_2/in
+ transmission_gate_3/en_b VSS transmission_gate
Xtransmission_gate_3 en VDD transmission_gate_3/nmos_tgate_0/w_n646_n262# in3 switch_5t_mux4_3/in
+ transmission_gate_3/en_b VSS transmission_gate
Xsky130_fd_sc_hd__nand2_1_0 s0 s1 VSS VDD switch_5t_mux4_3/en_b VSS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_1 s0 sky130_fd_sc_hd__inv_1_0/Y VSS VDD switch_5t_mux4_2/en_b
+ VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_2 s1 sky130_fd_sc_hd__inv_1_1/Y VSS VDD switch_5t_mux4_1/en_b
+ VSS VDD sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/Y
+ VSS VDD switch_5t_mux4_0/en_b VSS VDD sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/Y s0 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y s1 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_mux4_0 switch_5t_mux4_0/in out switch_5t_mux4_0/en switch_5t_mux4_0/en_b
+ switch_5t_mux4_0/a_300_216# VDD VSS switch_5t_mux4_flat
Xswitch_5t_mux4_1 switch_5t_mux4_1/in out switch_5t_mux4_1/en switch_5t_mux4_1/en_b
+ switch_5t_mux4_1/a_300_216# VDD VSS switch_5t_mux4_flat
Xswitch_5t_mux4_2 switch_5t_mux4_2/in out switch_5t_mux4_2/en switch_5t_mux4_2/en_b
+ switch_5t_mux4_2/a_300_216# VDD VSS switch_5t_mux4_flat
Xsky130_fd_sc_hd__inv_1_3 switch_5t_mux4_1/en switch_5t_mux4_1/en_b VSS VDD VSS VDD
+ sky130_fd_sc_hd__inv_1
C0 switch_5t_mux4_0/in transmission_gate_3/en_b 0.39fF
C1 out switch_5t_mux4_2/en 0.04fF
C2 switch_5t_mux4_0/en_b transmission_gate_3/en_b 0.05fF
C3 in1 VDD 0.10fF
C4 switch_5t_mux4_3/en switch_5t_mux4_3/a_300_216# -0.00fF
C5 switch_5t_mux4_1/en VDD 0.35fF
C6 s1 sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C7 switch_5t_mux4_1/in VDD 0.80fF
C8 s1 VDD 0.65fF
C9 switch_5t_mux4_1/en_b sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.01fF
C10 switch_5t_mux4_3/en_b switch_5t_mux4_2/in 0.09fF
C11 switch_5t_mux4_3/en_b switch_5t_mux4_2/en_b 0.38fF
C12 switch_5t_mux4_1/en_b VDD 0.34fF
C13 switch_5t_mux4_1/a_300_216# sky130_fd_sc_hd__inv_1_1/Y 0.02fF
C14 switch_5t_mux4_2/a_300_216# switch_5t_mux4_1/a_300_216# 0.30fF
C15 switch_5t_mux4_0/a_300_216# transmission_gate_3/en_b 0.02fF
C16 switch_5t_mux4_3/a_300_216# VDD 0.28fF
C17 sky130_fd_sc_hd__inv_1_0/Y VDD 0.88fF
C18 switch_5t_mux4_3/en VDD 0.34fF
C19 in0 in1 0.24fF
C20 switch_5t_mux4_0/in sky130_fd_sc_hd__inv_1_1/Y 0.02fF
C21 switch_5t_mux4_0/in s0 0.04fF
C22 in1 transmission_gate_3/en_b 0.31fF
C23 switch_5t_mux4_0/in en 0.23fF
C24 sky130_fd_sc_hd__inv_1_1/Y switch_5t_mux4_0/en_b 0.00fF
C25 out switch_5t_mux4_2/a_300_216# 0.34fF
C26 switch_5t_mux4_0/en_b s0 0.08fF
C27 switch_5t_mux4_2/in switch_5t_mux4_2/en_b 0.22fF
C28 in0 switch_5t_mux4_1/in 0.06fF
C29 switch_5t_mux4_1/en transmission_gate_3/en_b 0.01fF
C30 switch_5t_mux4_0/en_b en 0.07fF
C31 switch_5t_mux4_1/in transmission_gate_3/en_b 0.47fF
C32 s1 transmission_gate_3/en_b 1.15fF
C33 switch_5t_mux4_2/en switch_5t_mux4_1/en 0.17fF
C34 in2 switch_5t_mux4_2/in 0.00fF
C35 switch_5t_mux4_2/en switch_5t_mux4_1/in 0.02fF
C36 switch_5t_mux4_2/en s1 0.03fF
C37 switch_5t_mux4_1/en_b transmission_gate_3/en_b 0.04fF
C38 switch_5t_mux4_2/en switch_5t_mux4_1/en_b 0.44fF
C39 in3 VDD -0.11fF
C40 s0 sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C41 sky130_fd_sc_hd__inv_1_0/Y transmission_gate_3/en_b 0.10fF
C42 switch_5t_mux4_3/en transmission_gate_3/en_b 0.00fF
C43 switch_5t_mux4_2/en switch_5t_mux4_3/a_300_216# 0.01fF
C44 switch_5t_mux4_0/a_300_216# en 0.00fF
C45 switch_5t_mux4_2/en sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C46 switch_5t_mux4_3/en switch_5t_mux4_2/en 0.29fF
C47 out switch_5t_mux4_3/en_b 0.01fF
C48 sky130_fd_sc_hd__inv_1_1/Y in1 0.01fF
C49 in1 s0 0.01fF
C50 in1 en 0.31fF
C51 switch_5t_mux4_1/en sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C52 switch_5t_mux4_1/en s0 0.02fF
C53 switch_5t_mux4_3/en_b switch_5t_mux4_0/en_b 0.00fF
C54 switch_5t_mux4_1/in sky130_fd_sc_hd__inv_1_1/Y 0.07fF
C55 s1 sky130_fd_sc_hd__inv_1_1/Y 0.30fF
C56 switch_5t_mux4_1/in s0 0.07fF
C57 s1 s0 2.16fF
C58 switch_5t_mux4_1/in en 0.20fF
C59 s1 en 0.66fF
C60 s1 switch_5t_mux4_3/in 0.02fF
C61 switch_5t_mux4_2/in switch_5t_mux4_1/a_300_216# 0.06fF
C62 switch_5t_mux4_2/a_300_216# switch_5t_mux4_1/en 0.01fF
C63 switch_5t_mux4_2/en_b switch_5t_mux4_1/a_300_216# 0.01fF
C64 in0 VDD 0.03fF
C65 sky130_fd_sc_hd__inv_1_1/Y switch_5t_mux4_1/en_b 0.15fF
C66 switch_5t_mux4_2/a_300_216# switch_5t_mux4_1/in 0.07fF
C67 switch_5t_mux4_1/en_b s0 0.10fF
C68 switch_5t_mux4_2/a_300_216# s1 0.01fF
C69 switch_5t_mux4_1/en_b en 0.03fF
C70 VDD transmission_gate_3/en_b 0.93fF
C71 in3 transmission_gate_3/en_b 0.29fF
C72 switch_5t_mux4_2/a_300_216# switch_5t_mux4_1/en_b 0.05fF
C73 switch_5t_mux4_2/en VDD 0.32fF
C74 out switch_5t_mux4_2/en_b 0.04fF
C75 switch_5t_mux4_0/en switch_5t_mux4_1/a_300_216# 0.01fF
C76 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/Y 0.42fF
C77 sky130_fd_sc_hd__inv_1_0/Y s0 0.97fF
C78 switch_5t_mux4_2/in switch_5t_mux4_0/en_b 0.00fF
C79 switch_5t_mux4_3/a_300_216# switch_5t_mux4_3/in 0.02fF
C80 switch_5t_mux4_3/en s0 0.01fF
C81 switch_5t_mux4_2/en_b switch_5t_mux4_0/en_b 0.01fF
C82 sky130_fd_sc_hd__inv_1_0/Y en 0.07fF
C83 switch_5t_mux4_3/en switch_5t_mux4_3/in 0.11fF
C84 switch_5t_mux4_3/a_300_216# switch_5t_mux4_2/a_300_216# 0.30fF
C85 out switch_5t_mux4_0/en 0.01fF
C86 switch_5t_mux4_2/a_300_216# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C87 switch_5t_mux4_3/en switch_5t_mux4_2/a_300_216# 0.04fF
C88 switch_5t_mux4_0/in switch_5t_mux4_0/en 0.11fF
C89 switch_5t_mux4_0/en switch_5t_mux4_0/en_b 0.15fF
C90 in0 transmission_gate_3/en_b 0.23fF
C91 switch_5t_mux4_3/en_b s1 0.03fF
C92 switch_5t_mux4_2/en_b sky130_fd_sc_hd__nand2_1_1/a_113_47# -0.00fF
C93 sky130_fd_sc_hd__inv_1_1/Y VDD 0.72fF
C94 switch_5t_mux4_3/en_b switch_5t_mux4_1/en_b 0.01fF
C95 s0 VDD 0.85fF
C96 switch_5t_mux4_2/en transmission_gate_3/en_b 0.04fF
C97 en VDD 2.11fF
C98 switch_5t_mux4_3/in VDD 0.27fF
C99 en in3 0.28fF
C100 switch_5t_mux4_3/en_b sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.01fF
C101 switch_5t_mux4_3/in in3 0.00fF
C102 switch_5t_mux4_2/a_300_216# VDD 0.50fF
C103 switch_5t_mux4_2/in in1 0.06fF
C104 switch_5t_mux4_3/en_b switch_5t_mux4_3/a_300_216# 0.02fF
C105 switch_5t_mux4_0/en switch_5t_mux4_0/a_300_216# 0.07fF
C106 switch_5t_mux4_3/en_b sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C107 out switch_5t_mux4_1/a_300_216# 0.34fF
C108 switch_5t_mux4_2/in switch_5t_mux4_1/en 0.01fF
C109 switch_5t_mux4_3/en switch_5t_mux4_3/en_b 0.15fF
C110 switch_5t_mux4_2/en_b switch_5t_mux4_1/en 0.00fF
C111 switch_5t_mux4_0/in switch_5t_mux4_1/a_300_216# 0.07fF
C112 switch_5t_mux4_2/in switch_5t_mux4_1/in 0.30fF
C113 switch_5t_mux4_2/en_b switch_5t_mux4_1/in 0.01fF
C114 switch_5t_mux4_2/in s1 0.30fF
C115 switch_5t_mux4_2/en_b s1 0.07fF
C116 in2 in1 0.22fF
C117 switch_5t_mux4_1/a_300_216# switch_5t_mux4_0/en_b 0.07fF
C118 switch_5t_mux4_2/in switch_5t_mux4_1/en_b 0.03fF
C119 switch_5t_mux4_2/en_b switch_5t_mux4_1/en_b 0.23fF
C120 in2 switch_5t_mux4_1/in 0.07fF
C121 switch_5t_mux4_0/en switch_5t_mux4_1/en 0.20fF
C122 in2 s1 0.01fF
C123 switch_5t_mux4_0/en switch_5t_mux4_1/in 0.01fF
C124 switch_5t_mux4_0/en s1 0.03fF
C125 in0 en 0.18fF
C126 out switch_5t_mux4_0/en_b 0.03fF
C127 sky130_fd_sc_hd__inv_1_1/Y transmission_gate_3/en_b 0.04fF
C128 s0 transmission_gate_3/en_b 0.48fF
C129 switch_5t_mux4_0/in switch_5t_mux4_0/en_b 0.11fF
C130 switch_5t_mux4_0/en switch_5t_mux4_1/en_b 0.02fF
C131 en transmission_gate_3/en_b 2.59fF
C132 switch_5t_mux4_3/in transmission_gate_3/en_b 0.16fF
C133 switch_5t_mux4_2/in switch_5t_mux4_3/a_300_216# 0.07fF
C134 switch_5t_mux4_2/en_b switch_5t_mux4_3/a_300_216# 0.05fF
C135 switch_5t_mux4_2/in sky130_fd_sc_hd__inv_1_0/Y 0.08fF
C136 switch_5t_mux4_2/en s0 0.09fF
C137 switch_5t_mux4_2/en_b sky130_fd_sc_hd__inv_1_0/Y 0.04fF
C138 switch_5t_mux4_3/en switch_5t_mux4_2/in 0.04fF
C139 switch_5t_mux4_3/en switch_5t_mux4_2/en_b 0.56fF
C140 switch_5t_mux4_3/en_b VDD 0.19fF
C141 switch_5t_mux4_2/en en 0.03fF
C142 switch_5t_mux4_2/en switch_5t_mux4_3/in 0.04fF
C143 switch_5t_mux4_2/en switch_5t_mux4_2/a_300_216# 0.02fF
C144 in2 sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C145 switch_5t_mux4_1/a_300_216# switch_5t_mux4_0/a_300_216# 0.32fF
C146 switch_5t_mux4_0/en sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C147 switch_5t_mux4_0/en_b sky130_fd_sc_hd__nand2_1_3/a_113_47# -0.00fF
C148 out switch_5t_mux4_0/a_300_216# 0.20fF
C149 switch_5t_mux4_1/en switch_5t_mux4_1/a_300_216# 0.02fF
C150 switch_5t_mux4_0/in switch_5t_mux4_0/a_300_216# 0.10fF
C151 switch_5t_mux4_1/in switch_5t_mux4_1/a_300_216# 0.06fF
C152 switch_5t_mux4_2/in VDD 1.21fF
C153 switch_5t_mux4_2/en_b VDD 0.48fF
C154 switch_5t_mux4_2/in in3 0.07fF
C155 switch_5t_mux4_0/a_300_216# switch_5t_mux4_0/en_b 0.07fF
C156 switch_5t_mux4_1/a_300_216# switch_5t_mux4_1/en_b 0.08fF
C157 sky130_fd_sc_hd__inv_1_1/Y s0 0.29fF
C158 switch_5t_mux4_0/in in1 0.07fF
C159 sky130_fd_sc_hd__inv_1_1/Y en 0.03fF
C160 out switch_5t_mux4_1/en 0.04fF
C161 in2 VDD 0.07fF
C162 s0 en 0.55fF
C163 s0 switch_5t_mux4_3/in 0.01fF
C164 switch_5t_mux4_3/en_b transmission_gate_3/en_b 0.04fF
C165 in2 in3 0.22fF
C166 switch_5t_mux4_0/in switch_5t_mux4_1/en 0.09fF
C167 switch_5t_mux4_0/en VDD 0.23fF
C168 en switch_5t_mux4_3/in 0.17fF
C169 switch_5t_mux4_2/a_300_216# s0 0.02fF
C170 switch_5t_mux4_0/in switch_5t_mux4_1/in 0.45fF
C171 switch_5t_mux4_0/in s1 0.06fF
C172 switch_5t_mux4_2/en switch_5t_mux4_3/en_b 0.18fF
C173 switch_5t_mux4_1/en switch_5t_mux4_0/en_b 0.64fF
C174 switch_5t_mux4_2/a_300_216# switch_5t_mux4_3/in 0.06fF
C175 switch_5t_mux4_1/in switch_5t_mux4_0/en_b 0.10fF
C176 out switch_5t_mux4_1/en_b 0.04fF
C177 s1 switch_5t_mux4_0/en_b 0.07fF
C178 switch_5t_mux4_0/in switch_5t_mux4_1/en_b 0.04fF
C179 switch_5t_mux4_1/a_300_216# sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C180 switch_5t_mux4_0/en_b switch_5t_mux4_1/en_b 0.47fF
C181 out switch_5t_mux4_3/a_300_216# 0.14fF
C182 out switch_5t_mux4_3/en 0.03fF
C183 switch_5t_mux4_2/in transmission_gate_3/en_b 0.25fF
C184 switch_5t_mux4_2/en_b transmission_gate_3/en_b 0.04fF
C185 switch_5t_mux4_0/in sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C186 switch_5t_mux4_2/en switch_5t_mux4_2/in 0.09fF
C187 switch_5t_mux4_2/en switch_5t_mux4_2/en_b 0.60fF
C188 sky130_fd_sc_hd__inv_1_0/Y switch_5t_mux4_0/en_b 0.10fF
C189 in2 transmission_gate_3/en_b 0.32fF
C190 switch_5t_mux4_1/en switch_5t_mux4_0/a_300_216# 0.05fF
C191 switch_5t_mux4_1/in switch_5t_mux4_0/a_300_216# 0.06fF
C192 switch_5t_mux4_0/en transmission_gate_3/en_b 0.07fF
C193 switch_5t_mux4_1/a_300_216# VDD 0.54fF
C194 switch_5t_mux4_3/en_b s0 0.10fF
C195 switch_5t_mux4_3/en_b en 0.06fF
C196 switch_5t_mux4_3/en_b switch_5t_mux4_3/in 0.10fF
C197 switch_5t_mux4_0/a_300_216# switch_5t_mux4_1/en_b 0.02fF
C198 switch_5t_mux4_1/in in1 0.15fF
C199 switch_5t_mux4_3/en_b switch_5t_mux4_2/a_300_216# 0.05fF
C200 switch_5t_mux4_1/en switch_5t_mux4_1/in 0.11fF
C201 out VDD 1.58fF
C202 switch_5t_mux4_1/en s1 0.02fF
C203 switch_5t_mux4_1/in s1 0.08fF
C204 switch_5t_mux4_0/in VDD 1.07fF
C205 switch_5t_mux4_1/en switch_5t_mux4_1/en_b 0.22fF
C206 switch_5t_mux4_0/en_b VDD 0.13fF
C207 switch_5t_mux4_1/in switch_5t_mux4_1/en_b 0.31fF
C208 s1 switch_5t_mux4_1/en_b 0.27fF
C209 switch_5t_mux4_2/in sky130_fd_sc_hd__inv_1_1/Y 0.02fF
C210 switch_5t_mux4_2/en_b sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C211 switch_5t_mux4_2/in s0 0.46fF
C212 switch_5t_mux4_2/en_b s0 0.32fF
C213 switch_5t_mux4_2/in en 0.18fF
C214 switch_5t_mux4_2/en_b en 0.03fF
C215 switch_5t_mux4_2/in switch_5t_mux4_3/in 0.34fF
C216 switch_5t_mux4_2/en_b switch_5t_mux4_3/in 0.07fF
C217 switch_5t_mux4_2/in switch_5t_mux4_2/a_300_216# 0.02fF
C218 switch_5t_mux4_2/en_b switch_5t_mux4_2/a_300_216# 0.09fF
C219 switch_5t_mux4_1/en sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C220 in2 s0 0.00fF
C221 switch_5t_mux4_1/in sky130_fd_sc_hd__inv_1_0/Y 0.08fF
C222 sky130_fd_sc_hd__inv_1_0/Y s1 0.46fF
C223 in2 en 0.32fF
C224 switch_5t_mux4_0/en s0 0.03fF
C225 in2 switch_5t_mux4_3/in 0.06fF
C226 switch_5t_mux4_2/en switch_5t_mux4_1/a_300_216# 0.04fF
C227 switch_5t_mux4_0/en en 0.07fF
C228 sky130_fd_sc_hd__inv_1_0/Y switch_5t_mux4_1/en_b 0.19fF
C229 switch_5t_mux4_0/in in0 0.02fF
C230 switch_5t_mux4_0/a_300_216# VDD 0.45fF
C231 switch_5t_mux4_2/a_300_216# VSS 1.97fF
C232 switch_5t_mux4_1/en VSS 8.85fF
C233 switch_5t_mux4_1/a_300_216# VSS 1.97fF
C234 switch_5t_mux4_0/a_300_216# VSS 1.96fF
C235 sky130_fd_sc_hd__inv_1_0/Y VSS 42.07fF
C236 s1 VSS 46.15fF
C237 sky130_fd_sc_hd__inv_1_1/Y VSS 14.58fF
C238 switch_5t_mux4_0/en_b VSS 16.89fF
C239 sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS 0.01fF
C240 switch_5t_mux4_1/en_b VSS 16.29fF
C241 sky130_fd_sc_hd__nand2_1_2/a_113_47# VSS -0.00fF
C242 s0 VSS 46.08fF
C243 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.01fF
C244 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS -0.00fF
C245 en VSS 36.88fF
C246 switch_5t_mux4_3/in VSS 2.43fF
C247 in3 VSS 1.22fF
C248 VDD VSS -228.89fF
C249 switch_5t_mux4_2/in VSS 3.47fF
C250 in2 VSS 1.80fF
C251 transmission_gate_3/en_b VSS -3.38fF
C252 switch_5t_mux4_1/in VSS 2.26fF
C253 in1 VSS 1.81fF
C254 switch_5t_mux4_0/in VSS 3.65fF
C255 in0 VSS 1.89fF
C256 switch_5t_mux4_3/en VSS 4.74fF
C257 switch_5t_mux4_3/en_b VSS 6.22fF
C258 switch_5t_mux4_2/en VSS 9.63fF
C259 switch_5t_mux4_2/en_b VSS 12.63fF
C260 switch_5t_mux4_0/en VSS 4.31fF
C261 out VSS 6.86fF
C262 switch_5t_mux4_3/a_300_216# VSS 1.90fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TABSMU c1_n1210_n1160# m3_n1310_n1260# VSUBS
X0 c1_n1210_n1160# m3_n1310_n1260# sky130_fd_pr__cap_mim_m3_1 l=1.16e+07u w=1.16e+07u
C0 c1_n1210_n1160# m3_n1310_n1260# 13.72fF
C1 m3_n1310_n1260# VSUBS 4.03fF
.ends

.subckt sky130_fd_pr__pfet_01v8_VCQUSW a_n2818_n633# a_n4080_n100# a_n976_n730# a_2640_n100#
+ a_2010_n100# a_3852_131# a_2594_n401# a_1802_n633# a_n2866_n401# a_n2912_n100# a_n810_n633#
+ a_3600_n633# a_2548_n100# a_n182_n100# a_3644_n730# a_n3750_n633# a_n3120_n633#
+ a_n718_n633# a_n88_n633# a_n3916_n730# a_n3658_n633# a_n3028_n633# a_n1140_n100#
+ a_n1770_n100# a_n1398_n197# a_2172_131# a_n812_n100# a_n4128_131# a_n766_n401# a_3480_n100#
+ a_n3122_n100# a_n3752_n100# a_2012_n633# a_2642_n633# a_n2448_131# a_3388_n100#
+ a_3434_n401# a_240_n633# a_870_n633# a_284_n730# a_n3706_n401# a_492_131# a_n768_131#
+ a_3482_n633# a_n2238_n197# a_n1650_n633# a_n1020_n633# a_1500_n633# a_n2610_n100#
+ a_1544_n730# a_n1816_n730# a_n1558_n633# a_750_n100# a_120_n100# a_1380_n100# a_658_n100#
+ a_n510_n100# a_n1022_n100# a_n1652_n100# a_n138_n197# w_n4520_n852# a_2340_n633#
+ a_2970_n633# a_1288_n100# a_n3450_n100# a_n3078_n197# a_2384_n730# a_n2490_n633#
+ a_1334_n401# a_74_n401# a_702_n197# a_n2656_n730# a_n2398_n633# a_n1606_n401# a_1962_n197#
+ a_3012_131# a_1918_n100# a_28_n100# a_122_n633# a_752_n633# a_n2492_n100# a_1332_131#
+ a_n390_n633# a_1382_n633# a_n556_n730# a_3180_n633# a_2850_n100# a_2220_n100# a_n298_n633#
+ a_n3496_n730# a_2174_n401# a_n1608_131# a_n2446_n401# a_n3960_n633# a_n3330_n633#
+ a_3810_n633# a_2758_n100# a_2128_n100# a_n392_n100# a_3224_n730# a_n928_n633# a_2802_n197#
+ a_n3868_n633# a_n3238_n633# a_n1350_n100# a_n1980_n100# a_n346_n401# a_3690_n100#
+ a_3060_n100# a_2222_n633# a_2852_n633# a_n3332_n100# a_n3962_n100# a_2592_131# a_n3286_n401#
+ a_4020_n633# a_3598_n100# a_4064_n730# a_n4170_n633# a_3014_n401# a_n2868_131# a_450_n633#
+ a_n4078_n633# a_n2190_n100# a_3642_n197# a_1080_n633# a_n1396_n730# a_3062_n633#
+ a_3692_n633# a_n4172_n100# a_n2820_n100# a_1124_n730# a_n1860_n633# a_n1230_n633#
+ a_1710_n633# a_n1188_131# a_n4126_n401# a_960_n100# a_330_n100# a_n1768_n633# a_n1138_n633#
+ a_1590_n100# a_282_n197# a_n90_n100# a_n978_n197# a_n1186_n401# a_868_n100# a_238_n100#
+ a_n720_n100# a_n1232_n100# a_n1862_n100# a_n2070_n633# a_2550_n633# a_914_n401#
+ a_1498_n100# a_n3030_n100# a_n3660_n100# a_n2236_n730# a_1542_n197# a_n3918_n197#
+ a_n2700_n633# a_332_n633# a_962_n633# a_n2072_n100# a_3432_131# a_1592_n633# a_n2608_n633#
+ a_n136_n730# a_3390_n633# a_1752_131# a_2430_n100# a_n3076_n730# a_n2702_n100# a_n3708_131#
+ a_n600_n633# a_n2026_n401# a_2382_n197# a_2968_n100# a_2338_n100# a_n3540_n633#
+ a_n508_n633# a_n1560_n100# a_n3448_n633# a_3270_n100# a_n602_n100# a_n2028_131#
+ a_2432_n633# a_n3542_n100# a_n1818_n197# a_3178_n100# a_3900_n100# a_660_n633# a_3854_n401#
+ a_3222_n197# a_1290_n633# a_n348_131# a_3808_n100# a_704_n730# a_3272_n633# a_n2658_n197#
+ a_30_n633# a_1920_n633# a_n2400_n100# a_1964_n730# a_n1440_n633# a_n3288_131# a_4110_n100#
+ a_n1978_n633# a_n1348_n633# a_3902_n633# a_494_n401# a_540_n100# a_4062_n197# a_4018_n100#
+ a_1170_n100# a_72_131# a_n300_n100# a_n930_n100# a_n1442_n100# a_n558_n197# a_448_n100#
+ a_n3240_n100# a_n3870_n100# a_n3498_n197# a_n2280_n633# a_2130_n633# a_2760_n633#
+ a_1078_n100# a_1754_n401# a_1800_n100# a_4112_n633# a_1122_n197# a_n2188_n633# a_n2910_n633#
+ a_542_n633# a_1708_n100# a_912_131# a_2804_n730# VSUBS a_n180_n633# a_1172_n633#
+ a_n2282_n100#
X0 a_n90_n100# a_n138_n197# a_n182_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_330_n100# a_282_n197# a_238_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2 a_n88_n633# a_n136_n730# a_n180_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X3 a_1172_n633# a_1124_n730# a_1080_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X4 w_n4520_n852# w_n4520_n852# w_n4520_n852# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=2.48e+12p pd=2.096e+07u as=0p ps=0u w=1e+06u l=150000u
X5 a_n3450_n100# a_n3498_n197# a_n3542_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X6 a_3480_n100# a_3432_131# a_3388_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X7 a_3692_n633# a_3644_n730# a_3600_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X8 a_n1978_n633# a_n2026_n401# a_n2070_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X9 a_n1770_n100# a_n1818_n197# a_n1862_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X10 a_1800_n100# a_1752_131# a_1708_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X11 a_540_n100# a_492_131# a_448_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X12 a_2220_n100# a_2172_131# a_2128_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X13 a_n3658_n633# a_n3706_n401# a_n3750_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X14 a_n1138_n633# a_n1186_n401# a_n1230_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X15 a_n3660_n100# a_n3708_131# a_n3752_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X16 a_n300_n100# a_n348_131# a_n392_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X17 a_3690_n100# a_3642_n197# a_3598_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X18 a_4110_n100# a_4062_n197# a_4018_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X19 a_332_n633# a_284_n730# a_240_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X20 a_n298_n633# a_n346_n401# a_n390_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X21 a_1382_n633# a_1334_n401# a_1290_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X22 a_3902_n633# a_3854_n401# a_3810_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X23 a_n1980_n100# a_n2028_131# a_n2072_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X24 a_2010_n100# a_1962_n197# a_1918_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X25 a_n510_n100# a_n558_n197# a_n602_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X26 a_750_n100# a_702_n197# a_658_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X27 a_n2188_n633# a_n2236_n730# a_n2280_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X28 a_n3870_n100# a_n3918_n197# a_n3962_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X29 a_3900_n100# a_3852_131# a_3808_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X30 w_n4520_n852# w_n4520_n852# w_n4520_n852# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n3868_n633# a_n3916_n730# a_n3960_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X32 a_n1348_n633# a_n1396_n730# a_n1440_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X33 a_3062_n633# a_3014_n401# a_2970_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X34 a_n2190_n100# a_n2238_n197# a_n2282_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X35 a_542_n633# a_494_n401# a_450_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X36 a_2432_n633# a_2384_n730# a_2340_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X37 a_n720_n100# a_n768_131# a_n812_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X38 a_960_n100# a_912_131# a_868_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X39 a_n508_n633# a_n556_n730# a_n600_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X40 a_1592_n633# a_1544_n730# a_1500_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X41 a_2222_n633# a_2174_n401# a_2130_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X42 a_n4080_n100# a_n4128_131# a_n4172_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X43 a_n3028_n633# a_n3076_n730# a_n3120_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X44 a_n2398_n633# a_n2446_n401# a_n2490_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X45 a_n2400_n100# a_n2448_131# a_n2492_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X46 a_2430_n100# a_2382_n197# a_2338_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X47 a_n1558_n633# a_n1606_n401# a_n1650_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X48 w_n4520_n852# w_n4520_n852# w_n4520_n852# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_n930_n100# a_n978_n197# a_n1022_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X50 a_2642_n633# a_2594_n401# a_2550_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X51 a_3272_n633# a_3224_n730# a_3180_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X52 a_752_n633# a_704_n730# a_660_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X53 a_n1140_n100# a_n1188_131# a_n1232_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X54 a_1170_n100# a_1122_n197# a_1078_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X55 a_n4078_n633# a_n4126_n401# a_n4170_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X56 a_n718_n633# a_n766_n401# a_n810_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X57 a_1802_n633# a_1754_n401# a_1710_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X58 a_n2610_n100# a_n2658_n197# a_n2702_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X59 a_2640_n100# a_2592_131# a_2548_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X60 a_n3238_n633# a_n3286_n401# a_n3330_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X61 a_n3030_n100# a_n3078_n197# a_n3122_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X62 a_3060_n100# a_3012_131# a_2968_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X63 a_n2608_n633# a_n2656_n730# a_n2700_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X64 a_n1768_n633# a_n1816_n730# a_n1860_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X65 a_4112_n633# a_4064_n730# a_4020_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X66 a_n1350_n100# a_n1398_n197# a_n1442_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X67 a_1380_n100# a_1332_131# a_1288_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X68 a_962_n633# a_914_n401# a_870_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X69 a_2852_n633# a_2804_n730# a_2760_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X70 a_3482_n633# a_3434_n401# a_3390_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X71 a_n2820_n100# a_n2868_131# a_n2912_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X72 a_2850_n100# a_2802_n197# a_2758_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X73 a_n928_n633# a_n976_n730# a_n1020_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X74 a_n3240_n100# a_n3288_131# a_n3332_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X75 a_3270_n100# a_3222_n197# a_3178_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X76 w_n4520_n852# w_n4520_n852# w_n4520_n852# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_122_n633# a_74_n401# a_30_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X78 a_2012_n633# a_1964_n730# a_1920_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X79 a_n3448_n633# a_n3496_n730# a_n3540_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X80 a_n1560_n100# a_n1608_131# a_n1652_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X81 a_120_n100# a_72_131# a_28_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X82 a_1590_n100# a_1542_n197# a_1498_n100# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X83 a_n2818_n633# a_n2866_n401# a_n2910_n633# w_n4520_n852# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
C0 a_n3076_n730# a_n3496_n730# 0.01fF
C1 a_282_n197# a_n978_n197# 0.00fF
C2 a_2430_n100# a_1498_n100# 0.01fF
C3 a_3690_n100# a_2850_n100# 0.01fF
C4 a_3902_n633# a_2760_n633# 0.01fF
C5 a_3810_n633# a_2852_n633# 0.01fF
C6 a_n2700_n633# a_n3868_n633# 0.01fF
C7 a_n1230_n633# a_n1860_n633# 0.01fF
C8 a_n2026_n401# a_n2866_n401# 0.01fF
C9 a_n1860_n633# a_n2910_n633# 0.01fF
C10 a_1382_n633# a_962_n633# 0.02fF
C11 a_n3540_n633# a_n3658_n633# 0.07fF
C12 a_n3658_n633# w_n4520_n852# 0.04fF
C13 a_n1770_n100# a_n1980_n100# 0.03fF
C14 a_332_n633# a_330_n100# 0.00fF
C15 a_1920_n633# a_1918_n100# 0.00fF
C16 a_n2658_n197# a_n4128_131# 0.00fF
C17 a_2338_n100# a_1498_n100# 0.01fF
C18 a_n3540_n633# w_n4520_n852# 0.03fF
C19 a_3690_n100# a_2758_n100# 0.01fF
C20 a_3810_n633# a_2760_n633# 0.01fF
C21 a_3600_n633# a_2970_n633# 0.01fF
C22 a_3692_n633# a_2852_n633# 0.01fF
C23 a_n2818_n633# a_n3868_n633# 0.01fF
C24 a_1498_n100# a_868_n100# 0.01fF
C25 a_n2446_n401# a_n2866_n401# 0.01fF
C26 a_n1860_n633# a_n3028_n633# 0.01fF
C27 a_1290_n633# a_962_n633# 0.02fF
C28 a_1752_131# a_492_131# 0.00fF
C29 a_n1862_n100# a_n1980_n100# 0.07fF
C30 a_n1022_n100# a_n2610_n100# 0.00fF
C31 a_n3078_n197# a_n4128_131# 0.00fF
C32 a_n2700_n633# a_n2658_n197# 0.00fF
C33 a_2220_n100# a_1498_n100# 0.01fF
C34 a_3690_n100# a_2640_n100# 0.01fF
C35 a_1590_n100# a_540_n100# 0.01fF
C36 a_3692_n633# a_2760_n633# 0.01fF
C37 a_n2910_n633# a_n3868_n633# 0.01fF
C38 a_1498_n100# a_750_n100# 0.01fF
C39 a_n1860_n633# a_n3120_n633# 0.00fF
C40 a_1172_n633# a_962_n633# 0.03fF
C41 a_3272_n633# a_2432_n633# 0.01fF
C42 a_914_n401# w_n4520_n852# 0.10fF
C43 a_1288_n100# a_960_n100# 0.02fF
C44 a_240_n633# a_238_n100# 0.00fF
C45 a_n3498_n197# a_n4128_131# 0.00fF
C46 a_2128_n100# a_1498_n100# 0.01fF
C47 a_2804_n730# a_2174_n401# 0.00fF
C48 a_3690_n100# a_2548_n100# 0.01fF
C49 a_3900_n100# a_3598_n100# 0.02fF
C50 a_n1140_n100# a_n1770_n100# 0.01fF
C51 a_n3028_n633# a_n3868_n633# 0.01fF
C52 a_2548_n100# a_960_n100# 0.00fF
C53 a_2432_n633# a_962_n633# 0.00fF
C54 a_n1652_n100# a_n1608_131# 0.00fF
C55 a_n1768_n633# a_n3330_n633# 0.00fF
C56 a_n1860_n633# a_n3238_n633# 0.00fF
C57 a_3272_n633# a_2340_n633# 0.01fF
C58 a_n508_n633# a_n1138_n633# 0.01fF
C59 a_1382_n633# a_1334_n401# 0.00fF
C60 a_1498_n100# a_330_n100# 0.01fF
C61 a_n2702_n100# a_n3870_n100# 0.01fF
C62 a_n3918_n197# a_n4128_131# 0.01fF
C63 a_2010_n100# a_1498_n100# 0.01fF
C64 a_2804_n730# a_1754_n401# 0.00fF
C65 a_2384_n730# a_2174_n401# 0.01fF
C66 a_3690_n100# a_2430_n100# 0.00fF
C67 a_2642_n633# a_1592_n633# 0.01fF
C68 a_3808_n100# a_3598_n100# 0.03fF
C69 a_n1140_n100# a_n1862_n100# 0.01fF
C70 a_3900_n100# a_3480_n100# 0.02fF
C71 a_n558_n197# a_n1608_131# 0.00fF
C72 a_n3120_n633# a_n3868_n633# 0.01fF
C73 a_n1606_n401# a_n1608_131# 0.01fF
C74 a_2430_n100# a_960_n100# 0.00fF
C75 a_2340_n633# a_962_n633# 0.00fF
C76 a_n600_n633# a_n1138_n633# 0.01fF
C77 a_1290_n633# a_1334_n401# 0.00fF
C78 a_1498_n100# a_238_n100# 0.00fF
C79 a_n2820_n100# a_n3870_n100# 0.01fF
C80 a_1964_n730# a_2174_n401# 0.01fF
C81 a_n346_n401# a_n300_n100# 0.00fF
C82 a_1918_n100# a_1498_n100# 0.02fF
C83 a_2384_n730# a_1754_n401# 0.00fF
C84 a_1334_n401# a_1332_131# 0.01fF
C85 a_3690_n100# a_2338_n100# 0.00fF
C86 a_2550_n633# w_n4520_n852# 0.01fF
C87 a_2642_n633# a_1500_n633# 0.01fF
C88 a_n90_n100# a_n1652_n100# 0.00fF
C89 a_3900_n100# a_3388_n100# 0.01fF
C90 a_1288_n100# a_448_n100# 0.01fF
C91 a_3808_n100# a_3480_n100# 0.02fF
C92 a_n3238_n633# a_n3868_n633# 0.01fF
C93 a_n1560_n100# a_n2400_n100# 0.01fF
C94 a_2338_n100# a_960_n100# 0.00fF
C95 a_2852_n633# a_2804_n730# 0.00fF
C96 a_n2656_n730# a_n3916_n730# 0.00fF
C97 a_n2188_n633# a_n2236_n730# 0.00fF
C98 a_n718_n633# a_n1138_n633# 0.02fF
C99 a_30_n633# a_72_131# 0.00fF
C100 a_4112_n633# a_3482_n633# 0.01fF
C101 a_960_n100# a_868_n100# 0.09fF
C102 a_n2912_n100# a_n3870_n100# 0.01fF
C103 a_n138_n197# a_n768_131# 0.00fF
C104 a_1964_n730# a_1754_n401# 0.01fF
C105 a_1544_n730# a_2174_n401# 0.00fF
C106 a_3642_n197# w_n4520_n852# 0.09fF
C107 a_3690_n100# a_2220_n100# 0.00fF
C108 a_2642_n633# a_1382_n633# 0.00fF
C109 a_n3238_n633# a_n3286_n401# 0.00fF
C110 a_n182_n100# a_n1652_n100# 0.00fF
C111 a_3270_n100# a_2850_n100# 0.02fF
C112 a_3808_n100# a_3388_n100# 0.02fF
C113 a_2220_n100# a_960_n100# 0.00fF
C114 a_2760_n633# a_2804_n730# 0.00fF
C115 a_n88_n633# a_n508_n633# 0.02fF
C116 a_n2280_n633# a_n2236_n730# 0.00fF
C117 a_n2190_n100# a_n2400_n100# 0.03fF
C118 a_2222_n633# a_2174_n401# 0.00fF
C119 a_n2610_n100# a_n3752_n100# 0.01fF
C120 a_n810_n633# a_n1138_n633# 0.02fF
C121 a_4020_n633# a_3482_n633# 0.01fF
C122 a_960_n100# a_750_n100# 0.03fF
C123 a_4112_n633# a_3390_n633# 0.01fF
C124 a_n3030_n100# a_n3870_n100# 0.01fF
C125 a_702_n197# w_n4520_n852# 0.10fF
C126 a_n138_n197# a_n1188_131# 0.00fF
C127 a_n3120_n633# a_n3078_n197# 0.00fF
C128 a_1544_n730# a_1754_n401# 0.01fF
C129 a_3690_n100# a_2128_n100# 0.00fF
C130 a_4062_n197# a_3012_131# 0.00fF
C131 a_n2070_n633# a_n2072_n100# 0.00fF
C132 a_2642_n633# a_1290_n633# 0.00fF
C133 a_3180_n633# a_3178_n100# 0.00fF
C134 a_n300_n100# a_n1652_n100# 0.00fF
C135 a_3270_n100# a_2758_n100# 0.01fF
C136 a_2128_n100# a_960_n100# 0.01fF
C137 a_n180_n633# a_n508_n633# 0.02fF
C138 a_n88_n633# a_n600_n633# 0.01fF
C139 a_n1770_n100# w_n4520_n852# 0.02fF
C140 a_n2866_n401# a_n4126_n401# 0.00fF
C141 a_2130_n633# a_2174_n401# 0.00fF
C142 a_n928_n633# a_n1138_n633# 0.03fF
C143 a_962_n633# a_542_n633# 0.02fF
C144 a_3902_n633# a_3482_n633# 0.02fF
C145 a_4020_n633# a_3390_n633# 0.01fF
C146 a_n3122_n100# a_n3870_n100# 0.01fF
C147 a_1288_n100# a_658_n100# 0.01fF
C148 a_n390_n633# a_n348_131# 0.00fF
C149 a_2642_n633# a_1172_n633# 0.00fF
C150 a_960_n100# a_330_n100# 0.01fF
C151 a_868_n100# a_448_n100# 0.02fF
C152 a_3270_n100# a_2640_n100# 0.01fF
C153 a_3854_n401# a_3014_n401# 0.01fF
C154 a_n2400_n100# a_n2492_n100# 0.09fF
C155 a_n392_n100# a_n1652_n100# 0.00fF
C156 a_n3750_n633# a_n3960_n633# 0.03fF
C157 a_n978_n197# w_n4520_n852# 0.10fF
C158 a_1592_n633# a_752_n633# 0.01fF
C159 a_3012_131# a_2592_131# 0.01fF
C160 a_2010_n100# a_960_n100# 0.01fF
C161 a_704_n730# a_750_n100# 0.00fF
C162 a_n298_n633# a_n508_n633# 0.03fF
C163 a_n180_n633# a_n600_n633# 0.02fF
C164 a_n88_n633# a_n718_n633# 0.01fF
C165 a_n1862_n100# w_n4520_n852# 0.02fF
C166 a_28_n100# a_n1022_n100# 0.01fF
C167 a_n1020_n633# a_n1138_n633# 0.07fF
C168 a_962_n633# a_450_n633# 0.01fF
C169 a_n1860_n633# w_n4520_n852# 0.01fF
C170 a_3810_n633# a_3482_n633# 0.02fF
C171 a_3902_n633# a_3390_n633# 0.01fF
C172 a_n1652_n100# a_n2702_n100# 0.01fF
C173 a_1380_n100# a_120_n100# 0.00fF
C174 a_n3240_n100# a_n3870_n100# 0.01fF
C175 a_2642_n633# a_2432_n633# 0.03fF
C176 a_4064_n730# a_3854_n401# 0.01fF
C177 a_2852_n633# a_2222_n633# 0.01fF
C178 a_1800_n100# a_1380_n100# 0.02fF
C179 a_750_n100# a_448_n100# 0.02fF
C180 a_1078_n100# a_120_n100# 0.01fF
C181 a_960_n100# a_238_n100# 0.01fF
C182 a_3270_n100# a_2548_n100# 0.01fF
C183 a_n510_n100# a_n1652_n100# 0.01fF
C184 a_3854_n401# a_2594_n401# 0.00fF
C185 a_3434_n401# a_3014_n401# 0.01fF
C186 a_n1398_n197# w_n4520_n852# 0.10fF
C187 a_660_n633# w_n4520_n852# 0.01fF
C188 a_1500_n633# a_752_n633# 0.01fF
C189 a_1918_n100# a_960_n100# 0.01fF
C190 a_1800_n100# a_1078_n100# 0.01fF
C191 a_n180_n633# a_n718_n633# 0.01fF
C192 a_n298_n633# a_n600_n633# 0.02fF
C193 a_n390_n633# a_n508_n633# 0.07fF
C194 a_n88_n633# a_n810_n633# 0.01fF
C195 a_n90_n100# a_n1022_n100# 0.01fF
C196 a_2592_131# a_1332_131# 0.00fF
C197 a_3854_n401# a_3900_n100# 0.00fF
C198 a_3692_n633# a_3482_n633# 0.03fF
C199 a_3810_n633# a_3390_n633# 0.02fF
C200 a_n1652_n100# a_n2820_n100# 0.01fF
C201 a_n3332_n100# a_n3870_n100# 0.01fF
C202 a_n510_n100# a_n558_n197# 0.00fF
C203 a_2760_n633# a_2802_n197# 0.00fF
C204 a_4064_n730# a_3434_n401# 0.00fF
C205 a_2852_n633# a_2130_n633# 0.01fF
C206 a_2642_n633# a_2340_n633# 0.02fF
C207 a_2760_n633# a_2222_n633# 0.01fF
C208 a_3644_n730# a_3854_n401# 0.01fF
C209 a_n766_n401# a_n720_n100# 0.00fF
C210 a_n3658_n633# a_n3868_n633# 0.03fF
C211 a_2850_n100# a_1590_n100# 0.00fF
C212 a_1708_n100# a_1380_n100# 0.02fF
C213 a_n602_n100# a_n1652_n100# 0.01fF
C214 a_3270_n100# a_2430_n100# 0.01fF
C215 a_3434_n401# a_2594_n401# 0.01fF
C216 a_n1818_n197# w_n4520_n852# 0.10fF
C217 a_1382_n633# a_752_n633# 0.01fF
C218 a_n3540_n633# a_n3868_n633# 0.02fF
C219 a_1708_n100# a_1078_n100# 0.01fF
C220 a_448_n100# a_330_n100# 0.07fF
C221 a_n298_n633# a_n718_n633# 0.02fF
C222 a_n180_n633# a_n810_n633# 0.01fF
C223 a_n88_n633# a_n928_n633# 0.01fF
C224 a_n390_n633# a_n600_n633# 0.03fF
C225 a_n3868_n633# w_n4520_n852# 0.05fF
C226 a_122_n633# a_n1138_n633# 0.00fF
C227 a_n182_n100# a_n1022_n100# 0.01fF
C228 a_2010_n100# a_448_n100# 0.00fF
C229 a_284_n730# a_330_n100# 0.00fF
C230 a_3692_n633# a_3390_n633# 0.02fF
C231 a_n1652_n100# a_n2912_n100# 0.00fF
C232 a_n3330_n633# a_n3448_n633# 0.07fF
C233 a_4062_n197# a_3222_n197# 0.01fF
C234 a_868_n100# a_658_n100# 0.03fF
C235 a_n3450_n100# a_n3870_n100# 0.02fF
C236 a_n602_n100# a_n558_n197# 0.00fF
C237 a_n508_n633# a_n1440_n633# 0.01fF
C238 a_2852_n633# a_2012_n633# 0.01fF
C239 a_3644_n730# a_3434_n401# 0.01fF
C240 a_2760_n633# a_2130_n633# 0.01fF
C241 a_2758_n100# a_1590_n100# 0.01fF
C242 a_n720_n100# a_n1652_n100# 0.01fF
C243 a_3270_n100# a_2338_n100# 0.01fF
C244 a_n768_131# a_n2028_131# 0.00fF
C245 a_n2238_n197# w_n4520_n852# 0.10fF
C246 a_3690_n100# a_3178_n100# 0.01fF
C247 a_1290_n633# a_752_n633# 0.01fF
C248 a_n3286_n401# w_n4520_n852# 0.10fF
C249 a_n1980_n100# a_n2400_n100# 0.02fF
C250 a_2220_n100# a_658_n100# 0.00fF
C251 a_448_n100# a_238_n100# 0.03fF
C252 a_n1348_n633# a_n1978_n633# 0.01fF
C253 a_n298_n633# a_n810_n633# 0.01fF
C254 a_30_n633# a_n1138_n633# 0.01fF
C255 a_n390_n633# a_n718_n633# 0.02fF
C256 a_n180_n633# a_n928_n633# 0.01fF
C257 a_542_n633# a_494_n401# 0.00fF
C258 a_n88_n633# a_n1020_n633# 0.01fF
C259 a_1802_n633# a_1754_n401# 0.00fF
C260 a_n300_n100# a_n1022_n100# 0.01fF
C261 a_2382_n197# a_2592_131# 0.01fF
C262 a_n2610_n100# a_n2702_n100# 0.09fF
C263 a_870_n633# a_912_131# 0.00fF
C264 a_1918_n100# a_448_n100# 0.00fF
C265 a_n1652_n100# a_n3030_n100# 0.00fF
C266 a_750_n100# a_658_n100# 0.09fF
C267 a_n3542_n100# a_n3870_n100# 0.02fF
C268 a_n3658_n633# a_n3706_n401# 0.00fF
C269 a_n600_n633# a_n1440_n633# 0.01fF
C270 a_2760_n633# a_2012_n633# 0.01fF
C271 a_2852_n633# a_1920_n633# 0.01fF
C272 a_2640_n100# a_1590_n100# 0.01fF
C273 a_3222_n197# a_2592_131# 0.00fF
C274 a_3270_n100# a_2220_n100# 0.01fF
C275 a_n812_n100# a_n1652_n100# 0.01fF
C276 a_n1188_131# a_n2028_131# 0.01fF
C277 a_n2658_n197# w_n4520_n852# 0.10fF
C278 a_1080_n633# a_870_n633# 0.03fF
C279 a_1172_n633# a_752_n633# 0.02fF
C280 a_n3706_n401# w_n4520_n852# 0.10fF
C281 a_2128_n100# a_658_n100# 0.00fF
C282 a_n180_n633# a_n1020_n633# 0.01fF
C283 a_450_n633# a_494_n401# 0.00fF
C284 a_n390_n633# a_n810_n633# 0.02fF
C285 a_n298_n633# a_n928_n633# 0.01fF
C286 a_n1232_n100# a_n2282_n100# 0.01fF
C287 a_1288_n100# a_1590_n100# 0.02fF
C288 a_3062_n633# a_3014_n401# 0.00fF
C289 a_n392_n100# a_n1022_n100# 0.01fF
C290 a_1962_n197# a_2592_131# 0.00fF
C291 a_1710_n633# a_1754_n401# 0.00fF
C292 a_n2610_n100# a_n2820_n100# 0.03fF
C293 a_1122_n197# a_282_n197# 0.01fF
C294 a_n1652_n100# a_n3122_n100# 0.00fF
C295 a_n3660_n100# a_n3870_n100# 0.03fF
C296 a_284_n730# a_n976_n730# 0.00fF
C297 a_n718_n633# a_n1440_n633# 0.01fF
C298 a_2760_n633# a_1920_n633# 0.01fF
C299 a_2852_n633# a_1802_n633# 0.01fF
C300 a_2548_n100# a_1590_n100# 0.01fF
C301 a_3900_n100# a_2850_n100# 0.01fF
C302 a_n930_n100# a_n1652_n100# 0.01fF
C303 a_3270_n100# a_2128_n100# 0.01fF
C304 a_658_n100# a_330_n100# 0.02fF
C305 a_n3078_n197# w_n4520_n852# 0.10fF
C306 a_4112_n633# w_n4520_n852# 0.14fF
C307 a_122_n633# a_n88_n633# 0.03fF
C308 a_2010_n100# a_658_n100# 0.00fF
C309 a_n390_n633# a_n928_n633# 0.01fF
C310 a_n2448_131# a_n3708_131# 0.00fF
C311 a_n298_n633# a_n1020_n633# 0.01fF
C312 a_n510_n100# a_n1022_n100# 0.01fF
C313 a_n2610_n100# a_n2912_n100# 0.02fF
C314 a_n2866_n401# a_n2820_n100# 0.00fF
C315 a_n1652_n100# a_n3240_n100# 0.00fF
C316 a_n1140_n100# a_n2400_n100# 0.00fF
C317 a_n136_n730# a_n976_n730# 0.01fF
C318 a_n810_n633# a_n1440_n633# 0.01fF
C319 a_2852_n633# a_1710_n633# 0.01fF
C320 a_2760_n633# a_1802_n633# 0.01fF
C321 a_2430_n100# a_1590_n100# 0.01fF
C322 a_n3540_n633# a_n3498_n197# 0.00fF
C323 a_3900_n100# a_2758_n100# 0.01fF
C324 a_3808_n100# a_2850_n100# 0.01fF
C325 a_3270_n100# a_2010_n100# 0.00fF
C326 a_1170_n100# a_1122_n197# 0.00fF
C327 a_2340_n633# a_752_n633# 0.00fF
C328 a_658_n100# a_238_n100# 0.02fF
C329 a_2222_n633# a_870_n633# 0.00fF
C330 a_n3498_n197# w_n4520_n852# 0.11fF
C331 a_4020_n633# w_n4520_n852# 0.08fF
C332 a_122_n633# a_n180_n633# 0.02fF
C333 a_30_n633# a_n88_n633# 0.07fF
C334 a_282_n197# a_912_131# 0.00fF
C335 a_1918_n100# a_658_n100# 0.00fF
C336 a_n390_n633# a_n1020_n633# 0.01fF
C337 a_n602_n100# a_n1022_n100# 0.02fF
C338 a_28_n100# a_n90_n100# 0.07fF
C339 a_2594_n401# a_2640_n100# 0.00fF
C340 a_n2610_n100# a_n3030_n100# 0.02fF
C341 a_3600_n633# a_3272_n633# 0.02fF
C342 a_n1770_n100# a_n1862_n100# 0.09fF
C343 a_540_n100# a_120_n100# 0.02fF
C344 a_n556_n730# a_n976_n730# 0.01fF
C345 a_n928_n633# a_n1440_n633# 0.01fF
C346 a_n136_n730# a_n1396_n730# 0.00fF
C347 a_2760_n633# a_1710_n633# 0.01fF
C348 a_2338_n100# a_1590_n100# 0.01fF
C349 a_660_n633# a_702_n197# 0.00fF
C350 a_4018_n100# a_3598_n100# 0.02fF
C351 a_3808_n100# a_2758_n100# 0.01fF
C352 a_3900_n100# a_2640_n100# 0.00fF
C353 a_3388_n100# a_1800_n100# 0.00fF
C354 a_1800_n100# a_540_n100# 0.00fF
C355 a_3270_n100# a_1918_n100# 0.00fF
C356 a_2130_n633# a_870_n633# 0.00fF
C357 a_n1558_n633# a_n2070_n633# 0.01fF
C358 a_n3918_n197# w_n4520_n852# 0.11fF
C359 a_3598_n100# a_3060_n100# 0.01fF
C360 a_n766_n401# a_n768_131# 0.01fF
C361 a_3902_n633# w_n4520_n852# 0.06fF
C362 a_30_n633# a_n180_n633# 0.03fF
C363 a_122_n633# a_n298_n633# 0.02fF
C364 a_1590_n100# a_868_n100# 0.01fF
C365 a_n720_n100# a_n1022_n100# 0.02fF
C366 a_28_n100# a_n182_n100# 0.03fF
C367 a_n2610_n100# a_n3122_n100# 0.01fF
C368 a_n556_n730# a_n1396_n730# 0.01fF
C369 a_n1020_n633# a_n1440_n633# 0.02fF
C370 a_n1860_n633# a_n1862_n100# 0.00fF
C371 a_3062_n633# a_2970_n633# 0.09fF
C372 a_3180_n633# a_2852_n633# 0.02fF
C373 a_2220_n100# a_1590_n100# 0.01fF
C374 a_4018_n100# a_3480_n100# 0.01fF
C375 a_3808_n100# a_2640_n100# 0.01fF
C376 a_3900_n100# a_2548_n100# 0.00fF
C377 a_1708_n100# a_540_n100# 0.01fF
C378 a_2012_n633# a_870_n633# 0.01fF
C379 a_n1558_n633# a_n2188_n633# 0.01fF
C380 a_n1768_n633# a_n1978_n633# 0.03fF
C381 a_n1442_n100# a_n2282_n100# 0.01fF
C382 a_n1650_n633# a_n2070_n633# 0.02fF
C383 a_n978_n197# a_n1398_n197# 0.01fF
C384 a_3480_n100# a_3060_n100# 0.02fF
C385 a_122_n633# a_n390_n633# 0.01fF
C386 a_30_n633# a_n298_n633# 0.02fF
C387 a_3810_n633# w_n4520_n852# 0.05fF
C388 a_2220_n100# a_2172_131# 0.00fF
C389 a_1590_n100# a_750_n100# 0.01fF
C390 a_n1350_n100# a_n2282_n100# 0.01fF
C391 a_n812_n100# a_n1022_n100# 0.03fF
C392 a_28_n100# a_n300_n100# 0.02fF
C393 a_n90_n100# a_n182_n100# 0.09fF
C394 a_n2070_n633# a_n2608_n633# 0.01fF
C395 a_n1770_n100# a_n1818_n197# 0.00fF
C396 a_n2610_n100# a_n3240_n100# 0.01fF
C397 a_n1978_n633# a_n2026_n401# 0.00fF
C398 a_n556_n730# a_n1816_n730# 0.00fF
C399 a_3180_n633# a_2760_n633# 0.02fF
C400 a_3224_n730# a_2174_n401# 0.00fF
C401 a_2128_n100# a_1590_n100# 0.01fF
C402 a_4018_n100# a_3388_n100# 0.01fF
C403 a_3808_n100# a_2548_n100# 0.00fF
C404 a_3900_n100# a_2430_n100# 0.00fF
C405 a_1920_n633# a_870_n633# 0.01fF
C406 a_4112_n633# a_2550_n633# 0.00fF
C407 a_n2188_n633# a_n2190_n100# 0.00fF
C408 a_n1650_n633# a_n2188_n633# 0.01fF
C409 a_n1558_n633# a_n2280_n633# 0.01fF
C410 a_n558_n197# a_n768_131# 0.01fF
C411 a_n978_n197# a_n1818_n197# 0.01fF
C412 a_3270_n100# a_3178_n100# 0.09fF
C413 a_3388_n100# a_3060_n100# 0.02fF
C414 a_n1186_n401# a_n1188_131# 0.01fF
C415 a_30_n633# a_n390_n633# 0.02fF
C416 a_3692_n633# w_n4520_n852# 0.04fF
C417 a_752_n633# a_542_n633# 0.03fF
C418 a_2128_n100# a_2172_131# 0.00fF
C419 a_n930_n100# a_n1022_n100# 0.09fF
C420 a_n2070_n633# a_n2700_n633# 0.01fF
C421 a_n2188_n633# a_n2608_n633# 0.02fF
C422 a_28_n100# a_n392_n100# 0.02fF
C423 a_n90_n100# a_n300_n100# 0.03fF
C424 a_n1862_n100# a_n1818_n197# 0.00fF
C425 a_3482_n633# a_2222_n633# 0.00fF
C426 a_n2610_n100# a_n3332_n100# 0.01fF
C427 a_1590_n100# a_330_n100# 0.00fF
C428 a_n1860_n633# a_n1818_n197# 0.00fF
C429 a_122_n633# a_n1440_n633# 0.00fF
C430 a_n138_n197# a_n348_131# 0.01fF
C431 a_n2702_n100# a_n3752_n100# 0.01fF
C432 a_3224_n730# a_1754_n401# 0.00fF
C433 a_2010_n100# a_1590_n100# 0.02fF
C434 a_3808_n100# a_2430_n100# 0.00fF
C435 a_3900_n100# a_2338_n100# 0.00fF
C436 a_n2400_n100# w_n4520_n852# 0.02fF
C437 a_1802_n633# a_870_n633# 0.01fF
C438 a_n1650_n633# a_n2280_n633# 0.01fF
C439 a_4020_n633# a_2550_n633# 0.00fF
C440 a_n1558_n633# a_n2398_n633# 0.01fF
C441 a_n558_n197# a_n1188_131# 0.00fF
C442 a_n1398_n197# a_n1818_n197# 0.01fF
C443 a_n978_n197# a_n2238_n197# 0.00fF
C444 a_n2608_n633# a_n4078_n633# 0.00fF
C445 a_870_n633# a_332_n633# 0.01fF
C446 a_n138_n197# a_492_131# 0.00fF
C447 a_752_n633# a_450_n633# 0.02fF
C448 a_28_n100# a_n510_n100# 0.01fF
C449 a_n2280_n633# a_n2608_n633# 0.02fF
C450 a_3390_n633# a_2222_n633# 0.01fF
C451 a_3482_n633# a_2130_n633# 0.00fF
C452 a_n2070_n633# a_n2818_n633# 0.01fF
C453 a_n90_n100# a_n392_n100# 0.02fF
C454 a_n182_n100# a_n300_n100# 0.07fF
C455 a_n2188_n633# a_n2700_n633# 0.01fF
C456 a_1124_n730# a_2174_n401# 0.00fF
C457 a_n2610_n100# a_n3450_n100# 0.01fF
C458 a_1334_n401# a_1380_n100# 0.00fF
C459 a_1590_n100# a_238_n100# 0.00fF
C460 a_30_n633# a_n1440_n633# 0.00fF
C461 a_n2820_n100# a_n3752_n100# 0.01fF
C462 a_1918_n100# a_1590_n100# 0.02fF
C463 a_3808_n100# a_2338_n100# 0.00fF
C464 a_1710_n633# a_870_n633# 0.01fF
C465 a_3902_n633# a_2550_n633# 0.00fF
C466 a_n1558_n633# a_n2490_n633# 0.01fF
C467 a_n1650_n633# a_n2398_n633# 0.01fF
C468 a_1592_n633# a_1500_n633# 0.09fF
C469 a_n1398_n197# a_n2238_n197# 0.01fF
C470 a_n2700_n633# a_n4078_n633# 0.00fF
C471 a_870_n633# a_240_n633# 0.01fF
C472 a_n1230_n633# a_n2070_n633# 0.01fF
C473 a_n182_n100# a_n392_n100# 0.03fF
C474 a_3390_n633# a_2130_n633# 0.00fF
C475 a_n2188_n633# a_n2818_n633# 0.01fF
C476 a_3482_n633# a_2012_n633# 0.00fF
C477 a_n90_n100# a_n510_n100# 0.02fF
C478 a_n2070_n633# a_n2910_n633# 0.01fF
C479 a_28_n100# a_n602_n100# 0.01fF
C480 a_n2280_n633# a_n2700_n633# 0.02fF
C481 a_n2398_n633# a_n2608_n633# 0.03fF
C482 a_704_n730# a_2174_n401# 0.00fF
C483 a_1124_n730# a_1754_n401# 0.00fF
C484 a_n2610_n100# a_n3542_n100# 0.01fF
C485 a_n2912_n100# a_n3752_n100# 0.01fF
C486 a_4062_n197# a_3852_131# 0.01fF
C487 a_3808_n100# a_2220_n100# 0.00fF
C488 a_3810_n633# a_2550_n633# 0.00fF
C489 a_n1650_n633# a_n2490_n633# 0.01fF
C490 a_n1398_n197# a_n2658_n197# 0.00fF
C491 a_n1818_n197# a_n2238_n197# 0.01fF
C492 a_4110_n100# a_3690_n100# 0.02fF
C493 a_1592_n633# a_1382_n633# 0.03fF
C494 a_n2818_n633# a_n4078_n633# 0.00fF
C495 a_n1230_n633# a_n2188_n633# 0.01fF
C496 a_n90_n100# a_n602_n100# 0.01fF
C497 a_n2280_n633# a_n2818_n633# 0.01fF
C498 a_n2188_n633# a_n2910_n633# 0.01fF
C499 a_n2398_n633# a_n2700_n633# 0.02fF
C500 a_n2490_n633# a_n2608_n633# 0.07fF
C501 a_n300_n100# a_n392_n100# 0.09fF
C502 a_28_n100# a_n720_n100# 0.01fF
C503 a_3482_n633# a_1920_n633# 0.00fF
C504 a_n2070_n633# a_n3028_n633# 0.01fF
C505 a_n182_n100# a_n510_n100# 0.02fF
C506 a_3390_n633# a_2012_n633# 0.00fF
C507 a_704_n730# a_1754_n401# 0.00fF
C508 a_n2610_n100# a_n3660_n100# 0.01fF
C509 a_n3030_n100# a_n3752_n100# 0.01fF
C510 a_1122_n197# w_n4520_n852# 0.10fF
C511 a_332_n633# a_n1230_n633# 0.00fF
C512 a_4062_n197# a_3432_131# 0.00fF
C513 a_3692_n633# a_2550_n633# 0.01fF
C514 a_3600_n633# a_2642_n633# 0.01fF
C515 a_3178_n100# a_1590_n100# 0.00fF
C516 a_1592_n633# a_1290_n633# 0.02fF
C517 a_n1818_n197# a_n2658_n197# 0.01fF
C518 a_1500_n633# a_1382_n633# 0.07fF
C519 a_3852_131# a_2592_131# 0.00fF
C520 a_n2910_n633# a_n4078_n633# 0.01fF
C521 a_n1230_n633# a_n2280_n633# 0.01fF
C522 a_n90_n100# a_n720_n100# 0.01fF
C523 a_n2280_n633# a_n2910_n633# 0.01fF
C524 a_n2490_n633# a_n2700_n633# 0.03fF
C525 a_n300_n100# a_n510_n100# 0.03fF
C526 a_3390_n633# a_1920_n633# 0.00fF
C527 a_n182_n100# a_n602_n100# 0.02fF
C528 a_28_n100# a_n812_n100# 0.01fF
C529 a_n2188_n633# a_n3028_n633# 0.01fF
C530 a_n2398_n633# a_n2818_n633# 0.02fF
C531 a_n2070_n633# a_n3120_n633# 0.01fF
C532 a_284_n730# a_1754_n401# 0.00fF
C533 a_2804_n730# w_n4520_n852# 0.12fF
C534 a_n2490_n633# a_n2492_n100# 0.00fF
C535 a_962_n633# a_n508_n633# 0.00fF
C536 a_n3122_n100# a_n3752_n100# 0.01fF
C537 a_122_n633# a_120_n100# 0.00fF
C538 a_240_n633# a_n1230_n633# 0.00fF
C539 a_240_n633# a_282_n197# 0.00fF
C540 a_n2238_n197# a_n2658_n197# 0.01fF
C541 a_n1818_n197# a_n3078_n197# 0.00fF
C542 a_1500_n633# a_1290_n633# 0.03fF
C543 a_1592_n633# a_1172_n633# 0.02fF
C544 a_n3028_n633# a_n4078_n633# 0.01fF
C545 a_3432_131# a_2592_131# 0.01fF
C546 a_n3330_n633# a_n3332_n100# 0.00fF
C547 a_330_n100# a_n1232_n100# 0.00fF
C548 a_n1230_n633# a_n2398_n633# 0.01fF
C549 a_n3286_n401# a_n3706_n401# 0.01fF
C550 a_n2280_n633# a_n3028_n633# 0.01fF
C551 a_3390_n633# a_1802_n633# 0.00fF
C552 a_n182_n100# a_n720_n100# 0.01fF
C553 a_28_n100# a_n930_n100# 0.01fF
C554 a_n392_n100# a_n510_n100# 0.07fF
C555 a_n2490_n633# a_n2818_n633# 0.02fF
C556 a_n2188_n633# a_n3120_n633# 0.01fF
C557 a_n300_n100# a_n602_n100# 0.02fF
C558 a_n2398_n633# a_n2910_n633# 0.01fF
C559 a_n90_n100# a_n812_n100# 0.01fF
C560 a_n2070_n633# a_n3238_n633# 0.01fF
C561 a_n1978_n633# a_n3330_n633# 0.00fF
C562 a_2384_n730# w_n4520_n852# 0.12fF
C563 a_912_131# w_n4520_n852# 0.12fF
C564 a_962_n633# a_n600_n633# 0.00fF
C565 a_n3240_n100# a_n3752_n100# 0.01fF
C566 a_2850_n100# a_1800_n100# 0.01fF
C567 a_2432_n633# a_1592_n633# 0.01fF
C568 a_n2238_n197# a_n3078_n197# 0.01fF
C569 a_1382_n633# a_1290_n633# 0.09fF
C570 a_1500_n633# a_1172_n633# 0.02fF
C571 a_1080_n633# w_n4520_n852# 0.01fF
C572 a_n3120_n633# a_n4078_n633# 0.01fF
C573 a_238_n100# a_n1232_n100# 0.00fF
C574 a_n1230_n633# a_n2490_n633# 0.00fF
C575 a_n182_n100# a_n812_n100# 0.01fF
C576 a_n1978_n633# a_n3448_n633# 0.00fF
C577 a_n2280_n633# a_n3120_n633# 0.01fF
C578 a_n2490_n633# a_n2910_n633# 0.02fF
C579 a_n2188_n633# a_n3238_n633# 0.01fF
C580 a_n300_n100# a_n720_n100# 0.02fF
C581 a_n90_n100# a_n930_n100# 0.01fF
C582 a_n2398_n633# a_n3028_n633# 0.01fF
C583 a_n392_n100# a_n602_n100# 0.03fF
C584 a_1964_n730# w_n4520_n852# 0.12fF
C585 a_n3332_n100# a_n3752_n100# 0.02fF
C586 a_n2702_n100# a_n2820_n100# 0.07fF
C587 a_2850_n100# a_1708_n100# 0.01fF
C588 a_2758_n100# a_1800_n100# 0.01fF
C589 a_914_n401# a_912_131# 0.01fF
C590 a_2384_n730# a_914_n401# 0.00fF
C591 a_2340_n633# a_1592_n633# 0.01fF
C592 a_2432_n633# a_1500_n633# 0.01fF
C593 a_n3750_n633# a_n3708_131# 0.00fF
C594 a_3900_n100# a_3178_n100# 0.01fF
C595 a_n2658_n197# a_n3078_n197# 0.01fF
C596 a_1382_n633# a_1172_n633# 0.03fF
C597 a_n2238_n197# a_n3498_n197# 0.00fF
C598 a_n3238_n633# a_n4078_n633# 0.01fF
C599 a_n3330_n633# a_n3960_n633# 0.01fF
C600 a_n3448_n633# a_n3450_n100# 0.00fF
C601 a_n1770_n100# a_n2400_n100# 0.01fF
C602 a_n2398_n633# a_n3120_n633# 0.01fF
C603 a_n182_n100# a_n930_n100# 0.01fF
C604 a_n2280_n633# a_n3238_n633# 0.01fF
C605 a_n300_n100# a_n812_n100# 0.01fF
C606 a_n2490_n633# a_n3028_n633# 0.01fF
C607 a_n510_n100# a_n602_n100# 0.09fF
C608 a_n392_n100# a_n720_n100# 0.02fF
C609 a_3482_n633# a_3180_n633# 0.02fF
C610 a_1544_n730# w_n4520_n852# 0.12fF
C611 a_1290_n633# a_1332_131# 0.00fF
C612 a_494_n401# a_492_131# 0.01fF
C613 a_n3450_n100# a_n3752_n100# 0.02fF
C614 a_n2702_n100# a_n2912_n100# 0.03fF
C615 a_4018_n100# a_2850_n100# 0.01fF
C616 a_n1816_n730# a_n3076_n730# 0.00fF
C617 a_2640_n100# a_1800_n100# 0.01fF
C618 a_2758_n100# a_1708_n100# 0.01fF
C619 a_1964_n730# a_914_n401# 0.00fF
C620 a_2802_n197# w_n4520_n852# 0.10fF
C621 a_2340_n633# a_1500_n633# 0.01fF
C622 a_2432_n633# a_1382_n633# 0.01fF
C623 a_2222_n633# w_n4520_n852# 0.01fF
C624 a_3060_n100# a_2850_n100# 0.03fF
C625 a_n768_131# a_n1608_131# 0.01fF
C626 a_3808_n100# a_3178_n100# 0.01fF
C627 a_n2658_n197# a_n3498_n197# 0.01fF
C628 a_1288_n100# a_120_n100# 0.01fF
C629 a_1290_n633# a_1172_n633# 0.07fF
C630 a_n3448_n633# a_n3960_n633# 0.01fF
C631 a_n1862_n100# a_n2400_n100# 0.01fF
C632 a_1498_n100# a_1170_n100# 0.02fF
C633 a_494_n401# a_540_n100# 0.00fF
C634 a_2382_n197# a_3012_131# 0.00fF
C635 a_n2398_n633# a_n3238_n633# 0.01fF
C636 a_n300_n100# a_n930_n100# 0.01fF
C637 a_1288_n100# a_1800_n100# 0.01fF
C638 a_n510_n100# a_n720_n100# 0.03fF
C639 a_n392_n100# a_n812_n100# 0.02fF
C640 a_n2490_n633# a_n3120_n633# 0.01fF
C641 a_3390_n633# a_3180_n633# 0.03fF
C642 a_n3542_n100# a_n3752_n100# 0.03fF
C643 a_n2820_n100# a_n2912_n100# 0.09fF
C644 a_n2702_n100# a_n3030_n100# 0.02fF
C645 a_4018_n100# a_2758_n100# 0.00fF
C646 a_n2236_n730# a_n3076_n730# 0.01fF
C647 a_2640_n100# a_1708_n100# 0.01fF
C648 a_2548_n100# a_1800_n100# 0.01fF
C649 a_1544_n730# a_914_n401# 0.00fF
C650 a_3222_n197# a_3012_131# 0.01fF
C651 a_2432_n633# a_1290_n633# 0.01fF
C652 a_2340_n633# a_1382_n633# 0.01fF
C653 a_2130_n633# w_n4520_n852# 0.01fF
C654 a_n3496_n730# a_n2026_n401# 0.00fF
C655 a_3062_n633# a_3060_n100# 0.00fF
C656 a_n346_n401# a_n348_131# 0.01fF
C657 a_3060_n100# a_2758_n100# 0.02fF
C658 a_2968_n100# a_1498_n100# 0.00fF
C659 a_n508_n633# a_n1348_n633# 0.01fF
C660 a_n1188_131# a_n1608_131# 0.01fF
C661 a_n3078_n197# a_n3498_n197# 0.01fF
C662 a_n2658_n197# a_n3918_n197# 0.00fF
C663 a_4110_n100# a_3270_n100# 0.01fF
C664 a_n2448_131# a_n2868_131# 0.01fF
C665 a_4112_n633# a_4020_n633# 0.09fF
C666 a_1962_n197# a_3012_131# 0.00fF
C667 a_1288_n100# a_1708_n100# 0.02fF
C668 a_n602_n100# a_n720_n100# 0.07fF
C669 a_n510_n100# a_n812_n100# 0.02fF
C670 a_n2490_n633# a_n3238_n633# 0.01fF
C671 a_n392_n100# a_n930_n100# 0.01fF
C672 a_1122_n197# a_702_n197# 0.01fF
C673 a_1542_n197# a_282_n197# 0.00fF
C674 a_2382_n197# a_1332_131# 0.00fF
C675 a_n3660_n100# a_n3752_n100# 0.09fF
C676 a_n2820_n100# a_n3030_n100# 0.03fF
C677 a_n2702_n100# a_n3122_n100# 0.02fF
C678 a_4018_n100# a_2640_n100# 0.00fF
C679 a_n2656_n730# a_n3076_n730# 0.01fF
C680 a_2548_n100# a_1708_n100# 0.01fF
C681 a_2430_n100# a_1800_n100# 0.01fF
C682 a_2340_n633# a_1290_n633# 0.01fF
C683 a_2550_n633# a_1080_n633# 0.00fF
C684 a_2432_n633# a_1172_n633# 0.00fF
C685 a_n3496_n730# a_n2446_n401# 0.00fF
C686 a_2012_n633# w_n4520_n852# 0.01fF
C687 a_3060_n100# a_2640_n100# 0.02fF
C688 a_n600_n633# a_n1348_n633# 0.01fF
C689 a_n3078_n197# a_n3918_n197# 0.01fF
C690 a_n3750_n633# a_n4170_n633# 0.02fF
C691 a_n2070_n633# a_n3658_n633# 0.00fF
C692 a_n4080_n100# a_n4172_n100# 0.09fF
C693 a_1592_n633# a_542_n633# 0.01fF
C694 a_238_n100# a_n1350_n100# 0.00fF
C695 a_n2448_131# a_n3288_131# 0.01fF
C696 a_4112_n633# a_3902_n633# 0.03fF
C697 a_n602_n100# a_n812_n100# 0.03fF
C698 a_n510_n100# a_n930_n100# 0.02fF
C699 a_n2070_n633# a_n3540_n633# 0.00fF
C700 a_n3962_n100# a_n4172_n100# 0.03fF
C701 a_n3916_n730# w_n4520_n852# 0.13fF
C702 a_n2070_n633# w_n4520_n852# 0.01fF
C703 a_1962_n197# a_1332_131# 0.00fF
C704 a_n2702_n100# a_n3240_n100# 0.01fF
C705 a_n2820_n100# a_n3122_n100# 0.02fF
C706 a_n2912_n100# a_n3030_n100# 0.07fF
C707 a_4018_n100# a_2548_n100# 0.00fF
C708 a_2430_n100# a_1708_n100# 0.01fF
C709 a_2338_n100# a_1800_n100# 0.01fF
C710 a_2174_n401# a_2172_131# 0.01fF
C711 a_2340_n633# a_1172_n633# 0.01fF
C712 a_1920_n633# w_n4520_n852# 0.01fF
C713 a_n3496_n730# a_n2866_n401# 0.00fF
C714 a_3060_n100# a_2548_n100# 0.01fF
C715 a_868_n100# a_120_n100# 0.01fF
C716 a_n718_n633# a_n1348_n633# 0.01fF
C717 a_n3498_n197# a_n3918_n197# 0.01fF
C718 a_n2188_n633# a_n3658_n633# 0.00fF
C719 a_702_n197# a_912_131# 0.01fF
C720 a_1592_n633# a_450_n633# 0.01fF
C721 a_1500_n633# a_542_n633# 0.01fF
C722 a_1800_n100# a_868_n100# 0.01fF
C723 a_4112_n633# a_3810_n633# 0.02fF
C724 a_4020_n633# a_3902_n633# 0.07fF
C725 a_n602_n100# a_n930_n100# 0.02fF
C726 a_n720_n100# a_n812_n100# 0.09fF
C727 a_n2188_n633# a_n3540_n633# 0.00fF
C728 a_962_n633# a_122_n633# 0.01fF
C729 a_1754_n401# a_1752_131# 0.01fF
C730 a_n2188_n633# w_n4520_n852# 0.01fF
C731 a_n2702_n100# a_n3332_n100# 0.01fF
C732 a_n2820_n100# a_n3240_n100# 0.02fF
C733 a_n2912_n100# a_n3122_n100# 0.03fF
C734 a_4018_n100# a_2430_n100# 0.00fF
C735 a_2338_n100# a_1708_n100# 0.01fF
C736 a_2220_n100# a_1800_n100# 0.02fF
C737 a_2432_n633# a_2340_n633# 0.09fF
C738 a_2550_n633# a_2222_n633# 0.02fF
C739 a_n558_n197# a_n348_131# 0.01fF
C740 a_n3658_n633# a_n4078_n633# 0.02fF
C741 a_1802_n633# w_n4520_n852# 0.01fF
C742 a_3060_n100# a_2430_n100# 0.01fF
C743 a_750_n100# a_120_n100# 0.01fF
C744 a_3014_n401# a_2174_n401# 0.01fF
C745 a_n810_n633# a_n1348_n633# 0.01fF
C746 a_n2280_n633# a_n3658_n633# 0.00fF
C747 a_3222_n197# a_2382_n197# 0.01fF
C748 a_332_n633# w_n4520_n852# 0.01fF
C749 a_1500_n633# a_450_n633# 0.01fF
C750 a_1382_n633# a_542_n633# 0.01fF
C751 a_n3540_n633# a_n4078_n633# 0.01fF
C752 a_2340_n633# a_2382_n197# 0.00fF
C753 a_1708_n100# a_868_n100# 0.01fF
C754 a_1800_n100# a_750_n100# 0.01fF
C755 a_4020_n633# a_3810_n633# 0.03fF
C756 a_4112_n633# a_3692_n633# 0.02fF
C757 a_n720_n100# a_n930_n100# 0.03fF
C758 a_n4078_n633# w_n4520_n852# 0.08fF
C759 a_n1440_n633# a_n1396_n730# 0.00fF
C760 a_n2280_n633# a_n3540_n633# 0.00fF
C761 a_3272_n633# a_3062_n633# 0.03fF
C762 a_n558_n197# a_492_131# 0.00fF
C763 a_n1396_n730# a_n1350_n100# 0.00fF
C764 a_962_n633# a_30_n633# 0.01fF
C765 a_2382_n197# a_1962_n197# 0.01fF
C766 a_n2280_n633# w_n4520_n852# 0.01fF
C767 a_1170_n100# a_960_n100# 0.03fF
C768 a_n2820_n100# a_n3332_n100# 0.01fF
C769 a_n2912_n100# a_n3240_n100# 0.02fF
C770 a_n2702_n100# a_n3450_n100# 0.01fF
C771 a_n3030_n100# a_n3122_n100# 0.09fF
C772 a_3642_n197# a_2802_n197# 0.01fF
C773 a_2550_n633# a_2130_n633# 0.02fF
C774 a_2128_n100# a_1800_n100# 0.02fF
C775 a_2220_n100# a_1708_n100# 0.01fF
C776 a_1710_n633# w_n4520_n852# 0.01fF
C777 a_3060_n100# a_2338_n100# 0.01fF
C778 a_2594_n401# a_2174_n401# 0.01fF
C779 a_n928_n633# a_n1348_n633# 0.02fF
C780 a_3014_n401# a_1754_n401# 0.00fF
C781 a_n1232_n100# a_n2072_n100# 0.01fF
C782 a_n2398_n633# a_n3658_n633# 0.00fF
C783 a_3690_n100# a_2968_n100# 0.01fF
C784 a_1290_n633# a_542_n633# 0.01fF
C785 a_1382_n633# a_450_n633# 0.01fF
C786 a_n2282_n100# a_n3870_n100# 0.00fF
C787 a_n4080_n100# a_n4128_131# 0.00fF
C788 a_3222_n197# a_1962_n197# 0.00fF
C789 a_240_n633# w_n4520_n852# 0.01fF
C790 a_1124_n730# a_1170_n100# 0.00fF
C791 a_1708_n100# a_750_n100# 0.01fF
C792 a_3902_n633# a_3810_n633# 0.09fF
C793 a_4020_n633# a_3692_n633# 0.02fF
C794 a_330_n100# a_120_n100# 0.03fF
C795 a_n812_n100# a_n930_n100# 0.07fF
C796 a_n2398_n633# a_n3540_n633# 0.01fF
C797 a_n718_n633# a_n766_n401# 0.00fF
C798 a_1800_n100# a_330_n100# 0.00fF
C799 a_n2398_n633# w_n4520_n852# 0.01fF
C800 a_n2702_n100# a_n3542_n100# 0.01fF
C801 a_284_n730# a_282_n197# 0.01fF
C802 a_n2912_n100# a_n3332_n100# 0.02fF
C803 a_n3030_n100# a_n3240_n100# 0.03fF
C804 a_n2820_n100# a_n3450_n100# 0.01fF
C805 a_n508_n633# a_n1768_n633# 0.00fF
C806 a_2128_n100# a_1708_n100# 0.02fF
C807 a_2550_n633# a_2012_n633# 0.01fF
C808 a_2010_n100# a_1800_n100# 0.03fF
C809 a_3644_n730# a_2174_n401# 0.00fF
C810 a_3060_n100# a_2220_n100# 0.01fF
C811 a_n1020_n633# a_n1348_n633# 0.02fF
C812 a_2594_n401# a_1754_n401# 0.01fF
C813 a_n2490_n633# a_n3658_n633# 0.01fF
C814 a_1172_n633# a_542_n633# 0.01fF
C815 a_1080_n633# a_660_n633# 0.02fF
C816 a_1290_n633# a_450_n633# 0.01fF
C817 a_3902_n633# a_3692_n633# 0.03fF
C818 a_n600_n633# a_n558_n197# 0.00fF
C819 a_238_n100# a_120_n100# 0.07fF
C820 a_752_n633# a_n508_n633# 0.00fF
C821 a_n2490_n633# a_n3540_n633# 0.01fF
C822 a_n810_n633# a_n766_n401# 0.00fF
C823 a_n2492_n100# a_n4080_n100# 0.00fF
C824 a_n2490_n633# w_n4520_n852# 0.01fF
C825 a_1708_n100# a_330_n100# 0.00fF
C826 a_1800_n100# a_238_n100# 0.00fF
C827 a_n3030_n100# a_n3332_n100# 0.02fF
C828 a_n2912_n100# a_n3450_n100# 0.01fF
C829 a_n2702_n100# a_n3660_n100# 0.01fF
C830 a_n2820_n100# a_n3542_n100# 0.01fF
C831 a_n3122_n100# a_n3240_n100# 0.07fF
C832 a_n2492_n100# a_n3962_n100# 0.00fF
C833 a_2010_n100# a_1708_n100# 0.02fF
C834 a_1918_n100# a_1800_n100# 0.07fF
C835 a_n600_n633# a_n1768_n633# 0.01fF
C836 a_2550_n633# a_1920_n633# 0.01fF
C837 a_3180_n633# w_n4520_n852# 0.03fF
C838 a_1170_n100# a_448_n100# 0.01fF
C839 a_3060_n100# a_2128_n100# 0.01fF
C840 a_1498_n100# w_n4520_n852# 0.02fF
C841 a_1172_n633# a_450_n633# 0.01fF
C842 a_3810_n633# a_3692_n633# 0.07fF
C843 a_752_n633# a_n600_n633# 0.00fF
C844 a_4064_n730# a_4110_n100# 0.00fF
C845 a_1708_n100# a_238_n100# 0.00fF
C846 a_n3448_n633# a_n3496_n730# 0.00fF
C847 a_n3122_n100# a_n3332_n100# 0.03fF
C848 a_n2912_n100# a_n3542_n100# 0.01fF
C849 a_n2820_n100# a_n3660_n100# 0.01fF
C850 a_n720_n100# a_n768_131# 0.00fF
C851 a_n3030_n100# a_n3450_n100# 0.02fF
C852 a_1380_n100# a_28_n100# 0.00fF
C853 a_n718_n633# a_n1768_n633# 0.01fF
C854 a_2550_n633# a_1802_n633# 0.01fF
C855 a_1918_n100# a_1708_n100# 0.03fF
C856 a_122_n633# a_n1348_n633# 0.00fF
C857 a_3060_n100# a_2010_n100# 0.01fF
C858 a_n3496_n730# a_n4126_n401# 0.00fF
C859 a_2222_n633# a_660_n633# 0.00fF
C860 a_1078_n100# a_28_n100# 0.01fF
C861 a_4110_n100# a_3900_n100# 0.03fF
C862 a_282_n197# a_72_131# 0.01fF
C863 a_122_n633# a_74_n401# 0.00fF
C864 a_752_n633# a_n718_n633# 0.00fF
C865 a_n3240_n100# a_n3332_n100# 0.09fF
C866 a_n3030_n100# a_n3542_n100# 0.01fF
C867 a_n2912_n100# a_n3660_n100# 0.01fF
C868 a_n3122_n100# a_n3450_n100# 0.02fF
C869 a_n812_n100# a_n768_131# 0.00fF
C870 a_n1442_n100# a_n2072_n100# 0.01fF
C871 a_1380_n100# a_n90_n100# 0.00fF
C872 a_n810_n633# a_n1768_n633# 0.01fF
C873 a_2550_n633# a_1710_n633# 0.01fF
C874 a_540_n100# a_n1022_n100# 0.00fF
C875 a_30_n633# a_n1348_n633# 0.00fF
C876 a_3178_n100# a_1800_n100# 0.00fF
C877 a_3060_n100# a_1918_n100# 0.01fF
C878 a_2130_n633# a_660_n633# 0.00fF
C879 a_n1350_n100# a_n2072_n100# 0.01fF
C880 a_1078_n100# a_n90_n100# 0.01fF
C881 a_4110_n100# a_3808_n100# 0.02fF
C882 a_30_n633# a_74_n401# 0.00fF
C883 a_752_n633# a_n810_n633# 0.00fF
C884 a_448_n100# a_n1140_n100# 0.00fF
C885 a_n3030_n100# a_n3660_n100# 0.01fF
C886 a_n3240_n100# a_n3450_n100# 0.03fF
C887 a_n3122_n100# a_n3542_n100# 0.02fF
C888 a_1170_n100# a_658_n100# 0.01fF
C889 a_1542_n197# w_n4520_n852# 0.10fF
C890 a_1380_n100# a_n182_n100# 0.00fF
C891 a_n1138_n633# a_n1558_n633# 0.02fF
C892 a_n928_n633# a_n1768_n633# 0.01fF
C893 a_2970_n633# a_2852_n633# 0.07fF
C894 a_3178_n100# a_1708_n100# 0.00fF
C895 a_2012_n633# a_660_n633# 0.00fF
C896 a_1078_n100# a_n182_n100# 0.00fF
C897 a_n1652_n100# a_n2282_n100# 0.01fF
C898 a_n1860_n633# a_n2070_n633# 0.03fF
C899 a_3852_131# a_3012_131# 0.01fF
C900 a_3224_n730# w_n4520_n852# 0.12fF
C901 a_n3122_n100# a_n3660_n100# 0.01fF
C902 a_n3332_n100# a_n3450_n100# 0.07fF
C903 a_n3240_n100# a_n3542_n100# 0.02fF
C904 a_n1020_n633# a_n1768_n633# 0.01fF
C905 a_n1138_n633# a_n1650_n633# 0.01fF
C906 a_2970_n633# a_2760_n633# 0.03fF
C907 a_3180_n633# a_2550_n633# 0.01fF
C908 a_3062_n633# a_2642_n633# 0.02fF
C909 a_4018_n100# a_3178_n100# 0.01fF
C910 a_1920_n633# a_660_n633# 0.00fF
C911 a_1078_n100# a_n300_n100# 0.00fF
C912 a_n1860_n633# a_n2188_n633# 0.02fF
C913 a_3690_n100# w_n4520_n852# 0.04fF
C914 a_3432_131# a_3012_131# 0.01fF
C915 a_n1138_n633# a_n2608_n633# 0.00fF
C916 a_3178_n100# a_3060_n100# 0.07fF
C917 a_3270_n100# a_2968_n100# 0.02fF
C918 a_960_n100# w_n4520_n852# 0.02fF
C919 a_n3332_n100# a_n3542_n100# 0.03fF
C920 a_n3240_n100# a_n3660_n100# 0.02fF
C921 a_n3868_n633# a_n3916_n730# 0.00fF
C922 a_n348_131# a_n1608_131# 0.00fF
C923 a_2642_n633# a_2640_n100# 0.00fF
C924 a_1124_n730# w_n4520_n852# 0.12fF
C925 a_1802_n633# a_660_n633# 0.01fF
C926 a_1078_n100# a_n392_n100# 0.00fF
C927 a_n1860_n633# a_n2280_n633# 0.02fF
C928 a_1382_n633# a_1380_n100# 0.00fF
C929 a_n1138_n633# a_n2700_n633# 0.00fF
C930 a_660_n633# a_332_n633# 0.02fF
C931 a_542_n633# a_450_n633# 0.09fF
C932 a_n3450_n100# a_n3542_n100# 0.09fF
C933 a_n3332_n100# a_n3660_n100# 0.02fF
C934 a_n88_n633# a_n1558_n633# 0.00fF
C935 a_n3916_n730# a_n3286_n401# 0.00fF
C936 a_n2282_n100# a_n2610_n100# 0.02fF
C937 a_282_n197# a_1752_131# 0.00fF
C938 a_914_n401# a_960_n100# 0.00fF
C939 a_704_n730# w_n4520_n852# 0.12fF
C940 a_n1232_n100# a_n1560_n100# 0.02fF
C941 a_1710_n633# a_660_n633# 0.01fF
C942 a_1078_n100# a_n510_n100# 0.00fF
C943 a_n1860_n633# a_n2398_n633# 0.01fF
C944 a_660_n633# a_240_n633# 0.02fF
C945 a_752_n633# a_122_n633# 0.01fF
C946 a_2382_n197# a_3852_131# 0.00fF
C947 a_1124_n730# a_914_n401# 0.01fF
C948 a_1380_n100# a_1332_131# 0.00fF
C949 a_n3868_n633# a_n4078_n633# 0.03fF
C950 a_n3450_n100# a_n3660_n100# 0.03fF
C951 a_n180_n633# a_n1558_n633# 0.00fF
C952 a_n88_n633# a_n1650_n633# 0.00fF
C953 a_n3916_n730# a_n3706_n401# 0.01fF
C954 a_448_n100# w_n4520_n852# 0.02fF
C955 a_540_n100# a_28_n100# 0.01fF
C956 a_n2280_n633# a_n3868_n633# 0.00fF
C957 a_3222_n197# a_3852_131# 0.00fF
C958 a_284_n730# w_n4520_n852# 0.12fF
C959 a_n1020_n633# a_n1022_n100# 0.00fF
C960 a_n768_131# a_n1188_131# 0.01fF
C961 a_n1138_n633# a_n1230_n633# 0.09fF
C962 a_n1860_n633# a_n2490_n633# 0.01fF
C963 a_2640_n100# a_2592_131# 0.00fF
C964 a_n1232_n100# a_n2190_n100# 0.01fF
C965 a_752_n633# a_30_n633# 0.01fF
C966 a_1590_n100# a_1170_n100# 0.02fF
C967 a_870_n633# a_n88_n633# 0.01fF
C968 a_2382_n197# a_3432_131# 0.00fF
C969 a_704_n730# a_914_n401# 0.01fF
C970 a_n1022_n100# a_n2282_n100# 0.00fF
C971 a_n2280_n633# a_n2238_n197# 0.00fF
C972 a_n3542_n100# a_n3660_n100# 0.07fF
C973 a_n298_n633# a_n1558_n633# 0.00fF
C974 a_n180_n633# a_n1650_n633# 0.00fF
C975 a_540_n100# a_n90_n100# 0.01fF
C976 a_n2398_n633# a_n3868_n633# 0.00fF
C977 a_3222_n197# a_3432_131# 0.01fF
C978 a_n136_n730# w_n4520_n852# 0.12fF
C979 a_2968_n100# a_1590_n100# 0.00fF
C980 a_3600_n633# a_2432_n633# 0.01fF
C981 a_2548_n100# a_2592_131# 0.00fF
C982 a_3810_n633# a_2222_n633# 0.00fF
C983 a_870_n633# a_n180_n633# 0.01fF
C984 a_n2028_131# a_n2868_131# 0.01fF
C985 a_1962_n197# a_3432_131# 0.00fF
C986 a_284_n730# a_914_n401# 0.00fF
C987 a_1542_n197# a_702_n197# 0.01fF
C988 a_n300_n100# a_n348_131# 0.00fF
C989 a_n298_n633# a_n1650_n633# 0.00fF
C990 a_n390_n633# a_n1558_n633# 0.01fF
C991 a_n1232_n100# a_n2492_n100# 0.00fF
C992 a_540_n100# a_n182_n100# 0.01fF
C993 a_n2490_n633# a_n3868_n633# 0.00fF
C994 a_3690_n100# a_3642_n197# 0.00fF
C995 a_n556_n730# w_n4520_n852# 0.12fF
C996 a_3600_n633# a_2340_n633# 0.00fF
C997 a_3692_n633# a_2222_n633# 0.00fF
C998 a_870_n633# a_n298_n633# 0.01fF
C999 a_n2028_131# a_n3288_131# 0.00fF
C1000 a_n4080_n100# w_n4520_n852# 0.08fF
C1001 a_n136_n730# a_914_n401# 0.00fF
C1002 a_658_n100# w_n4520_n852# 0.02fF
C1003 a_1754_n401# a_1800_n100# 0.00fF
C1004 a_72_131# w_n4520_n852# 0.12fF
C1005 a_n392_n100# a_n348_131# 0.00fF
C1006 a_n3752_n100# a_n3708_131# 0.00fF
C1007 a_n3916_n730# a_n3918_n197# 0.01fF
C1008 a_n390_n633# a_n1650_n633# 0.00fF
C1009 a_n1442_n100# a_n1560_n100# 0.07fF
C1010 a_n3962_n100# w_n4520_n852# 0.06fF
C1011 a_n3028_n633# a_n3076_n730# 0.00fF
C1012 a_540_n100# a_n300_n100# 0.01fF
C1013 a_n88_n633# a_n1230_n633# 0.01fF
C1014 a_n1350_n100# a_n1560_n100# 0.03fF
C1015 a_3692_n633# a_2130_n633# 0.00fF
C1016 a_n1440_n633# a_n1558_n633# 0.07fF
C1017 a_1122_n197# a_912_131# 0.01fF
C1018 a_3270_n100# w_n4520_n852# 0.03fF
C1019 a_870_n633# a_n390_n633# 0.00fF
C1020 a_n556_n730# a_914_n401# 0.00fF
C1021 a_n1230_n633# a_n1232_n100# 0.00fF
C1022 a_1080_n633# a_1122_n197# 0.00fF
C1023 a_n3120_n633# a_n3076_n730# 0.00fF
C1024 a_2804_n730# a_2384_n730# 0.01fF
C1025 a_540_n100# a_n392_n100# 0.01fF
C1026 a_n1442_n100# a_n2190_n100# 0.01fF
C1027 a_n180_n633# a_n1230_n633# 0.01fF
C1028 a_n1138_n633# a_n1140_n100# 0.00fF
C1029 a_3900_n100# a_2968_n100# 0.01fF
C1030 a_n976_n730# a_494_n401# 0.00fF
C1031 a_n1440_n633# a_n1650_n633# 0.03fF
C1032 a_n1350_n100# a_n2190_n100# 0.01fF
C1033 a_n3330_n633# a_n4170_n633# 0.01fF
C1034 a_3482_n633# a_2970_n633# 0.01fF
C1035 a_n1440_n633# a_n2608_n633# 0.01fF
C1036 a_704_n730# a_702_n197# 0.01fF
C1037 a_540_n100# a_n510_n100# 0.01fF
C1038 a_2804_n730# a_1964_n730# 0.01fF
C1039 a_1332_131# a_492_131# 0.01fF
C1040 a_n298_n633# a_n1230_n633# 0.01fF
C1041 a_n508_n633# a_n510_n100# 0.00fF
C1042 a_n1232_n100# a_n1980_n100# 0.01fF
C1043 a_n976_n730# a_74_n401# 0.00fF
C1044 a_4112_n633# a_3180_n633# 0.01fF
C1045 a_n2282_n100# a_n3752_n100# 0.00fF
C1046 a_3808_n100# a_2968_n100# 0.01fF
C1047 a_n3448_n633# a_n4170_n633# 0.01fF
C1048 a_n2492_n100# a_n2448_131# 0.00fF
C1049 a_3390_n633# a_2970_n633# 0.02fF
C1050 a_n1440_n633# a_n2700_n633# 0.00fF
C1051 a_n1442_n100# a_n2492_n100# 0.01fF
C1052 a_n4170_n633# a_n4126_n401# 0.00fF
C1053 a_n1348_n633# a_n1396_n730# 0.00fF
C1054 a_n1350_n100# a_n2492_n100# 0.01fF
C1055 a_2804_n730# a_1544_n730# 0.00fF
C1056 a_2384_n730# a_1964_n730# 0.01fF
C1057 a_540_n100# a_n602_n100# 0.01fF
C1058 a_n390_n633# a_n1230_n633# 0.01fF
C1059 a_4110_n100# a_4018_n100# 0.09fF
C1060 a_2970_n633# a_2968_n100# 0.00fF
C1061 a_4020_n633# a_3180_n633# 0.01fF
C1062 a_n1396_n730# a_74_n401# 0.00fF
C1063 a_n976_n730# a_n346_n401# 0.00fF
C1064 a_n3496_n730# a_n3450_n100# 0.00fF
C1065 a_4110_n100# a_3060_n100# 0.01fF
C1066 a_2804_n730# a_2802_n197# 0.01fF
C1067 a_n1440_n633# a_n2818_n633# 0.00fF
C1068 a_752_n633# a_750_n100# 0.00fF
C1069 a_2384_n730# a_1544_n730# 0.01fF
C1070 a_540_n100# a_n720_n100# 0.00fF
C1071 a_n600_n633# a_n602_n100# 0.00fF
C1072 a_1590_n100# w_n4520_n852# 0.02fF
C1073 a_660_n633# a_704_n730# 0.00fF
C1074 a_n976_n730# a_n766_n401# 0.01fF
C1075 a_n1396_n730# a_n346_n401# 0.00fF
C1076 a_3902_n633# a_3180_n633# 0.01fF
C1077 a_1752_131# w_n4520_n852# 0.12fF
C1078 a_n1230_n633# a_n1440_n633# 0.03fF
C1079 a_2172_131# w_n4520_n852# 0.12fF
C1080 a_n1140_n100# a_n1232_n100# 0.09fF
C1081 a_n1440_n633# a_n2910_n633# 0.00fF
C1082 a_1962_n197# a_492_131# 0.00fF
C1083 a_1964_n730# a_1544_n730# 0.01fF
C1084 a_540_n100# a_n812_n100# 0.00fF
C1085 a_30_n633# a_28_n100# 0.00fF
C1086 a_2222_n633# a_1080_n633# 0.01fF
C1087 a_n1816_n730# a_n346_n401# 0.00fF
C1088 a_n1396_n730# a_n766_n401# 0.00fF
C1089 a_3810_n633# a_3180_n633# 0.01fF
C1090 a_n976_n730# a_n1186_n401# 0.01fF
C1091 a_658_n100# a_702_n197# 0.00fF
C1092 a_702_n197# a_72_131# 0.00fF
C1093 a_n1138_n633# w_n4520_n852# 0.01fF
C1094 a_n1440_n633# a_n3028_n633# 0.00fF
C1095 a_n2398_n633# a_n2400_n100# 0.00fF
C1096 a_n2072_n100# a_n2028_131# 0.00fF
C1097 a_3014_n401# w_n4520_n852# 0.10fF
C1098 a_n1442_n100# a_n1980_n100# 0.01fF
C1099 a_540_n100# a_n930_n100# 0.00fF
C1100 a_n718_n633# a_n720_n100# 0.00fF
C1101 a_2130_n633# a_1080_n633# 0.01fF
C1102 a_n1350_n100# a_n1980_n100# 0.01fF
C1103 a_n976_n730# a_n1606_n401# 0.00fF
C1104 a_3692_n633# a_3180_n633# 0.01fF
C1105 a_n1396_n730# a_n1186_n401# 0.01fF
C1106 a_n1816_n730# a_n766_n401# 0.00fF
C1107 a_1592_n633# a_122_n633# 0.00fF
C1108 a_4064_n730# w_n4520_n852# 0.11fF
C1109 a_3272_n633# a_2852_n633# 0.02fF
C1110 a_n978_n197# a_72_131# 0.00fF
C1111 a_2594_n401# w_n4520_n852# 0.10fF
C1112 a_2012_n633# a_1080_n633# 0.01fF
C1113 a_n3076_n730# w_n4520_n852# 0.12fF
C1114 a_3900_n100# w_n4520_n852# 0.06fF
C1115 a_n1816_n730# a_n1186_n401# 0.00fF
C1116 a_n2236_n730# a_n766_n401# 0.00fF
C1117 a_n976_n730# a_n2026_n401# 0.00fF
C1118 a_n1396_n730# a_n1606_n401# 0.01fF
C1119 a_3852_131# a_3432_131# 0.01fF
C1120 a_n2282_n100# a_n2702_n100# 0.02fF
C1121 a_1288_n100# a_28_n100# 0.00fF
C1122 a_1592_n633# a_30_n633# 0.00fF
C1123 a_1500_n633# a_122_n633# 0.00fF
C1124 a_2012_n633# a_1964_n730# 0.00fF
C1125 a_n2866_n401# a_n2868_131# 0.01fF
C1126 a_3644_n730# w_n4520_n852# 0.10fF
C1127 a_330_n100# a_n1022_n100# 0.00fF
C1128 a_3272_n633# a_2760_n633# 0.01fF
C1129 a_n1398_n197# a_72_131# 0.00fF
C1130 a_660_n633# a_658_n100# 0.00fF
C1131 a_n508_n633# a_n1978_n633# 0.00fF
C1132 a_2222_n633# a_2130_n633# 0.09fF
C1133 a_n348_131# a_n768_131# 0.01fF
C1134 a_n810_n633# a_n812_n100# 0.00fF
C1135 a_1920_n633# a_1080_n633# 0.01fF
C1136 a_3062_n633# a_1592_n633# 0.00fF
C1137 a_2174_n401# a_1334_n401# 0.01fF
C1138 a_3808_n100# w_n4520_n852# 0.05fF
C1139 a_n1396_n730# a_n2026_n401# 0.00fF
C1140 a_n2236_n730# a_n1186_n401# 0.00fF
C1141 a_n1816_n730# a_n1606_n401# 0.01fF
C1142 a_n976_n730# a_n2446_n401# 0.00fF
C1143 a_n2282_n100# a_n2820_n100# 0.01fF
C1144 a_n1140_n100# a_n1442_n100# 0.02fF
C1145 a_1288_n100# a_n90_n100# 0.00fF
C1146 a_1500_n633# a_30_n633# 0.00fF
C1147 a_1382_n633# a_122_n633# 0.00fF
C1148 a_n88_n633# w_n4520_n852# 0.01fF
C1149 a_542_n633# a_540_n100# 0.00fF
C1150 a_1920_n633# a_1964_n730# 0.00fF
C1151 a_238_n100# a_n1022_n100# 0.00fF
C1152 a_n1140_n100# a_n1350_n100# 0.03fF
C1153 a_542_n633# a_n508_n633# 0.01fF
C1154 a_n1768_n633# a_n1816_n730# 0.00fF
C1155 a_492_131# a_n768_131# 0.00fF
C1156 a_450_n633# a_492_131# 0.00fF
C1157 a_n1232_n100# w_n4520_n852# 0.02fF
C1158 a_n600_n633# a_n1978_n633# 0.00fF
C1159 a_n348_131# a_n1188_131# 0.01fF
C1160 a_2222_n633# a_2012_n633# 0.03fF
C1161 a_1802_n633# a_1080_n633# 0.01fF
C1162 a_3062_n633# a_1500_n633# 0.00fF
C1163 a_2970_n633# w_n4520_n852# 0.03fF
C1164 a_1754_n401# a_1334_n401# 0.01fF
C1165 a_n1816_n730# a_n2026_n401# 0.01fF
C1166 a_n2656_n730# a_n1186_n401# 0.00fF
C1167 a_n1396_n730# a_n2446_n401# 0.00fF
C1168 a_n2236_n730# a_n1606_n401# 0.00fF
C1169 a_n2282_n100# a_n2912_n100# 0.01fF
C1170 a_1288_n100# a_n182_n100# 0.00fF
C1171 a_n180_n633# w_n4520_n852# 0.01fF
C1172 a_1080_n633# a_332_n633# 0.01fF
C1173 a_1382_n633# a_30_n633# 0.00fF
C1174 a_1290_n633# a_122_n633# 0.01fF
C1175 a_3642_n197# a_2172_131# 0.00fF
C1176 a_542_n633# a_n600_n633# 0.01fF
C1177 a_450_n633# a_n508_n633# 0.01fF
C1178 a_n720_n100# a_n2282_n100# 0.00fF
C1179 a_1754_n401# a_494_n401# 0.00fF
C1180 a_n718_n633# a_n1978_n633# 0.00fF
C1181 a_702_n197# a_1752_131# 0.00fF
C1182 a_2222_n633# a_1920_n633# 0.02fF
C1183 a_2130_n633# a_2012_n633# 0.07fF
C1184 a_n928_n633# a_n930_n100# 0.00fF
C1185 a_1170_n100# a_120_n100# 0.01fF
C1186 a_1710_n633# a_1080_n633# 0.01fF
C1187 a_n2236_n730# a_n2026_n401# 0.01fF
C1188 a_n1396_n730# a_n2866_n401# 0.00fF
C1189 a_n1816_n730# a_n2446_n401# 0.00fF
C1190 a_868_n100# a_28_n100# 0.01fF
C1191 a_n2656_n730# a_n1606_n401# 0.00fF
C1192 a_n2282_n100# a_n3030_n100# 0.01fF
C1193 a_702_n197# a_2172_131# 0.00fF
C1194 a_1288_n100# a_n300_n100# 0.00fF
C1195 a_n298_n633# w_n4520_n852# 0.01fF
C1196 a_1172_n633# a_122_n633# 0.01fF
C1197 a_1290_n633# a_30_n633# 0.00fF
C1198 a_1080_n633# a_240_n633# 0.01fF
C1199 a_1800_n100# a_1170_n100# 0.01fF
C1200 a_3692_n633# a_3690_n100# 0.00fF
C1201 a_1380_n100# a_1078_n100# 0.02fF
C1202 a_450_n633# a_n600_n633# 0.01fF
C1203 a_542_n633# a_n718_n633# 0.00fF
C1204 a_n812_n100# a_n2282_n100# 0.00fF
C1205 a_2550_n633# a_2594_n401# 0.00fF
C1206 a_n1652_n100# a_n2072_n100# 0.02fF
C1207 a_n810_n633# a_n1978_n633# 0.01fF
C1208 a_2222_n633# a_1802_n633# 0.02fF
C1209 a_2130_n633# a_1920_n633# 0.03fF
C1210 a_2968_n100# a_1800_n100# 0.01fF
C1211 a_n1816_n730# a_n2866_n401# 0.00fF
C1212 a_868_n100# a_n90_n100# 0.01fF
C1213 a_n2656_n730# a_n2026_n401# 0.00fF
C1214 a_n2236_n730# a_n2446_n401# 0.01fF
C1215 a_750_n100# a_28_n100# 0.01fF
C1216 a_n2282_n100# a_n3122_n100# 0.01fF
C1217 a_n390_n633# w_n4520_n852# 0.01fF
C1218 a_1172_n633# a_30_n633# 0.01fF
C1219 a_1708_n100# a_1170_n100# 0.01fF
C1220 a_450_n633# a_n718_n633# 0.01fF
C1221 a_542_n633# a_n810_n633# 0.00fF
C1222 a_n930_n100# a_n2282_n100# 0.00fF
C1223 a_n2608_n633# a_n3750_n633# 0.01fF
C1224 a_n928_n633# a_n1978_n633# 0.01fF
C1225 a_2222_n633# a_1710_n633# 0.01fF
C1226 a_2012_n633# a_1920_n633# 0.09fF
C1227 a_2130_n633# a_1802_n633# 0.02fF
C1228 a_n3330_n633# a_n3288_131# 0.00fF
C1229 a_2968_n100# a_1708_n100# 0.00fF
C1230 a_n2656_n730# a_n2610_n100# 0.00fF
C1231 a_n2236_n730# a_n2866_n401# 0.00fF
C1232 a_868_n100# a_n182_n100# 0.01fF
C1233 a_n2656_n730# a_n2446_n401# 0.01fF
C1234 a_750_n100# a_n90_n100# 0.01fF
C1235 a_n2282_n100# a_n3240_n100# 0.01fF
C1236 a_n2448_131# w_n4520_n852# 0.12fF
C1237 a_3644_n730# a_3642_n197# 0.01fF
C1238 a_n1608_131# a_n2868_131# 0.00fF
C1239 a_n810_n633# a_n768_131# 0.00fF
C1240 a_n3870_n100# a_n4172_n100# 0.02fF
C1241 a_330_n100# a_28_n100# 0.02fF
C1242 a_542_n633# a_n928_n633# 0.00fF
C1243 a_1542_n197# a_1122_n197# 0.01fF
C1244 a_450_n633# a_n810_n633# 0.00fF
C1245 a_n1442_n100# w_n4520_n852# 0.02fF
C1246 a_120_n100# a_n1140_n100# 0.00fF
C1247 a_1288_n100# a_1290_n633# 0.00fF
C1248 a_962_n633# a_870_n633# 0.09fF
C1249 a_n1440_n633# w_n4520_n852# 0.01fF
C1250 a_282_n197# a_n138_n197# 0.01fF
C1251 a_n1350_n100# w_n4520_n852# 0.02fF
C1252 a_n2700_n633# a_n3750_n633# 0.01fF
C1253 a_n1020_n633# a_n1978_n633# 0.01fF
C1254 a_n1138_n633# a_n1860_n633# 0.01fF
C1255 a_2012_n633# a_1802_n633# 0.03fF
C1256 a_2130_n633# a_1710_n633# 0.02fF
C1257 a_1288_n100# a_1332_131# 0.00fF
C1258 a_2970_n633# a_2550_n633# 0.02fF
C1259 a_2852_n633# a_2642_n633# 0.03fF
C1260 a_3062_n633# a_2432_n633# 0.01fF
C1261 a_4018_n100# a_2968_n100# 0.01fF
C1262 a_750_n100# a_n182_n100# 0.01fF
C1263 a_n2656_n730# a_n2866_n401# 0.01fF
C1264 a_868_n100# a_n300_n100# 0.01fF
C1265 a_n2070_n633# a_n2188_n633# 0.07fF
C1266 a_n2282_n100# a_n3332_n100# 0.01fF
C1267 a_3060_n100# a_2968_n100# 0.09fF
C1268 a_450_n633# a_n928_n633# 0.00fF
C1269 a_542_n633# a_n1020_n633# 0.00fF
C1270 a_330_n100# a_n90_n100# 0.02fF
C1271 a_238_n100# a_28_n100# 0.03fF
C1272 a_n3660_n100# a_n3708_131# 0.00fF
C1273 a_n2072_n100# a_n2610_n100# 0.01fF
C1274 a_n2818_n633# a_n3750_n633# 0.01fF
C1275 a_n3962_n100# a_n3918_n197# 0.00fF
C1276 a_3224_n730# a_2804_n730# 0.01fF
C1277 a_2012_n633# a_1710_n633# 0.02fF
C1278 a_1920_n633# a_1802_n633# 0.07fF
C1279 a_3062_n633# a_2340_n633# 0.01fF
C1280 a_3180_n633# a_2222_n633# 0.01fF
C1281 a_2760_n633# a_2642_n633# 0.07fF
C1282 a_4110_n100# a_4062_n197# 0.00fF
C1283 a_868_n100# a_n392_n100# 0.00fF
C1284 a_1920_n633# a_332_n633# 0.00fF
C1285 a_750_n100# a_n300_n100# 0.01fF
C1286 a_n2282_n100# a_n3450_n100# 0.01fF
C1287 a_1542_n197# a_912_131# 0.00fF
C1288 a_n2070_n633# a_n2280_n633# 0.03fF
C1289 a_3480_n100# a_3432_131# 0.00fF
C1290 a_3600_n633# a_3598_n100# 0.00fF
C1291 a_330_n100# a_n182_n100# 0.01fF
C1292 a_238_n100# a_n90_n100# 0.02fF
C1293 a_450_n633# a_n1020_n633# 0.00fF
C1294 a_n2910_n633# a_n3750_n633# 0.01fF
C1295 a_1124_n730# a_1122_n197# 0.01fF
C1296 a_3224_n730# a_2384_n730# 0.01fF
C1297 a_1920_n633# a_1710_n633# 0.03fF
C1298 a_3180_n633# a_2130_n633# 0.01fF
C1299 a_n1232_n100# a_n1770_n100# 0.01fF
C1300 a_3482_n633# a_3272_n633# 0.03fF
C1301 a_1802_n633# a_332_n633# 0.00fF
C1302 a_868_n100# a_n510_n100# 0.00fF
C1303 a_750_n100# a_n392_n100# 0.01fF
C1304 a_n2282_n100# a_n3542_n100# 0.00fF
C1305 a_n2188_n633# a_n2280_n633# 0.09fF
C1306 a_n2070_n633# a_n2398_n633# 0.02fF
C1307 a_n1022_n100# a_n2072_n100# 0.01fF
C1308 a_3388_n100# a_3432_131# 0.00fF
C1309 a_542_n633# a_122_n633# 0.02fF
C1310 a_n1348_n633# a_n1558_n633# 0.03fF
C1311 a_330_n100# a_n300_n100# 0.01fF
C1312 a_238_n100# a_n182_n100# 0.02fF
C1313 a_n3028_n633# a_n3750_n633# 0.01fF
C1314 a_n3960_n633# a_n4170_n633# 0.03fF
C1315 a_3224_n730# a_1964_n730# 0.00fF
C1316 a_960_n100# a_912_131# 0.00fF
C1317 a_1802_n633# a_1710_n633# 0.09fF
C1318 a_3180_n633# a_2012_n633# 0.01fF
C1319 a_2432_n633# a_2430_n100# 0.00fF
C1320 a_n1232_n100# a_n1862_n100# 0.01fF
C1321 a_868_n100# a_n602_n100# 0.00fF
C1322 a_1802_n633# a_240_n633# 0.00fF
C1323 a_1710_n633# a_332_n633# 0.00fF
C1324 a_750_n100# a_n510_n100# 0.00fF
C1325 a_3390_n633# a_3272_n633# 0.07fF
C1326 a_n2070_n633# a_n2490_n633# 0.02fF
C1327 a_n2188_n633# a_n2398_n633# 0.03fF
C1328 a_n2282_n100# a_n3660_n100# 0.00fF
C1329 a_1544_n730# a_1542_n197# 0.01fF
C1330 a_1380_n100# a_540_n100# 0.01fF
C1331 a_2430_n100# a_2382_n197# 0.00fF
C1332 a_332_n633# a_240_n633# 0.09fF
C1333 a_660_n633# a_n88_n633# 0.01fF
C1334 a_542_n633# a_30_n633# 0.01fF
C1335 a_450_n633# a_122_n633# 0.02fF
C1336 a_n1348_n633# a_n1650_n633# 0.02fF
C1337 a_2384_n730# a_1124_n730# 0.00fF
C1338 a_238_n100# a_n300_n100# 0.01fF
C1339 a_330_n100# a_n392_n100# 0.01fF
C1340 a_1078_n100# a_540_n100# 0.01fF
C1341 a_2802_n197# a_1542_n197# 0.00fF
C1342 a_n2492_n100# a_n3870_n100# 0.00fF
C1343 a_n2400_n100# a_n3962_n100# 0.00fF
C1344 a_n3120_n633# a_n3750_n633# 0.01fF
C1345 a_n1348_n633# a_n2608_n633# 0.00fF
C1346 a_120_n100# w_n4520_n852# 0.02fF
C1347 a_3180_n633# a_1920_n633# 0.00fF
C1348 a_1080_n633# a_1124_n730# 0.00fF
C1349 a_1800_n100# w_n4520_n852# 0.02fF
C1350 a_750_n100# a_n602_n100# 0.00fF
C1351 a_1710_n633# a_240_n633# 0.00fF
C1352 a_868_n100# a_n720_n100# 0.00fF
C1353 a_n2188_n633# a_n2490_n633# 0.02fF
C1354 a_n2280_n633# a_n2398_n633# 0.07fF
C1355 a_n3076_n730# a_n3286_n401# 0.01fF
C1356 a_2338_n100# a_2382_n197# 0.00fF
C1357 a_450_n633# a_30_n633# 0.02fF
C1358 a_660_n633# a_n180_n633# 0.01fF
C1359 a_1964_n730# a_1124_n730# 0.01fF
C1360 a_238_n100# a_n392_n100# 0.01fF
C1361 a_330_n100# a_n510_n100# 0.01fF
C1362 a_n3238_n633# a_n3750_n633# 0.01fF
C1363 a_n298_n633# a_n1860_n633# 0.00fF
C1364 a_n1348_n633# a_n2700_n633# 0.00fF
C1365 a_3180_n633# a_1802_n633# 0.00fF
C1366 a_n2490_n633# a_n4078_n633# 0.00fF
C1367 a_2340_n633# a_2338_n100# 0.00fF
C1368 a_1708_n100# w_n4520_n852# 0.02fF
C1369 a_750_n100# a_n720_n100# 0.00fF
C1370 a_n2280_n633# a_n2490_n633# 0.03fF
C1371 a_n2656_n730# a_n4126_n401# 0.00fF
C1372 a_n3076_n730# a_n3706_n401# 0.00fF
C1373 a_660_n633# a_n298_n633# 0.01fF
C1374 a_1544_n730# a_1124_n730# 0.01fF
C1375 a_1964_n730# a_704_n730# 0.00fF
C1376 a_330_n100# a_n602_n100# 0.01fF
C1377 a_238_n100# a_n510_n100# 0.01fF
C1378 a_4112_n633# a_4064_n730# 0.00fF
C1379 a_n2820_n100# a_n2868_131# 0.00fF
C1380 a_3854_n401# a_3852_131# 0.01fF
C1381 a_n390_n633# a_n1860_n633# 0.00fF
C1382 a_n1442_n100# a_n1770_n100# 0.02fF
C1383 a_n1560_n100# a_n1652_n100# 0.09fF
C1384 a_n1348_n633# a_n2818_n633# 0.00fF
C1385 a_3180_n633# a_1710_n633# 0.00fF
C1386 a_4018_n100# w_n4520_n852# 0.08fF
C1387 a_n1350_n100# a_n1770_n100# 0.02fF
C1388 a_n3076_n730# a_n3078_n197# 0.01fF
C1389 a_750_n100# a_n812_n100# 0.00fF
C1390 a_n2398_n633# a_n2490_n633# 0.09fF
C1391 a_1122_n197# a_72_131# 0.00fF
C1392 a_3598_n100# a_3480_n100# 0.07fF
C1393 a_3060_n100# w_n4520_n852# 0.03fF
C1394 a_n978_n197# a_n2448_131# 0.00fF
C1395 a_660_n633# a_n390_n633# 0.01fF
C1396 a_1544_n730# a_704_n730# 0.01fF
C1397 a_238_n100# a_n602_n100# 0.01fF
C1398 a_330_n100# a_n720_n100# 0.01fF
C1399 a_n1980_n100# a_n2028_131# 0.00fF
C1400 a_4020_n633# a_4064_n730# 0.00fF
C1401 a_n2912_n100# a_n2868_131# 0.00fF
C1402 a_n1606_n401# a_n1560_n100# 0.00fF
C1403 a_n1230_n633# a_n1348_n633# 0.07fF
C1404 a_n1442_n100# a_n1862_n100# 0.02fF
C1405 a_n1348_n633# a_n2910_n633# 0.00fF
C1406 a_n1558_n633# a_n1606_n401# 0.00fF
C1407 a_n1652_n100# a_n2190_n100# 0.01fF
C1408 a_n1650_n633# a_n1652_n100# 0.00fF
C1409 a_n1350_n100# a_n1862_n100# 0.01fF
C1410 a_n2610_n100# a_n4172_n100# 0.00fF
C1411 a_n1558_n633# a_n1768_n633# 0.03fF
C1412 a_n1440_n633# a_n1860_n633# 0.02fF
C1413 a_3598_n100# a_3388_n100# 0.03fF
C1414 a_n1398_n197# a_n2448_131# 0.00fF
C1415 a_492_131# a_n348_131# 0.01fF
C1416 a_1544_n730# a_284_n730# 0.00fF
C1417 a_238_n100# a_n720_n100# 0.01fF
C1418 a_330_n100# a_n812_n100# 0.01fF
C1419 a_n1442_n100# a_n1398_n197# 0.00fF
C1420 a_3434_n401# a_3432_131# 0.01fF
C1421 a_n1440_n633# a_n1398_n197# 0.00fF
C1422 a_n1350_n100# a_n1398_n197# 0.00fF
C1423 a_n1650_n633# a_n1606_n401# 0.00fF
C1424 a_912_131# a_72_131# 0.01fF
C1425 a_n138_n197# w_n4520_n852# 0.10fF
C1426 a_4112_n633# a_2970_n633# 0.01fF
C1427 a_n1650_n633# a_n1768_n633# 0.07fF
C1428 a_3480_n100# a_3388_n100# 0.09fF
C1429 a_3902_n633# a_3900_n100# 0.00fF
C1430 a_2010_n100# a_1962_n197# 0.00fF
C1431 a_n1818_n197# a_n2448_131# 0.00fF
C1432 a_238_n100# a_n812_n100# 0.01fF
C1433 a_330_n100# a_n930_n100# 0.00fF
C1434 a_n1768_n633# a_n2608_n633# 0.01fF
C1435 a_3482_n633# a_2642_n633# 0.01fF
C1436 a_n1652_n100# a_n2492_n100# 0.01fF
C1437 a_n1560_n100# a_n2610_n100# 0.01fF
C1438 a_540_n100# a_492_131# 0.00fF
C1439 a_4020_n633# a_2970_n633# 0.01fF
C1440 a_n2238_n197# a_n2448_131# 0.01fF
C1441 a_1918_n100# a_1962_n197# 0.00fF
C1442 a_870_n633# a_752_n633# 0.07fF
C1443 a_238_n100# a_n930_n100# 0.01fF
C1444 a_n3658_n633# a_n3750_n633# 0.09fF
C1445 a_3390_n633# a_2642_n633# 0.01fF
C1446 a_n1768_n633# a_n2700_n633# 0.01fF
C1447 a_3272_n633# w_n4520_n852# 0.03fF
C1448 a_n2190_n100# a_n2610_n100# 0.02fF
C1449 a_n3540_n633# a_n3750_n633# 0.03fF
C1450 a_n3750_n633# w_n4520_n852# 0.04fF
C1451 a_n1230_n633# a_n1186_n401# 0.00fF
C1452 a_n2608_n633# a_n2610_n100# 0.00fF
C1453 a_n1022_n100# a_n1560_n100# 0.01fF
C1454 a_3902_n633# a_2970_n633# 0.01fF
C1455 a_3810_n633# a_3808_n100# 0.00fF
C1456 a_n2658_n197# a_n2448_131# 0.01fF
C1457 a_n1768_n633# a_n2818_n633# 0.01fF
C1458 a_3692_n633# a_3644_n730# 0.00fF
C1459 a_962_n633# w_n4520_n852# 0.01fF
C1460 a_n3240_n100# a_n3288_131# 0.00fF
C1461 a_n976_n730# a_n930_n100# 0.00fF
C1462 a_n508_n633# a_n600_n633# 0.09fF
C1463 a_1498_n100# a_1542_n197# 0.00fF
C1464 a_1122_n197# a_1752_131# 0.00fF
C1465 a_282_n197# a_n558_n197# 0.01fF
C1466 a_3178_n100# a_3222_n197# 0.00fF
C1467 a_2850_n100# a_1380_n100# 0.00fF
C1468 a_1122_n197# a_2172_131# 0.00fF
C1469 a_3810_n633# a_2970_n633# 0.01fF
C1470 a_n3078_n197# a_n2448_131# 0.00fF
C1471 a_n1022_n100# a_n2190_n100# 0.01fF
C1472 a_3180_n633# a_3224_n730# 0.00fF
C1473 a_n2492_n100# a_n2610_n100# 0.07fF
C1474 a_n1230_n633# a_n1768_n633# 0.01fF
C1475 a_n1768_n633# a_n2910_n633# 0.01fF
C1476 a_n3332_n100# a_n3288_131# 0.00fF
C1477 a_n508_n633# a_n718_n633# 0.03fF
C1478 a_n1652_n100# a_n1980_n100# 0.02fF
C1479 a_n2072_n100# a_n2702_n100# 0.01fF
C1480 a_962_n633# a_914_n401# 0.00fF
C1481 a_2758_n100# a_1380_n100# 0.00fF
C1482 a_332_n633# a_284_n730# 0.00fF
C1483 a_3692_n633# a_2970_n633# 0.01fF
C1484 a_3600_n633# a_3062_n633# 0.01fF
C1485 a_n510_n100# a_n2072_n100# 0.00fF
C1486 a_n3498_n197# a_n2448_131# 0.00fF
C1487 a_1498_n100# a_960_n100# 0.01fF
C1488 a_n1768_n633# a_n3028_n633# 0.00fF
C1489 a_1752_131# a_912_131# 0.01fF
C1490 a_n1232_n100# a_n2400_n100# 0.01fF
C1491 a_n508_n633# a_n810_n633# 0.02fF
C1492 a_n600_n633# a_n718_n633# 0.07fF
C1493 a_2172_131# a_912_131# 0.00fF
C1494 a_n2072_n100# a_n2820_n100# 0.01fF
C1495 a_n1022_n100# a_n2492_n100# 0.00fF
C1496 a_2804_n730# a_3014_n401# 0.01fF
C1497 a_2640_n100# a_1380_n100# 0.00fF
C1498 a_240_n633# a_284_n730# 0.00fF
C1499 a_n2818_n633# a_n2866_n401# 0.00fF
C1500 a_n602_n100# a_n2072_n100# 0.00fF
C1501 a_n2028_131# w_n4520_n852# 0.12fF
C1502 a_n3918_n197# a_n2448_131# 0.00fF
C1503 a_n3752_n100# a_n4172_n100# 0.02fF
C1504 a_2640_n100# a_1078_n100# 0.00fF
C1505 a_n1768_n633# a_n3120_n633# 0.00fF
C1506 a_n3870_n100# w_n4520_n852# 0.05fF
C1507 a_3272_n633# a_2550_n633# 0.01fF
C1508 a_1288_n100# a_1380_n100# 0.09fF
C1509 a_n600_n633# a_n810_n633# 0.03fF
C1510 a_n508_n633# a_n928_n633# 0.02fF
C1511 a_1334_n401# w_n4520_n852# 0.10fF
C1512 a_n2026_n401# a_n1980_n100# 0.00fF
C1513 a_702_n197# a_n138_n197# 0.01fF
C1514 a_3434_n401# a_3480_n100# 0.00fF
C1515 a_4064_n730# a_2804_n730# 0.00fF
C1516 a_n2072_n100# a_n2912_n100# 0.01fF
C1517 a_1288_n100# a_1078_n100# 0.03fF
C1518 a_2804_n730# a_2594_n401# 0.01fF
C1519 a_n1186_n401# a_n1140_n100# 0.00fF
C1520 a_2384_n730# a_3014_n401# 0.00fF
C1521 a_2548_n100# a_1380_n100# 0.01fF
C1522 a_2852_n633# a_1592_n633# 0.00fF
C1523 a_n2910_n633# a_n2866_n401# 0.00fF
C1524 a_n720_n100# a_n2072_n100# 0.00fF
C1525 a_n1140_n100# a_n1652_n100# 0.01fF
C1526 a_494_n401# w_n4520_n852# 0.10fF
C1527 a_2548_n100# a_1078_n100# 0.00fF
C1528 a_2550_n633# a_962_n633# 0.00fF
C1529 a_1544_n730# a_1590_n100# 0.00fF
C1530 a_n1768_n633# a_n3238_n633# 0.00fF
C1531 a_n1560_n100# a_n1608_131# 0.00fF
C1532 a_n1980_n100# a_n2610_n100# 0.01fF
C1533 a_n600_n633# a_n928_n633# 0.02fF
C1534 a_n718_n633# a_n810_n633# 0.09fF
C1535 a_n508_n633# a_n1020_n633# 0.01fF
C1536 a_n4078_n633# a_n4080_n100# 0.00fF
C1537 a_1498_n100# a_448_n100# 0.01fF
C1538 a_n2608_n633# a_n3330_n633# 0.01fF
C1539 a_3644_n730# a_2804_n730# 0.01fF
C1540 a_n2072_n100# a_n3030_n100# 0.01fF
C1541 a_n1348_n633# w_n4520_n852# 0.01fF
C1542 a_n138_n197# a_n978_n197# 0.01fF
C1543 a_1964_n730# a_3014_n401# 0.00fF
C1544 a_2384_n730# a_2594_n401# 0.01fF
C1545 a_2802_n197# a_1752_131# 0.00fF
C1546 a_2430_n100# a_1380_n100# 0.01fF
C1547 a_2760_n633# a_1592_n633# 0.01fF
C1548 a_2852_n633# a_1500_n633# 0.00fF
C1549 a_3598_n100# a_2850_n100# 0.01fF
C1550 a_28_n100# a_n1560_n100# 0.00fF
C1551 a_1334_n401# a_914_n401# 0.01fF
C1552 a_n812_n100# a_n2072_n100# 0.00fF
C1553 a_2802_n197# a_2172_131# 0.00fF
C1554 a_74_n401# w_n4520_n852# 0.10fF
C1555 a_2430_n100# a_1078_n100# 0.00fF
C1556 a_n600_n633# a_n1020_n633# 0.02fF
C1557 a_n718_n633# a_n928_n633# 0.03fF
C1558 a_n1650_n633# a_n1608_131# 0.00fF
C1559 a_3644_n730# a_2384_n730# 0.00fF
C1560 a_n2608_n633# a_n3448_n633# 0.01fF
C1561 a_n2700_n633# a_n3330_n633# 0.01fF
C1562 a_n2072_n100# a_n3122_n100# 0.01fF
C1563 a_914_n401# a_494_n401# 0.01fF
C1564 a_n2190_n100# a_n3752_n100# 0.00fF
C1565 a_1544_n730# a_3014_n401# 0.00fF
C1566 a_n138_n197# a_n1398_n197# 0.00fF
C1567 a_1964_n730# a_2594_n401# 0.00fF
C1568 a_2338_n100# a_1380_n100# 0.01fF
C1569 a_2760_n633# a_1500_n633# 0.00fF
C1570 a_2642_n633# w_n4520_n852# 0.02fF
C1571 a_2852_n633# a_1382_n633# 0.00fF
C1572 a_n4126_n401# a_n4128_131# 0.01fF
C1573 a_3480_n100# a_2850_n100# 0.01fF
C1574 a_3598_n100# a_2758_n100# 0.01fF
C1575 a_n90_n100# a_n1560_n100# 0.00fF
C1576 a_n2400_n100# a_n2448_131# 0.00fF
C1577 a_n1022_n100# a_n1980_n100# 0.01fF
C1578 a_n930_n100# a_n2072_n100# 0.01fF
C1579 a_n1442_n100# a_n2400_n100# 0.01fF
C1580 a_2338_n100# a_1078_n100# 0.00fF
C1581 a_n346_n401# w_n4520_n852# 0.10fF
C1582 a_2130_n633# a_2172_131# 0.00fF
C1583 a_1380_n100# a_868_n100# 0.01fF
C1584 a_122_n633# a_n508_n633# 0.01fF
C1585 a_n1350_n100# a_n2400_n100# 0.01fF
C1586 a_n718_n633# a_n1020_n633# 0.02fF
C1587 a_n810_n633# a_n928_n633# 0.07fF
C1588 a_n2700_n633# a_n3448_n633# 0.01fF
C1589 a_n2818_n633# a_n3330_n633# 0.01fF
C1590 a_1078_n100# a_868_n100# 0.03fF
C1591 a_n2072_n100# a_n3240_n100# 0.01fF
C1592 a_914_n401# a_74_n401# 0.01fF
C1593 a_n1140_n100# a_n2610_n100# 0.00fF
C1594 a_4062_n197# w_n4520_n852# 0.10fF
C1595 a_1544_n730# a_2594_n401# 0.00fF
C1596 a_2220_n100# a_1380_n100# 0.01fF
C1597 a_2852_n633# a_1290_n633# 0.00fF
C1598 a_2760_n633# a_1382_n633# 0.00fF
C1599 a_3480_n100# a_2758_n100# 0.01fF
C1600 a_n182_n100# a_n1560_n100# 0.00fF
C1601 a_3598_n100# a_2640_n100# 0.01fF
C1602 a_3388_n100# a_2850_n100# 0.01fF
C1603 a_1080_n633# a_n88_n633# 0.01fF
C1604 a_2220_n100# a_1078_n100# 0.01fF
C1605 a_n766_n401# w_n4520_n852# 0.10fF
C1606 a_1380_n100# a_750_n100# 0.01fF
C1607 a_122_n633# a_n600_n633# 0.01fF
C1608 a_30_n633# a_n508_n633# 0.01fF
C1609 a_1498_n100# a_658_n100# 0.01fF
C1610 a_n2492_n100# a_n3752_n100# 0.00fF
C1611 a_n810_n633# a_n1020_n633# 0.03fF
C1612 a_n2910_n633# a_n3330_n633# 0.02fF
C1613 a_1078_n100# a_750_n100# 0.02fF
C1614 a_n2818_n633# a_n3448_n633# 0.01fF
C1615 a_n2072_n100# a_n3332_n100# 0.00fF
C1616 a_914_n401# a_n346_n401# 0.00fF
C1617 a_2128_n100# a_1380_n100# 0.01fF
C1618 a_2760_n633# a_1290_n633# 0.00fF
C1619 a_3598_n100# a_2548_n100# 0.01fF
C1620 a_3480_n100# a_2640_n100# 0.01fF
C1621 a_3388_n100# a_2758_n100# 0.01fF
C1622 a_n300_n100# a_n1560_n100# 0.00fF
C1623 a_1080_n633# a_n180_n633# 0.00fF
C1624 a_2592_131# w_n4520_n852# 0.12fF
C1625 a_n1186_n401# w_n4520_n852# 0.10fF
C1626 a_2128_n100# a_1078_n100# 0.01fF
C1627 a_n2702_n100# a_n4172_n100# 0.00fF
C1628 a_30_n633# a_n600_n633# 0.01fF
C1629 a_n1652_n100# w_n4520_n852# 0.02fF
C1630 a_122_n633# a_n718_n633# 0.01fF
C1631 a_n1022_n100# a_n1140_n100# 0.07fF
C1632 a_n928_n633# a_n1020_n633# 0.09fF
C1633 a_962_n633# a_660_n633# 0.02fF
C1634 a_n3028_n633# a_n3330_n633# 0.02fF
C1635 a_n2910_n633# a_n3448_n633# 0.01fF
C1636 a_n2072_n100# a_n3450_n100# 0.00fF
C1637 a_1380_n100# a_330_n100# 0.01fF
C1638 a_n1138_n633# a_n2070_n633# 0.01fF
C1639 a_1124_n730# a_704_n730# 0.01fF
C1640 a_2852_n633# a_2432_n633# 0.02fF
C1641 a_2010_n100# a_1380_n100# 0.01fF
C1642 a_2760_n633# a_1172_n633# 0.00fF
C1643 a_4020_n633# a_4018_n100# 0.00fF
C1644 a_3598_n100# a_2430_n100# 0.01fF
C1645 a_3480_n100# a_2548_n100# 0.01fF
C1646 a_960_n100# a_448_n100# 0.01fF
C1647 a_n392_n100# a_n1560_n100# 0.01fF
C1648 a_3388_n100# a_2640_n100# 0.01fF
C1649 a_1078_n100# a_330_n100# 0.01fF
C1650 a_3854_n401# a_3434_n401# 0.01fF
C1651 a_n3750_n633# a_n3868_n633# 0.07fF
C1652 a_1080_n633# a_n298_n633# 0.00fF
C1653 a_n558_n197# w_n4520_n852# 0.10fF
C1654 a_1592_n633# a_870_n633# 0.01fF
C1655 a_n2820_n100# a_n4172_n100# 0.00fF
C1656 a_2010_n100# a_1078_n100# 0.01fF
C1657 a_n1606_n401# w_n4520_n852# 0.10fF
C1658 a_30_n633# a_n718_n633# 0.01fF
C1659 a_122_n633# a_n810_n633# 0.01fF
C1660 a_1288_n100# a_540_n100# 0.01fF
C1661 a_n1768_n633# w_n4520_n852# 0.01fF
C1662 a_n1560_n100# a_n2702_n100# 0.01fF
C1663 a_n3120_n633# a_n3330_n633# 0.03fF
C1664 a_n3028_n633# a_n3448_n633# 0.02fF
C1665 a_1380_n100# a_238_n100# 0.01fF
C1666 a_n2072_n100# a_n3542_n100# 0.00fF
C1667 a_n1138_n633# a_n2188_n633# 0.01fF
C1668 a_1124_n730# a_284_n730# 0.01fF
C1669 a_2970_n633# a_2222_n633# 0.01fF
C1670 a_2852_n633# a_2340_n633# 0.01fF
C1671 a_2760_n633# a_2432_n633# 0.02fF
C1672 a_2642_n633# a_2550_n633# 0.09fF
C1673 a_1710_n633# a_1752_131# 0.00fF
C1674 a_1918_n100# a_1380_n100# 0.01fF
C1675 a_3598_n100# a_2338_n100# 0.00fF
C1676 a_3480_n100# a_2430_n100# 0.01fF
C1677 a_1078_n100# a_238_n100# 0.01fF
C1678 a_n510_n100# a_n1560_n100# 0.01fF
C1679 a_3388_n100# a_2548_n100# 0.01fF
C1680 a_1542_n197# a_72_131# 0.00fF
C1681 a_1080_n633# a_n390_n633# 0.00fF
C1682 a_1500_n633# a_870_n633# 0.01fF
C1683 a_752_n633# w_n4520_n852# 0.01fF
C1684 a_n978_n197# a_n2028_131# 0.00fF
C1685 a_n2912_n100# a_n4172_n100# 0.00fF
C1686 a_1918_n100# a_1078_n100# 0.01fF
C1687 a_n2026_n401# w_n4520_n852# 0.10fF
C1688 a_30_n633# a_n810_n633# 0.01fF
C1689 a_122_n633# a_n928_n633# 0.01fF
C1690 a_332_n633# a_n1138_n633# 0.00fF
C1691 a_n3076_n730# a_n3916_n730# 0.01fF
C1692 a_n3238_n633# a_n3330_n633# 0.09fF
C1693 a_n1560_n100# a_n2820_n100# 0.00fF
C1694 a_n3120_n633# a_n3448_n633# 0.02fF
C1695 a_n2072_n100# a_n3660_n100# 0.00fF
C1696 a_n1138_n633# a_n2280_n633# 0.01fF
C1697 a_1124_n730# a_n136_n730# 0.00fF
C1698 a_704_n730# a_284_n730# 0.01fF
C1699 a_2760_n633# a_2340_n633# 0.02fF
C1700 a_2970_n633# a_2130_n633# 0.01fF
C1701 a_n2190_n100# a_n2702_n100# 0.01fF
C1702 a_n3750_n633# a_n3706_n401# 0.00fF
C1703 a_3598_n100# a_2220_n100# 0.00fF
C1704 a_n602_n100# a_n1560_n100# 0.01fF
C1705 a_1170_n100# a_28_n100# 0.01fF
C1706 a_3480_n100# a_2338_n100# 0.01fF
C1707 a_3388_n100# a_2430_n100# 0.01fF
C1708 a_n1398_n197# a_n2028_131# 0.00fF
C1709 a_1382_n633# a_870_n633# 0.01fF
C1710 a_n3030_n100# a_n4172_n100# 0.01fF
C1711 a_n2610_n100# w_n4520_n852# 0.02fF
C1712 a_n2446_n401# w_n4520_n852# 0.10fF
C1713 a_122_n633# a_n1020_n633# 0.01fF
C1714 a_240_n633# a_n1138_n633# 0.00fF
C1715 a_30_n633# a_n928_n633# 0.01fF
C1716 a_3224_n730# a_3270_n100# 0.00fF
C1717 a_n1560_n100# a_n2912_n100# 0.00fF
C1718 a_n3238_n633# a_n3448_n633# 0.03fF
C1719 a_4112_n633# a_3272_n633# 0.01fF
C1720 a_4062_n197# a_3642_n197# 0.01fF
C1721 a_960_n100# a_658_n100# 0.02fF
C1722 a_704_n730# a_n136_n730# 0.01fF
C1723 a_n1138_n633# a_n2398_n633# 0.00fF
C1724 a_2970_n633# a_2012_n633# 0.01fF
C1725 a_n2190_n100# a_n2820_n100# 0.01fF
C1726 a_1590_n100# a_1498_n100# 0.09fF
C1727 a_n720_n100# a_n1560_n100# 0.01fF
C1728 a_3480_n100# a_2220_n100# 0.00fF
C1729 a_3598_n100# a_2128_n100# 0.00fF
C1730 a_1170_n100# a_n90_n100# 0.00fF
C1731 a_3388_n100# a_2338_n100# 0.01fF
C1732 a_2550_n633# a_2592_131# 0.00fF
C1733 a_3690_n100# a_3270_n100# 0.02fF
C1734 a_n1818_n197# a_n2028_131# 0.01fF
C1735 a_1290_n633# a_870_n633# 0.02fF
C1736 a_n3122_n100# a_n4172_n100# 0.01fF
C1737 a_n602_n100# a_n2190_n100# 0.00fF
C1738 a_n2700_n633# a_n2702_n100# 0.00fF
C1739 a_n2866_n401# w_n4520_n852# 0.10fF
C1740 a_30_n633# a_n1020_n633# 0.01fF
C1741 a_n1348_n633# a_n1860_n633# 0.01fF
C1742 a_868_n100# a_540_n100# 0.02fF
C1743 a_n2492_n100# a_n2702_n100# 0.03fF
C1744 a_n1560_n100# a_n3030_n100# 0.00fF
C1745 a_4020_n633# a_3272_n633# 0.01fF
C1746 a_n3868_n633# a_n3870_n100# 0.00fF
C1747 a_n1022_n100# w_n4520_n852# 0.02fF
C1748 a_n1138_n633# a_n2490_n633# 0.00fF
C1749 a_704_n730# a_n556_n730# 0.00fF
C1750 a_284_n730# a_n136_n730# 0.01fF
C1751 a_2970_n633# a_1920_n633# 0.01fF
C1752 a_n2190_n100# a_n2912_n100# 0.01fF
C1753 a_3598_n100# a_2010_n100# 0.00fF
C1754 a_3480_n100# a_2128_n100# 0.00fF
C1755 a_3388_n100# a_2220_n100# 0.01fF
C1756 a_3642_n197# a_2592_131# 0.00fF
C1757 a_n812_n100# a_n1560_n100# 0.01fF
C1758 a_1170_n100# a_n182_n100# 0.00fF
C1759 a_n2238_n197# a_n2028_131# 0.01fF
C1760 a_1172_n633# a_870_n633# 0.02fF
C1761 a_n3240_n100# a_n4172_n100# 0.01fF
C1762 a_n720_n100# a_n2190_n100# 0.00fF
C1763 a_332_n633# a_n88_n633# 0.02fF
C1764 a_750_n100# a_540_n100# 0.03fF
C1765 a_n2492_n100# a_n2820_n100# 0.02fF
C1766 a_28_n100# a_n1140_n100# 0.01fF
C1767 a_n1560_n100# a_n3122_n100# 0.00fF
C1768 a_3902_n633# a_3272_n633# 0.01fF
C1769 a_284_n730# a_n556_n730# 0.01fF
C1770 a_2970_n633# a_1802_n633# 0.01fF
C1771 a_n2190_n100# a_n3030_n100# 0.01fF
C1772 a_2128_n100# a_540_n100# 0.00fF
C1773 a_1170_n100# a_n300_n100# 0.00fF
C1774 a_3480_n100# a_2010_n100# 0.00fF
C1775 a_n930_n100# a_n1560_n100# 0.01fF
C1776 a_3388_n100# a_2128_n100# 0.00fF
C1777 a_2432_n633# a_870_n633# 0.00fF
C1778 a_658_n100# a_448_n100# 0.03fF
C1779 a_n2658_n197# a_n2028_131# 0.00fF
C1780 a_n812_n100# a_n2190_n100# 0.00fF
C1781 a_n3332_n100# a_n4172_n100# 0.01fF
C1782 a_332_n633# a_n180_n633# 0.01fF
C1783 a_240_n633# a_n88_n633# 0.02fF
C1784 a_n2818_n633# a_n2820_n100# 0.00fF
C1785 a_122_n633# a_30_n633# 0.09fF
C1786 a_n2492_n100# a_n2912_n100# 0.02fF
C1787 a_n90_n100# a_n1140_n100# 0.01fF
C1788 a_1590_n100# a_1542_n197# 0.00fF
C1789 a_n1652_n100# a_n1770_n100# 0.07fF
C1790 a_n2236_n730# a_n3496_n730# 0.00fF
C1791 a_3810_n633# a_3272_n633# 0.01fF
C1792 a_1542_n197# a_1752_131# 0.01fF
C1793 a_n136_n730# a_n556_n730# 0.01fF
C1794 a_540_n100# a_330_n100# 0.03fF
C1795 a_2970_n633# a_1710_n633# 0.00fF
C1796 a_n2190_n100# a_n3122_n100# 0.01fF
C1797 a_702_n197# a_n558_n197# 0.00fF
C1798 a_3480_n100# a_1918_n100# 0.00fF
C1799 a_1170_n100# a_n392_n100# 0.00fF
C1800 a_3388_n100# a_2010_n100# 0.00fF
C1801 a_2010_n100# a_540_n100# 0.00fF
C1802 a_2340_n633# a_870_n633# 0.00fF
C1803 a_1542_n197# a_2172_131# 0.00fF
C1804 a_n392_n100# a_n1980_n100# 0.00fF
C1805 a_n3078_n197# a_n2028_131# 0.00fF
C1806 a_n3450_n100# a_n4172_n100# 0.01fF
C1807 a_n930_n100# a_n2190_n100# 0.00fF
C1808 a_332_n633# a_n298_n633# 0.01fF
C1809 a_282_n197# a_1332_131# 0.00fF
C1810 a_240_n633# a_n180_n633# 0.02fF
C1811 a_n3330_n633# a_n3658_n633# 0.02fF
C1812 a_n182_n100# a_n1140_n100# 0.01fF
C1813 a_n2492_n100# a_n3030_n100# 0.01fF
C1814 a_n2656_n730# a_n3496_n730# 0.01fF
C1815 a_n1652_n100# a_n1862_n100# 0.03fF
C1816 a_3692_n633# a_3272_n633# 0.02fF
C1817 a_n3330_n633# a_n3540_n633# 0.03fF
C1818 a_n1980_n100# a_n2702_n100# 0.01fF
C1819 a_540_n100# a_238_n100# 0.02fF
C1820 a_n2190_n100# a_n3240_n100# 0.01fF
C1821 a_n1768_n633# a_n1770_n100# 0.00fF
C1822 a_n3330_n633# w_n4520_n852# 0.03fF
C1823 a_2850_n100# a_2758_n100# 0.09fF
C1824 a_3388_n100# a_1918_n100# 0.00fF
C1825 a_1918_n100# a_540_n100# 0.00fF
C1826 a_n510_n100# a_n1980_n100# 0.00fF
C1827 a_n1558_n633# a_n1978_n633# 0.02fF
C1828 a_n1440_n633# a_n2070_n633# 0.01fF
C1829 a_n3498_n197# a_n2028_131# 0.00fF
C1830 a_3598_n100# a_3178_n100# 0.02fF
C1831 a_n3542_n100# a_n4172_n100# 0.01fF
C1832 a_2968_n100# a_3012_131# 0.00fF
C1833 a_n558_n197# a_n978_n197# 0.01fF
C1834 a_332_n633# a_n390_n633# 0.01fF
C1835 a_240_n633# a_n298_n633# 0.01fF
C1836 a_n2910_n633# a_n2912_n100# 0.00fF
C1837 a_1590_n100# a_960_n100# 0.01fF
C1838 a_n3448_n633# a_n3658_n633# 0.03fF
C1839 a_n300_n100# a_n1140_n100# 0.01fF
C1840 a_n2492_n100# a_n3122_n100# 0.01fF
C1841 a_n1980_n100# a_n2820_n100# 0.01fF
C1842 a_n3448_n633# a_n3540_n633# 0.09fF
C1843 a_n930_n100# a_n2492_n100# 0.00fF
C1844 a_3180_n633# a_2970_n633# 0.03fF
C1845 a_n2190_n100# a_n3332_n100# 0.01fF
C1846 a_3224_n730# a_3014_n401# 0.01fF
C1847 a_n3448_n633# w_n4520_n852# 0.03fF
C1848 a_2850_n100# a_2640_n100# 0.03fF
C1849 a_n3962_n100# a_n4080_n100# 0.07fF
C1850 a_n602_n100# a_n1980_n100# 0.00fF
C1851 a_n1768_n633# a_n1860_n633# 0.09fF
C1852 a_n1440_n633# a_n2188_n633# 0.01fF
C1853 a_n1650_n633# a_n1978_n633# 0.02fF
C1854 a_n1608_131# w_n4520_n852# 0.12fF
C1855 a_n558_n197# a_n1398_n197# 0.01fF
C1856 a_3480_n100# a_3178_n100# 0.02fF
C1857 a_n3660_n100# a_n4172_n100# 0.01fF
C1858 a_240_n633# a_n390_n633# 0.01fF
C1859 a_n4126_n401# w_n4520_n852# 0.12fF
C1860 a_1172_n633# a_1170_n100# 0.00fF
C1861 a_1288_n100# a_2850_n100# 0.00fF
C1862 a_n3752_n100# w_n4520_n852# 0.04fF
C1863 a_n1978_n633# a_n2608_n633# 0.01fF
C1864 a_3482_n633# a_2432_n633# 0.01fF
C1865 a_n2492_n100# a_n3240_n100# 0.01fF
C1866 a_n1770_n100# a_n2610_n100# 0.01fF
C1867 a_n392_n100# a_n1140_n100# 0.01fF
C1868 a_n3870_n100# a_n3918_n197# 0.00fF
C1869 a_1122_n197# a_n138_n197# 0.00fF
C1870 a_4064_n730# a_3224_n730# 0.01fF
C1871 a_n1980_n100# a_n2912_n100# 0.01fF
C1872 a_28_n100# w_n4520_n852# 0.02fF
C1873 a_n2190_n100# a_n3450_n100# 0.00fF
C1874 a_3224_n730# a_2594_n401# 0.00fF
C1875 a_2850_n100# a_2548_n100# 0.02fF
C1876 a_2758_n100# a_2640_n100# 0.07fF
C1877 a_n720_n100# a_n1980_n100# 0.00fF
C1878 a_n1440_n633# a_n2280_n633# 0.01fF
C1879 a_4112_n633# a_2642_n633# 0.00fF
C1880 a_n1140_n100# a_n2702_n100# 0.00fF
C1881 a_n558_n197# a_n1818_n197# 0.00fF
C1882 a_3388_n100# a_3178_n100# 0.03fF
C1883 a_n3028_n633# a_n3030_n100# 0.00fF
C1884 a_752_n633# a_660_n633# 0.09fF
C1885 a_870_n633# a_542_n633# 0.02fF
C1886 a_n2868_131# a_n3708_131# 0.01fF
C1887 a_1288_n100# a_2758_n100# 0.00fF
C1888 a_n1978_n633# a_n2700_n633# 0.01fF
C1889 a_3482_n633# a_2340_n633# 0.01fF
C1890 a_3390_n633# a_2432_n633# 0.01fF
C1891 a_n510_n100# a_n1140_n100# 0.01fF
C1892 a_n1862_n100# a_n2610_n100# 0.01fF
C1893 a_n2492_n100# a_n3332_n100# 0.01fF
C1894 a_1590_n100# a_448_n100# 0.01fF
C1895 a_3644_n730# a_3224_n730# 0.01fF
C1896 a_n1980_n100# a_n3030_n100# 0.01fF
C1897 a_n90_n100# w_n4520_n852# 0.02fF
C1898 a_n2190_n100# a_n3542_n100# 0.00fF
C1899 a_2850_n100# a_2430_n100# 0.02fF
C1900 a_2758_n100# a_2548_n100# 0.03fF
C1901 a_3900_n100# a_3690_n100# 0.03fF
C1902 a_n812_n100# a_n1980_n100# 0.01fF
C1903 a_n1022_n100# a_n1770_n100# 0.01fF
C1904 a_n1440_n633# a_n2398_n633# 0.01fF
C1905 a_4020_n633# a_2642_n633# 0.00fF
C1906 a_n2608_n633# a_n3960_n633# 0.00fF
C1907 a_870_n633# a_450_n633# 0.02fF
C1908 a_n138_n197# a_912_131# 0.00fF
C1909 a_3644_n730# a_3690_n100# 0.00fF
C1910 a_1288_n100# a_2640_n100# 0.00fF
C1911 a_n3288_131# a_n3708_131# 0.01fF
C1912 a_n1978_n633# a_n2818_n633# 0.01fF
C1913 a_1124_n730# a_2594_n401# 0.00fF
C1914 a_3390_n633# a_2340_n633# 0.01fF
C1915 a_n2492_n100# a_n3450_n100# 0.01fF
C1916 a_n602_n100# a_n1140_n100# 0.01fF
C1917 a_n2490_n633# a_n2448_131# 0.00fF
C1918 a_n1980_n100# a_n3122_n100# 0.01fF
C1919 a_n182_n100# w_n4520_n852# 0.02fF
C1920 a_n1022_n100# a_n978_n197# 0.00fF
C1921 a_n2190_n100# a_n3660_n100# 0.00fF
C1922 a_2640_n100# a_2548_n100# 0.09fF
C1923 a_2850_n100# a_2338_n100# 0.01fF
C1924 a_2758_n100# a_2430_n100# 0.02fF
C1925 a_4020_n633# a_4062_n197# 0.00fF
C1926 a_3808_n100# a_3690_n100# 0.07fF
C1927 a_n1022_n100# a_n1862_n100# 0.01fF
C1928 a_n930_n100# a_n1980_n100# 0.01fF
C1929 a_3902_n633# a_2642_n633# 0.00fF
C1930 a_n1440_n633# a_n2490_n633# 0.01fF
C1931 a_1592_n633# w_n4520_n852# 0.01fF
C1932 a_n2700_n633# a_n3960_n633# 0.00fF
C1933 a_n3120_n633# a_n3122_n100# 0.00fF
C1934 a_n1230_n633# a_n1978_n633# 0.01fF
C1935 a_n2400_n100# a_n3870_n100# 0.00fF
C1936 a_n2026_n401# a_n3286_n401# 0.00fF
C1937 a_1288_n100# a_2548_n100# 0.00fF
C1938 a_n1978_n633# a_n2910_n633# 0.01fF
C1939 a_n2492_n100# a_n3542_n100# 0.01fF
C1940 a_n720_n100# a_n1140_n100# 0.02fF
C1941 a_n1980_n100# a_n3240_n100# 0.00fF
C1942 a_n300_n100# w_n4520_n852# 0.02fF
C1943 a_2640_n100# a_2430_n100# 0.03fF
C1944 a_2850_n100# a_2220_n100# 0.01fF
C1945 a_2758_n100# a_2338_n100# 0.02fF
C1946 a_3600_n633# a_2852_n633# 0.01fF
C1947 a_3810_n633# a_2642_n633# 0.01fF
C1948 a_1500_n633# w_n4520_n852# 0.01fF
C1949 a_n928_n633# a_n976_n730# 0.00fF
C1950 a_n2818_n633# a_n3960_n633# 0.01fF
C1951 a_1590_n100# a_658_n100# 0.01fF
C1952 a_n2446_n401# a_n3286_n401# 0.01fF
C1953 a_1288_n100# a_2430_n100# 0.01fF
C1954 a_n1978_n633# a_n3028_n633# 0.01fF
C1955 a_n2492_n100# a_n3660_n100# 0.01fF
C1956 a_n812_n100# a_n1140_n100# 0.02fF
C1957 a_n1980_n100# a_n3332_n100# 0.00fF
C1958 a_n392_n100# w_n4520_n852# 0.02fF
C1959 a_1802_n633# a_1800_n100# 0.00fF
C1960 a_282_n197# a_n768_131# 0.00fF
C1961 a_2548_n100# a_2430_n100# 0.07fF
C1962 a_2640_n100# a_2338_n100# 0.02fF
C1963 a_2850_n100# a_2128_n100# 0.01fF
C1964 a_2758_n100# a_2220_n100# 0.01fF
C1965 a_n1978_n633# a_n1980_n100# 0.00fF
C1966 a_3692_n633# a_2642_n633# 0.01fF
C1967 a_3600_n633# a_2760_n633# 0.01fF
C1968 a_1382_n633# w_n4520_n852# 0.01fF
C1969 a_n1020_n633# a_n976_n730# 0.00fF
C1970 a_3012_131# w_n4520_n852# 0.13fF
C1971 a_n3238_n633# a_n3240_n100# 0.00fF
C1972 a_n2910_n633# a_n3960_n633# 0.01fF
C1973 a_n2610_n100# a_n2658_n197# 0.00fF
C1974 a_n2446_n401# a_n3706_n401# 0.00fF
C1975 a_n2866_n401# a_n3286_n401# 0.01fF
C1976 a_1288_n100# a_2338_n100# 0.01fF
C1977 a_n1978_n633# a_n3120_n633# 0.01fF
C1978 a_n2702_n100# w_n4520_n852# 0.02fF
C1979 a_1080_n633# a_962_n633# 0.07fF
C1980 a_n930_n100# a_n1140_n100# 0.03fF
C1981 a_n1980_n100# a_n3450_n100# 0.00fF
C1982 a_n510_n100# w_n4520_n852# 0.02fF
C1983 a_1288_n100# a_868_n100# 0.02fF
C1984 a_n1230_n633# a_n1188_131# 0.00fF
C1985 a_282_n197# a_n1188_131# 0.00fF
C1986 a_2758_n100# a_2128_n100# 0.01fF
C1987 a_2640_n100# a_2220_n100# 0.02fF
C1988 a_2548_n100# a_2338_n100# 0.03fF
C1989 a_2850_n100# a_2010_n100# 0.01fF
C1990 a_1290_n633# w_n4520_n852# 0.01fF
C1991 a_n3028_n633# a_n3960_n633# 0.01fF
C1992 a_n2866_n401# a_n3706_n401# 0.01fF
C1993 a_n1860_n633# a_n3330_n633# 0.00fF
C1994 a_1288_n100# a_2220_n100# 0.01fF
C1995 a_n1978_n633# a_n3238_n633# 0.00fF
C1996 a_n2820_n100# w_n4520_n852# 0.02fF
C1997 a_3272_n633# a_2222_n633# 0.01fF
C1998 a_1332_131# w_n4520_n852# 0.12fF
C1999 a_n1980_n100# a_n3542_n100# 0.00fF
C2000 a_n602_n100# w_n4520_n852# 0.02fF
C2001 a_1288_n100# a_750_n100# 0.01fF
C2002 a_1710_n633# a_1708_n100# 0.00fF
C2003 a_2548_n100# a_2220_n100# 0.02fF
C2004 a_2430_n100# a_2338_n100# 0.09fF
C2005 a_2640_n100# a_2128_n100# 0.01fF
C2006 a_2758_n100# a_2010_n100# 0.01fF
C2007 a_2850_n100# a_1918_n100# 0.01fF
C2008 a_2804_n730# a_1334_n401# 0.00fF
C2009 a_2550_n633# a_1592_n633# 0.01fF
C2010 a_n88_n633# a_n136_n730# 0.00fF
C2011 a_1172_n633# w_n4520_n852# 0.01fF
C2012 a_n978_n197# a_n1608_131# 0.00fF
C2013 a_n3120_n633# a_n3960_n633# 0.01fF
C2014 a_2430_n100# a_868_n100# 0.00fF
C2015 a_2222_n633# a_962_n633# 0.00fF
C2016 a_n1860_n633# a_n3448_n633# 0.00fF
C2017 a_1288_n100# a_2128_n100# 0.01fF
C2018 a_n2912_n100# w_n4520_n852# 0.03fF
C2019 a_3272_n633# a_2130_n633# 0.01fF
C2020 a_1498_n100# a_120_n100# 0.00fF
C2021 a_n720_n100# w_n4520_n852# 0.02fF
C2022 a_2640_n100# a_2010_n100# 0.01fF
C2023 a_2548_n100# a_2128_n100# 0.02fF
C2024 a_2758_n100# a_1918_n100# 0.01fF
C2025 a_2430_n100# a_2220_n100# 0.03fF
C2026 a_1800_n100# a_1498_n100# 0.02fF
C2027 a_2384_n730# a_1334_n401# 0.00fF
C2028 a_2550_n633# a_1500_n633# 0.01fF
C2029 a_n180_n633# a_n136_n730# 0.00fF
C2030 a_2432_n633# w_n4520_n852# 0.01fF
C2031 a_3900_n100# a_3270_n100# 0.01fF
C2032 a_1288_n100# a_330_n100# 0.01fF
C2033 a_n1398_n197# a_n1608_131# 0.01fF
C2034 a_n3330_n633# a_n3868_n633# 0.01fF
C2035 a_n3238_n633# a_n3960_n633# 0.01fF
C2036 a_4110_n100# a_3598_n100# 0.01fF
C2037 a_n1652_n100# a_n2400_n100# 0.01fF
C2038 a_2338_n100# a_868_n100# 0.00fF
C2039 a_2130_n633# a_962_n633# 0.01fF
C2040 a_1288_n100# a_2010_n100# 0.01fF
C2041 a_2382_n197# w_n4520_n852# 0.10fF
C2042 a_n3030_n100# w_n4520_n852# 0.03fF
C2043 a_3272_n633# a_2012_n633# 0.00fF
C2044 a_n812_n100# w_n4520_n852# 0.02fF
C2045 a_2338_n100# a_2220_n100# 0.07fF
C2046 a_2548_n100# a_2010_n100# 0.01fF
C2047 a_2430_n100# a_2128_n100# 0.02fF
C2048 a_2640_n100# a_1918_n100# 0.01fF
C2049 a_1964_n730# a_1334_n401# 0.00fF
C2050 a_1708_n100# a_1498_n100# 0.03fF
C2051 a_3222_n197# w_n4520_n852# 0.10fF
C2052 a_2340_n633# w_n4520_n852# 0.01fF
C2053 a_2550_n633# a_1382_n633# 0.01fF
C2054 a_n3330_n633# a_n3286_n401# 0.00fF
C2055 a_n182_n100# a_n1770_n100# 0.00fF
C2056 a_3178_n100# a_2850_n100# 0.02fF
C2057 a_1288_n100# a_238_n100# 0.01fF
C2058 a_3808_n100# a_3270_n100# 0.01fF
C2059 a_n1818_n197# a_n1608_131# 0.01fF
C2060 a_n3448_n633# a_n3868_n633# 0.02fF
C2061 a_4110_n100# a_3480_n100# 0.01fF
C2062 a_2338_n100# a_750_n100# 0.00fF
C2063 a_2220_n100# a_868_n100# 0.00fF
C2064 a_2012_n633# a_962_n633# 0.01fF
C2065 a_1962_n197# w_n4520_n852# 0.10fF
C2066 a_1288_n100# a_1918_n100# 0.01fF
C2067 a_n3122_n100# w_n4520_n852# 0.03fF
C2068 a_2172_131# a_1752_131# 0.01fF
C2069 a_3272_n633# a_1920_n633# 0.00fF
C2070 a_1964_n730# a_494_n401# 0.00fF
C2071 a_868_n100# a_750_n100# 0.07fF
C2072 a_n930_n100# w_n4520_n852# 0.02fF
C2073 a_n1140_n100# a_n1188_131# 0.00fF
C2074 a_2430_n100# a_2010_n100# 0.02fF
C2075 a_2338_n100# a_2128_n100# 0.03fF
C2076 a_2548_n100# a_1918_n100# 0.01fF
C2077 a_1544_n730# a_1334_n401# 0.01fF
C2078 a_3642_n197# a_3012_131# 0.00fF
C2079 a_2550_n633# a_1290_n633# 0.00fF
C2080 a_n300_n100# a_n1770_n100# 0.00fF
C2081 a_3178_n100# a_2758_n100# 0.02fF
C2082 a_3060_n100# a_1498_n100# 0.00fF
C2083 a_n2238_n197# a_n1608_131# 0.00fF
C2084 a_4110_n100# a_3388_n100# 0.01fF
C2085 a_2128_n100# a_868_n100# 0.00fF
C2086 a_2220_n100# a_750_n100# 0.00fF
C2087 a_1920_n633# a_962_n633# 0.01fF
C2088 a_n2188_n633# a_n3750_n633# 0.00fF
C2089 a_n3240_n100# w_n4520_n852# 0.03fF
C2090 a_n3286_n401# a_n4126_n401# 0.01fF
C2091 a_3272_n633# a_1802_n633# 0.00fF
C2092 a_1544_n730# a_494_n401# 0.00fF
C2093 a_1122_n197# a_2592_131# 0.00fF
C2094 a_2338_n100# a_2010_n100# 0.02fF
C2095 a_2220_n100# a_2128_n100# 0.09fF
C2096 a_2430_n100# a_1918_n100# 0.01fF
C2097 a_2642_n633# a_1080_n633# 0.00fF
C2098 a_2550_n633# a_1172_n633# 0.00fF
C2099 a_n300_n100# a_n1862_n100# 0.00fF
C2100 a_n392_n100# a_n1770_n100# 0.00fF
C2101 a_868_n100# a_330_n100# 0.01fF
C2102 a_3178_n100# a_2640_n100# 0.01fF
C2103 a_n2400_n100# a_n2610_n100# 0.03fF
C2104 a_n2446_n401# a_n2400_n100# 0.00fF
C2105 a_n3750_n633# a_n4078_n633# 0.02fF
C2106 a_n2658_n197# a_n1608_131# 0.00fF
C2107 a_n2072_n100# a_n2282_n100# 0.03fF
C2108 a_1592_n633# a_660_n633# 0.01fF
C2109 a_2128_n100# a_750_n100# 0.00fF
C2110 a_2010_n100# a_868_n100# 0.01fF
C2111 a_n2280_n633# a_n3750_n633# 0.00fF
C2112 a_1802_n633# a_962_n633# 0.01fF
C2113 a_n3332_n100# w_n4520_n852# 0.03fF
C2114 a_n3706_n401# a_n4126_n401# 0.01fF
C2115 a_n1978_n633# a_n3540_n633# 0.00fF
C2116 a_3272_n633# a_1710_n633# 0.00fF
C2117 a_962_n633# a_332_n633# 0.01fF
C2118 a_n1978_n633# w_n4520_n852# 0.01fF
C2119 a_1544_n730# a_74_n401# 0.00fF
C2120 a_n1770_n100# a_n2702_n100# 0.01fF
C2121 a_2220_n100# a_2010_n100# 0.03fF
C2122 a_2550_n633# a_2432_n633# 0.07fF
C2123 a_2338_n100# a_1918_n100# 0.02fF
C2124 a_960_n100# a_120_n100# 0.01fF
C2125 a_n510_n100# a_n1770_n100# 0.00fF
C2126 a_868_n100# a_238_n100# 0.01fF
C2127 a_n392_n100# a_n1862_n100# 0.00fF
C2128 a_750_n100# a_330_n100# 0.02fF
C2129 a_3178_n100# a_2548_n100# 0.01fF
C2130 a_n3078_n197# a_n1608_131# 0.00fF
C2131 a_702_n197# a_1332_131# 0.00fF
C2132 a_1500_n633# a_660_n633# 0.01fF
C2133 a_542_n633# w_n4520_n852# 0.01fF
C2134 a_1800_n100# a_960_n100# 0.01fF
C2135 a_2010_n100# a_750_n100# 0.00fF
C2136 a_1918_n100# a_868_n100# 0.01fF
C2137 a_n2398_n633# a_n3750_n633# 0.00fF
C2138 a_1710_n633# a_962_n633# 0.01fF
C2139 a_n3450_n100# w_n4520_n852# 0.03fF
C2140 a_962_n633# a_240_n633# 0.01fF
C2141 a_3390_n633# a_3432_131# 0.00fF
C2142 a_n1022_n100# a_n2400_n100# 0.00fF
C2143 a_n2070_n633# a_n2028_131# 0.00fF
C2144 a_3600_n633# a_3482_n633# 0.07fF
C2145 a_n1770_n100# a_n2820_n100# 0.01fF
C2146 a_n1862_n100# a_n2702_n100# 0.01fF
C2147 a_2550_n633# a_2340_n633# 0.03fF
C2148 a_2642_n633# a_2222_n633# 0.02fF
C2149 a_2128_n100# a_2010_n100# 0.07fF
C2150 a_2220_n100# a_1918_n100# 0.02fF
C2151 a_4064_n730# a_3014_n401# 0.00fF
C2152 a_n3916_n730# a_n3870_n100# 0.00fF
C2153 a_n3658_n633# a_n3960_n633# 0.02fF
C2154 a_n602_n100# a_n1770_n100# 0.01fF
C2155 a_750_n100# a_238_n100# 0.01fF
C2156 a_n510_n100# a_n1862_n100# 0.00fF
C2157 a_3014_n401# a_2594_n401# 0.01fF
C2158 a_3178_n100# a_2430_n100# 0.01fF
C2159 a_3434_n401# a_2174_n401# 0.00fF
C2160 a_n768_131# w_n4520_n852# 0.12fF
C2161 a_3642_n197# a_2382_n197# 0.00fF
C2162 a_450_n633# w_n4520_n852# 0.01fF
C2163 a_1382_n633# a_660_n633# 0.01fF
C2164 a_n3540_n633# a_n3542_n100# 0.00fF
C2165 a_n3540_n633# a_n3960_n633# 0.02fF
C2166 a_1708_n100# a_960_n100# 0.01fF
C2167 a_1918_n100# a_750_n100# 0.01fF
C2168 a_n2490_n633# a_n3750_n633# 0.00fF
C2169 a_1380_n100# a_1170_n100# 0.03fF
C2170 a_n3960_n633# w_n4520_n852# 0.06fF
C2171 a_n3542_n100# w_n4520_n852# 0.04fF
C2172 a_3272_n633# a_3180_n633# 0.09fF
C2173 a_n558_n197# a_912_131# 0.00fF
C2174 a_1170_n100# a_1078_n100# 0.09fF
C2175 a_3600_n633# a_3390_n633# 0.03fF
C2176 a_n1770_n100# a_n2912_n100# 0.01fF
C2177 a_n1862_n100# a_n2820_n100# 0.01fF
C2178 a_4062_n197# a_2802_n197# 0.00fF
C2179 a_3642_n197# a_3222_n197# 0.01fF
C2180 a_n508_n633# a_n1558_n633# 0.01fF
C2181 a_2642_n633# a_2130_n633# 0.01fF
C2182 a_2128_n100# a_1918_n100# 0.03fF
C2183 a_4018_n100# a_3690_n100# 0.02fF
C2184 a_3644_n730# a_3014_n401# 0.00fF
C2185 a_4064_n730# a_2594_n401# 0.00fF
C2186 a_n3658_n633# a_n3660_n100# 0.00fF
C2187 a_n720_n100# a_n1770_n100# 0.01fF
C2188 a_n602_n100# a_n1862_n100# 0.00fF
C2189 a_3178_n100# a_2338_n100# 0.01fF
C2190 a_n1188_131# w_n4520_n852# 0.12fF
C2191 a_3690_n100# a_3060_n100# 0.01fF
C2192 a_2968_n100# a_1380_n100# 0.00fF
C2193 a_1290_n633# a_660_n633# 0.01fF
C2194 a_330_n100# a_238_n100# 0.09fF
C2195 a_448_n100# a_120_n100# 0.02fF
C2196 a_n1348_n633# a_n2070_n633# 0.01fF
C2197 a_n3660_n100# w_n4520_n852# 0.04fF
C2198 a_n88_n633# a_n1138_n633# 0.01fF
C2199 a_1918_n100# a_330_n100# 0.00fF
C2200 a_1800_n100# a_448_n100# 0.00fF
C2201 a_4064_n730# a_3644_n730# 0.01fF
C2202 a_n1862_n100# a_n2912_n100# 0.01fF
C2203 a_n1770_n100# a_n3030_n100# 0.00fF
C2204 a_n600_n633# a_n1558_n633# 0.01fF
C2205 a_n508_n633# a_n1650_n633# 0.01fF
C2206 a_3644_n730# a_2594_n401# 0.00fF
C2207 a_2642_n633# a_2012_n633# 0.01fF
C2208 a_2010_n100# a_1918_n100# 0.09fF
C2209 a_2802_n197# a_2592_131# 0.01fF
C2210 a_n812_n100# a_n1770_n100# 0.01fF
C2211 a_n720_n100# a_n1862_n100# 0.01fF
C2212 a_3178_n100# a_2220_n100# 0.01fF
C2213 a_1962_n197# a_702_n197# 0.00fF
C2214 a_1172_n633# a_660_n633# 0.01fF
C2215 a_1080_n633# a_752_n633# 0.02fF
C2216 a_n1348_n633# a_n2188_n633# 0.01fF
C2217 a_n180_n633# a_n1138_n633# 0.01fF
C2218 a_n2868_131# a_n3288_131# 0.01fF
C2219 a_870_n633# a_n508_n633# 0.00fF
C2220 a_2970_n633# a_3014_n401# 0.00fF
C2221 a_1708_n100# a_448_n100# 0.00fF
C2222 a_n1862_n100# a_n3030_n100# 0.01fF
C2223 a_n1770_n100# a_n3122_n100# 0.00fF
C2224 a_2642_n633# a_1920_n633# 0.01fF
C2225 a_n718_n633# a_n1558_n633# 0.01fF
C2226 a_n600_n633# a_n1650_n633# 0.01fF
C2227 a_n812_n100# a_n1862_n100# 0.01fF
C2228 a_n930_n100# a_n1770_n100# 0.01fF
C2229 a_3900_n100# a_3808_n100# 0.09fF
C2230 a_3178_n100# a_2128_n100# 0.01fF
C2231 a_n1348_n633# a_n2280_n633# 0.01fF
C2232 a_n298_n633# a_n1138_n633# 0.01fF
C2233 a_870_n633# a_n600_n633# 0.00fF
C2234 a_n2702_n100# a_n2658_n197# 0.00fF
C2235 a_282_n197# a_n348_131# 0.00fF
C2236 a_n1862_n100# a_n3122_n100# 0.00fF
C2237 a_n1770_n100# a_n3240_n100# 0.00fF
C2238 a_n930_n100# a_n978_n197# 0.00fF
C2239 a_2642_n633# a_1802_n633# 0.01fF
C2240 a_n810_n633# a_n1558_n633# 0.01fF
C2241 a_n718_n633# a_n1650_n633# 0.01fF
C2242 a_3272_n633# a_3224_n730# 0.00fF
C2243 a_240_n633# a_n1348_n633# 0.00fF
C2244 a_n930_n100# a_n1862_n100# 0.01fF
C2245 a_3178_n100# a_2010_n100# 0.01fF
C2246 a_658_n100# a_120_n100# 0.01fF
C2247 a_2222_n633# a_752_n633# 0.00fF
C2248 a_120_n100# a_72_131# 0.00fF
C2249 a_282_n197# a_492_131# 0.01fF
C2250 a_n2400_n100# a_n3752_n100# 0.00fF
C2251 a_n1348_n633# a_n2398_n633# 0.01fF
C2252 a_1800_n100# a_658_n100# 0.01fF
C2253 a_n390_n633# a_n1138_n633# 0.01fF
C2254 a_870_n633# a_n718_n633# 0.00fF
C2255 a_3482_n633# a_3480_n100# 0.00fF
C2256 a_n1770_n100# a_n3332_n100# 0.00fF
C2257 a_n1862_n100# a_n3240_n100# 0.00fF
C2258 a_n810_n633# a_n1650_n633# 0.01fF
C2259 a_n928_n633# a_n1558_n633# 0.01fF
C2260 a_2642_n633# a_1710_n633# 0.01fF
C2261 a_2852_n633# a_2850_n100# 0.00fF
C2262 a_3270_n100# a_1800_n100# 0.00fF
C2263 a_3178_n100# a_1918_n100# 0.00fF
C2264 a_n3708_131# a_n4128_131# 0.01fF
C2265 a_n508_n633# a_n1230_n633# 0.01fF
C2266 a_2130_n633# a_752_n633# 0.00fF
C2267 a_4110_n100# a_2850_n100# 0.00fF
C2268 a_3852_131# w_n4520_n852# 0.11fF
C2269 a_3598_n100# a_2968_n100# 0.01fF
C2270 a_n4170_n633# a_n4172_n100# 0.00fF
C2271 a_n88_n633# a_n180_n633# 0.09fF
C2272 a_1708_n100# a_658_n100# 0.01fF
C2273 a_n1348_n633# a_n2490_n633# 0.01fF
C2274 a_n1862_n100# a_n3332_n100# 0.00fF
C2275 a_962_n633# a_960_n100# 0.00fF
C2276 a_702_n197# a_n768_131# 0.00fF
C2277 a_n928_n633# a_n1650_n633# 0.01fF
C2278 a_n976_n730# a_n1396_n730# 0.01fF
C2279 a_n1020_n633# a_n1558_n633# 0.01fF
C2280 a_n1138_n633# a_n1440_n633# 0.02fF
C2281 a_3062_n633# a_2852_n633# 0.03fF
C2282 a_3270_n100# a_1708_n100# 0.00fF
C2283 a_4110_n100# a_2758_n100# 0.00fF
C2284 a_n1560_n100# a_n2282_n100# 0.01fF
C2285 a_2012_n633# a_752_n633# 0.00fF
C2286 a_n600_n633# a_n1230_n633# 0.01fF
C2287 a_n1768_n633# a_n2070_n633# 0.02fF
C2288 a_n1860_n633# a_n1978_n633# 0.07fF
C2289 a_3432_131# w_n4520_n852# 0.12fF
C2290 a_3480_n100# a_2968_n100# 0.01fF
C2291 a_n88_n633# a_n298_n633# 0.03fF
C2292 a_1170_n100# a_540_n100# 0.01fF
C2293 a_3390_n633# a_3388_n100# 0.00fF
C2294 a_n1862_n100# a_n3450_n100# 0.00fF
C2295 a_n136_n730# a_n138_n197# 0.01fF
C2296 a_n2070_n633# a_n2026_n401# 0.00fF
C2297 a_n976_n730# a_n1816_n730# 0.01fF
C2298 a_n1020_n633# a_n1650_n633# 0.01fF
C2299 a_3180_n633# a_2642_n633# 0.01fF
C2300 a_3062_n633# a_2760_n633# 0.02fF
C2301 a_2760_n633# a_2758_n100# 0.00fF
C2302 a_4018_n100# a_3270_n100# 0.01fF
C2303 a_n718_n633# a_n1230_n633# 0.01fF
C2304 a_1920_n633# a_752_n633# 0.01fF
C2305 a_4110_n100# a_2640_n100# 0.00fF
C2306 a_n978_n197# a_n768_131# 0.01fF
C2307 a_n1768_n633# a_n2188_n633# 0.02fF
C2308 a_1380_n100# w_n4520_n852# 0.02fF
C2309 a_n1020_n633# a_n2608_n633# 0.00fF
C2310 a_3270_n100# a_3060_n100# 0.03fF
C2311 a_3388_n100# a_2968_n100# 0.02fF
C2312 a_3600_n633# w_n4520_n852# 0.04fF
C2313 a_n88_n633# a_n390_n633# 0.02fF
C2314 a_n2190_n100# a_n2282_n100# 0.09fF
C2315 a_n180_n633# a_n298_n633# 0.07fF
C2316 a_660_n633# a_542_n633# 0.07fF
C2317 a_n3030_n100# a_n3078_n197# 0.00fF
C2318 a_1078_n100# w_n4520_n852# 0.02fF
C2319 a_n3286_n401# a_n3240_n100# 0.00fF
C2320 a_n3540_n633# a_n3496_n730# 0.00fF
C2321 a_n3916_n730# a_n2446_n401# 0.00fF
C2322 a_n976_n730# a_n2236_n730# 0.00fF
C2323 a_n1396_n730# a_n1816_n730# 0.01fF
C2324 a_n3496_n730# w_n4520_n852# 0.12fF
C2325 a_n810_n633# a_n1230_n633# 0.02fF
C2326 a_4110_n100# a_2548_n100# 0.00fF
C2327 a_1802_n633# a_752_n633# 0.01fF
C2328 a_n978_n197# a_n1188_131# 0.01fF
C2329 a_n1398_n197# a_n768_131# 0.00fF
C2330 a_4020_n633# a_2432_n633# 0.00fF
C2331 a_n1768_n633# a_n2280_n633# 0.01fF
C2332 a_n4170_n633# a_n4128_131# 0.00fF
C2333 a_n2608_n633# a_n4170_n633# 0.00fF
C2334 a_n180_n633# a_n390_n633# 0.03fF
C2335 a_n138_n197# a_72_131# 0.01fF
C2336 a_660_n633# a_450_n633# 0.03fF
C2337 a_752_n633# a_332_n633# 0.02fF
C2338 a_n3122_n100# a_n3078_n197# 0.00fF
C2339 a_2174_n401# a_2220_n100# 0.00fF
C2340 a_1590_n100# a_120_n100# 0.00fF
C2341 a_n88_n633# a_n1440_n633# 0.00fF
C2342 a_30_n633# a_n1558_n633# 0.00fF
C2343 a_n3916_n730# a_n2866_n401# 0.00fF
C2344 a_n1396_n730# a_n2236_n730# 0.01fF
C2345 a_1800_n100# a_1590_n100# 0.03fF
C2346 a_n2282_n100# a_n2492_n100# 0.03fF
C2347 a_1800_n100# a_1752_131# 0.00fF
C2348 a_n1232_n100# a_n1442_n100# 0.03fF
C2349 a_1710_n633# a_752_n633# 0.01fF
C2350 a_n928_n633# a_n1230_n633# 0.02fF
C2351 a_n1818_n197# a_n768_131# 0.00fF
C2352 a_3902_n633# a_2432_n633# 0.00fF
C2353 a_n1768_n633# a_n2398_n633# 0.01fF
C2354 a_n1398_n197# a_n1188_131# 0.01fF
C2355 a_n2700_n633# a_n4170_n633# 0.00fF
C2356 a_n298_n633# a_n390_n633# 0.09fF
C2357 a_752_n633# a_240_n633# 0.01fF
C2358 a_870_n633# a_122_n633# 0.01fF
C2359 a_n1232_n100# a_n1350_n100# 0.07fF
C2360 a_n2400_n100# a_n2702_n100# 0.02fF
C2361 a_1124_n730# a_1334_n401# 0.01fF
C2362 a_n3868_n633# a_n3960_n633# 0.09fF
C2363 a_n180_n633# a_n1440_n633# 0.00fF
C2364 a_n1816_n730# a_n2236_n730# 0.01fF
C2365 a_n1396_n730# a_n2656_n730# 0.00fF
C2366 a_1708_n100# a_1590_n100# 0.07fF
C2367 a_3642_n197# a_3852_131# 0.01fF
C2368 a_1708_n100# a_1752_131# 0.00fF
C2369 a_n1020_n633# a_n1230_n633# 0.03fF
C2370 a_n2238_n197# a_n768_131# 0.00fF
C2371 a_n1768_n633# a_n2490_n633# 0.01fF
C2372 a_n1818_n197# a_n1188_131# 0.00fF
C2373 a_3810_n633# a_2432_n633# 0.00fF
C2374 a_3902_n633# a_2340_n633# 0.00fF
C2375 a_1124_n730# a_494_n401# 0.00fF
C2376 a_n2818_n633# a_n4170_n633# 0.00fF
C2377 a_n2400_n100# a_n2820_n100# 0.02fF
C2378 a_870_n633# a_30_n633# 0.01fF
C2379 a_704_n730# a_1334_n401# 0.00fF
C2380 a_3272_n633# a_3270_n100# 0.00fF
C2381 a_n298_n633# a_n1440_n633# 0.01fF
C2382 a_n2398_n633# a_n2446_n401# 0.00fF
C2383 a_n1816_n730# a_n2656_n730# 0.01fF
C2384 a_3642_n197# a_3432_131# 0.01fF
C2385 a_3482_n633# a_3434_n401# 0.00fF
C2386 a_3060_n100# a_1590_n100# 0.00fF
C2387 a_3810_n633# a_2340_n633# 0.00fF
C2388 a_3692_n633# a_2432_n633# 0.00fF
C2389 a_3600_n633# a_2550_n633# 0.01fF
C2390 a_n2238_n197# a_n1188_131# 0.00fF
C2391 a_704_n730# a_494_n401# 0.01fF
C2392 a_3598_n100# w_n4520_n852# 0.04fF
C2393 a_1124_n730# a_74_n401# 0.00fF
C2394 a_n2910_n633# a_n4170_n633# 0.00fF
C2395 a_n2400_n100# a_n2912_n100# 0.01fF
C2396 a_284_n730# a_1334_n401# 0.00fF
C2397 a_n390_n633# a_n1440_n633# 0.01fF
C2398 a_n2490_n633# a_n2446_n401# 0.00fF
C2399 a_n2236_n730# a_n2656_n730# 0.01fF
C2400 a_1542_n197# a_2592_131# 0.00fF
C2401 a_n348_131# w_n4520_n852# 0.12fF
C2402 a_122_n633# a_n1230_n633# 0.00fF
C2403 a_3600_n633# a_3642_n197# 0.00fF
C2404 a_3390_n633# a_3434_n401# 0.00fF
C2405 a_n2658_n197# a_n1188_131# 0.00fF
C2406 a_3692_n633# a_2340_n633# 0.00fF
C2407 a_n1980_n100# a_n2282_n100# 0.02fF
C2408 a_1592_n633# a_1080_n633# 0.01fF
C2409 a_1124_n730# a_n346_n401# 0.00fF
C2410 a_284_n730# a_494_n401# 0.01fF
C2411 a_704_n730# a_74_n401# 0.00fF
C2412 a_3480_n100# w_n4520_n852# 0.04fF
C2413 a_n3028_n633# a_n4170_n633# 0.01fF
C2414 a_n2400_n100# a_n3030_n100# 0.01fF
C2415 a_n2070_n633# a_n3330_n633# 0.00fF
C2416 a_n3450_n100# a_n3498_n197# 0.00fF
C2417 a_n136_n730# a_1334_n401# 0.00fF
C2418 a_492_131# w_n4520_n852# 0.12fF
C2419 a_n3706_n401# a_n3660_n100# 0.00fF
C2420 a_n812_n100# a_n2400_n100# 0.00fF
C2421 a_3014_n401# a_3060_n100# 0.00fF
C2422 a_n1440_n633# a_n1442_n100# 0.00fF
C2423 a_30_n633# a_n1230_n633# 0.00fF
C2424 a_n1350_n100# a_n1442_n100# 0.09fF
C2425 a_1500_n633# a_1080_n633# 0.02fF
C2426 a_1122_n197# a_1332_131# 0.01fF
C2427 a_n136_n730# a_494_n401# 0.00fF
C2428 a_3388_n100# w_n4520_n852# 0.03fF
C2429 a_704_n730# a_n346_n401# 0.00fF
C2430 a_284_n730# a_74_n401# 0.01fF
C2431 a_540_n100# w_n4520_n852# 0.02fF
C2432 a_n3120_n633# a_n4170_n633# 0.01fF
C2433 a_n2400_n100# a_n3122_n100# 0.01fF
C2434 a_120_n100# a_n1232_n100# 0.00fF
C2435 a_n508_n633# w_n4520_n852# 0.01fF
C2436 a_n2070_n633# a_n3448_n633# 0.00fF
C2437 a_n2188_n633# a_n3330_n633# 0.01fF
C2438 a_n3542_n100# a_n3498_n197# 0.00fF
C2439 a_1592_n633# a_1544_n730# 0.00fF
C2440 a_n930_n100# a_n2400_n100# 0.00fF
C2441 a_n3916_n730# a_n4126_n401# 0.01fF
C2442 a_n3870_n100# a_n4080_n100# 0.03fF
C2443 a_4018_n100# a_3900_n100# 0.07fF
C2444 a_2222_n633# a_1592_n633# 0.01fF
C2445 a_n3870_n100# a_n3962_n100# 0.09fF
C2446 a_1382_n633# a_1080_n633# 0.02fF
C2447 a_3900_n100# a_3060_n100# 0.01fF
C2448 a_n556_n730# a_494_n401# 0.00fF
C2449 a_704_n730# a_n766_n401# 0.00fF
C2450 a_284_n730# a_n346_n401# 0.00fF
C2451 a_n136_n730# a_74_n401# 0.01fF
C2452 a_n3330_n633# a_n4078_n633# 0.01fF
C2453 a_n3238_n633# a_n4170_n633# 0.01fF
C2454 a_n2400_n100# a_n3240_n100# 0.01fF
C2455 a_n600_n633# w_n4520_n852# 0.01fF
C2456 a_n2188_n633# a_n3448_n633# 0.00fF
C2457 a_n3960_n633# a_n3918_n197# 0.00fF
C2458 a_n2280_n633# a_n3330_n633# 0.01fF
C2459 a_3482_n633# a_3062_n633# 0.02fF
C2460 a_1500_n633# a_1544_n730# 0.00fF
C2461 a_n1140_n100# a_n2282_n100# 0.01fF
C2462 a_4018_n100# a_3808_n100# 0.03fF
C2463 a_1332_131# a_912_131# 0.01fF
C2464 a_2130_n633# a_1592_n633# 0.01fF
C2465 a_2222_n633# a_1500_n633# 0.01fF
C2466 a_2382_n197# a_1122_n197# 0.00fF
C2467 a_2968_n100# a_2850_n100# 0.07fF
C2468 a_3808_n100# a_3060_n100# 0.01fF
C2469 a_1290_n633# a_1080_n633# 0.03fF
C2470 a_n136_n730# a_n346_n401# 0.01fF
C2471 a_284_n730# a_n766_n401# 0.00fF
C2472 a_n556_n730# a_74_n401# 0.00fF
C2473 a_n3448_n633# a_n4078_n633# 0.01fF
C2474 a_2758_n100# a_1170_n100# 0.00fF
C2475 a_n2400_n100# a_n3332_n100# 0.01fF
C2476 a_n718_n633# w_n4520_n852# 0.01fF
C2477 a_n2398_n633# a_n3330_n633# 0.01fF
C2478 a_n2280_n633# a_n3448_n633# 0.01fF
C2479 a_3390_n633# a_3062_n633# 0.02fF
C2480 a_870_n633# a_868_n100# 0.00fF
C2481 a_n4078_n633# a_n4126_n401# 0.00fF
C2482 a_74_n401# a_72_131# 0.01fF
C2483 a_2012_n633# a_1592_n633# 0.02fF
C2484 a_3598_n100# a_3642_n197# 0.00fF
C2485 a_2222_n633# a_1382_n633# 0.01fF
C2486 a_2130_n633# a_1500_n633# 0.01fF
C2487 a_2802_n197# a_3012_131# 0.01fF
C2488 a_1962_n197# a_1122_n197# 0.01fF
C2489 a_2968_n100# a_2758_n100# 0.03fF
C2490 a_1172_n633# a_1080_n633# 0.09fF
C2491 a_n136_n730# a_n766_n401# 0.00fF
C2492 a_n556_n730# a_n346_n401# 0.01fF
C2493 a_284_n730# a_n1186_n401# 0.00fF
C2494 a_4110_n100# a_3178_n100# 0.01fF
C2495 a_n2400_n100# a_n3450_n100# 0.01fF
C2496 a_2640_n100# a_1170_n100# 0.00fF
C2497 a_n3708_131# w_n4520_n852# 0.13fF
C2498 a_n810_n633# w_n4520_n852# 0.01fF
C2499 a_2432_n633# a_2384_n730# 0.00fF
C2500 a_n2398_n633# a_n3448_n633# 0.01fF
C2501 a_n2490_n633# a_n3330_n633# 0.01fF
C2502 a_2384_n730# a_2382_n197# 0.01fF
C2503 a_2382_n197# a_912_131# 0.00fF
C2504 a_1288_n100# a_1170_n100# 0.07fF
C2505 a_2222_n633# a_1290_n633# 0.01fF
C2506 a_2432_n633# a_1080_n633# 0.00fF
C2507 a_2130_n633# a_1382_n633# 0.01fF
C2508 a_2012_n633# a_1500_n633# 0.01fF
C2509 a_1920_n633# a_1592_n633# 0.02fF
C2510 a_120_n100# a_n1442_n100# 0.00fF
C2511 a_752_n633# a_704_n730# 0.00fF
C2512 a_2968_n100# a_2640_n100# 0.02fF
C2513 a_n136_n730# a_n1186_n401# 0.00fF
C2514 a_n556_n730# a_n766_n401# 0.01fF
C2515 a_n2400_n100# a_n3542_n100# 0.01fF
C2516 a_2548_n100# a_1170_n100# 0.00fF
C2517 a_120_n100# a_n1350_n100# 0.00fF
C2518 a_2802_n197# a_1332_131# 0.00fF
C2519 a_n928_n633# w_n4520_n852# 0.01fF
C2520 a_2340_n633# a_2384_n730# 0.00fF
C2521 a_n2490_n633# a_n3448_n633# 0.01fF
C2522 a_702_n197# a_n348_131# 0.00fF
C2523 a_3854_n401# w_n4520_n852# 0.09fF
C2524 a_1962_n197# a_912_131# 0.00fF
C2525 a_2222_n633# a_1172_n633# 0.01fF
C2526 a_n180_n633# a_n138_n197# 0.00fF
C2527 a_1802_n633# a_1592_n633# 0.03fF
C2528 a_1920_n633# a_1500_n633# 0.02fF
C2529 a_2340_n633# a_1080_n633# 0.00fF
C2530 a_2130_n633# a_1290_n633# 0.01fF
C2531 a_2012_n633# a_1382_n633# 0.01fF
C2532 a_n3496_n730# a_n3286_n401# 0.01fF
C2533 a_n2868_131# a_n4128_131# 0.00fF
C2534 a_2968_n100# a_2548_n100# 0.02fF
C2535 a_n556_n730# a_n1186_n401# 0.00fF
C2536 a_n136_n730# a_n1606_n401# 0.00fF
C2537 a_1592_n633# a_332_n633# 0.00fF
C2538 a_702_n197# a_492_131# 0.01fF
C2539 a_n2400_n100# a_n3660_n100# 0.00fF
C2540 a_2430_n100# a_1170_n100# 0.00fF
C2541 a_n1020_n633# w_n4520_n852# 0.01fF
C2542 a_3434_n401# w_n4520_n852# 0.09fF
C2543 a_1964_n730# a_1962_n197# 0.01fF
C2544 a_1498_n100# a_28_n100# 0.00fF
C2545 a_n2282_n100# w_n4520_n852# 0.02fF
C2546 a_2432_n633# a_2222_n633# 0.03fF
C2547 a_n978_n197# a_n348_131# 0.00fF
C2548 a_n3658_n633# a_n4170_n633# 0.01fF
C2549 a_1920_n633# a_1382_n633# 0.01fF
C2550 a_1710_n633# a_1592_n633# 0.07fF
C2551 a_2012_n633# a_1290_n633# 0.01fF
C2552 a_1802_n633# a_1500_n633# 0.02fF
C2553 a_2130_n633# a_1172_n633# 0.01fF
C2554 a_n3496_n730# a_n3706_n401# 0.01fF
C2555 a_n556_n730# a_n558_n197# 0.01fF
C2556 a_n3288_131# a_n4128_131# 0.01fF
C2557 a_2968_n100# a_2430_n100# 0.01fF
C2558 a_n556_n730# a_n1606_n401# 0.00fF
C2559 a_1500_n633# a_332_n633# 0.01fF
C2560 a_1592_n633# a_240_n633# 0.00fF
C2561 a_2802_n197# a_2382_n197# 0.01fF
C2562 a_n3540_n633# a_n4170_n633# 0.01fF
C2563 a_2338_n100# a_1170_n100# 0.01fF
C2564 a_4112_n633# a_3600_n633# 0.01fF
C2565 a_n4170_n633# w_n4520_n852# 0.14fF
C2566 a_3272_n633# a_2970_n633# 0.02fF
C2567 a_n558_n197# a_72_131# 0.00fF
C2568 a_962_n633# a_n88_n633# 0.01fF
C2569 a_n978_n197# a_492_131# 0.00fF
C2570 a_1170_n100# a_868_n100# 0.02fF
C2571 a_1498_n100# a_n90_n100# 0.00fF
C2572 a_3222_n197# a_2802_n197# 0.01fF
C2573 a_2340_n633# a_2222_n633# 0.07fF
C2574 a_2432_n633# a_2130_n633# 0.02fF
C2575 a_n1398_n197# a_n348_131# 0.00fF
C2576 a_1802_n633# a_1382_n633# 0.02fF
C2577 a_1710_n633# a_1500_n633# 0.03fF
C2578 a_2012_n633# a_1172_n633# 0.01fF
C2579 a_1920_n633# a_1290_n633# 0.01fF
C2580 a_2968_n100# a_2338_n100# 0.01fF
C2581 a_n556_n730# a_n2026_n401# 0.00fF
C2582 a_122_n633# w_n4520_n852# 0.01fF
C2583 a_1382_n633# a_332_n633# 0.01fF
C2584 a_2802_n197# a_1962_n197# 0.01fF
C2585 a_1500_n633# a_240_n633# 0.00fF
C2586 a_3810_n633# a_3852_131# 0.00fF
C2587 a_2220_n100# a_1170_n100# 0.01fF
C2588 a_4020_n633# a_3600_n633# 0.02fF
C2589 a_448_n100# a_n1022_n100# 0.00fF
C2590 a_330_n100# a_282_n197# 0.00fF
C2591 a_962_n633# a_n180_n633# 0.01fF
C2592 a_1170_n100# a_750_n100# 0.02fF
C2593 a_2340_n633# a_2130_n633# 0.03fF
C2594 a_n508_n633# a_n1860_n633# 0.00fF
C2595 a_2432_n633# a_2012_n633# 0.02fF
C2596 a_n3496_n730# a_n3498_n197# 0.01fF
C2597 a_n1818_n197# a_n348_131# 0.00fF
C2598 a_1710_n633# a_1382_n633# 0.02fF
C2599 a_1802_n633# a_1290_n633# 0.01fF
C2600 a_1920_n633# a_1172_n633# 0.01fF
C2601 a_3180_n633# a_1592_n633# 0.00fF
C2602 a_2968_n100# a_2220_n100# 0.01fF
C2603 a_2850_n100# w_n4520_n852# 0.03fF
C2604 a_2594_n401# a_1334_n401# 0.00fF
C2605 a_2174_n401# a_1754_n401# 0.01fF
C2606 a_n2910_n633# a_n2868_131# 0.00fF
C2607 a_n1138_n633# a_n1348_n633# 0.03fF
C2608 a_1080_n633# a_542_n633# 0.01fF
C2609 a_30_n633# w_n4520_n852# 0.01fF
C2610 a_1290_n633# a_332_n633# 0.01fF
C2611 a_1382_n633# a_240_n633# 0.01fF
C2612 a_2128_n100# a_1170_n100# 0.01fF
C2613 a_3902_n633# a_3600_n633# 0.02fF
C2614 a_660_n633# a_n508_n633# 0.01fF
C2615 a_n2610_n100# a_n4080_n100# 0.00fF
C2616 a_238_n100# a_282_n197# 0.00fF
C2617 a_962_n633# a_n298_n633# 0.00fF
C2618 a_n2610_n100# a_n3962_n100# 0.00fF
C2619 a_2340_n633# a_2012_n633# 0.02fF
C2620 a_n600_n633# a_n1860_n633# 0.00fF
C2621 a_2432_n633# a_1920_n633# 0.01fF
C2622 a_1710_n633# a_1290_n633# 0.02fF
C2623 a_1802_n633# a_1172_n633# 0.01fF
C2624 a_3062_n633# w_n4520_n852# 0.03fF
C2625 a_1170_n100# a_330_n100# 0.01fF
C2626 a_2758_n100# w_n4520_n852# 0.02fF
C2627 a_2968_n100# a_2128_n100# 0.01fF
C2628 a_1500_n633# a_1498_n100# 0.00fF
C2629 a_1290_n633# a_240_n633# 0.01fF
C2630 a_1172_n633# a_332_n633# 0.01fF
C2631 a_1080_n633# a_450_n633# 0.01fF
C2632 a_2010_n100# a_1170_n100# 0.01fF
C2633 a_3810_n633# a_3600_n633# 0.03fF
C2634 a_660_n633# a_n600_n633# 0.00fF
C2635 a_n2236_n730# a_n2190_n100# 0.00fF
C2636 a_962_n633# a_n390_n633# 0.00fF
C2637 a_1708_n100# a_120_n100# 0.00fF
C2638 a_2340_n633# a_1920_n633# 0.02fF
C2639 a_n718_n633# a_n1860_n633# 0.01fF
C2640 a_1800_n100# a_1708_n100# 0.09fF
C2641 a_2432_n633# a_1802_n633# 0.01fF
C2642 a_1170_n100# a_238_n100# 0.01fF
C2643 a_1710_n633# a_1172_n633# 0.01fF
C2644 a_2968_n100# a_2010_n100# 0.01fF
C2645 a_2640_n100# w_n4520_n852# 0.02fF
C2646 a_960_n100# a_28_n100# 0.01fF
C2647 a_1172_n633# a_240_n633# 0.01fF
C2648 a_1920_n633# a_1962_n197# 0.00fF
C2649 a_2592_131# a_1752_131# 0.01fF
C2650 a_1918_n100# a_1170_n100# 0.01fF
C2651 a_3692_n633# a_3600_n633# 0.09fF
C2652 a_660_n633# a_n718_n633# 0.00fF
C2653 a_2642_n633# a_2594_n401# 0.00fF
C2654 a_2592_131# a_2172_131# 0.01fF
C2655 a_1288_n100# w_n4520_n852# 0.02fF
C2656 a_n2608_n633# a_n2656_n730# 0.00fF
C2657 a_n1560_n100# a_n2072_n100# 0.01fF
C2658 a_n810_n633# a_n1860_n633# 0.01fF
C2659 a_2340_n633# a_1802_n633# 0.01fF
C2660 a_2432_n633# a_1710_n633# 0.01fF
C2661 a_n88_n633# a_n1348_n633# 0.00fF
C2662 a_2968_n100# a_1918_n100# 0.01fF
C2663 a_3060_n100# a_1800_n100# 0.00fF
C2664 a_2548_n100# w_n4520_n852# 0.02fF
C2665 a_2130_n633# a_542_n633# 0.00fF
C2666 a_960_n100# a_n90_n100# 0.01fF
C2667 a_4064_n730# a_4062_n197# 0.01fF
C2668 a_660_n633# a_n810_n633# 0.00fF
C2669 a_n1138_n633# a_n1186_n401# 0.00fF
C2670 a_330_n100# a_n1140_n100# 0.00fF
C2671 a_n2700_n633# a_n2656_n730# 0.00fF
C2672 a_1500_n633# a_1542_n197# 0.00fF
C2673 a_n928_n633# a_n1860_n633# 0.01fF
C2674 a_2340_n633# a_1710_n633# 0.01fF
C2675 a_n180_n633# a_n1348_n633# 0.01fF
C2676 a_n2072_n100# a_n2190_n100# 0.07fF
C2677 a_3060_n100# a_1708_n100# 0.00fF
C2678 a_2430_n100# w_n4520_n852# 0.02fF
C2679 a_2012_n633# a_542_n633# 0.00fF
C2680 a_n1770_n100# a_n2282_n100# 0.01fF
C2681 a_960_n100# a_n182_n100# 0.01fF
C2682 a_n1978_n633# a_n2070_n633# 0.09fF
C2683 a_n1020_n633# a_n978_n197# 0.00fF
C2684 a_660_n633# a_n928_n633# 0.00fF
C2685 a_448_n100# a_28_n100# 0.02fF
C2686 a_238_n100# a_n1140_n100# 0.00fF
C2687 a_2594_n401# a_2592_131# 0.01fF
C2688 a_1542_n197# a_3012_131# 0.00fF
C2689 a_n1138_n633# a_n1768_n633# 0.01fF
C2690 a_n1020_n633# a_n1860_n633# 0.01fF
C2691 a_3180_n633# a_2432_n633# 0.01fF
C2692 a_2852_n633# a_2760_n633# 0.09fF
C2693 a_3062_n633# a_2550_n633# 0.01fF
C2694 a_2970_n633# a_2642_n633# 0.02fF
C2695 a_n298_n633# a_n1348_n633# 0.01fF
C2696 a_4018_n100# a_3060_n100# 0.01fF
C2697 a_2338_n100# w_n4520_n852# 0.02fF
C2698 a_1920_n633# a_542_n633# 0.00fF
C2699 a_960_n100# a_n300_n100# 0.00fF
C2700 a_2012_n633# a_450_n633# 0.00fF
C2701 a_n1862_n100# a_n2282_n100# 0.02fF
C2702 a_n1978_n633# a_n2188_n633# 0.03fF
C2703 a_3178_n100# a_2968_n100# 0.03fF
C2704 a_n2028_131# a_n2448_131# 0.01fF
C2705 a_n2238_n197# a_n3708_131# 0.00fF
C2706 a_448_n100# a_n90_n100# 0.01fF
C2707 a_868_n100# w_n4520_n852# 0.02fF
C2708 a_n2072_n100# a_n2492_n100# 0.02fF
C2709 a_3180_n633# a_3222_n197# 0.00fF
C2710 a_3180_n633# a_2340_n633# 0.01fF
C2711 a_n3960_n633# a_n3916_n730# 0.00fF
C2712 a_n390_n633# a_n1348_n633# 0.01fF
C2713 a_2220_n100# w_n4520_n852# 0.02fF
C2714 a_1802_n633# a_542_n633# 0.00fF
C2715 a_960_n100# a_n392_n100# 0.00fF
C2716 a_1920_n633# a_450_n633# 0.00fF
C2717 a_1078_n100# a_1122_n197# 0.00fF
C2718 a_n3076_n730# a_n1606_n401# 0.00fF
C2719 a_1542_n197# a_1332_131# 0.01fF
C2720 a_n1978_n633# a_n2280_n633# 0.02fF
C2721 a_542_n633# a_332_n633# 0.03fF
C2722 a_n2658_n197# a_n3708_131# 0.00fF
C2723 a_n298_n633# a_n346_n401# 0.00fF
C2724 a_n3706_n401# a_n3708_131# 0.01fF
C2725 a_448_n100# a_n182_n100# 0.01fF
C2726 a_750_n100# w_n4520_n852# 0.02fF
C2727 a_n4126_n401# a_n4080_n100# 0.00fF
C2728 a_n136_n730# a_n90_n100# 0.00fF
C2729 a_n3752_n100# a_n4080_n100# 0.02fF
C2730 a_2550_n633# a_2548_n100# 0.00fF
C2731 a_n3752_n100# a_n3962_n100# 0.03fF
C2732 a_2128_n100# w_n4520_n852# 0.02fF
C2733 a_n1232_n100# a_n1652_n100# 0.02fF
C2734 a_960_n100# a_n510_n100# 0.00fF
C2735 a_1802_n633# a_450_n633# 0.00fF
C2736 a_1710_n633# a_542_n633# 0.01fF
C2737 a_n3076_n730# a_n2026_n401# 0.00fF
C2738 a_n1978_n633# a_n2398_n633# 0.02fF
C2739 a_658_n100# a_28_n100# 0.01fF
C2740 a_28_n100# a_72_131# 0.00fF
C2741 a_450_n633# a_332_n633# 0.07fF
C2742 a_542_n633# a_240_n633# 0.02fF
C2743 a_660_n633# a_122_n633# 0.01fF
C2744 a_n3078_n197# a_n3708_131# 0.00fF
C2745 a_n1348_n633# a_n1440_n633# 0.09fF
C2746 a_n390_n633# a_n346_n401# 0.00fF
C2747 a_448_n100# a_n300_n100# 0.01fF
C2748 a_n1348_n633# a_n1350_n100# 0.00fF
C2749 a_n3868_n633# a_n4170_n633# 0.02fF
C2750 a_n3960_n633# a_n4078_n633# 0.07fF
C2751 a_330_n100# w_n4520_n852# 0.02fF
C2752 a_n2282_n100# a_n2238_n197# 0.00fF
C2753 a_2802_n197# a_3852_131# 0.00fF
C2754 a_2382_n197# a_1542_n197# 0.01fF
C2755 a_2010_n100# w_n4520_n852# 0.02fF
C2756 a_960_n100# a_n602_n100# 0.00fF
C2757 a_1710_n633# a_450_n633# 0.00fF
C2758 a_658_n100# a_n90_n100# 0.01fF
C2759 a_n1978_n633# a_n2490_n633# 0.01fF
C2760 a_n3076_n730# a_n2446_n401# 0.00fF
C2761 a_660_n633# a_30_n633# 0.01fF
C2762 a_450_n633# a_240_n633# 0.03fF
C2763 a_752_n633# a_n88_n633# 0.01fF
C2764 a_n2868_131# w_n4520_n852# 0.12fF
C2765 a_n3498_n197# a_n3708_131# 0.01fF
C2766 a_448_n100# a_n392_n100# 0.01fF
C2767 a_1080_n633# a_1078_n100# 0.00fF
C2768 a_n180_n633# a_n1768_n633# 0.00fF
C2769 a_238_n100# w_n4520_n852# 0.02fF
C2770 a_n1980_n100# a_n2072_n100# 0.09fF
C2771 a_n2398_n633# a_n3960_n633# 0.00fF
C2772 a_2802_n197# a_3432_131# 0.00fF
C2773 a_1962_n197# a_1542_n197# 0.01fF
C2774 a_1172_n633# a_1124_n730# 0.00fF
C2775 a_1918_n100# w_n4520_n852# 0.02fF
C2776 a_658_n100# a_n182_n100# 0.01fF
C2777 a_n3076_n730# a_n2866_n401# 0.01fF
C2778 a_752_n633# a_n180_n633# 0.01fF
C2779 a_3224_n730# a_3222_n197# 0.01fF
C2780 a_n3288_131# w_n4520_n852# 0.13fF
C2781 a_n3918_n197# a_n3708_131# 0.01fF
C2782 a_448_n100# a_n510_n100# 0.01fF
C2783 a_n298_n633# a_n1768_n633# 0.00fF
C2784 a_n1232_n100# a_n2610_n100# 0.00fF
C2785 a_n2490_n633# a_n3960_n633# 0.00fF
C2786 a_n976_n730# w_n4520_n852# 0.12fF
C2787 a_658_n100# a_n300_n100# 0.01fF
C2788 a_3600_n633# a_2222_n633# 0.00fF
C2789 a_752_n633# a_n298_n633# 0.01fF
C2790 a_448_n100# a_n602_n100# 0.01fF
C2791 a_1122_n197# a_n348_131# 0.00fF
C2792 a_n390_n633# a_n1768_n633# 0.00fF
C2793 a_n1442_n100# a_n1652_n100# 0.03fF
C2794 a_3902_n633# a_3854_n401# 0.00fF
C2795 a_n4172_n100# a_n4128_131# 0.00fF
C2796 a_n1558_n633# a_n1560_n100# 0.00fF
C2797 a_n1396_n730# w_n4520_n852# 0.12fF
C2798 a_n1350_n100# a_n1652_n100# 0.02fF
C2799 a_658_n100# a_n392_n100# 0.01fF
C2800 a_3600_n633# a_2130_n633# 0.00fF
C2801 a_1122_n197# a_492_131# 0.00fF
C2802 a_3178_n100# w_n4520_n852# 0.03fF
C2803 a_n1140_n100# a_n2072_n100# 0.01fF
C2804 a_752_n633# a_n390_n633# 0.01fF
C2805 a_448_n100# a_n720_n100# 0.01fF
C2806 a_n1022_n100# a_n1232_n100# 0.03fF
C2807 a_n556_n730# a_n510_n100# 0.00fF
C2808 a_1590_n100# a_28_n100# 0.00fF
C2809 a_3810_n633# a_3854_n401# 0.00fF
C2810 a_n2702_n100# a_n4080_n100# 0.00fF
C2811 a_n1560_n100# a_n2190_n100# 0.01fF
C2812 a_74_n401# a_120_n100# 0.00fF
C2813 a_n1816_n730# w_n4520_n852# 0.12fF
C2814 a_n2702_n100# a_n3962_n100# 0.00fF
C2815 a_3600_n633# a_2012_n633# 0.00fF
C2816 a_n1558_n633# a_n1650_n633# 0.09fF
C2817 a_n1440_n633# a_n1768_n633# 0.02fF
C2818 a_658_n100# a_n510_n100# 0.01fF
C2819 a_750_n100# a_702_n197# 0.00fF
C2820 a_912_131# a_n348_131# 0.00fF
C2821 a_448_n100# a_n812_n100# 0.00fF
C2822 a_n1558_n633# a_n2608_n633# 0.01fF
C2823 a_3482_n633# a_2852_n633# 0.01fF
C2824 a_n2820_n100# a_n4080_n100# 0.00fF
C2825 a_912_131# a_492_131# 0.01fF
C2826 a_1332_131# a_72_131# 0.00fF
C2827 a_n2236_n730# w_n4520_n852# 0.12fF
C2828 a_n2820_n100# a_n3962_n100# 0.01fF
C2829 a_4112_n633# a_3062_n633# 0.01fF
C2830 a_658_n100# a_n602_n100# 0.00fF
C2831 a_448_n100# a_n930_n100# 0.00fF
C2832 a_n2446_n401# a_n2448_131# 0.01fF
C2833 a_n3496_n730# a_n3916_n730# 0.01fF
C2834 a_n1650_n633# a_n2608_n633# 0.01fF
C2835 a_n1558_n633# a_n2700_n633# 0.01fF
C2836 a_3482_n633# a_2760_n633# 0.01fF
C2837 a_3390_n633# a_2852_n633# 0.01fF
C2838 a_n1560_n100# a_n2492_n100# 0.01fF
C2839 a_n1442_n100# a_n2610_n100# 0.01fF
C2840 a_n2912_n100# a_n4080_n100# 0.01fF
C2841 a_n1350_n100# a_n2610_n100# 0.00fF
C2842 a_n2656_n730# w_n4520_n852# 0.12fF
C2843 a_n2912_n100# a_n3962_n100# 0.01fF
C2844 a_1592_n633# a_1590_n100# 0.00fF
C2845 a_4020_n633# a_3062_n633# 0.01fF
C2846 a_658_n100# a_n720_n100# 0.00fF
C2847 a_n3076_n730# a_n4126_n401# 0.00fF
C2848 a_4110_n100# a_2968_n100# 0.01fF
C2849 a_1080_n633# a_n508_n633# 0.00fF
C2850 a_n1650_n633# a_n2700_n633# 0.01fF
C2851 a_n1558_n633# a_n2818_n633# 0.00fF
C2852 a_3390_n633# a_2760_n633# 0.01fF
C2853 a_n2190_n100# a_n2492_n100# 0.02fF
C2854 a_n2282_n100# a_n2400_n100# 0.07fF
C2855 a_n3030_n100# a_n4080_n100# 0.01fF
C2856 a_n2608_n633# a_n2700_n633# 0.09fF
C2857 a_n3030_n100# a_n3962_n100# 0.01fF
C2858 a_n1022_n100# a_n1442_n100# 0.02fF
C2859 a_3902_n633# a_3062_n633# 0.01fF
C2860 a_658_n100# a_n812_n100# 0.00fF
C2861 a_n1230_n633# a_n1558_n633# 0.02fF
C2862 a_n1022_n100# a_n1350_n100# 0.02fF
C2863 a_n1558_n633# a_n2910_n633# 0.00fF
C2864 a_n1650_n633# a_n2818_n633# 0.01fF
C2865 a_n2072_n100# w_n4520_n852# 0.02fF
C2866 a_4018_n100# a_4062_n197# 0.00fF
C2867 a_n3122_n100# a_n4080_n100# 0.01fF
C2868 a_n2608_n633# a_n2818_n633# 0.03fF
C2869 a_3270_n100# a_3222_n197# 0.00fF
C2870 a_n3122_n100# a_n3962_n100# 0.01fF
C2871 a_658_n100# a_n930_n100# 0.00fF
C2872 a_3810_n633# a_3062_n633# 0.01fF
C2873 a_3012_131# a_1752_131# 0.00fF
C2874 a_n1398_n197# a_n2868_131# 0.00fF
C2875 a_n1230_n633# a_n1650_n633# 0.02fF
C2876 a_28_n100# a_n1232_n100# 0.00fF
C2877 a_n1558_n633# a_n3028_n633# 0.00fF
C2878 a_n1650_n633# a_n2910_n633# 0.00fF
C2879 a_3012_131# a_2172_131# 0.01fF
C2880 a_n1230_n633# a_n2608_n633# 0.00fF
C2881 a_n3240_n100# a_n4080_n100# 0.01fF
C2882 a_n2700_n633# a_n2818_n633# 0.07fF
C2883 a_n2608_n633# a_n2910_n633# 0.02fF
C2884 a_n1560_n100# a_n1980_n100# 0.02fF
C2885 a_450_n633# a_448_n100# 0.00fF
C2886 a_n88_n633# a_n90_n100# 0.00fF
C2887 a_2804_n730# a_3854_n401# 0.00fF
C2888 a_n3240_n100# a_n3962_n100# 0.01fF
C2889 a_n976_n730# a_n978_n197# 0.01fF
C2890 a_3692_n633# a_3062_n633# 0.01fF
C2891 a_1498_n100# a_1380_n100# 0.07fF
C2892 a_3600_n633# a_3180_n633# 0.02fF
C2893 a_n1818_n197# a_n2868_131# 0.00fF
C2894 a_1498_n100# a_1078_n100# 0.02fF
C2895 a_n90_n100# a_n1232_n100# 0.01fF
C2896 a_n1558_n633# a_n3120_n633# 0.00fF
C2897 a_n1650_n633# a_n3028_n633# 0.00fF
C2898 a_1752_131# a_1332_131# 0.01fF
C2899 a_2174_n401# w_n4520_n852# 0.10fF
C2900 a_3014_n401# a_3012_131# 0.01fF
C2901 a_n1230_n633# a_n2700_n633# 0.00fF
C2902 a_n3332_n100# a_n4080_n100# 0.01fF
C2903 a_n2700_n633# a_n2910_n633# 0.03fF
C2904 a_n2608_n633# a_n3028_n633# 0.02fF
C2905 a_2172_131# a_1332_131# 0.01fF
C2906 a_n1980_n100# a_n2190_n100# 0.03fF
C2907 a_2804_n730# a_3434_n401# 0.00fF
C2908 a_2384_n730# a_3854_n401# 0.00fF
C2909 a_n3332_n100# a_n3962_n100# 0.01fF
C2910 a_n1816_n730# a_n1770_n100# 0.00fF
C2911 a_n1818_n197# a_n3288_131# 0.00fF
C2912 a_n2238_n197# a_n2868_131# 0.00fF
C2913 a_n182_n100# a_n1232_n100# 0.01fF
C2914 a_n1650_n633# a_n3120_n633# 0.00fF
C2915 a_3272_n633# a_2642_n633# 0.01fF
C2916 a_1754_n401# w_n4520_n852# 0.10fF
C2917 a_n1230_n633# a_n2818_n633# 0.00fF
C2918 a_n3450_n100# a_n4080_n100# 0.01fF
C2919 a_n2700_n633# a_n3028_n633# 0.02fF
C2920 a_n2818_n633# a_n2910_n633# 0.09fF
C2921 a_n2608_n633# a_n3120_n633# 0.01fF
C2922 a_n508_n633# a_n2070_n633# 0.00fF
C2923 a_n180_n633# a_n182_n100# 0.00fF
C2924 a_2384_n730# a_3434_n401# 0.00fF
C2925 a_n3450_n100# a_n3962_n100# 0.01fF
C2926 a_n1396_n730# a_n1398_n197# 0.01fF
C2927 a_2970_n633# a_1592_n633# 0.00fF
C2928 a_2174_n401# a_914_n401# 0.00fF
C2929 a_n1140_n100# a_n1560_n100# 0.02fF
C2930 a_n1608_131# a_n2448_131# 0.01fF
C2931 a_1500_n633# a_n88_n633# 0.00fF
C2932 a_n2658_n197# a_n2868_131# 0.01fF
C2933 a_n2238_n197# a_n3288_131# 0.00fF
C2934 a_n300_n100# a_n1232_n100# 0.01fF
C2935 a_n3286_n401# a_n3288_131# 0.01fF
C2936 a_2382_n197# a_1752_131# 0.00fF
C2937 a_120_n100# a_n1022_n100# 0.01fF
C2938 a_n1650_n633# a_n3238_n633# 0.00fF
C2939 a_n1860_n633# a_n1816_n730# 0.00fF
C2940 a_72_131# a_n768_131# 0.01fF
C2941 a_n1980_n100# a_n2492_n100# 0.01fF
C2942 a_2382_n197# a_2172_131# 0.01fF
C2943 a_n3542_n100# a_n4080_n100# 0.01fF
C2944 a_n2700_n633# a_n3120_n633# 0.02fF
C2945 a_n2818_n633# a_n3028_n633# 0.03fF
C2946 a_n2608_n633# a_n3238_n633# 0.01fF
C2947 a_n600_n633# a_n2070_n633# 0.00fF
C2948 a_n138_n197# a_n558_n197# 0.01fF
C2949 a_1964_n730# a_3434_n401# 0.00fF
C2950 a_3222_n197# a_1752_131# 0.00fF
C2951 a_n3542_n100# a_n3962_n100# 0.02fF
C2952 a_2970_n633# a_1500_n633# 0.00fF
C2953 a_n3960_n633# a_n3962_n100# 0.00fF
C2954 a_2852_n633# w_n4520_n852# 0.03fF
C2955 a_1754_n401# a_914_n401# 0.01fF
C2956 a_28_n100# a_n1442_n100# 0.00fF
C2957 a_4110_n100# w_n4520_n852# 0.14fF
C2958 a_1382_n633# a_n88_n633# 0.00fF
C2959 a_3222_n197# a_2172_131# 0.00fF
C2960 a_n3078_n197# a_n2868_131# 0.01fF
C2961 a_n1140_n100# a_n2190_n100# 0.01fF
C2962 a_n2658_n197# a_n3288_131# 0.00fF
C2963 a_28_n100# a_n1350_n100# 0.00fF
C2964 a_n392_n100# a_n1232_n100# 0.01fF
C2965 a_1962_n197# a_1752_131# 0.01fF
C2966 a_2804_n730# a_2850_n100# 0.00fF
C2967 a_332_n633# a_n508_n633# 0.01fF
C2968 a_72_131# a_n1188_131# 0.00fF
C2969 a_1962_n197# a_2172_131# 0.01fF
C2970 a_n3660_n100# a_n4080_n100# 0.02fF
C2971 a_n2818_n633# a_n3120_n633# 0.02fF
C2972 a_n2700_n633# a_n3238_n633# 0.01fF
C2973 a_n2910_n633# a_n3028_n633# 0.07fF
C2974 a_1334_n401# a_494_n401# 0.01fF
C2975 a_n298_n633# a_n300_n100# 0.00fF
C2976 a_n718_n633# a_n2070_n633# 0.00fF
C2977 a_n600_n633# a_n2188_n633# 0.00fF
C2978 a_2970_n633# a_1382_n633# 0.00fF
C2979 a_n1816_n730# a_n1818_n197# 0.01fF
C2980 a_n3660_n100# a_n3962_n100# 0.02fF
C2981 a_2760_n633# w_n4520_n852# 0.02fF
C2982 a_2970_n633# a_3012_131# 0.00fF
C2983 a_n1232_n100# a_n2702_n100# 0.00fF
C2984 a_n90_n100# a_n1442_n100# 0.00fF
C2985 a_1080_n633# a_122_n633# 0.01fF
C2986 a_1382_n633# a_n180_n633# 0.00fF
C2987 a_1290_n633# a_n88_n633# 0.00fF
C2988 a_n3498_n197# a_n2868_131# 0.00fF
C2989 a_n3078_n197# a_n3288_131# 0.01fF
C2990 a_n510_n100# a_n1232_n100# 0.01fF
C2991 a_n90_n100# a_n1350_n100# 0.00fF
C2992 a_240_n633# a_n508_n633# 0.01fF
C2993 a_332_n633# a_n600_n633# 0.01fF
C2994 a_1380_n100# a_960_n100# 0.02fF
C2995 a_1078_n100# a_960_n100# 0.07fF
C2996 a_n2910_n633# a_n3120_n633# 0.03fF
C2997 a_n2818_n633# a_n3238_n633# 0.02fF
C2998 a_1334_n401# a_74_n401# 0.00fF
C2999 a_n1770_n100# a_n2072_n100# 0.02fF
C3000 a_n718_n633# a_n2188_n633# 0.00fF
C3001 a_n810_n633# a_n2070_n633# 0.00fF
C3002 a_n1140_n100# a_n2492_n100# 0.00fF
C3003 a_n4172_n100# w_n4520_n852# 0.14fF
C3004 a_n1232_n100# a_n2820_n100# 0.00fF
C3005 a_3482_n633# a_3390_n633# 0.09fF
C3006 a_n182_n100# a_n1442_n100# 0.00fF
C3007 a_n1816_n730# a_n3286_n401# 0.00fF
C3008 a_1172_n633# a_n88_n633# 0.00fF
C3009 a_1290_n633# a_n180_n633# 0.00fF
C3010 a_1080_n633# a_30_n633# 0.01fF
C3011 a_n3498_n197# a_n3288_131# 0.01fF
C3012 a_n3918_n197# a_n2868_131# 0.00fF
C3013 a_n3076_n730# a_n3030_n100# 0.00fF
C3014 a_n602_n100# a_n1232_n100# 0.01fF
C3015 a_n182_n100# a_n1350_n100# 0.01fF
C3016 a_332_n633# a_n718_n633# 0.01fF
C3017 a_240_n633# a_n600_n633# 0.01fF
C3018 a_494_n401# a_74_n401# 0.01fF
C3019 a_n3028_n633# a_n3120_n633# 0.09fF
C3020 a_n2910_n633# a_n3238_n633# 0.02fF
C3021 a_n1862_n100# a_n2072_n100# 0.03fF
C3022 a_n810_n633# a_n2188_n633# 0.00fF
C3023 a_n390_n633# a_n392_n100# 0.00fF
C3024 a_n718_n633# a_n2280_n633# 0.00fF
C3025 a_n928_n633# a_n2070_n633# 0.01fF
C3026 a_n2236_n730# a_n2238_n197# 0.01fF
C3027 a_n300_n100# a_n1442_n100# 0.01fF
C3028 a_n2236_n730# a_n3286_n401# 0.00fF
C3029 a_1498_n100# a_540_n100# 0.01fF
C3030 a_1290_n633# a_n298_n633# 0.00fF
C3031 a_1172_n633# a_n180_n633# 0.00fF
C3032 a_n3918_n197# a_n3288_131# 0.00fF
C3033 a_n720_n100# a_n1232_n100# 0.01fF
C3034 a_n300_n100# a_n1350_n100# 0.01fF
C3035 a_240_n633# a_n718_n633# 0.01fF
C3036 a_332_n633# a_n810_n633# 0.01fF
C3037 a_n1560_n100# w_n4520_n852# 0.02fF
C3038 a_494_n401# a_n346_n401# 0.01fF
C3039 a_962_n633# a_752_n633# 0.03fF
C3040 a_n1558_n633# w_n4520_n852# 0.01fF
C3041 a_n3028_n633# a_n3238_n633# 0.03fF
C3042 a_1380_n100# a_448_n100# 0.01fF
C3043 a_n1138_n633# a_n1978_n633# 0.01fF
C3044 a_n1020_n633# a_n2070_n633# 0.01fF
C3045 a_n928_n633# a_n2188_n633# 0.00fF
C3046 a_n810_n633# a_n2280_n633# 0.00fF
C3047 a_2852_n633# a_2550_n633# 0.02fF
C3048 a_2970_n633# a_2432_n633# 0.01fF
C3049 a_2850_n100# a_2802_n197# 0.00fF
C3050 a_1078_n100# a_448_n100# 0.01fF
C3051 a_n392_n100# a_n1442_n100# 0.01fF
C3052 a_n2656_n730# a_n3286_n401# 0.00fF
C3053 a_n2236_n730# a_n3706_n401# 0.00fF
C3054 a_1172_n633# a_n298_n633# 0.00fF
C3055 a_n392_n100# a_n1350_n100# 0.01fF
C3056 a_n812_n100# a_n1232_n100# 0.02fF
C3057 a_240_n633# a_n810_n633# 0.01fF
C3058 a_120_n100# a_28_n100# 0.09fF
C3059 a_332_n633# a_n928_n633# 0.00fF
C3060 a_494_n401# a_n766_n401# 0.00fF
C3061 a_74_n401# a_n346_n401# 0.01fF
C3062 a_n2608_n633# a_n3658_n633# 0.01fF
C3063 a_n2190_n100# w_n4520_n852# 0.02fF
C3064 a_n1650_n633# w_n4520_n852# 0.01fF
C3065 a_n1442_n100# a_n2702_n100# 0.00fF
C3066 a_n3120_n633# a_n3238_n633# 0.07fF
C3067 a_n2608_n633# a_n3540_n633# 0.01fF
C3068 a_n1020_n633# a_n2188_n633# 0.01fF
C3069 a_n928_n633# a_n2280_n633# 0.00fF
C3070 a_n810_n633# a_n2398_n633# 0.00fF
C3071 a_3062_n633# a_2222_n633# 0.01fF
C3072 a_2760_n633# a_2550_n633# 0.03fF
C3073 a_2970_n633# a_2340_n633# 0.01fF
C3074 a_2758_n100# a_2802_n197# 0.00fF
C3075 a_n4128_131# w_n4520_n852# 0.14fF
C3076 a_n2608_n633# w_n4520_n852# 0.01fF
C3077 a_n2656_n730# a_n2658_n197# 0.01fF
C3078 a_n1350_n100# a_n2702_n100# 0.00fF
C3079 a_n510_n100# a_n1442_n100# 0.01fF
C3080 a_n2656_n730# a_n3706_n401# 0.00fF
C3081 a_1542_n197# a_492_131# 0.00fF
C3082 a_3690_n100# a_3598_n100# 0.09fF
C3083 a_n1140_n100# a_n1980_n100# 0.01fF
C3084 a_n558_n197# a_n2028_131# 0.00fF
C3085 a_1172_n633# a_n390_n633# 0.00fF
C3086 a_870_n633# w_n4520_n852# 0.01fF
C3087 a_n510_n100# a_n1350_n100# 0.01fF
C3088 a_n930_n100# a_n1232_n100# 0.02fF
C3089 a_2384_n730# a_2430_n100# 0.00fF
C3090 a_120_n100# a_n90_n100# 0.03fF
C3091 a_332_n633# a_n1020_n633# 0.00fF
C3092 a_240_n633# a_n928_n633# 0.01fF
C3093 a_450_n633# a_n1138_n633# 0.00fF
C3094 a_74_n401# a_n766_n401# 0.01fF
C3095 a_n2700_n633# a_n3658_n633# 0.01fF
C3096 a_n1442_n100# a_n2820_n100# 0.00fF
C3097 a_n2700_n633# a_n3540_n633# 0.01fF
C3098 a_n1020_n633# a_n2280_n633# 0.00fF
C3099 a_n928_n633# a_n2398_n633# 0.00fF
C3100 a_3062_n633# a_2130_n633# 0.01fF
C3101 a_n2700_n633# w_n4520_n852# 0.02fF
C3102 a_n1350_n100# a_n2820_n100# 0.00fF
C3103 a_n602_n100# a_n1442_n100# 0.01fF
C3104 a_3690_n100# a_3480_n100# 0.03fF
C3105 a_n2492_n100# w_n4520_n852# 0.02fF
C3106 a_n2280_n633# a_n2282_n100# 0.00fF
C3107 a_n2026_n401# a_n2028_131# 0.01fF
C3108 a_n602_n100# a_n1350_n100# 0.01fF
C3109 a_240_n633# a_n1020_n633# 0.00fF
C3110 a_120_n100# a_n182_n100# 0.02fF
C3111 a_n346_n401# a_n766_n401# 0.01fF
C3112 a_74_n401# a_n1186_n401# 0.00fF
C3113 a_n2818_n633# a_n3658_n633# 0.01fF
C3114 a_1380_n100# a_658_n100# 0.01fF
C3115 a_n4078_n633# a_n4170_n633# 0.09fF
C3116 a_870_n633# a_914_n401# 0.00fF
C3117 a_n1442_n100# a_n2912_n100# 0.00fF
C3118 a_n2818_n633# a_n3540_n633# 0.01fF
C3119 a_1078_n100# a_658_n100# 0.02fF
C3120 a_868_n100# a_912_131# 0.00fF
C3121 a_n928_n633# a_n2490_n633# 0.00fF
C3122 a_n1020_n633# a_n2398_n633# 0.00fF
C3123 a_3062_n633# a_2012_n633# 0.01fF
C3124 a_n2818_n633# w_n4520_n852# 0.02fF
C3125 a_n1350_n100# a_n2912_n100# 0.00fF
C3126 a_n720_n100# a_n1442_n100# 0.01fF
C3127 a_3690_n100# a_3388_n100# 0.02fF
C3128 a_542_n633# a_n88_n633# 0.01fF
C3129 a_332_n633# a_122_n633# 0.03fF
C3130 a_n720_n100# a_n1350_n100# 0.01fF
C3131 a_n1348_n633# a_n1768_n633# 0.02fF
C3132 a_120_n100# a_n300_n100# 0.02fF
C3133 a_n346_n401# a_n1186_n401# 0.01fF
C3134 a_n2910_n633# a_n3658_n633# 0.01fF
C3135 a_960_n100# a_540_n100# 0.02fF
C3136 a_n2610_n100# a_n3870_n100# 0.00fF
C3137 a_n1442_n100# a_n3030_n100# 0.00fF
C3138 a_n2910_n633# a_n3540_n633# 0.01fF
C3139 a_n1020_n633# a_n2490_n633# 0.00fF
C3140 a_3062_n633# a_1920_n633# 0.01fF
C3141 a_282_n197# w_n4520_n852# 0.10fF
C3142 a_n1230_n633# w_n4520_n852# 0.01fF
C3143 a_n138_n197# a_n1608_131# 0.00fF
C3144 a_n2910_n633# w_n4520_n852# 0.03fF
C3145 a_4062_n197# a_2592_131# 0.00fF
C3146 a_n812_n100# a_n1442_n100# 0.01fF
C3147 a_1710_n633# a_122_n633# 0.00fF
C3148 a_332_n633# a_30_n633# 0.02fF
C3149 a_240_n633# a_122_n633# 0.07fF
C3150 a_542_n633# a_n180_n633# 0.01fF
C3151 a_450_n633# a_n88_n633# 0.01fF
C3152 a_n812_n100# a_n1350_n100# 0.01fF
C3153 a_120_n100# a_n392_n100# 0.01fF
C3154 a_n766_n401# a_n1186_n401# 0.01fF
C3155 a_n346_n401# a_n1606_n401# 0.00fF
C3156 a_n3028_n633# a_n3658_n633# 0.01fF
C3157 a_3482_n633# w_n4520_n852# 0.03fF
C3158 a_n3330_n633# a_n3750_n633# 0.02fF
C3159 a_n3028_n633# a_n3540_n633# 0.01fF
C3160 a_3062_n633# a_1802_n633# 0.00fF
C3161 a_n3028_n633# w_n4520_n852# 0.03fF
C3162 a_n930_n100# a_n1442_n100# 0.01fF
C3163 a_448_n100# a_492_131# 0.00fF
C3164 a_240_n633# a_30_n633# 0.03fF
C3165 a_450_n633# a_n180_n633# 0.01fF
C3166 a_542_n633# a_n298_n633# 0.01fF
C3167 a_n930_n100# a_n1350_n100# 0.02fF
C3168 a_120_n100# a_n510_n100# 0.01fF
C3169 a_1170_n100# w_n4520_n852# 0.02fF
C3170 a_n766_n401# a_n1606_n401# 0.01fF
C3171 a_n1980_n100# w_n4520_n852# 0.02fF
C3172 a_n3120_n633# a_n3658_n633# 0.01fF
C3173 a_n90_n100# a_n138_n197# 0.00fF
C3174 a_3390_n633# w_n4520_n852# 0.03fF
C3175 a_n3448_n633# a_n3750_n633# 0.02fF
C3176 a_n390_n633# a_n1978_n633# 0.00fF
C3177 a_n1232_n100# a_n1188_131# 0.00fF
C3178 a_n1560_n100# a_n1770_n100# 0.03fF
C3179 a_n3120_n633# a_n3540_n633# 0.02fF
C3180 a_540_n100# a_448_n100# 0.09fF
C3181 a_3062_n633# a_1710_n633# 0.00fF
C3182 a_2222_n633# a_2220_n100# 0.00fF
C3183 a_n3120_n633# w_n4520_n852# 0.03fF
C3184 a_2968_n100# w_n4520_n852# 0.03fF
C3185 a_n3750_n633# a_n3752_n100# 0.00fF
C3186 a_542_n633# a_n390_n633# 0.01fF
C3187 a_450_n633# a_n298_n633# 0.01fF
C3188 a_1964_n730# a_2010_n100# 0.00fF
C3189 a_120_n100# a_n602_n100# 0.01fF
C3190 a_3432_131# a_2172_131# 0.00fF
C3191 a_n1186_n401# a_n1606_n401# 0.01fF
C3192 a_n766_n401# a_n2026_n401# 0.00fF
C3193 a_n3238_n633# a_n3658_n633# 0.02fF
C3194 a_n182_n100# a_n138_n197# 0.00fF
C3195 a_n1560_n100# a_n1862_n100# 0.02fF
C3196 a_n3238_n633# a_n3540_n633# 0.02fF
C3197 a_n1770_n100# a_n2190_n100# 0.02fF
C3198 a_3224_n730# a_3854_n401# 0.00fF
C3199 a_n3238_n633# w_n4520_n852# 0.03fF
C3200 a_2850_n100# a_1498_n100# 0.00fF
C3201 a_1590_n100# a_1380_n100# 0.03fF
C3202 a_n1558_n633# a_n1860_n633# 0.02fF
C3203 a_n1440_n633# a_n1978_n633# 0.01fF
C3204 a_3598_n100# a_3270_n100# 0.02fF
C3205 a_3060_n100# a_3012_131# 0.00fF
C3206 a_72_131# a_n348_131# 0.01fF
C3207 a_450_n633# a_n390_n633# 0.01fF
C3208 a_1590_n100# a_1078_n100# 0.01fF
C3209 a_120_n100# a_n720_n100# 0.01fF
C3210 a_n1186_n401# a_n2026_n401# 0.01fF
C3211 a_3180_n633# a_3062_n633# 0.07fF
C3212 a_2130_n633# a_2128_n100# 0.00fF
C3213 a_n1140_n100# w_n4520_n852# 0.02fF
C3214 a_n1862_n100# a_n2190_n100# 0.02fF
C3215 a_492_131# a_72_131# 0.01fF
C3216 a_3224_n730# a_3434_n401# 0.01fF
C3217 a_2758_n100# a_1498_n100# 0.00fF
C3218 a_3900_n100# a_3852_131# 0.00fF
C3219 a_4112_n633# a_2852_n633# 0.00fF
C3220 a_n1650_n633# a_n1860_n633# 0.03fF
C3221 a_n508_n633# a_n556_n730# 0.00fF
C3222 a_3480_n100# a_3270_n100# 0.03fF
C3223 a_4112_n633# a_4110_n100# 0.00fF
C3224 a_n2072_n100# a_n2400_n100# 0.02fF
C3225 a_120_n100# a_n812_n100# 0.01fF
C3226 a_n1606_n401# a_n2026_n401# 0.01fF
C3227 a_n1186_n401# a_n2446_n401# 0.00fF
C3228 a_3482_n633# a_2550_n633# 0.01fF
C3229 a_n1860_n633# a_n2608_n633# 0.01fF
C3230 a_n1770_n100# a_n2492_n100# 0.01fF
C3231 a_n1652_n100# a_n2610_n100# 0.01fF
C3232 a_658_n100# a_540_n100# 0.07fF
C3233 a_2640_n100# a_1498_n100# 0.01fF
C3234 a_3808_n100# a_3852_131# 0.00fF
C3235 a_4112_n633# a_2760_n633# 0.00fF
C3236 a_4020_n633# a_2852_n633# 0.01fF
C3237 a_n1188_131# a_n2448_131# 0.00fF
C3238 a_n1608_131# a_n2028_131# 0.01fF
C3239 a_n600_n633# a_n556_n730# 0.00fF
C3240 a_3388_n100# a_3270_n100# 0.07fF
C3241 a_870_n633# a_660_n633# 0.03fF
C3242 a_120_n100# a_n930_n100# 0.01fF
C3243 a_n1606_n401# a_n2446_n401# 0.01fF
C3244 a_n1860_n633# a_n2700_n633# 0.01fF
C3245 a_1288_n100# a_1498_n100# 0.03fF
C3246 a_3390_n633# a_2550_n633# 0.01fF
C3247 a_n1862_n100# a_n2492_n100# 0.01fF
C3248 a_1592_n633# a_962_n633# 0.01fF
C3249 a_702_n197# a_282_n197# 0.01fF
C3250 a_n3752_n100# a_n3870_n100# 0.07fF
C3251 a_2012_n633# a_2010_n100# 0.00fF
C3252 a_2548_n100# a_1498_n100# 0.01fF
C3253 a_n1022_n100# a_n1652_n100# 0.01fF
C3254 a_3902_n633# a_2852_n633# 0.01fF
C3255 a_4020_n633# a_2760_n633# 0.00fF
C3256 a_n2608_n633# a_n3868_n633# 0.00fF
C3257 a_n138_n197# a_1332_131# 0.00fF
C3258 a_n1606_n401# a_n2866_n401# 0.00fF
C3259 a_n2026_n401# a_n2446_n401# 0.01fF
C3260 a_n1860_n633# a_n2818_n633# 0.01fF
C3261 a_1500_n633# a_962_n633# 0.01fF
C3262 a_3600_n633# a_3644_n730# 0.00fF
C3263 a_n2190_n100# a_n2238_n197# 0.00fF
C3264 w_n4520_n852# VSUBS 31.76fF
.ends

.subckt latch_pmos_pair sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n852# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n633#
+ VSUBS sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
Xsky130_fd_pr__pfet_01v8_VCQUSW_0 sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n852# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n730# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n730#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n730#
+ VSUBS sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n633# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n633#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100# sky130_fd_pr__pfet_01v8_VCQUSW
C0 sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n852# VSUBS 31.76fF
.ends

.subckt sky130_fd_pr__pfet_01v8_VCG74W a_543_n100# a_159_n100# a_n609_n100# a_495_n197#
+ a_n705_n100# a_255_n100# a_n657_n197# a_n369_131# a_351_n100# a_n417_n100# a_n801_n100#
+ a_303_n197# a_n129_n100# a_n513_n100# a_n465_n197# a_n561_131# a_63_n100# a_n225_n100#
+ a_399_131# a_111_n197# a_n321_n100# a_n273_n197# a_15_131# a_n753_131# a_639_n100#
+ w_n1031_n319# a_591_131# a_207_131# a_735_n100# a_n33_n100# a_687_n197# a_447_n100#
+ a_n81_n197# a_n177_131# VSUBS
X0 a_63_n100# a_15_131# a_n33_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n129_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_255_n100# a_207_131# a_159_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_351_n100# a_303_n197# a_255_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_543_n100# a_495_n197# a_447_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 w_n1031_n319# w_n1031_n319# a_735_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=5.24e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_159_n100# a_111_n197# a_63_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_447_n100# a_399_131# a_351_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_639_n100# a_591_131# a_543_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_735_n100# a_687_n197# a_639_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n801_n100# w_n1031_n319# w_n1031_n319# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_n513_n100# a_n561_131# a_n609_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_n321_n100# a_n369_131# a_n417_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_n225_n100# a_n273_n197# a_n321_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_n705_n100# a_n753_131# a_n801_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_n609_n100# a_n657_n197# a_n705_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n417_n100# a_n465_n197# a_n513_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n129_n100# a_n177_131# a_n225_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_351_n100# a_n705_n100# 0.01fF
C1 a_255_n100# a_n609_n100# 0.01fF
C2 a_639_n100# a_255_n100# 0.02fF
C3 a_159_n100# a_n129_n100# 0.02fF
C4 a_255_n100# a_n705_n100# 0.01fF
C5 a_543_n100# a_495_n197# 0.00fF
C6 a_351_n100# a_n801_n100# 0.01fF
C7 a_n657_n197# a_n81_n197# 0.01fF
C8 a_399_131# a_111_n197# 0.00fF
C9 a_399_131# a_303_n197# 0.01fF
C10 a_n177_131# a_n657_n197# 0.00fF
C11 a_n561_131# a_111_n197# 0.00fF
C12 a_n561_131# a_303_n197# 0.00fF
C13 w_n1031_n319# a_447_n100# 0.05fF
C14 a_255_n100# a_n801_n100# 0.01fF
C15 a_15_131# a_n33_n100# 0.00fF
C16 w_n1031_n319# a_543_n100# 0.06fF
C17 w_n1031_n319# a_351_n100# 0.05fF
C18 a_n273_n197# a_111_n197# 0.01fF
C19 a_n273_n197# a_303_n197# 0.01fF
C20 w_n1031_n319# a_255_n100# 0.05fF
C21 a_63_n100# a_111_n197# 0.00fF
C22 a_n753_131# a_399_131# 0.00fF
C23 a_n561_131# a_n753_131# 0.04fF
C24 a_n657_n197# a_n609_n100# 0.00fF
C25 a_n561_131# a_n513_n100# 0.00fF
C26 a_n657_n197# a_n705_n100# 0.00fF
C27 a_447_n100# a_n33_n100# 0.01fF
C28 a_447_n100# a_735_n100# 0.02fF
C29 a_n273_n197# a_n225_n100# 0.00fF
C30 a_n465_n197# a_n657_n197# 0.04fF
C31 a_n657_n197# a_687_n197# 0.00fF
C32 a_n273_n197# a_n321_n100# 0.00fF
C33 a_63_n100# a_n225_n100# 0.02fF
C34 a_n273_n197# a_n753_131# 0.00fF
C35 a_543_n100# a_n33_n100# 0.01fF
C36 a_n657_n197# a_495_n197# 0.00fF
C37 a_543_n100# a_735_n100# 0.04fF
C38 a_63_n100# a_n321_n100# 0.02fF
C39 a_63_n100# a_n417_n100# 0.01fF
C40 a_351_n100# a_n33_n100# 0.02fF
C41 a_351_n100# a_735_n100# 0.02fF
C42 a_63_n100# a_n513_n100# 0.01fF
C43 a_207_131# a_399_131# 0.04fF
C44 a_591_131# a_n81_n197# 0.00fF
C45 a_255_n100# a_n33_n100# 0.02fF
C46 a_255_n100# a_735_n100# 0.01fF
C47 a_n657_n197# w_n1031_n319# 0.16fF
C48 a_n561_131# a_207_131# 0.01fF
C49 a_n177_131# a_591_131# 0.01fF
C50 a_n369_131# a_399_131# 0.01fF
C51 a_n369_131# a_n561_131# 0.04fF
C52 a_n273_n197# a_207_131# 0.00fF
C53 a_15_131# a_399_131# 0.01fF
C54 a_n561_131# a_15_131# 0.01fF
C55 a_159_n100# a_n609_n100# 0.01fF
C56 a_639_n100# a_159_n100# 0.01fF
C57 a_n273_n197# a_n369_131# 0.01fF
C58 a_159_n100# a_n705_n100# 0.01fF
C59 a_303_n197# a_111_n197# 0.04fF
C60 a_159_n100# a_n801_n100# 0.01fF
C61 a_591_131# a_639_n100# 0.00fF
C62 a_n273_n197# a_15_131# 0.00fF
C63 a_n465_n197# a_591_131# 0.00fF
C64 a_591_131# a_687_n197# 0.01fF
C65 a_15_131# a_63_n100# 0.00fF
C66 a_591_131# a_495_n197# 0.01fF
C67 a_n129_n100# a_n81_n197# 0.00fF
C68 a_399_131# a_447_n100# 0.00fF
C69 w_n1031_n319# a_159_n100# 0.04fF
C70 a_n177_131# a_n129_n100# 0.00fF
C71 a_n753_131# a_111_n197# 0.00fF
C72 a_n753_131# a_303_n197# 0.00fF
C73 w_n1031_n319# a_591_131# 0.12fF
C74 a_399_131# a_351_n100# 0.00fF
C75 a_447_n100# a_63_n100# 0.02fF
C76 a_n225_n100# a_n321_n100# 0.09fF
C77 a_n225_n100# a_n417_n100# 0.04fF
C78 a_n129_n100# a_n609_n100# 0.01fF
C79 a_639_n100# a_n129_n100# 0.01fF
C80 a_n225_n100# a_n513_n100# 0.02fF
C81 a_n321_n100# a_n417_n100# 0.09fF
C82 a_543_n100# a_63_n100# 0.01fF
C83 a_n321_n100# a_n513_n100# 0.04fF
C84 a_n129_n100# a_n705_n100# 0.01fF
C85 a_207_131# a_111_n197# 0.01fF
C86 a_159_n100# a_n33_n100# 0.04fF
C87 a_159_n100# a_735_n100# 0.01fF
C88 a_207_131# a_303_n197# 0.01fF
C89 a_351_n100# a_63_n100# 0.02fF
C90 a_n129_n100# a_n801_n100# 0.01fF
C91 a_n417_n100# a_n513_n100# 0.09fF
C92 a_n369_131# a_111_n197# 0.00fF
C93 a_255_n100# a_63_n100# 0.04fF
C94 a_n369_131# a_303_n197# 0.00fF
C95 a_n177_131# a_n81_n197# 0.01fF
C96 a_n657_n197# a_399_131# 0.00fF
C97 a_15_131# a_111_n197# 0.01fF
C98 a_n657_n197# a_n561_131# 0.01fF
C99 a_15_131# a_303_n197# 0.00fF
C100 w_n1031_n319# a_n129_n100# 0.04fF
C101 a_n753_131# a_207_131# 0.01fF
C102 a_n369_131# a_n321_n100# 0.00fF
C103 a_n369_131# a_n753_131# 0.01fF
C104 a_n369_131# a_n417_n100# 0.00fF
C105 a_n273_n197# a_n657_n197# 0.01fF
C106 a_n753_131# a_15_131# 0.01fF
C107 a_n465_n197# a_n81_n197# 0.01fF
C108 a_n33_n100# a_n129_n100# 0.09fF
C109 a_n129_n100# a_735_n100# 0.01fF
C110 a_687_n197# a_n81_n197# 0.01fF
C111 a_n465_n197# a_n177_131# 0.00fF
C112 a_n177_131# a_687_n197# 0.00fF
C113 a_495_n197# a_n81_n197# 0.01fF
C114 a_n369_131# a_207_131# 0.01fF
C115 a_n177_131# a_495_n197# 0.00fF
C116 a_351_n100# a_303_n197# 0.00fF
C117 a_255_n100# a_303_n197# 0.00fF
C118 a_447_n100# a_n225_n100# 0.01fF
C119 w_n1031_n319# a_n81_n197# 0.13fF
C120 a_447_n100# a_n321_n100# 0.01fF
C121 a_n177_131# w_n1031_n319# 0.13fF
C122 a_591_131# a_399_131# 0.04fF
C123 a_207_131# a_15_131# 0.04fF
C124 a_n561_131# a_591_131# 0.00fF
C125 a_447_n100# a_n417_n100# 0.01fF
C126 a_543_n100# a_n225_n100# 0.01fF
C127 a_639_n100# a_n609_n100# 0.00fF
C128 a_543_n100# a_n321_n100# 0.01fF
C129 a_n609_n100# a_n705_n100# 0.09fF
C130 a_639_n100# a_n705_n100# 0.00fF
C131 a_447_n100# a_n513_n100# 0.01fF
C132 a_n369_131# a_15_131# 0.01fF
C133 a_639_n100# a_n801_n100# 0.00fF
C134 a_351_n100# a_n225_n100# 0.01fF
C135 a_543_n100# a_n417_n100# 0.01fF
C136 a_n609_n100# a_n801_n100# 0.04fF
C137 a_n705_n100# a_n801_n100# 0.09fF
C138 a_543_n100# a_n513_n100# 0.01fF
C139 a_351_n100# a_n321_n100# 0.01fF
C140 a_255_n100# a_n225_n100# 0.01fF
C141 a_639_n100# a_687_n197# 0.00fF
C142 a_159_n100# a_63_n100# 0.09fF
C143 a_255_n100# a_n321_n100# 0.01fF
C144 a_351_n100# a_n417_n100# 0.01fF
C145 a_n273_n197# a_591_131# 0.00fF
C146 a_351_n100# a_n513_n100# 0.01fF
C147 a_255_n100# a_n417_n100# 0.01fF
C148 a_n465_n197# a_687_n197# 0.00fF
C149 a_255_n100# a_n513_n100# 0.01fF
C150 a_n465_n197# a_495_n197# 0.01fF
C151 w_n1031_n319# a_n609_n100# 0.06fF
C152 a_687_n197# a_495_n197# 0.04fF
C153 w_n1031_n319# a_639_n100# 0.08fF
C154 a_n657_n197# a_111_n197# 0.01fF
C155 a_n657_n197# a_303_n197# 0.01fF
C156 a_n33_n100# a_n81_n197# 0.00fF
C157 w_n1031_n319# a_n705_n100# 0.08fF
C158 w_n1031_n319# a_n801_n100# 0.15fF
C159 a_n465_n197# w_n1031_n319# 0.14fF
C160 w_n1031_n319# a_687_n197# 0.13fF
C161 w_n1031_n319# a_495_n197# 0.11fF
C162 a_207_131# a_255_n100# 0.00fF
C163 a_n657_n197# a_n753_131# 0.01fF
C164 a_n33_n100# a_n609_n100# 0.01fF
C165 a_n609_n100# a_735_n100# 0.00fF
C166 a_639_n100# a_n33_n100# 0.01fF
C167 a_639_n100# a_735_n100# 0.09fF
C168 a_n33_n100# a_n705_n100# 0.01fF
C169 a_n705_n100# a_735_n100# 0.00fF
C170 a_n33_n100# a_n801_n100# 0.01fF
C171 a_n801_n100# a_735_n100# 0.00fF
C172 a_63_n100# a_n129_n100# 0.04fF
C173 a_687_n197# a_735_n100# 0.00fF
C174 a_159_n100# a_111_n197# 0.00fF
C175 a_n657_n197# a_207_131# 0.00fF
C176 a_591_131# a_111_n197# 0.00fF
C177 a_591_131# a_303_n197# 0.00fF
C178 a_447_n100# a_543_n100# 0.09fF
C179 w_n1031_n319# a_n33_n100# 0.04fF
C180 w_n1031_n319# a_735_n100# 0.15fF
C181 a_n657_n197# a_n369_131# 0.00fF
C182 a_447_n100# a_351_n100# 0.09fF
C183 a_159_n100# a_n225_n100# 0.02fF
C184 a_447_n100# a_255_n100# 0.04fF
C185 a_399_131# a_n81_n197# 0.00fF
C186 a_n561_131# a_n81_n197# 0.00fF
C187 a_n177_131# a_399_131# 0.01fF
C188 a_159_n100# a_n321_n100# 0.01fF
C189 a_543_n100# a_351_n100# 0.04fF
C190 a_n177_131# a_n561_131# 0.01fF
C191 a_n657_n197# a_15_131# 0.00fF
C192 a_159_n100# a_n417_n100# 0.01fF
C193 a_543_n100# a_255_n100# 0.02fF
C194 a_159_n100# a_n513_n100# 0.01fF
C195 a_n753_131# a_591_131# 0.00fF
C196 a_351_n100# a_255_n100# 0.09fF
C197 a_n273_n197# a_n81_n197# 0.04fF
C198 a_n273_n197# a_n177_131# 0.01fF
C199 a_n33_n100# a_735_n100# 0.01fF
C200 a_n561_131# a_n609_n100# 0.00fF
C201 a_207_131# a_159_n100# 0.00fF
C202 a_207_131# a_591_131# 0.01fF
C203 a_n465_n197# a_399_131# 0.00fF
C204 a_399_131# a_687_n197# 0.00fF
C205 a_n465_n197# a_n561_131# 0.01fF
C206 a_n561_131# a_687_n197# 0.00fF
C207 a_399_131# a_495_n197# 0.01fF
C208 a_n561_131# a_495_n197# 0.00fF
C209 a_n369_131# a_591_131# 0.01fF
C210 a_63_n100# a_n609_n100# 0.01fF
C211 a_639_n100# a_63_n100# 0.01fF
C212 a_n129_n100# a_n225_n100# 0.09fF
C213 w_n1031_n319# a_399_131# 0.12fF
C214 a_63_n100# a_n705_n100# 0.01fF
C215 w_n1031_n319# a_n561_131# 0.14fF
C216 a_n129_n100# a_n321_n100# 0.04fF
C217 a_n273_n197# a_n465_n197# 0.04fF
C218 a_n273_n197# a_687_n197# 0.01fF
C219 a_15_131# a_591_131# 0.01fF
C220 a_63_n100# a_n801_n100# 0.01fF
C221 a_n129_n100# a_n417_n100# 0.02fF
C222 a_n273_n197# a_495_n197# 0.01fF
C223 a_n129_n100# a_n513_n100# 0.02fF
C224 a_n273_n197# w_n1031_n319# 0.13fF
C225 w_n1031_n319# a_63_n100# 0.04fF
C226 a_447_n100# a_159_n100# 0.02fF
C227 a_111_n197# a_n81_n197# 0.04fF
C228 a_303_n197# a_n81_n197# 0.01fF
C229 a_n177_131# a_111_n197# 0.00fF
C230 a_n177_131# a_303_n197# 0.00fF
C231 a_543_n100# a_159_n100# 0.02fF
C232 a_351_n100# a_159_n100# 0.04fF
C233 a_591_131# a_543_n100# 0.00fF
C234 a_255_n100# a_159_n100# 0.09fF
C235 a_n177_131# a_n225_n100# 0.00fF
C236 a_n753_131# a_n81_n197# 0.00fF
C237 a_n177_131# a_n753_131# 0.01fF
C238 a_63_n100# a_n33_n100# 0.09fF
C239 a_63_n100# a_735_n100# 0.01fF
C240 a_n465_n197# a_111_n197# 0.01fF
C241 a_687_n197# a_111_n197# 0.01fF
C242 a_n465_n197# a_303_n197# 0.01fF
C243 a_687_n197# a_303_n197# 0.01fF
C244 a_495_n197# a_111_n197# 0.01fF
C245 a_495_n197# a_303_n197# 0.04fF
C246 a_n225_n100# a_n609_n100# 0.02fF
C247 a_639_n100# a_n225_n100# 0.01fF
C248 a_447_n100# a_n129_n100# 0.01fF
C249 a_n321_n100# a_n609_n100# 0.02fF
C250 a_639_n100# a_n321_n100# 0.01fF
C251 a_207_131# a_n81_n197# 0.00fF
C252 a_n225_n100# a_n705_n100# 0.01fF
C253 w_n1031_n319# a_111_n197# 0.12fF
C254 a_n177_131# a_207_131# 0.01fF
C255 w_n1031_n319# a_303_n197# 0.11fF
C256 a_n417_n100# a_n609_n100# 0.04fF
C257 a_639_n100# a_n417_n100# 0.01fF
C258 a_n225_n100# a_n801_n100# 0.01fF
C259 a_n321_n100# a_n705_n100# 0.02fF
C260 a_n657_n197# a_591_131# 0.00fF
C261 a_n753_131# a_n705_n100# 0.00fF
C262 a_n369_131# a_n81_n197# 0.00fF
C263 a_n321_n100# a_n801_n100# 0.01fF
C264 a_n417_n100# a_n705_n100# 0.02fF
C265 a_543_n100# a_n129_n100# 0.01fF
C266 a_n513_n100# a_n609_n100# 0.09fF
C267 a_639_n100# a_n513_n100# 0.01fF
C268 a_n177_131# a_n369_131# 0.04fF
C269 a_n753_131# a_n801_n100# 0.00fF
C270 a_n417_n100# a_n801_n100# 0.02fF
C271 a_n513_n100# a_n705_n100# 0.04fF
C272 a_n465_n197# a_n753_131# 0.00fF
C273 a_n753_131# a_687_n197# 0.00fF
C274 a_n465_n197# a_n417_n100# 0.00fF
C275 a_n513_n100# a_n801_n100# 0.02fF
C276 a_351_n100# a_n129_n100# 0.01fF
C277 a_n753_131# a_495_n197# 0.00fF
C278 a_n465_n197# a_n513_n100# 0.00fF
C279 a_255_n100# a_n129_n100# 0.02fF
C280 a_15_131# a_n81_n197# 0.01fF
C281 a_n561_131# a_399_131# 0.01fF
C282 w_n1031_n319# a_n225_n100# 0.04fF
C283 a_n177_131# a_15_131# 0.04fF
C284 w_n1031_n319# a_n321_n100# 0.05fF
C285 w_n1031_n319# a_n753_131# 0.17fF
C286 w_n1031_n319# a_n417_n100# 0.05fF
C287 w_n1031_n319# a_n513_n100# 0.05fF
C288 a_n273_n197# a_399_131# 0.00fF
C289 a_n273_n197# a_n561_131# 0.00fF
C290 a_n465_n197# a_207_131# 0.00fF
C291 a_207_131# a_687_n197# 0.00fF
C292 a_207_131# a_495_n197# 0.00fF
C293 a_n465_n197# a_n369_131# 0.01fF
C294 a_n369_131# a_687_n197# 0.00fF
C295 a_n369_131# a_495_n197# 0.00fF
C296 a_n33_n100# a_n225_n100# 0.04fF
C297 a_n225_n100# a_735_n100# 0.01fF
C298 w_n1031_n319# a_207_131# 0.12fF
C299 a_n33_n100# a_n321_n100# 0.02fF
C300 a_n321_n100# a_735_n100# 0.01fF
C301 a_n465_n197# a_15_131# 0.00fF
C302 a_15_131# a_687_n197# 0.00fF
C303 a_n33_n100# a_n417_n100# 0.02fF
C304 a_n369_131# w_n1031_n319# 0.13fF
C305 a_n417_n100# a_735_n100# 0.01fF
C306 a_15_131# a_495_n197# 0.00fF
C307 a_n33_n100# a_n513_n100# 0.01fF
C308 a_n513_n100# a_735_n100# 0.00fF
C309 w_n1031_n319# a_15_131# 0.12fF
C310 a_447_n100# a_n609_n100# 0.01fF
C311 a_639_n100# a_447_n100# 0.04fF
C312 a_447_n100# a_n705_n100# 0.01fF
C313 a_543_n100# a_n609_n100# 0.01fF
C314 a_639_n100# a_543_n100# 0.09fF
C315 a_447_n100# a_n801_n100# 0.00fF
C316 a_543_n100# a_n705_n100# 0.00fF
C317 a_447_n100# a_495_n197# 0.00fF
C318 a_639_n100# a_351_n100# 0.02fF
C319 a_543_n100# a_n801_n100# 0.00fF
C320 a_351_n100# a_n609_n100# 0.01fF
C321 w_n1031_n319# VSUBS 3.95fF
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
C0 VPB VPWR 0.24fF
C1 VPWR VGND 0.06fF
C2 VPB X 0.00fF
C3 VPWR X 0.30fF
C4 VGND X 0.19fF
C5 a_27_47# VPB 0.12fF
C6 a_27_47# VPWR 0.24fF
C7 a_27_47# VGND 0.19fF
C8 VPB A 0.10fF
C9 A VPWR 0.02fF
C10 a_27_47# X 0.26fF
C11 A VGND 0.02fF
C12 A X 0.01fF
C13 a_27_47# A 0.21fF
C14 VGND VNB 0.28fF
C15 X VNB 0.00fF
C16 VPWR VNB 0.08fF
C17 A VNB 0.13fF
C18 VPB VNB 0.43fF
C19 a_27_47# VNB 0.15fF
.ends

.subckt precharge_pmos sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131#
+ VSUBS
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ VSUBS sky130_fd_pr__pfet_01v8_VCG74W
C0 sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319# VSUBS 3.95fF
.ends

.subckt current_tail a_543_n100# a_159_n100# a_n609_n100# a_n1569_n100# a_n705_n100#
+ a_255_n100# a_1407_n100# a_351_n100# a_n417_n100# a_n801_n100# a_1503_n100# a_1119_n100#
+ a_n1377_n100# a_n129_n100# a_n513_n100# a_1215_n100# a_63_n100# a_n1089_n100# a_n1473_n100#
+ a_n225_n100# a_1311_n100# a_927_n100# a_n1185_n100# a_n321_n100# a_1023_n100# a_639_n100#
+ a_n1281_n100# a_735_n100# a_n33_n100# a_n897_n100# a_831_n100# a_447_n100# a_n1521_122#
+ a_n993_n100# a_n1763_n274#
X0 a_n801_n100# a_n1521_122# a_n897_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n513_n100# a_n1521_122# a_n609_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n321_n100# a_n1521_122# a_n417_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n225_n100# a_n1521_122# a_n321_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_n897_n100# a_n1521_122# a_n993_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 a_n705_n100# a_n1521_122# a_n801_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n609_n100# a_n1521_122# a_n705_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n417_n100# a_n1521_122# a_n513_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n129_n100# a_n1521_122# a_n225_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_63_n100# a_n1521_122# a_n33_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_927_n100# a_n1521_122# a_831_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11 a_1023_n100# a_n1521_122# a_927_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1569_n100# a_n1763_n274# a_n1763_n274# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=6.2e+11p ps=5.24e+06u w=1e+06u l=150000u
X13 a_1119_n100# a_n1521_122# a_1023_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_1215_n100# a_n1521_122# a_1119_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_1311_n100# a_n1521_122# a_1215_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_1407_n100# a_n1521_122# a_1311_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_1503_n100# a_n1521_122# a_1407_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1763_n274# a_n1763_n274# a_1503_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n33_n100# a_n1521_122# a_n129_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_351_n100# a_n1521_122# a_255_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X21 a_159_n100# a_n1521_122# a_63_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22 a_255_n100# a_n1521_122# a_159_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_447_n100# a_n1521_122# a_351_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X24 a_543_n100# a_n1521_122# a_447_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X25 a_639_n100# a_n1521_122# a_543_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_735_n100# a_n1521_122# a_639_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_831_n100# a_n1521_122# a_735_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n1473_n100# a_n1521_122# a_n1569_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X29 a_n1377_n100# a_n1521_122# a_n1473_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X30 a_n1281_n100# a_n1521_122# a_n1377_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X31 a_n1185_n100# a_n1521_122# a_n1281_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X32 a_n1089_n100# a_n1521_122# a_n1185_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X33 a_n993_n100# a_n1521_122# a_n1089_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_735_n100# a_543_n100# 0.04fF
C1 a_831_n100# a_543_n100# 0.02fF
C2 a_543_n100# a_n801_n100# 0.00fF
C3 a_351_n100# a_n609_n100# 0.01fF
C4 a_639_n100# a_n897_n100# 0.00fF
C5 a_447_n100# a_n705_n100# 0.01fF
C6 a_255_n100# a_n609_n100# 0.01fF
C7 a_159_n100# a_n609_n100# 0.01fF
C8 a_63_n100# a_n513_n100# 0.01fF
C9 a_n1089_n100# a_n1473_n100# 0.02fF
C10 a_447_n100# a_n129_n100# 0.01fF
C11 a_n33_n100# a_n513_n100# 0.01fF
C12 a_1503_n100# a_1215_n100# 0.02fF
C13 a_1215_n100# a_1023_n100# 0.04fF
C14 a_1215_n100# a_927_n100# 0.02fF
C15 a_735_n100# a_n609_n100# 0.00fF
C16 a_831_n100# a_n609_n100# 0.00fF
C17 a_n417_n100# a_n993_n100# 0.01fF
C18 a_n513_n100# a_n897_n100# 0.02fF
C19 a_n609_n100# a_n801_n100# 0.04fF
C20 a_n321_n100# a_n1089_n100# 0.01fF
C21 a_n129_n100# a_n705_n100# 0.01fF
C22 a_1407_n100# a_63_n100# 0.00fF
C23 a_1215_n100# a_543_n100# 0.01fF
C24 a_63_n100# a_n225_n100# 0.02fF
C25 a_1311_n100# a_63_n100# 0.00fF
C26 a_1407_n100# a_n33_n100# 0.00fF
C27 a_1311_n100# a_n33_n100# 0.00fF
C28 a_n33_n100# a_n225_n100# 0.04fF
C29 a_n417_n100# a_n1473_n100# 0.01fF
C30 a_n225_n100# a_n897_n100# 0.01fF
C31 a_n321_n100# a_n417_n100# 0.09fF
C32 a_1119_n100# a_351_n100# 0.01fF
C33 a_351_n100# a_255_n100# 0.09fF
C34 a_n1089_n100# a_n1281_n100# 0.04fF
C35 a_n1089_n100# a_n1185_n100# 0.09fF
C36 a_351_n100# a_159_n100# 0.04fF
C37 a_447_n100# a_63_n100# 0.02fF
C38 a_1119_n100# a_255_n100# 0.01fF
C39 a_n1089_n100# a_n1377_n100# 0.02fF
C40 a_n609_n100# a_n1569_n100# 0.01fF
C41 a_255_n100# a_159_n100# 0.09fF
C42 a_447_n100# a_n33_n100# 0.01fF
C43 a_1119_n100# a_159_n100# 0.01fF
C44 a_255_n100# a_n1521_122# 0.03fF
C45 a_735_n100# a_351_n100# 0.02fF
C46 a_831_n100# a_351_n100# 0.01fF
C47 a_543_n100# a_n993_n100# 0.00fF
C48 a_447_n100# a_n897_n100# 0.00fF
C49 a_351_n100# a_n801_n100# 0.01fF
C50 a_735_n100# a_255_n100# 0.01fF
C51 a_1119_n100# a_735_n100# 0.02fF
C52 a_831_n100# a_255_n100# 0.01fF
C53 a_1119_n100# a_831_n100# 0.02fF
C54 a_255_n100# a_n801_n100# 0.01fF
C55 a_735_n100# a_159_n100# 0.01fF
C56 a_831_n100# a_159_n100# 0.01fF
C57 a_831_n100# a_n1521_122# 0.03fF
C58 a_159_n100# a_n801_n100# 0.01fF
C59 a_63_n100# a_n705_n100# 0.01fF
C60 a_1023_n100# a_n321_n100# 0.00fF
C61 a_n33_n100# a_n705_n100# 0.01fF
C62 a_927_n100# a_n321_n100# 0.00fF
C63 a_831_n100# a_735_n100# 0.09fF
C64 a_735_n100# a_n801_n100# 0.00fF
C65 a_63_n100# a_n129_n100# 0.04fF
C66 a_831_n100# a_n801_n100# 0.00fF
C67 a_n417_n100# a_n1281_n100# 0.01fF
C68 a_n513_n100# a_n1089_n100# 0.01fF
C69 a_n609_n100# a_n993_n100# 0.02fF
C70 a_n417_n100# a_n1185_n100# 0.01fF
C71 a_n705_n100# a_n897_n100# 0.04fF
C72 a_n33_n100# a_n129_n100# 0.09fF
C73 a_n417_n100# a_n1377_n100# 0.01fF
C74 a_n129_n100# a_n897_n100# 0.01fF
C75 a_543_n100# a_n321_n100# 0.01fF
C76 a_639_n100# a_n417_n100# 0.01fF
C77 a_1215_n100# a_351_n100# 0.01fF
C78 a_1215_n100# a_255_n100# 0.01fF
C79 a_1215_n100# a_1119_n100# 0.09fF
C80 a_n609_n100# a_n1473_n100# 0.01fF
C81 a_1215_n100# a_159_n100# 0.01fF
C82 a_1215_n100# a_n1521_122# 0.03fF
C83 a_n225_n100# a_n1089_n100# 0.01fF
C84 a_n321_n100# a_n609_n100# 0.02fF
C85 a_n417_n100# a_n513_n100# 0.09fF
C86 a_1215_n100# a_735_n100# 0.01fF
C87 a_1215_n100# a_831_n100# 0.02fF
C88 a_1503_n100# a_639_n100# 0.01fF
C89 a_n801_n100# a_n1569_n100# 0.01fF
C90 a_1023_n100# a_639_n100# 0.02fF
C91 a_927_n100# a_639_n100# 0.02fF
C92 a_63_n100# a_n33_n100# 0.09fF
C93 a_447_n100# a_n1089_n100# 0.00fF
C94 a_351_n100# a_n993_n100# 0.00fF
C95 a_255_n100# a_n993_n100# 0.00fF
C96 a_159_n100# a_n993_n100# 0.01fF
C97 a_63_n100# a_n897_n100# 0.01fF
C98 a_1023_n100# a_n513_n100# 0.00fF
C99 a_n33_n100# a_n897_n100# 0.01fF
C100 a_n225_n100# a_n417_n100# 0.04fF
C101 a_927_n100# a_n513_n100# 0.00fF
C102 a_639_n100# a_543_n100# 0.09fF
C103 a_n609_n100# a_n1281_n100# 0.01fF
C104 a_n705_n100# a_n1089_n100# 0.02fF
C105 a_n609_n100# a_n1185_n100# 0.01fF
C106 a_n801_n100# a_n993_n100# 0.04fF
C107 a_n609_n100# a_n1377_n100# 0.01fF
C108 a_159_n100# a_n1473_n100# 0.00fF
C109 a_n1473_n100# a_n1521_122# 0.03fF
C110 a_n129_n100# a_n1089_n100# 0.01fF
C111 a_639_n100# a_n609_n100# 0.00fF
C112 a_1503_n100# a_1407_n100# 0.09fF
C113 a_543_n100# a_n513_n100# 0.01fF
C114 a_351_n100# a_n321_n100# 0.01fF
C115 a_447_n100# a_n417_n100# 0.01fF
C116 a_1407_n100# a_1023_n100# 0.02fF
C117 a_1503_n100# a_1311_n100# 0.04fF
C118 a_1119_n100# a_n321_n100# 0.00fF
C119 a_255_n100# a_n321_n100# 0.01fF
C120 a_1023_n100# a_n225_n100# 0.00fF
C121 a_1407_n100# a_927_n100# 0.01fF
C122 a_1311_n100# a_1023_n100# 0.02fF
C123 a_159_n100# a_n321_n100# 0.01fF
C124 a_927_n100# a_n225_n100# 0.01fF
C125 a_n801_n100# a_n1473_n100# 0.01fF
C126 a_1311_n100# a_927_n100# 0.02fF
C127 a_n321_n100# a_n1521_122# 0.03fF
C128 a_735_n100# a_n321_n100# 0.01fF
C129 a_831_n100# a_n321_n100# 0.01fF
C130 a_n321_n100# a_n801_n100# 0.01fF
C131 a_n513_n100# a_n609_n100# 0.09fF
C132 a_n417_n100# a_n705_n100# 0.02fF
C133 a_1407_n100# a_543_n100# 0.01fF
C134 a_1503_n100# a_447_n100# 0.01fF
C135 a_1023_n100# a_447_n100# 0.01fF
C136 a_n993_n100# a_n1569_n100# 0.01fF
C137 a_543_n100# a_n225_n100# 0.01fF
C138 a_1311_n100# a_543_n100# 0.01fF
C139 a_927_n100# a_447_n100# 0.01fF
C140 a_n129_n100# a_n417_n100# 0.02fF
C141 a_351_n100# a_n1281_n100# 0.00fF
C142 a_351_n100# a_n1185_n100# 0.00fF
C143 a_255_n100# a_n1281_n100# 0.00fF
C144 a_255_n100# a_n1185_n100# 0.00fF
C145 a_255_n100# a_n1377_n100# 0.00fF
C146 a_159_n100# a_n1281_n100# 0.00fF
C147 a_n1281_n100# a_n1521_122# 0.03fF
C148 a_63_n100# a_n1089_n100# 0.01fF
C149 a_159_n100# a_n1185_n100# 0.00fF
C150 a_159_n100# a_n1377_n100# 0.00fF
C151 a_n1473_n100# a_n1569_n100# 0.09fF
C152 a_n33_n100# a_n1089_n100# 0.01fF
C153 a_n225_n100# a_n609_n100# 0.02fF
C154 a_927_n100# a_n705_n100# 0.00fF
C155 a_543_n100# a_447_n100# 0.09fF
C156 a_639_n100# a_351_n100# 0.02fF
C157 a_639_n100# a_255_n100# 0.02fF
C158 a_1119_n100# a_639_n100# 0.01fF
C159 a_1503_n100# a_n129_n100# 0.00fF
C160 a_n801_n100# a_n1281_n100# 0.01fF
C161 a_1215_n100# a_n321_n100# 0.00fF
C162 a_1023_n100# a_n129_n100# 0.01fF
C163 a_n897_n100# a_n1089_n100# 0.04fF
C164 a_n801_n100# a_n1185_n100# 0.02fF
C165 a_639_n100# a_159_n100# 0.01fF
C166 a_639_n100# a_n1521_122# 0.03fF
C167 a_n801_n100# a_n1377_n100# 0.01fF
C168 a_n321_n100# a_n1569_n100# 0.00fF
C169 a_927_n100# a_n129_n100# 0.01fF
C170 a_735_n100# a_639_n100# 0.09fF
C171 a_831_n100# a_639_n100# 0.04fF
C172 a_351_n100# a_n513_n100# 0.01fF
C173 a_543_n100# a_n705_n100# 0.00fF
C174 a_447_n100# a_n609_n100# 0.01fF
C175 a_639_n100# a_n801_n100# 0.00fF
C176 a_255_n100# a_n513_n100# 0.01fF
C177 a_1119_n100# a_n513_n100# 0.00fF
C178 a_63_n100# a_n417_n100# 0.01fF
C179 a_159_n100# a_n513_n100# 0.01fF
C180 a_n513_n100# a_n1521_122# 0.03fF
C181 a_n993_n100# a_n1473_n100# 0.01fF
C182 a_543_n100# a_n129_n100# 0.01fF
C183 a_n33_n100# a_n417_n100# 0.02fF
C184 a_735_n100# a_n513_n100# 0.00fF
C185 a_831_n100# a_n513_n100# 0.00fF
C186 a_n513_n100# a_n801_n100# 0.02fF
C187 a_n609_n100# a_n705_n100# 0.09fF
C188 a_n321_n100# a_n993_n100# 0.01fF
C189 a_n417_n100# a_n897_n100# 0.01fF
C190 a_n1281_n100# a_n1569_n100# 0.02fF
C191 a_1407_n100# a_351_n100# 0.01fF
C192 a_n1185_n100# a_n1569_n100# 0.02fF
C193 a_351_n100# a_n225_n100# 0.01fF
C194 a_n1377_n100# a_n1569_n100# 0.04fF
C195 a_1407_n100# a_255_n100# 0.01fF
C196 a_1311_n100# a_351_n100# 0.01fF
C197 a_1407_n100# a_1119_n100# 0.02fF
C198 a_n129_n100# a_n609_n100# 0.01fF
C199 a_255_n100# a_n225_n100# 0.01fF
C200 a_1311_n100# a_255_n100# 0.01fF
C201 a_1119_n100# a_n225_n100# 0.00fF
C202 a_1407_n100# a_159_n100# 0.00fF
C203 a_1311_n100# a_1119_n100# 0.04fF
C204 a_1503_n100# a_63_n100# 0.00fF
C205 a_1023_n100# a_63_n100# 0.01fF
C206 a_1407_n100# a_n1521_122# 0.03fF
C207 a_159_n100# a_n225_n100# 0.02fF
C208 a_1215_n100# a_639_n100# 0.01fF
C209 a_1311_n100# a_159_n100# 0.01fF
C210 a_1503_n100# a_n33_n100# 0.00fF
C211 a_927_n100# a_63_n100# 0.01fF
C212 a_1023_n100# a_n33_n100# 0.01fF
C213 a_927_n100# a_n33_n100# 0.01fF
C214 a_n321_n100# a_n1473_n100# 0.01fF
C215 a_1407_n100# a_735_n100# 0.01fF
C216 a_1407_n100# a_831_n100# 0.01fF
C217 a_1311_n100# a_735_n100# 0.01fF
C218 a_735_n100# a_n225_n100# 0.01fF
C219 a_831_n100# a_n225_n100# 0.01fF
C220 a_1311_n100# a_831_n100# 0.01fF
C221 a_n225_n100# a_n801_n100# 0.01fF
C222 a_447_n100# a_351_n100# 0.09fF
C223 a_447_n100# a_255_n100# 0.04fF
C224 a_1119_n100# a_447_n100# 0.01fF
C225 a_n993_n100# a_n1281_n100# 0.02fF
C226 a_n993_n100# a_n1185_n100# 0.04fF
C227 a_447_n100# a_159_n100# 0.02fF
C228 a_543_n100# a_63_n100# 0.01fF
C229 a_447_n100# a_n1521_122# 0.03fF
C230 a_n993_n100# a_n1377_n100# 0.02fF
C231 a_n513_n100# a_n1569_n100# 0.01fF
C232 a_543_n100# a_n33_n100# 0.01fF
C233 a_735_n100# a_447_n100# 0.02fF
C234 a_831_n100# a_447_n100# 0.02fF
C235 a_543_n100# a_n897_n100# 0.00fF
C236 a_447_n100# a_n801_n100# 0.00fF
C237 a_639_n100# a_n993_n100# 0.00fF
C238 a_351_n100# a_n705_n100# 0.01fF
C239 a_255_n100# a_n705_n100# 0.01fF
C240 a_n1281_n100# a_n1473_n100# 0.04fF
C241 a_159_n100# a_n705_n100# 0.01fF
C242 a_63_n100# a_n609_n100# 0.01fF
C243 a_n705_n100# a_n1521_122# 0.03fF
C244 a_n1185_n100# a_n1473_n100# 0.02fF
C245 a_n1377_n100# a_n1473_n100# 0.09fF
C246 a_351_n100# a_n129_n100# 0.01fF
C247 a_1407_n100# a_1215_n100# 0.04fF
C248 a_n33_n100# a_n609_n100# 0.01fF
C249 a_255_n100# a_n129_n100# 0.02fF
C250 a_1215_n100# a_n225_n100# 0.00fF
C251 a_1119_n100# a_n129_n100# 0.00fF
C252 a_1311_n100# a_1215_n100# 0.09fF
C253 a_159_n100# a_n129_n100# 0.02fF
C254 a_735_n100# a_n705_n100# 0.00fF
C255 a_n225_n100# a_n1569_n100# 0.00fF
C256 a_831_n100# a_n705_n100# 0.00fF
C257 a_n129_n100# a_n1521_122# 0.03fF
C258 a_n321_n100# a_n1281_n100# 0.01fF
C259 a_n417_n100# a_n1089_n100# 0.01fF
C260 a_n513_n100# a_n993_n100# 0.01fF
C261 a_n609_n100# a_n897_n100# 0.02fF
C262 a_n321_n100# a_n1185_n100# 0.01fF
C263 a_n705_n100# a_n801_n100# 0.09fF
C264 a_n321_n100# a_n1377_n100# 0.01fF
C265 a_735_n100# a_n129_n100# 0.01fF
C266 a_831_n100# a_n129_n100# 0.01fF
C267 a_n129_n100# a_n801_n100# 0.01fF
C268 a_639_n100# a_n321_n100# 0.01fF
C269 a_1215_n100# a_447_n100# 0.01fF
C270 a_n513_n100# a_n1473_n100# 0.01fF
C271 a_n225_n100# a_n993_n100# 0.01fF
C272 a_n321_n100# a_n513_n100# 0.04fF
C273 a_n1185_n100# a_n1281_n100# 0.09fF
C274 a_n1281_n100# a_n1377_n100# 0.09fF
C275 a_351_n100# a_63_n100# 0.02fF
C276 a_n1185_n100# a_n1377_n100# 0.04fF
C277 a_n705_n100# a_n1569_n100# 0.01fF
C278 a_1119_n100# a_63_n100# 0.01fF
C279 a_255_n100# a_63_n100# 0.04fF
C280 a_351_n100# a_n33_n100# 0.02fF
C281 a_159_n100# a_63_n100# 0.09fF
C282 a_255_n100# a_n33_n100# 0.02fF
C283 a_63_n100# a_n1521_122# 0.03fF
C284 a_1119_n100# a_n33_n100# 0.01fF
C285 a_1215_n100# a_n129_n100# 0.00fF
C286 a_159_n100# a_n33_n100# 0.04fF
C287 a_n225_n100# a_n1473_n100# 0.00fF
C288 a_n129_n100# a_n1569_n100# 0.00fF
C289 a_543_n100# a_n1089_n100# 0.00fF
C290 a_351_n100# a_n897_n100# 0.00fF
C291 a_447_n100# a_n993_n100# 0.00fF
C292 a_255_n100# a_n897_n100# 0.01fF
C293 a_735_n100# a_63_n100# 0.01fF
C294 a_831_n100# a_63_n100# 0.01fF
C295 a_159_n100# a_n897_n100# 0.01fF
C296 a_63_n100# a_n801_n100# 0.01fF
C297 a_n897_n100# a_n1521_122# 0.03fF
C298 a_735_n100# a_n33_n100# 0.01fF
C299 a_1023_n100# a_n417_n100# 0.00fF
C300 a_831_n100# a_n33_n100# 0.01fF
C301 a_n225_n100# a_n321_n100# 0.09fF
C302 a_n33_n100# a_n801_n100# 0.01fF
C303 a_1311_n100# a_n321_n100# 0.00fF
C304 a_927_n100# a_n417_n100# 0.00fF
C305 a_735_n100# a_n897_n100# 0.00fF
C306 a_n513_n100# a_n1281_n100# 0.01fF
C307 a_n513_n100# a_n1185_n100# 0.01fF
C308 a_n609_n100# a_n1089_n100# 0.01fF
C309 a_n801_n100# a_n897_n100# 0.09fF
C310 a_n705_n100# a_n993_n100# 0.02fF
C311 a_n513_n100# a_n1377_n100# 0.01fF
C312 a_n129_n100# a_n993_n100# 0.01fF
C313 a_639_n100# a_n513_n100# 0.01fF
C314 a_543_n100# a_n417_n100# 0.01fF
C315 a_447_n100# a_n321_n100# 0.01fF
C316 a_1503_n100# a_1023_n100# 0.01fF
C317 a_1503_n100# a_927_n100# 0.01fF
C318 a_1023_n100# a_927_n100# 0.09fF
C319 a_n705_n100# a_n1473_n100# 0.01fF
C320 a_1215_n100# a_63_n100# 0.01fF
C321 a_n225_n100# a_n1281_n100# 0.01fF
C322 a_63_n100# a_n1569_n100# 0.00fF
C323 a_1215_n100# a_n33_n100# 0.00fF
C324 a_n225_n100# a_n1185_n100# 0.01fF
C325 a_n129_n100# a_n1473_n100# 0.00fF
C326 a_n33_n100# a_n1569_n100# 0.00fF
C327 a_n225_n100# a_n1377_n100# 0.01fF
C328 a_n417_n100# a_n609_n100# 0.04fF
C329 a_n321_n100# a_n705_n100# 0.02fF
C330 a_1503_n100# a_543_n100# 0.01fF
C331 a_1407_n100# a_639_n100# 0.01fF
C332 a_1023_n100# a_543_n100# 0.01fF
C333 a_n897_n100# a_n1569_n100# 0.01fF
C334 a_1311_n100# a_639_n100# 0.01fF
C335 a_639_n100# a_n225_n100# 0.01fF
C336 a_n129_n100# a_n321_n100# 0.04fF
C337 a_927_n100# a_543_n100# 0.02fF
C338 a_351_n100# a_n1089_n100# 0.00fF
C339 a_447_n100# a_n1185_n100# 0.00fF
C340 a_255_n100# a_n1089_n100# 0.00fF
C341 a_63_n100# a_n993_n100# 0.01fF
C342 a_159_n100# a_n1089_n100# 0.00fF
C343 a_n1089_n100# a_n1521_122# 0.03fF
C344 a_1023_n100# a_n609_n100# 0.00fF
C345 a_n33_n100# a_n993_n100# 0.01fF
C346 a_n225_n100# a_n513_n100# 0.02fF
C347 a_927_n100# a_n609_n100# 0.00fF
C348 a_639_n100# a_447_n100# 0.04fF
C349 a_n705_n100# a_n1281_n100# 0.01fF
C350 a_n801_n100# a_n1089_n100# 0.02fF
C351 a_n705_n100# a_n1185_n100# 0.01fF
C352 a_n897_n100# a_n993_n100# 0.09fF
C353 a_n705_n100# a_n1377_n100# 0.01fF
C354 a_n129_n100# a_n1281_n100# 0.01fF
C355 a_63_n100# a_n1473_n100# 0.00fF
C356 a_n129_n100# a_n1185_n100# 0.01fF
C357 a_n33_n100# a_n1473_n100# 0.00fF
C358 a_n129_n100# a_n1377_n100# 0.00fF
C359 a_543_n100# a_n609_n100# 0.01fF
C360 a_351_n100# a_n417_n100# 0.01fF
C361 a_447_n100# a_n513_n100# 0.01fF
C362 a_639_n100# a_n705_n100# 0.00fF
C363 a_1407_n100# a_n225_n100# 0.00fF
C364 a_1407_n100# a_1311_n100# 0.09fF
C365 a_255_n100# a_n417_n100# 0.01fF
C366 a_1119_n100# a_n417_n100# 0.00fF
C367 a_1311_n100# a_n225_n100# 0.00fF
C368 a_n897_n100# a_n1473_n100# 0.01fF
C369 a_159_n100# a_n417_n100# 0.01fF
C370 a_63_n100# a_n321_n100# 0.02fF
C371 a_639_n100# a_n129_n100# 0.01fF
C372 a_n33_n100# a_n321_n100# 0.02fF
C373 a_735_n100# a_n417_n100# 0.01fF
C374 a_831_n100# a_n417_n100# 0.00fF
C375 a_n513_n100# a_n705_n100# 0.04fF
C376 a_n321_n100# a_n897_n100# 0.01fF
C377 a_n417_n100# a_n801_n100# 0.02fF
C378 a_1407_n100# a_447_n100# 0.01fF
C379 a_1503_n100# a_351_n100# 0.01fF
C380 a_n1089_n100# a_n1569_n100# 0.01fF
C381 a_1023_n100# a_351_n100# 0.01fF
C382 a_1311_n100# a_447_n100# 0.01fF
C383 a_1503_n100# a_255_n100# 0.00fF
C384 a_447_n100# a_n225_n100# 0.01fF
C385 a_1503_n100# a_1119_n100# 0.02fF
C386 a_1119_n100# a_1023_n100# 0.09fF
C387 a_927_n100# a_351_n100# 0.01fF
C388 a_1023_n100# a_255_n100# 0.01fF
C389 a_n129_n100# a_n513_n100# 0.02fF
C390 a_1503_n100# a_159_n100# 0.00fF
C391 a_927_n100# a_255_n100# 0.01fF
C392 a_1023_n100# a_159_n100# 0.01fF
C393 a_1119_n100# a_927_n100# 0.04fF
C394 a_1023_n100# a_n1521_122# 0.03fF
C395 a_927_n100# a_159_n100# 0.01fF
C396 a_1503_n100# a_735_n100# 0.01fF
C397 a_1023_n100# a_735_n100# 0.02fF
C398 a_63_n100# a_n1281_n100# 0.00fF
C399 a_1503_n100# a_831_n100# 0.01fF
C400 a_1023_n100# a_831_n100# 0.04fF
C401 a_63_n100# a_n1185_n100# 0.00fF
C402 a_927_n100# a_735_n100# 0.04fF
C403 a_n33_n100# a_n1281_n100# 0.00fF
C404 a_63_n100# a_n1377_n100# 0.00fF
C405 a_n33_n100# a_n1185_n100# 0.01fF
C406 a_927_n100# a_831_n100# 0.09fF
C407 a_n225_n100# a_n705_n100# 0.01fF
C408 a_543_n100# a_351_n100# 0.04fF
C409 a_n33_n100# a_n1377_n100# 0.00fF
C410 a_543_n100# a_255_n100# 0.02fF
C411 a_1407_n100# a_n129_n100# 0.00fF
C412 a_1119_n100# a_543_n100# 0.01fF
C413 a_n897_n100# a_n1281_n100# 0.02fF
C414 a_1215_n100# a_n417_n100# 0.00fF
C415 a_n993_n100# a_n1089_n100# 0.09fF
C416 a_n897_n100# a_n1185_n100# 0.02fF
C417 a_n129_n100# a_n225_n100# 0.09fF
C418 a_639_n100# a_63_n100# 0.01fF
C419 a_543_n100# a_159_n100# 0.02fF
C420 a_1311_n100# a_n129_n100# 0.00fF
C421 a_n417_n100# a_n1569_n100# 0.01fF
C422 a_n897_n100# a_n1377_n100# 0.01fF
C423 a_639_n100# a_n33_n100# 0.01fF
C424 a_1503_n100# a_n1763_n274# 0.14fF
C425 a_1407_n100# a_n1763_n274# 0.07fF
C426 a_1311_n100# a_n1763_n274# 0.06fF
C427 a_1215_n100# a_n1763_n274# 0.05fF
C428 a_1119_n100# a_n1763_n274# 0.04fF
C429 a_1023_n100# a_n1763_n274# 0.04fF
C430 a_927_n100# a_n1763_n274# 0.03fF
C431 a_831_n100# a_n1763_n274# 0.03fF
C432 a_735_n100# a_n1763_n274# 0.03fF
C433 a_639_n100# a_n1763_n274# 0.03fF
C434 a_543_n100# a_n1763_n274# 0.03fF
C435 a_447_n100# a_n1763_n274# 0.03fF
C436 a_351_n100# a_n1763_n274# 0.03fF
C437 a_255_n100# a_n1763_n274# 0.03fF
C438 a_159_n100# a_n1763_n274# 0.03fF
C439 a_63_n100# a_n1763_n274# 0.02fF
C440 a_n33_n100# a_n1763_n274# 0.03fF
C441 a_n129_n100# a_n1763_n274# 0.02fF
C442 a_n225_n100# a_n1763_n274# 0.03fF
C443 a_n321_n100# a_n1763_n274# 0.03fF
C444 a_n417_n100# a_n1763_n274# 0.03fF
C445 a_n513_n100# a_n1763_n274# 0.03fF
C446 a_n609_n100# a_n1763_n274# 0.03fF
C447 a_n705_n100# a_n1763_n274# 0.03fF
C448 a_n801_n100# a_n1763_n274# 0.03fF
C449 a_n897_n100# a_n1763_n274# 0.03fF
C450 a_n993_n100# a_n1763_n274# 0.03fF
C451 a_n1089_n100# a_n1763_n274# 0.04fF
C452 a_n1185_n100# a_n1763_n274# 0.04fF
C453 a_n1281_n100# a_n1763_n274# 0.05fF
C454 a_n1377_n100# a_n1763_n274# 0.06fF
C455 a_n1473_n100# a_n1763_n274# 0.08fF
C456 a_n1569_n100# a_n1763_n274# 0.15fF
C457 a_n1521_122# a_n1763_n274# 3.88fF
.ends

.subckt sky130_fd_pr__nfet_01v8_J3WY8C a_n4080_n100# a_n1188_122# a_282_n188# a_n978_n188#
+ a_1542_n188# a_n3918_n188# a_3432_122# a_1752_122# a_n3708_122# a_2382_n188# a_4228_n100#
+ a_n2028_122# a_n1818_n188# a_3222_n188# a_n348_122# a_n2658_n188# a_n3288_122# a_4062_n188#
+ a_72_122# a_n558_n188# a_n3498_n188# a_1122_n188# a_912_122# a_n4172_n100# a_3852_122#
+ a_n1398_n188# a_2172_122# a_n4128_122# a_n2448_122# a_492_122# a_n768_122# a_n2238_n188#
+ a_n138_n188# a_n3078_n188# a_1962_n188# a_702_n188# a_3012_122# a_1332_122# a_n1608_122#
+ a_n4382_n100# a_2802_n188# a_2592_122# a_3642_n188# a_n2868_122# VSUBS
X0 a_n4080_n100# a_n1398_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=1.24e+13p pd=1.048e+08u as=1.24e+13p ps=1.048e+08u w=1e+06u l=150000u
X1 a_n4080_n100# a_1332_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n4080_n100# a_n2868_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n4080_n100# a_2802_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n4080_n100# a_n3288_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n4080_n100# a_3222_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n4080_n100# a_72_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n4080_n100# a_n1608_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n4080_n100# a_1542_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n4080_n100# a_n138_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n4080_n100# a_282_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n4080_n100# a_n3498_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n4080_n100# a_3432_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n4080_n100# a_n1818_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n4080_n100# a_1752_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n4080_n100# a_492_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n4080_n100# a_2172_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n4080_n100# a_n3708_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n4080_n100# a_n348_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n4080_n100# a_3642_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n4080_n100# a_4062_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n4080_n100# a_n2028_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n4080_n100# a_1962_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n4080_n100# a_702_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n4080_n100# a_n3918_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n4080_n100# a_n558_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n4080_n100# a_3852_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_4228_n100# a_4228_n100# a_4228_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X28 a_n4080_n100# a_n2238_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_n4080_n100# a_n768_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n4080_n100# a_912_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n4080_n100# a_n4128_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_n4080_n100# a_n2448_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_n4080_n100# a_2382_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_n4080_n100# a_n978_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n4382_n100# a_n4382_n100# a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X36 a_n4080_n100# a_n1188_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_n4080_n100# a_1122_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n4080_n100# a_n2658_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_n4080_n100# a_2592_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_n4080_n100# a_n3078_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_n4080_n100# a_3012_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_3642_n188# a_n4172_n100# 0.02fF
C1 a_702_n188# a_n558_n188# 0.00fF
C2 a_n2028_122# a_n3078_n188# 0.00fF
C3 a_n2238_n188# a_n2658_n188# 0.01fF
C4 a_n1608_122# a_n2448_122# 0.01fF
C5 a_3012_122# a_1542_n188# 0.00fF
C6 a_282_n188# a_n978_n188# 0.00fF
C7 a_3222_n188# a_3012_122# 0.00fF
C8 a_3432_122# a_2802_n188# 0.00fF
C9 a_n4080_n100# a_2802_n188# 0.06fF
C10 a_n2658_n188# a_n3498_n188# 0.01fF
C11 a_282_n188# a_n768_122# 0.00fF
C12 a_2382_n188# a_1752_122# 0.00fF
C13 a_2172_122# a_n4172_n100# 0.06fF
C14 a_2592_122# a_1752_122# 0.01fF
C15 a_1962_n188# a_912_122# 0.00fF
C16 a_3852_122# a_2802_n188# 0.00fF
C17 a_n3918_n188# a_n4172_n100# 0.02fF
C18 a_1752_122# a_282_n188# 0.00fF
C19 a_282_n188# a_n1188_122# 0.00fF
C20 a_1542_n188# a_1332_122# 0.00fF
C21 a_912_122# a_n138_n188# 0.00fF
C22 a_3012_122# a_3642_n188# 0.00fF
C23 a_1542_n188# a_72_122# 0.00fF
C24 a_n3918_n188# a_n3708_122# 0.00fF
C25 a_n3288_122# a_n4382_n100# 0.00fF
C26 a_n3498_n188# a_n4128_122# 0.00fF
C27 a_282_n188# a_492_122# 0.00fF
C28 a_n2448_122# a_n3918_n188# 0.00fF
C29 a_n558_n188# a_n978_n188# 0.01fF
C30 a_3432_122# a_1962_n188# 0.00fF
C31 a_n4080_n100# a_1962_n188# 0.06fF
C32 a_n558_n188# a_n768_122# 0.00fF
C33 a_n4080_n100# a_n138_n188# 0.06fF
C34 a_n558_n188# a_n1398_n188# 0.01fF
C35 a_1122_n188# a_1332_122# 0.00fF
C36 a_1122_n188# a_72_122# 0.00fF
C37 a_n558_n188# a_n1188_122# 0.00fF
C38 a_n1818_n188# a_n2658_n188# 0.01fF
C39 a_n2238_n188# a_n3078_n188# 0.01fF
C40 a_2802_n188# a_n4172_n100# 0.02fF
C41 a_n1608_122# a_n2658_n188# 0.00fF
C42 a_n2238_n188# a_n2028_122# 0.00fF
C43 a_492_122# a_n558_n188# 0.00fF
C44 a_3012_122# a_2172_122# 0.01fF
C45 a_n4080_n100# a_n4382_n100# 0.14fF
C46 a_n3078_n188# a_n3498_n188# 0.01fF
C47 a_n2028_122# a_n3498_n188# 0.00fF
C48 a_2382_n188# a_912_122# 0.00fF
C49 a_702_n188# a_n768_122# 0.00fF
C50 a_1962_n188# a_n4172_n100# 0.02fF
C51 a_n138_n188# a_n4172_n100# 0.02fF
C52 a_912_122# a_282_n188# 0.00fF
C53 a_1752_122# a_702_n188# 0.00fF
C54 a_2172_122# a_1332_122# 0.01fF
C55 a_2802_n188# a_3012_122# 0.00fF
C56 a_3432_122# a_2382_n188# 0.00fF
C57 a_702_n188# a_492_122# 0.00fF
C58 a_n4080_n100# a_2382_n188# 0.06fF
C59 a_n2658_n188# a_n3918_n188# 0.00fF
C60 a_3432_122# a_2592_122# 0.01fF
C61 a_n4080_n100# a_2592_122# 0.02fF
C62 a_n4080_n100# a_282_n188# 0.06fF
C63 a_3852_122# a_2382_n188# 0.00fF
C64 a_n1398_n188# a_n2868_122# 0.00fF
C65 a_n4382_n100# a_n4172_n100# 0.21fF
C66 a_n1818_n188# a_n3078_n188# 0.00fF
C67 a_3852_122# a_2592_122# 0.00fF
C68 a_912_122# a_n558_n188# 0.00fF
C69 a_n1818_n188# a_n2028_122# 0.00fF
C70 a_n1608_122# a_n3078_n188# 0.00fF
C71 a_n1608_122# a_n2028_122# 0.01fF
C72 a_n3918_n188# a_n4128_122# 0.00fF
C73 a_n3708_122# a_n4382_n100# 0.00fF
C74 a_3012_122# a_1962_n188# 0.00fF
C75 a_2802_n188# a_1332_122# 0.00fF
C76 a_n978_n188# a_n768_122# 0.00fF
C77 a_4062_n188# a_3432_122# 0.00fF
C78 a_n978_n188# a_n1398_n188# 0.01fF
C79 a_n4080_n100# a_4062_n188# 0.06fF
C80 a_n4080_n100# a_n558_n188# 0.06fF
C81 a_1122_n188# a_n348_122# 0.00fF
C82 a_n768_122# a_n1398_n188# 0.00fF
C83 a_n978_n188# a_n1188_122# 0.00fF
C84 a_n348_122# a_n1818_n188# 0.00fF
C85 a_n2238_n188# a_n3498_n188# 0.00fF
C86 a_2382_n188# a_n4172_n100# 0.02fF
C87 a_3852_122# a_4062_n188# 0.00fF
C88 a_n348_122# a_n1608_122# 0.00fF
C89 a_n768_122# a_n1188_122# 0.01fF
C90 a_2592_122# a_n4172_n100# 0.06fF
C91 a_n1398_n188# a_n1188_122# 0.00fF
C92 a_492_122# a_n978_n188# 0.00fF
C93 a_282_n188# a_n4172_n100# 0.02fF
C94 a_492_122# a_n768_122# 0.00fF
C95 a_702_n188# a_912_122# 0.00fF
C96 a_1962_n188# a_1332_122# 0.00fF
C97 a_1752_122# a_492_122# 0.00fF
C98 a_3222_n188# a_4228_n100# 0.00fF
C99 a_n2868_122# a_n3288_122# 0.01fF
C100 a_n3078_n188# a_n3918_n188# 0.01fF
C101 a_1332_122# a_n138_n188# 0.00fF
C102 a_n138_n188# a_72_122# 0.00fF
C103 a_n4080_n100# a_702_n188# 0.06fF
C104 a_4062_n188# a_n4172_n100# 0.02fF
C105 a_n558_n188# a_n4172_n100# 0.02fF
C106 a_n1818_n188# a_n2238_n188# 0.01fF
C107 a_4228_n100# a_3642_n188# 0.00fF
C108 a_n1608_122# a_n2238_n188# 0.00fF
C109 a_3012_122# a_2382_n188# 0.00fF
C110 a_n2658_n188# a_n4382_n100# 0.00fF
C111 a_3012_122# a_2592_122# 0.01fF
C112 a_n4080_n100# a_n2868_122# 0.02fF
C113 a_n4382_n100# a_n4128_122# 0.00fF
C114 a_1752_122# a_912_122# 0.01fF
C115 a_702_n188# a_n4172_n100# 0.02fF
C116 a_2382_n188# a_1332_122# 0.00fF
C117 a_1542_n188# a_1122_n188# 0.01fF
C118 a_4062_n188# a_3012_122# 0.00fF
C119 a_2592_122# a_1332_122# 0.00fF
C120 a_n4080_n100# a_n978_n188# 0.06fF
C121 a_1332_122# a_282_n188# 0.00fF
C122 a_912_122# a_492_122# 0.01fF
C123 a_n4080_n100# a_n768_122# 0.02fF
C124 a_282_n188# a_72_122# 0.00fF
C125 a_n4080_n100# a_n1398_n188# 0.06fF
C126 a_n4080_n100# a_1752_122# 0.02fF
C127 a_n4080_n100# a_n1188_122# 0.02fF
C128 a_n2868_122# a_n4172_n100# 0.06fF
C129 a_n4080_n100# a_492_122# 0.02fF
C130 a_n1818_n188# a_n1608_122# 0.00fF
C131 a_3222_n188# a_3642_n188# 0.01fF
C132 a_n3498_n188# a_n3918_n188# 0.01fF
C133 a_n3078_n188# a_n4382_n100# 0.00fF
C134 a_n2868_122# a_n3708_122# 0.01fF
C135 a_2802_n188# a_4228_n100# 0.00fF
C136 a_n2448_122# a_n2868_122# 0.01fF
C137 a_n138_n188# a_n348_122# 0.00fF
C138 a_72_122# a_n558_n188# 0.00fF
C139 a_n978_n188# a_n4172_n100# 0.02fF
C140 a_2172_122# a_1542_n188# 0.00fF
C141 a_n768_122# a_n4172_n100# 0.06fF
C142 a_n1398_n188# a_n4172_n100# 0.02fF
C143 a_1752_122# a_n4172_n100# 0.06fF
C144 a_n1188_122# a_n4172_n100# 0.06fF
C145 a_n978_n188# a_n2448_122# 0.00fF
C146 a_3222_n188# a_2172_122# 0.00fF
C147 a_n4080_n100# a_n3288_122# 0.02fF
C148 a_2172_122# a_1122_n188# 0.00fF
C149 a_492_122# a_n4172_n100# 0.06fF
C150 a_n1398_n188# a_n2448_122# 0.00fF
C151 a_1332_122# a_702_n188# 0.00fF
C152 a_n1188_122# a_n2448_122# 0.00fF
C153 a_702_n188# a_72_122# 0.00fF
C154 a_2172_122# a_3642_n188# 0.00fF
C155 a_n4080_n100# a_912_122# 0.02fF
C156 a_2802_n188# a_1542_n188# 0.00fF
C157 a_3222_n188# a_2802_n188# 0.01fF
C158 a_282_n188# a_n348_122# 0.00fF
C159 a_n4080_n100# a_3432_122# 0.02fF
C160 a_n2658_n188# a_n2868_122# 0.00fF
C161 a_n558_n188# a_n2028_122# 0.00fF
C162 a_3012_122# a_1752_122# 0.00fF
C163 a_3852_122# a_3432_122# 0.01fF
C164 a_n4080_n100# a_3852_122# 0.02fF
C165 a_n3288_122# a_n4172_n100# 0.06fF
C166 a_1962_n188# a_1542_n188# 0.01fF
C167 a_2802_n188# a_3642_n188# 0.01fF
C168 a_n3498_n188# a_n4382_n100# 0.00fF
C169 a_n2868_122# a_n4128_122# 0.00fF
C170 a_n3288_122# a_n3708_122# 0.01fF
C171 a_n2448_122# a_n3288_122# 0.01fF
C172 a_n558_n188# a_n348_122# 0.00fF
C173 a_72_122# a_n978_n188# 0.00fF
C174 a_2592_122# a_4228_n100# 0.00fF
C175 a_912_122# a_n4172_n100# 0.06fF
C176 a_3222_n188# a_1962_n188# 0.00fF
C177 a_72_122# a_n768_122# 0.01fF
C178 a_1962_n188# a_1122_n188# 0.01fF
C179 a_72_122# a_n1398_n188# 0.00fF
C180 a_1752_122# a_1332_122# 0.01fF
C181 a_n1398_n188# a_n2658_n188# 0.00fF
C182 a_1122_n188# a_n138_n188# 0.00fF
C183 a_72_122# a_n1188_122# 0.00fF
C184 a_n1188_122# a_n2658_n188# 0.00fF
C185 a_3432_122# a_n4172_n100# 0.06fF
C186 a_n138_n188# a_n1608_122# 0.00fF
C187 a_1332_122# a_492_122# 0.01fF
C188 a_n4080_n100# a_n4172_n100# 15.77fF
C189 a_492_122# a_72_122# 0.01fF
C190 a_2802_n188# a_2172_122# 0.00fF
C191 a_3852_122# a_n4172_n100# 0.06fF
C192 a_n4080_n100# a_n3708_122# 0.02fF
C193 a_4062_n188# a_4228_n100# 0.00fF
C194 a_n4080_n100# a_n2448_122# 0.02fF
C195 a_n3078_n188# a_n2868_122# 0.00fF
C196 a_702_n188# a_n348_122# 0.00fF
C197 a_n2028_122# a_n2868_122# 0.01fF
C198 a_2382_n188# a_1542_n188# 0.01fF
C199 a_2592_122# a_1542_n188# 0.00fF
C200 a_1962_n188# a_2172_122# 0.00fF
C201 a_1542_n188# a_282_n188# 0.00fF
C202 a_3432_122# a_3012_122# 0.01fF
C203 a_3222_n188# a_2382_n188# 0.01fF
C204 a_n4080_n100# a_3012_122# 0.02fF
C205 a_n2658_n188# a_n3288_122# 0.00fF
C206 a_n978_n188# a_n2028_122# 0.00fF
C207 a_3222_n188# a_2592_122# 0.00fF
C208 a_2382_n188# a_1122_n188# 0.00fF
C209 a_n768_122# a_n2028_122# 0.00fF
C210 a_2592_122# a_1122_n188# 0.00fF
C211 a_3852_122# a_3012_122# 0.01fF
C212 a_n3708_122# a_n4172_n100# 0.06fF
C213 a_n1398_n188# a_n2028_122# 0.00fF
C214 a_1122_n188# a_282_n188# 0.01fF
C215 a_1332_122# a_912_122# 0.01fF
C216 a_n2448_122# a_n4172_n100# 0.06fF
C217 a_912_122# a_72_122# 0.01fF
C218 a_n1188_122# a_n2028_122# 0.01fF
C219 a_2382_n188# a_3642_n188# 0.00fF
C220 a_n3288_122# a_n4128_122# 0.01fF
C221 a_n3918_n188# a_n4382_n100# 0.01fF
C222 a_n2448_122# a_n3708_122# 0.00fF
C223 a_2592_122# a_3642_n188# 0.00fF
C224 a_n348_122# a_n978_n188# 0.00fF
C225 a_2802_n188# a_1962_n188# 0.01fF
C226 a_n348_122# a_n768_122# 0.01fF
C227 a_n4080_n100# a_1332_122# 0.02fF
C228 a_4062_n188# a_3222_n188# 0.01fF
C229 a_n4080_n100# a_72_122# 0.02fF
C230 a_n348_122# a_n1398_n188# 0.00fF
C231 a_n4080_n100# a_n2658_n188# 0.06fF
C232 a_n348_122# a_n1188_122# 0.01fF
C233 a_n558_n188# a_n1818_n188# 0.00fF
C234 a_n2238_n188# a_n2868_122# 0.00fF
C235 a_3012_122# a_n4172_n100# 0.06fF
C236 a_n558_n188# a_n1608_122# 0.00fF
C237 a_492_122# a_n348_122# 0.01fF
C238 a_2382_n188# a_2172_122# 0.00fF
C239 a_4062_n188# a_3642_n188# 0.01fF
C240 a_2592_122# a_2172_122# 0.01fF
C241 a_n4080_n100# a_n4128_122# 0.02fF
C242 a_1542_n188# a_702_n188# 0.01fF
C243 a_n3078_n188# a_n3288_122# 0.00fF
C244 a_n2868_122# a_n3498_n188# 0.00fF
C245 a_n2028_122# a_n3288_122# 0.00fF
C246 a_n978_n188# a_n2238_n188# 0.00fF
C247 a_n768_122# a_n2238_n188# 0.00fF
C248 a_1332_122# a_n4172_n100# 0.06fF
C249 a_n1398_n188# a_n2238_n188# 0.01fF
C250 a_72_122# a_n4172_n100# 0.06fF
C251 a_n2658_n188# a_n4172_n100# 0.02fF
C252 a_1122_n188# a_702_n188# 0.01fF
C253 a_n1188_122# a_n2238_n188# 0.00fF
C254 a_2802_n188# a_2382_n188# 0.01fF
C255 a_n2658_n188# a_n3708_122# 0.00fF
C256 a_2802_n188# a_2592_122# 0.00fF
C257 a_n2658_n188# a_n2448_122# 0.00fF
C258 a_n4080_n100# a_n3078_n188# 0.06fF
C259 a_n4128_122# a_n4172_n100# 0.06fF
C260 a_n4080_n100# a_n2028_122# 0.02fF
C261 a_n1818_n188# a_n2868_122# 0.00fF
C262 a_912_122# a_n348_122# 0.00fF
C263 a_n1608_122# a_n2868_122# 0.00fF
C264 a_n3708_122# a_n4128_122# 0.01fF
C265 a_2382_n188# a_1962_n188# 0.01fF
C266 a_2592_122# a_1962_n188# 0.00fF
C267 a_1542_n188# a_1752_122# 0.00fF
C268 a_4062_n188# a_2802_n188# 0.00fF
C269 a_n4080_n100# a_n348_122# 0.02fF
C270 a_2172_122# a_702_n188# 0.00fF
C271 a_n978_n188# a_n1818_n188# 0.01fF
C272 a_282_n188# a_n138_n188# 0.01fF
C273 a_n2238_n188# a_n3288_122# 0.00fF
C274 a_1542_n188# a_492_122# 0.00fF
C275 a_n978_n188# a_n1608_122# 0.00fF
C276 a_n768_122# a_n1818_n188# 0.00fF
C277 a_3222_n188# a_1752_122# 0.00fF
C278 a_n1398_n188# a_n1818_n188# 0.01fF
C279 a_n768_122# a_n1608_122# 0.01fF
C280 a_1752_122# a_1122_n188# 0.00fF
C281 a_n3078_n188# a_n4172_n100# 0.02fF
C282 a_n1188_122# a_n1818_n188# 0.00fF
C283 a_n1398_n188# a_n1608_122# 0.00fF
C284 a_n2028_122# a_n4172_n100# 0.06fF
C285 a_n1188_122# a_n1608_122# 0.01fF
C286 a_1122_n188# a_492_122# 0.00fF
C287 a_n3078_n188# a_n3708_122# 0.00fF
C288 a_n3498_n188# a_n3288_122# 0.00fF
C289 a_n2868_122# a_n3918_n188# 0.00fF
C290 a_3432_122# a_4228_n100# 0.00fF
C291 a_1332_122# a_72_122# 0.00fF
C292 a_n4080_n100# a_4228_n100# 0.21fF
C293 a_n2448_122# a_n3078_n188# 0.00fF
C294 a_n138_n188# a_n558_n188# 0.01fF
C295 a_n2028_122# a_n2448_122# 0.01fF
C296 a_3852_122# a_4228_n100# 0.01fF
C297 a_n4080_n100# a_n2238_n188# 0.06fF
C298 a_n348_122# a_n4172_n100# 0.06fF
C299 a_n2658_n188# a_n4128_122# 0.00fF
C300 a_2382_n188# a_2592_122# 0.00fF
C301 a_n4080_n100# a_n3498_n188# 0.06fF
C302 a_2172_122# a_1752_122# 0.01fF
C303 a_1542_n188# a_912_122# 0.00fF
C304 a_1962_n188# a_702_n188# 0.00fF
C305 a_n1818_n188# a_n3288_122# 0.00fF
C306 a_702_n188# a_n138_n188# 0.01fF
C307 a_4228_n100# a_n4172_n100# 0.14fF
C308 a_n4080_n100# a_1542_n188# 0.06fF
C309 a_1122_n188# a_912_122# 0.00fF
C310 a_n2238_n188# a_n4172_n100# 0.02fF
C311 a_4062_n188# a_2592_122# 0.00fF
C312 a_3222_n188# a_3432_122# 0.00fF
C313 a_282_n188# a_n558_n188# 0.01fF
C314 a_n4080_n100# a_3222_n188# 0.06fF
C315 a_n2238_n188# a_n3708_122# 0.00fF
C316 a_n2658_n188# a_n3078_n188# 0.01fF
C317 a_n2238_n188# a_n2448_122# 0.00fF
C318 a_n2028_122# a_n2658_n188# 0.00fF
C319 a_2802_n188# a_1752_122# 0.00fF
C320 a_n4080_n100# a_1122_n188# 0.06fF
C321 a_n4080_n100# a_n1818_n188# 0.06fF
C322 a_3852_122# a_3222_n188# 0.00fF
C323 a_n3498_n188# a_n4172_n100# 0.02fF
C324 a_n4080_n100# a_n1608_122# 0.02fF
C325 a_3432_122# a_3642_n188# 0.00fF
C326 a_n3288_122# a_n3918_n188# 0.00fF
C327 a_n2868_122# a_n4382_n100# 0.00fF
C328 a_3012_122# a_4228_n100# 0.00fF
C329 a_n3078_n188# a_n4128_122# 0.00fF
C330 a_n3498_n188# a_n3708_122# 0.00fF
C331 a_n4080_n100# a_3642_n188# 0.06fF
C332 a_n2448_122# a_n3498_n188# 0.00fF
C333 a_n138_n188# a_n978_n188# 0.01fF
C334 a_72_122# a_n348_122# 0.01fF
C335 a_n138_n188# a_n768_122# 0.00fF
C336 a_1542_n188# a_n4172_n100# 0.02fF
C337 a_3852_122# a_3642_n188# 0.00fF
C338 a_1962_n188# a_1752_122# 0.00fF
C339 a_2172_122# a_912_122# 0.00fF
C340 a_n138_n188# a_n1398_n188# 0.00fF
C341 a_n138_n188# a_n1188_122# 0.00fF
C342 a_702_n188# a_282_n188# 0.01fF
C343 a_1962_n188# a_492_122# 0.00fF
C344 a_3222_n188# a_n4172_n100# 0.02fF
C345 a_492_122# a_n138_n188# 0.00fF
C346 a_1122_n188# a_n4172_n100# 0.02fF
C347 a_n1818_n188# a_n4172_n100# 0.02fF
C348 a_3432_122# a_2172_122# 0.00fF
C349 a_n4080_n100# a_2172_122# 0.02fF
C350 a_n1608_122# a_n4172_n100# 0.06fF
C351 a_n4080_n100# a_n3918_n188# 0.06fF
C352 a_n1818_n188# a_n2448_122# 0.00fF
C353 a_n4080_n100# VSUBS 1.08fF
C354 a_n4172_n100# VSUBS 1.03fF
C355 a_4062_n188# VSUBS 0.11fF
C356 a_4228_n100# VSUBS 0.17fF
C357 a_3642_n188# VSUBS 0.10fF
C358 a_3852_122# VSUBS 0.09fF
C359 a_3222_n188# VSUBS 0.11fF
C360 a_3432_122# VSUBS 0.11fF
C361 a_2802_n188# VSUBS 0.12fF
C362 a_3012_122# VSUBS 0.11fF
C363 a_2382_n188# VSUBS 0.12fF
C364 a_2592_122# VSUBS 0.12fF
C365 a_1962_n188# VSUBS 0.12fF
C366 a_2172_122# VSUBS 0.12fF
C367 a_1542_n188# VSUBS 0.12fF
C368 a_1752_122# VSUBS 0.12fF
C369 a_1122_n188# VSUBS 0.12fF
C370 a_1332_122# VSUBS 0.12fF
C371 a_702_n188# VSUBS 0.12fF
C372 a_912_122# VSUBS 0.12fF
C373 a_282_n188# VSUBS 0.12fF
C374 a_492_122# VSUBS 0.12fF
C375 a_n138_n188# VSUBS 0.12fF
C376 a_72_122# VSUBS 0.12fF
C377 a_n558_n188# VSUBS 0.12fF
C378 a_n348_122# VSUBS 0.12fF
C379 a_n978_n188# VSUBS 0.12fF
C380 a_n768_122# VSUBS 0.12fF
C381 a_n1398_n188# VSUBS 0.12fF
C382 a_n1188_122# VSUBS 0.12fF
C383 a_n1818_n188# VSUBS 0.12fF
C384 a_n1608_122# VSUBS 0.12fF
C385 a_n2238_n188# VSUBS 0.12fF
C386 a_n2028_122# VSUBS 0.12fF
C387 a_n2658_n188# VSUBS 0.12fF
C388 a_n2448_122# VSUBS 0.12fF
C389 a_n3078_n188# VSUBS 0.12fF
C390 a_n2868_122# VSUBS 0.12fF
C391 a_n3498_n188# VSUBS 0.12fF
C392 a_n3288_122# VSUBS 0.12fF
C393 a_n3918_n188# VSUBS 0.12fF
C394 a_n3708_122# VSUBS 0.12fF
C395 a_n4382_n100# VSUBS 0.20fF
C396 a_n4128_122# VSUBS 0.13fF
.ends

.subckt latch_nmos_pair sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
C0 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.01fF
C2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C4 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# -0.00fF
C5 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C6 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C7 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C8 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C9 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C10 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C11 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C12 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.57fF
C13 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C14 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C15 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C16 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C17 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C18 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C19 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C20 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C21 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C22 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C23 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C24 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C25 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C26 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C27 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C28 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C29 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C30 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C31 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C32 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C33 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C34 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C35 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C36 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C37 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C38 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C39 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.02fF
C40 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C41 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.02fF
C42 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# -0.00fF
C43 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C44 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C45 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C46 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C47 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C48 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C49 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C50 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C51 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C52 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C53 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.01fF
C54 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C55 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C56 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C57 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C58 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.02fF
C59 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C60 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C61 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C62 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C63 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C64 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C65 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C66 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.02fF
C67 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C68 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C69 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.27fF
C70 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C71 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C72 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# -0.00fF
C73 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C74 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C75 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C76 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C77 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C78 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C79 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C80 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C81 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.02fF
C82 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C83 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.42fF
C84 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C85 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C86 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C87 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C88 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C89 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C90 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.02fF
C91 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.02fF
C92 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C93 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C94 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C95 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C96 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C97 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C98 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C99 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# -0.00fF
C100 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C102 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C103 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C105 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C106 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C107 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C108 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# -0.00fF
C109 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C110 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C111 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C112 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C114 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C117 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C118 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C119 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# -0.01fF
C120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C121 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# -0.01fF
C122 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C124 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C125 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C126 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C127 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C128 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C131 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C132 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C133 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C134 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# -0.00fF
C135 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C136 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C137 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C138 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C140 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C141 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C142 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C143 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C144 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C145 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C147 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C148 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# -0.00fF
C149 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C152 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C153 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C154 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C155 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C156 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C158 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C161 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C162 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C163 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C164 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C165 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C167 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# -0.00fF
C168 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C169 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C170 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C172 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C173 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C174 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C175 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C176 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C177 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C178 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C180 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C181 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.02fF
C182 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C183 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C184 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# -0.00fF
C185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C186 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C190 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C191 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C192 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C193 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C194 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C196 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.02fF
C197 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# -0.00fF
C198 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C199 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C200 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# -0.00fF
C201 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C202 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C203 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C204 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C205 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C206 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# -0.00fF
C207 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.02fF
C208 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C209 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C210 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# -0.00fF
C211 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.57fF
C212 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.02fF
C213 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C214 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.02fF
C215 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C216 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C217 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.24fF
C218 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C219 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# -0.00fF
C220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C222 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C223 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C224 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C225 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C226 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C227 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C228 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C229 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C230 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C231 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.02fF
C232 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C233 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C235 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C236 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C237 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C238 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C239 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C240 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C241 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C242 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C243 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C244 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C245 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# -0.00fF
C246 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C247 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C248 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C249 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C250 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C251 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C252 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C253 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C254 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C255 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C256 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C257 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C258 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C259 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C260 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C261 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C262 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C264 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C265 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C266 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C267 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C268 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C269 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.01fF
C270 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C271 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C272 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C273 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C274 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C275 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C276 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C277 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.02fF
C278 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C279 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C280 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C281 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C282 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C283 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C284 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C285 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C286 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C287 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C288 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C289 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C291 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C292 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C293 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C294 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C295 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C296 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C297 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C298 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# -0.00fF
C299 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C300 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# -0.00fF
C301 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C302 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C304 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C305 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C306 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C307 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C308 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C309 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C310 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C311 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C312 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C313 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C314 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C315 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C316 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C317 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C318 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.01fF
C319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.01fF
C320 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C321 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C322 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C323 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C324 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C325 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C326 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C327 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C329 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C330 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.02fF
C331 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C332 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C333 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C334 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C335 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C336 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C337 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C338 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C339 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C340 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C341 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# -0.00fF
C342 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C343 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C344 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C345 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C346 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# -0.00fF
C347 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C348 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C350 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C352 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C353 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C354 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.02fF
C355 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C356 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C357 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C358 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C359 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C360 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C362 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# -0.00fF
C363 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C364 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C365 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C367 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# -0.01fF
C368 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# -0.00fF
C369 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C373 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C374 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C375 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C376 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C378 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C379 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C380 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C381 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C382 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C383 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C384 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C385 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C386 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C389 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C390 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C391 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C392 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.44fF
C393 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C394 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C395 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C396 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.02fF
C397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C398 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C399 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C400 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C401 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C402 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C403 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C405 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C406 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C407 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C408 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C409 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# -0.01fF
C410 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C411 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C412 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C413 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C414 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C415 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C416 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C417 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# -0.01fF
C418 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.02fF
C419 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C421 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C422 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C423 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C424 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C426 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C427 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C428 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C429 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C430 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C432 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C434 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# -0.00fF
C435 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C436 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C437 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.02fF
C438 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C440 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C441 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C442 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C443 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C444 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C445 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.02fF
C446 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C447 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C448 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.22fF
C449 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C450 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C451 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C452 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C453 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C454 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.02fF
C455 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C457 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C458 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C459 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C460 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C461 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C462 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.02fF
C463 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C464 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C466 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C467 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C468 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C469 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C470 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C471 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C472 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C473 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C474 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C475 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C476 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C477 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C478 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C479 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C480 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C481 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C484 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C485 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C486 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C488 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C489 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C490 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C491 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C492 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C493 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C494 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C495 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C496 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C497 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C498 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C499 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C500 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C501 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C502 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C503 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C504 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C505 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C506 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C507 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C508 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C509 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# -0.00fF
C510 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C511 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C512 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# -0.00fF
C513 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C514 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C515 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.02fF
C516 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C517 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.02fF
C519 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C520 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C521 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C522 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C523 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# -0.00fF
C524 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C525 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.02fF
C526 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C527 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C528 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# -0.00fF
C529 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C530 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C531 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C532 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C533 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C534 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C535 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C536 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.01fF
C537 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C538 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C541 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C542 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C543 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C544 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C545 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C546 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C547 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C548 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C549 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C550 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C551 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C552 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C553 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# -0.00fF
C554 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C555 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C556 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C557 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C558 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# -0.00fF
C559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C560 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C563 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C564 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C565 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# -0.00fF
C567 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C568 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C569 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C571 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C572 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.00fF
C574 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# -0.00fF
C576 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# -0.00fF
C577 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C579 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C581 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C582 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C585 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C586 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C587 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C588 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C590 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# -0.00fF
C591 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C592 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C593 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C594 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C595 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C597 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C598 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C599 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C600 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C601 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C602 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# -0.00fF
C603 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C605 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C606 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C607 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C608 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C609 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C611 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C613 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.02fF
C614 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C615 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C616 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C618 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C619 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C620 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# -0.00fF
C621 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C622 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C623 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.76fF
C624 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.30fF
C625 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C626 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C627 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C628 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C629 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C630 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C631 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# -0.00fF
C632 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C633 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C634 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C635 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C636 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C637 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C638 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.02fF
C639 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C640 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.02fF
C641 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C642 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C643 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C644 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C645 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C646 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.02fF
C647 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C649 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C650 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C652 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C653 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C654 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C655 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# -0.01fF
C656 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C657 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C658 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C659 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C660 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C661 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.02fF
C662 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# -0.00fF
C663 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C664 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C665 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C666 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C667 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C668 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C669 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C670 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C671 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C672 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C673 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C674 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C675 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C677 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C679 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C680 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C683 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C684 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C686 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C687 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C688 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C689 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C690 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C691 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C692 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.01fF
C693 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C694 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C695 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C696 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C697 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C698 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.02fF
C699 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C700 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C701 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C702 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C703 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C704 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C705 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C706 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C707 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C708 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C709 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C710 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C711 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C712 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C713 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C714 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C715 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C716 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C717 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.02fF
C718 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C719 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# -0.00fF
C720 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C721 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C722 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# -0.00fF
C723 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C724 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C726 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C727 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C728 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C729 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C730 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C731 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C732 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C733 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C734 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C735 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C736 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.42fF
C737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C738 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C739 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C740 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C741 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C742 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C743 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C744 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# -0.00fF
C745 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C746 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C747 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C748 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C749 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C750 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C751 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.02fF
C752 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# -0.00fF
C753 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C754 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C755 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.02fF
C756 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.42fF
C757 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# -0.00fF
C758 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C759 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C760 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C761 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C762 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C763 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C764 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C765 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C766 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C767 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C768 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C769 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.02fF
C770 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C771 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# -0.00fF
C772 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C773 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.42fF
C774 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C775 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.01fF
C776 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C777 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C778 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.02fF
C779 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C780 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C781 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C782 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C783 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C784 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C785 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C786 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C787 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C788 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C789 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C790 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C791 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# -0.00fF
C792 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C793 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C794 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C795 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C796 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C797 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C798 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.27fF
C800 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C801 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C802 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# -0.00fF
C803 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C805 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# -0.00fF
C806 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C807 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C808 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C809 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C810 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.02fF
C811 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C812 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C813 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C814 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C815 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C816 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C817 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C818 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C819 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C820 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C821 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C822 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C823 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C824 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C825 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C826 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C827 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C828 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C829 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C830 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.02fF
C831 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C832 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C833 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C834 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C835 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C836 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C837 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C838 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C839 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# -0.00fF
C840 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C841 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C842 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C843 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C844 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C845 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# -0.00fF
C846 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.00fF
C847 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C848 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C849 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C850 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# -0.00fF
C851 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C852 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C853 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C854 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C855 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C856 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C857 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C858 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C859 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# -0.00fF
C860 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C861 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C862 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C863 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C864 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.17fF
C866 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C867 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C868 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C869 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C870 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C871 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C872 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C873 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C874 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C875 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C876 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C877 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C878 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C879 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C880 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# -0.01fF
C881 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C882 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C883 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C884 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C885 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C886 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C887 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C888 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C889 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C890 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C891 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C892 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# -0.00fF
C893 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C894 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C895 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C896 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C897 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C898 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C899 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# -0.01fF
C900 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C901 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C902 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C903 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C904 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C905 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C906 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C907 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C908 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C909 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C910 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C911 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C912 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# -0.00fF
C913 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C914 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C915 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C916 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C917 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C918 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C919 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C920 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C921 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.93fF
C922 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C923 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C924 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C925 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C926 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# -0.01fF
C927 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C928 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C929 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C930 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C931 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C932 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C933 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C934 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C935 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C936 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.31fF
C937 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C938 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C939 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C940 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# -0.00fF
C941 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C942 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C943 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C944 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C945 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C946 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C947 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.02fF
C948 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# -0.01fF
C949 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C950 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C951 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C952 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C953 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C954 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C955 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C956 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# -0.00fF
C957 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C958 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C959 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C960 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C961 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C962 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C963 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C964 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# -0.00fF
C965 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C966 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C967 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C968 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# -0.00fF
C969 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C970 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C971 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C972 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C973 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# -0.00fF
C974 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C975 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C976 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C977 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C978 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C979 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.02fF
C980 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C981 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C982 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C983 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C984 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C985 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C986 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C987 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C988 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C989 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C990 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C991 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C992 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C993 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C994 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C995 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C996 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C997 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C998 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C999 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1000 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1001 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1002 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# -0.00fF
C1003 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1004 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C1005 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1006 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1007 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1008 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.02fF
C1009 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C1010 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1011 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1012 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C1013 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1014 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1015 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1016 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1017 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1018 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1019 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1020 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1021 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1022 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1023 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1024 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C1025 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1026 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1027 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C1028 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1029 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1030 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1031 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1032 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C1033 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1034 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C1035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C1036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1037 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C1038 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1039 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1040 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1041 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1042 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1043 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.02fF
C1044 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1045 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C1046 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1047 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C1048 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1049 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1050 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1052 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C1053 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1054 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.02fF
C1055 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# -0.00fF
C1056 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1057 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 1.18fF
C1058 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1059 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1060 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1061 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1062 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C1063 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1064 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1065 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1066 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C1067 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1068 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C1069 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C1070 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1072 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1073 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1074 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1075 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1077 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C1078 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C1079 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C1080 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1081 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C1082 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C1083 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C1084 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C1085 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# -0.01fF
C1086 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1087 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C1088 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C1089 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1090 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C1091 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1092 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1093 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1094 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C1095 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C1096 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1097 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1098 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C1099 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.00fF
C1100 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1101 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.31fF
C1102 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 1.18fF
C1103 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C1104 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C1105 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1106 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1107 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1108 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1109 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1110 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1111 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1112 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# -0.00fF
C1113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.02fF
C1114 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C1115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C1116 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C1117 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1118 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1119 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C1120 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1121 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C1122 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C1123 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C1125 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C1126 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# -0.00fF
C1128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1129 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C1130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# -0.00fF
C1131 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1132 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1133 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C1134 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1135 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1136 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# -0.00fF
C1138 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.02fF
C1140 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1141 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1142 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C1143 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# -0.00fF
C1144 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C1145 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.00fF
C1146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1147 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C1148 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C1149 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C1150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1151 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1152 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1153 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1154 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C1155 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C1156 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.27fF
C1157 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C1158 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C1159 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C1160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1162 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C1163 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C1164 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.02fF
C1165 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# -0.00fF
C1166 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C1167 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1168 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1169 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1170 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# -0.00fF
C1171 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1172 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C1173 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1174 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1175 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1176 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1177 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1178 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1182 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.02fF
C1183 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1184 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C1185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1186 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1187 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1188 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# -0.00fF
C1189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1190 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1191 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# -0.00fF
C1192 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1193 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1194 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1195 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1196 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1197 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C1198 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1199 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1201 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1202 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C1203 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1206 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1207 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.02fF
C1208 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1209 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C1210 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C1211 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C1212 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1213 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1214 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C1215 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1216 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1217 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1218 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1219 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1221 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1222 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1223 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1224 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1225 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1226 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C1227 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C1228 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# -0.00fF
C1229 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1230 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C1231 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C1232 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# -0.00fF
C1233 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1234 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1235 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1236 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C1237 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C1238 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1239 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C1240 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# -0.00fF
C1241 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1242 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C1243 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1244 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C1245 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1246 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1247 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# -0.00fF
C1248 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1249 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C1250 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1251 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C1252 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C1253 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C1254 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C1255 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1256 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1257 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C1258 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1259 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C1260 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1261 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1262 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1263 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C1264 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1265 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1266 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1268 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1269 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1270 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 1.18fF
C1271 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C1272 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1273 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# -0.00fF
C1274 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.01fF
C1275 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# -0.00fF
C1276 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1277 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1278 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C1279 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1281 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1283 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.02fF
C1284 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1285 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.02fF
C1286 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1287 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.57fF
C1288 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1289 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C1290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1291 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1292 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1293 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1294 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.02fF
C1295 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C1296 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1297 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# -0.00fF
C1298 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1299 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1300 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.02fF
C1301 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1302 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C1303 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1304 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1305 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C1306 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# -0.00fF
C1307 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1308 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1309 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.02fF
C1310 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C1311 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C1312 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.02fF
C1313 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1314 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1315 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1316 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# -0.00fF
C1317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# -0.00fF
C1318 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1319 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1320 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C1321 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1322 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1323 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1324 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C1325 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1326 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C1327 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1328 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1329 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C1330 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.02fF
C1331 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# -0.00fF
C1332 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1333 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# -0.00fF
C1334 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1335 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C1336 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1337 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# -0.01fF
C1338 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C1339 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# -0.00fF
C1340 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1341 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1342 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1343 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1344 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.00fF
C1345 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C1346 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1347 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C1348 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1349 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1350 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C1351 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1352 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1353 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1354 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1355 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.02fF
C1356 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1357 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1358 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C1359 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# -0.00fF
C1360 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# -0.00fF
C1361 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1362 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1363 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1364 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# -0.00fF
C1365 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.02fF
C1366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1367 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1368 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1369 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1371 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C1373 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1374 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C1375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1376 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1377 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C1378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C1379 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1380 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C1381 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C1382 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C1383 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C1384 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1385 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# -0.00fF
C1386 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C1388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1389 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1390 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1391 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1392 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1393 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1394 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1395 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C1396 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C1398 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C1399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1401 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C1404 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1405 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1406 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1407 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1408 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C1409 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1410 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1411 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1412 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1413 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1414 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1415 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C1416 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C1417 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1418 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1419 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C1420 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.02fF
C1421 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C1422 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1423 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1424 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C1425 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C1426 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1427 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.01fF
C1428 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1429 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1430 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C1431 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C1432 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# -0.00fF
C1433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C1434 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1435 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1436 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# -0.00fF
C1437 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.02fF
C1438 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C1439 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1440 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C1441 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1442 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1443 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1444 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1446 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1447 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C1448 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1449 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1450 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1451 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C1452 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1453 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1454 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C1455 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.44fF
C1456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1458 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C1459 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1460 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1462 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1463 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C1464 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.93fF
C1465 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1466 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1467 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C1468 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C1469 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1470 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1471 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C1472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1473 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1474 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C1475 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1476 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1477 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1478 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1479 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# -0.00fF
C1480 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C1481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C1482 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1483 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1484 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.02fF
C1485 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1486 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C1488 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1489 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1490 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1491 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1492 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1493 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1494 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1495 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1496 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1497 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1498 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1499 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C1500 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1501 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.00fF
C1503 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1504 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1505 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1506 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1507 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1508 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C1509 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1510 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C1511 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C1512 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C1513 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1514 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1515 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C1516 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1517 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# -0.00fF
C1518 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1519 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C1520 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C1521 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1522 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1523 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1524 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C1525 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# -0.00fF
C1526 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.01fF
C1527 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1528 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C1529 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1530 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C1531 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C1532 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1533 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C1534 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1535 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C1536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# -0.00fF
C1537 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C1538 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1539 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.02fF
C1540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C1541 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1542 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1543 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C1544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1545 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1546 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C1547 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1548 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.01fF
C1549 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# -0.00fF
C1550 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1551 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# -0.00fF
C1552 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.02fF
C1553 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1554 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1555 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.02fF
C1556 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C1557 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1558 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# -0.00fF
C1560 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# VSUBS 1.08fF
C1561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# VSUBS 1.03fF
C1562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# VSUBS 0.11fF
C1563 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# VSUBS 0.17fF
C1564 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# VSUBS 0.10fF
C1565 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# VSUBS 0.09fF
C1566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# VSUBS 0.11fF
C1567 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# VSUBS 0.11fF
C1568 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# VSUBS 0.12fF
C1569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# VSUBS 0.11fF
C1570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# VSUBS 0.12fF
C1571 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# VSUBS 0.12fF
C1572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# VSUBS 0.12fF
C1573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# VSUBS 0.12fF
C1574 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# VSUBS 0.12fF
C1575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# VSUBS 0.12fF
C1576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# VSUBS 0.12fF
C1577 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# VSUBS 0.12fF
C1578 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# VSUBS 0.12fF
C1579 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# VSUBS 0.12fF
C1580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# VSUBS 0.12fF
C1581 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# VSUBS 0.12fF
C1582 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# VSUBS 0.12fF
C1583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# VSUBS 0.12fF
C1584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# VSUBS 0.12fF
C1585 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# VSUBS 0.12fF
C1586 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# VSUBS 0.12fF
C1587 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# VSUBS 0.12fF
C1588 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# VSUBS 0.12fF
C1589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# VSUBS 0.12fF
C1590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# VSUBS 0.12fF
C1591 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# VSUBS 0.12fF
C1592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# VSUBS 0.12fF
C1593 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# VSUBS 0.12fF
C1594 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# VSUBS 0.12fF
C1595 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# VSUBS 0.12fF
C1596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# VSUBS 0.12fF
C1597 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# VSUBS 0.12fF
C1598 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# VSUBS 0.12fF
C1599 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# VSUBS 0.12fF
C1600 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# VSUBS 0.12fF
C1601 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# VSUBS 0.12fF
C1602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# VSUBS 0.20fF
C1603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# VSUBS 0.13fF
C1604 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# VSUBS 1.08fF
C1605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# VSUBS 1.03fF
C1606 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# VSUBS 0.11fF
C1607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# VSUBS 0.17fF
C1608 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# VSUBS 0.10fF
C1609 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# VSUBS 0.09fF
C1610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# VSUBS 0.11fF
C1611 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# VSUBS 0.11fF
C1612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# VSUBS 0.12fF
C1613 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# VSUBS 0.11fF
C1614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# VSUBS 0.12fF
C1615 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# VSUBS 0.12fF
C1616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# VSUBS 0.12fF
C1617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# VSUBS 0.12fF
C1618 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# VSUBS 0.12fF
C1619 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# VSUBS 0.12fF
C1620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# VSUBS 0.12fF
C1621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# VSUBS 0.12fF
C1622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# VSUBS 0.12fF
C1623 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# VSUBS 0.12fF
C1624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# VSUBS 0.12fF
C1625 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# VSUBS 0.12fF
C1626 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# VSUBS 0.12fF
C1627 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# VSUBS 0.12fF
C1628 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# VSUBS 0.12fF
C1629 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# VSUBS 0.12fF
C1630 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# VSUBS 0.12fF
C1631 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# VSUBS 0.12fF
C1632 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# VSUBS 0.12fF
C1633 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# VSUBS 0.12fF
C1634 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# VSUBS 0.12fF
C1635 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# VSUBS 0.12fF
C1636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# VSUBS 0.12fF
C1637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# VSUBS 0.12fF
C1638 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# VSUBS 0.12fF
C1639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# VSUBS 0.12fF
C1640 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# VSUBS 0.12fF
C1641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# VSUBS 0.12fF
C1642 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# VSUBS 0.12fF
C1643 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# VSUBS 0.12fF
C1644 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# VSUBS 0.12fF
C1645 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# VSUBS 0.12fF
C1646 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# VSUBS 0.20fF
C1647 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# VSUBS 0.13fF
C1648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# VSUBS 1.08fF
C1649 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# VSUBS 1.03fF
C1650 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# VSUBS 0.11fF
C1651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# VSUBS 0.17fF
C1652 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# VSUBS 0.10fF
C1653 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# VSUBS 0.09fF
C1654 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# VSUBS 0.11fF
C1655 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# VSUBS 0.11fF
C1656 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# VSUBS 0.12fF
C1657 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# VSUBS 0.11fF
C1658 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# VSUBS 0.12fF
C1659 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# VSUBS 0.12fF
C1660 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# VSUBS 0.12fF
C1661 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# VSUBS 0.12fF
C1662 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# VSUBS 0.12fF
C1663 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# VSUBS 0.12fF
C1664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# VSUBS 0.12fF
C1665 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# VSUBS 0.12fF
C1666 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# VSUBS 0.12fF
C1667 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# VSUBS 0.12fF
C1668 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# VSUBS 0.12fF
C1669 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# VSUBS 0.12fF
C1670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# VSUBS 0.12fF
C1671 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# VSUBS 0.12fF
C1672 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# VSUBS 0.12fF
C1673 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# VSUBS 0.12fF
C1674 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# VSUBS 0.12fF
C1675 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# VSUBS 0.12fF
C1676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# VSUBS 0.12fF
C1677 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# VSUBS 0.12fF
C1678 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# VSUBS 0.12fF
C1679 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# VSUBS 0.12fF
C1680 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# VSUBS 0.12fF
C1681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# VSUBS 0.12fF
C1682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# VSUBS 0.12fF
C1683 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# VSUBS 0.12fF
C1684 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# VSUBS 0.12fF
C1685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# VSUBS 0.12fF
C1686 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# VSUBS 0.12fF
C1687 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# VSUBS 0.12fF
C1688 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# VSUBS 0.12fF
C1689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# VSUBS 0.12fF
C1690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# VSUBS 0.20fF
C1691 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# VSUBS 0.13fF
C1692 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# VSUBS 1.08fF
C1693 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# VSUBS 1.03fF
C1694 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# VSUBS 0.11fF
C1695 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# VSUBS 0.17fF
C1696 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# VSUBS 0.10fF
C1697 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# VSUBS 0.09fF
C1698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# VSUBS 0.11fF
C1699 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# VSUBS 0.11fF
C1700 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# VSUBS 0.12fF
C1701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# VSUBS 0.11fF
C1702 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# VSUBS 0.12fF
C1703 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# VSUBS 0.12fF
C1704 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# VSUBS 0.12fF
C1705 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# VSUBS 0.12fF
C1706 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# VSUBS 0.12fF
C1707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# VSUBS 0.12fF
C1708 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# VSUBS 0.12fF
C1709 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# VSUBS 0.12fF
C1710 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# VSUBS 0.12fF
C1711 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# VSUBS 0.12fF
C1712 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# VSUBS 0.12fF
C1713 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# VSUBS 0.12fF
C1714 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# VSUBS 0.12fF
C1715 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# VSUBS 0.12fF
C1716 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# VSUBS 0.12fF
C1717 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# VSUBS 0.12fF
C1718 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# VSUBS 0.12fF
C1719 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# VSUBS 0.12fF
C1720 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# VSUBS 0.12fF
C1721 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# VSUBS 0.12fF
C1722 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# VSUBS 0.12fF
C1723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# VSUBS 0.12fF
C1724 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# VSUBS 0.12fF
C1725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# VSUBS 0.12fF
C1726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# VSUBS 0.12fF
C1727 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# VSUBS 0.12fF
C1728 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# VSUBS 0.12fF
C1729 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# VSUBS 0.12fF
C1730 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# VSUBS 0.12fF
C1731 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# VSUBS 0.12fF
C1732 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# VSUBS 0.12fF
C1733 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# VSUBS 0.12fF
C1734 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# VSUBS 0.20fF
C1735 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# VSUBS 0.13fF
.ends

.subckt input_diff_pair sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_4 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_5 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_6 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_7 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
C0 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C2 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C4 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C5 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C6 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C7 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C8 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C9 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C10 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.44fF
C11 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C12 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C13 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C14 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C15 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C16 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C17 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C18 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C19 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C20 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C21 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C22 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C23 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.01fF
C24 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C25 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C26 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C27 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.01fF
C28 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# -0.00fF
C29 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C30 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.24fF
C31 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C32 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C33 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.02fF
C34 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C35 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C36 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C37 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C38 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C39 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C40 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C41 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C42 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C43 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C44 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C45 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C46 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C47 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C48 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C49 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C50 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C51 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C52 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C53 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.02fF
C54 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C55 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.02fF
C56 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C57 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C58 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C59 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.02fF
C60 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C61 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C62 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C63 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C64 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C65 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C66 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C67 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C68 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C69 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C70 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C71 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C72 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.02fF
C73 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C74 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C75 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.02fF
C76 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C77 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C78 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.01fF
C79 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C80 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C81 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.02fF
C82 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C83 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C84 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C85 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C86 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C87 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C88 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C89 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C90 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.01fF
C91 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C92 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C93 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C94 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C95 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C96 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C97 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# -0.00fF
C98 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# -0.00fF
C99 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# 0.00fF
C100 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 1.18fF
C101 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C103 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C104 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C106 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C107 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C108 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C109 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C111 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C112 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C114 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C116 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# -0.00fF
C118 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C119 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C121 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C122 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.00fF
C124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C125 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C126 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C127 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C128 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C129 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C131 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.02fF
C132 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C133 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C134 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C135 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C136 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C137 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C138 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C139 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C140 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C142 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C143 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C144 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C146 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.19fF
C147 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C148 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C149 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C150 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C151 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C152 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C153 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C154 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C155 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C156 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C157 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C158 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.02fF
C159 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C160 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.02fF
C161 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C162 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C163 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.44fF
C164 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C165 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C166 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.01fF
C167 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C168 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C169 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C170 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C171 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.02fF
C172 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C173 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# 0.02fF
C174 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.02fF
C175 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C176 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C177 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C178 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C179 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C182 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C183 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.01fF
C184 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C186 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C187 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C188 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.02fF
C189 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C190 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C191 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C192 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C193 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.01fF
C194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C195 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C196 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C197 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C199 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C200 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C201 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.02fF
C202 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C203 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.02fF
C204 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C205 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C206 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C207 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C208 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.02fF
C209 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C210 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C211 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C212 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C213 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C214 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C215 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C216 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C217 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C218 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C219 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C222 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.02fF
C223 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C224 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C225 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C226 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.01fF
C227 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C228 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C229 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C230 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C231 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.00fF
C232 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C233 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C234 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.01fF
C235 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C236 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# -0.00fF
C237 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C238 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.93fF
C239 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.02fF
C240 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C241 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C242 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C243 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C244 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.01fF
C245 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C246 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C247 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C249 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C250 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C251 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C252 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# -0.00fF
C253 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C254 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C255 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C256 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C257 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C258 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C259 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C260 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.01fF
C261 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C262 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C263 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C264 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C265 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C266 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C268 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C269 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C270 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# -0.00fF
C271 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C272 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C273 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C274 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C275 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C276 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C277 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C278 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C279 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C280 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C281 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C282 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C283 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C284 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C285 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C286 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C287 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C288 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.02fF
C289 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C290 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C291 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C292 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C293 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C294 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C295 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C296 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C297 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C298 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C299 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C300 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C301 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C302 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# -0.00fF
C303 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C304 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C305 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C306 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C307 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C308 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C309 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C310 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C311 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C312 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# -0.00fF
C313 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C314 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C315 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C316 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C317 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C318 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C319 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C320 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.01fF
C321 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C322 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C323 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C324 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.01fF
C325 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C326 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# -0.00fF
C327 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C328 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.01fF
C329 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C330 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C331 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.01fF
C332 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C333 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C334 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C335 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.01fF
C336 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C337 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C338 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C339 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C340 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C341 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C342 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C343 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.02fF
C344 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.01fF
C345 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C346 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C347 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C348 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C349 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.02fF
C350 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C351 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C352 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C353 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C354 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C355 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.02fF
C356 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C357 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C358 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C359 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C360 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C361 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C362 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C363 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C364 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C365 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C367 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.02fF
C368 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C369 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C370 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C372 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C373 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C374 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C375 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C376 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# -0.00fF
C377 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C378 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C379 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C380 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# -0.00fF
C381 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C382 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C383 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C384 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C385 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C386 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C387 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C388 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C389 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C390 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C391 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C392 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C393 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C394 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C395 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.00fF
C396 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C397 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C398 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# -0.00fF
C401 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C402 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C403 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C405 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C406 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C407 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.02fF
C408 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C409 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C410 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C411 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C412 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C413 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C414 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C415 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C416 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C417 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C418 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C419 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C420 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C421 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.02fF
C422 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C423 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C424 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C425 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C426 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C427 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C428 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C429 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C430 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C432 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C433 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C434 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C435 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C436 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C437 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C438 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C440 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C441 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C442 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C443 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# -0.00fF
C444 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C446 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C447 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C448 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C449 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C450 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C451 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C452 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C453 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C454 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C455 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C456 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.02fF
C458 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C459 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C460 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C462 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C463 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C464 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C465 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C466 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C467 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C468 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C469 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.01fF
C470 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C471 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C472 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C473 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C474 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# -0.00fF
C475 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C476 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.02fF
C477 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C478 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C479 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C480 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.01fF
C481 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C482 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.00fF
C483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C484 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C485 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.01fF
C486 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C487 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C488 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C489 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C490 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C491 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C492 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C493 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C494 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C495 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C496 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C497 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C498 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C499 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C500 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C501 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C502 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.02fF
C503 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C504 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C505 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C506 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.02fF
C507 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C508 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C509 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.01fF
C510 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C511 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C512 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C513 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C515 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C516 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C517 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C519 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.02fF
C520 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C521 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C522 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C523 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C524 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C525 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C526 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C527 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C528 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.02fF
C529 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C530 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C531 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C532 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C533 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C534 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C535 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C537 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C538 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C541 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C542 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C543 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C544 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C545 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C546 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.01fF
C547 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C548 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C549 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C550 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C551 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C552 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C553 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C554 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C555 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C556 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C557 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C558 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C559 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.00fF
C560 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C562 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C563 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C564 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C565 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C566 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C567 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.02fF
C568 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C569 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.01fF
C570 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C571 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C572 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C573 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C574 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C575 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C576 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C577 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C578 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C579 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.02fF
C581 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C582 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C583 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C584 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C585 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C586 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# -0.00fF
C587 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C588 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C590 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C591 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# -0.00fF
C592 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C593 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C594 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C595 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C596 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C597 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C598 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C599 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.02fF
C600 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C601 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C602 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C603 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C604 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C605 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C606 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.01fF
C607 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C608 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C609 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.02fF
C610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C611 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C613 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C614 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C615 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C617 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C618 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.02fF
C619 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.02fF
C620 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C621 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C622 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C623 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C624 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C625 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.02fF
C626 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C627 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C628 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C629 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C630 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# -0.01fF
C631 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.93fF
C632 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C633 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C634 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C635 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C636 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C638 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C640 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C642 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C643 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C644 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C645 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C646 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C647 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C648 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# -0.00fF
C649 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C650 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C651 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C652 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C653 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C654 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C655 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C656 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C657 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# -0.00fF
C658 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C659 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.02fF
C660 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C661 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C662 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C663 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.01fF
C664 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C665 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C666 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C667 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.42fF
C668 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C669 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# -0.00fF
C670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C671 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C672 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C673 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C674 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C675 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# -0.00fF
C676 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C677 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C678 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C679 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C680 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C681 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C683 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C684 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C685 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C686 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C687 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C688 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C689 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C690 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C691 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C692 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C693 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C694 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C695 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C696 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C697 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.02fF
C698 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C699 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.02fF
C700 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C702 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C703 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# -0.00fF
C704 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C705 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.57fF
C706 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C707 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C708 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C709 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C710 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C711 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C712 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C713 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C714 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C715 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C716 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C717 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C718 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C719 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C720 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C721 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.00fF
C722 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.02fF
C723 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C724 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C725 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C727 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C728 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.44fF
C729 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C730 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C731 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C732 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C733 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C734 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C735 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C736 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C737 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C738 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C739 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C740 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C741 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C742 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C743 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# 0.00fF
C744 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C745 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C746 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C747 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C748 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C749 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C750 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C751 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.22fF
C752 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C753 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.02fF
C754 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.02fF
C755 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# -0.00fF
C756 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C757 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C758 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C759 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C760 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C761 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.01fF
C762 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C763 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C764 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C765 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.02fF
C766 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C767 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C768 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C769 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C770 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C771 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# -0.00fF
C772 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.22fF
C773 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C774 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C775 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C776 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C777 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C778 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C779 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C780 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C781 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C782 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.93fF
C783 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C784 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C785 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.02fF
C786 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C787 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C788 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.02fF
C789 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C790 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C791 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C792 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C793 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C794 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C795 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# -0.00fF
C796 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C797 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C798 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C799 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C800 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C801 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C802 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# -0.00fF
C803 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C804 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C805 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C806 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C807 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C808 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C809 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C810 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C811 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# -0.00fF
C812 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C813 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C814 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C815 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C816 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C817 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.02fF
C818 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C819 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C820 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C821 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C822 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C823 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.02fF
C824 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C825 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C826 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C827 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.01fF
C828 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C829 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C830 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.01fF
C831 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C832 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C833 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C834 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C835 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C836 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C837 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C838 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C839 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C840 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.01fF
C841 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C842 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C843 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C844 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C845 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.02fF
C846 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C847 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C848 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C849 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C850 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C851 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C852 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C853 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C854 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C855 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C856 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C857 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C858 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C859 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# -0.00fF
C860 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# -0.00fF
C861 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C862 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# -0.00fF
C863 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C864 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C865 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.19fF
C866 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C867 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# -0.00fF
C868 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C869 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C870 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C871 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C872 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C873 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C874 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.01fF
C875 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.01fF
C876 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C877 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C878 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C879 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C880 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C881 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C882 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C883 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C884 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C885 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C886 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C887 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C888 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C889 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C890 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C891 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C892 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C893 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.02fF
C894 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C896 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C897 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C898 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C899 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.01fF
C900 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.42fF
C901 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C902 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C903 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C904 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C905 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C906 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C907 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C908 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C909 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C910 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.01fF
C911 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C912 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C913 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C914 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.27fF
C915 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C916 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C917 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C918 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# 0.01fF
C919 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C920 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C921 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C922 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C923 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C924 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.93fF
C925 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C926 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C927 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C928 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C929 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C930 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C931 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C932 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C933 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C934 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C935 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C936 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C937 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C938 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# -0.00fF
C939 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C940 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C941 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C942 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.02fF
C943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# -0.00fF
C944 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C945 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C946 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C947 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.93fF
C948 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# -0.00fF
C949 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C950 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C951 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C952 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C953 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.02fF
C954 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C955 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C956 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C957 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C958 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C959 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C960 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C961 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C962 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# -0.00fF
C963 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.01fF
C964 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C965 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C966 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C967 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C968 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C969 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C970 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C971 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C972 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C973 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C974 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C975 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C976 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C978 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C979 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C980 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C981 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C982 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C983 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C984 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C985 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C986 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C987 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C988 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C989 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C990 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C991 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C993 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C994 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.02fF
C995 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C996 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C997 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C998 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.46fF
C999 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1000 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C1001 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C1002 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C1003 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.02fF
C1004 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C1005 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C1006 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1007 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1008 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1009 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C1010 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C1011 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C1012 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C1013 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1014 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1015 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1016 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1017 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C1018 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C1019 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1020 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C1021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C1022 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1023 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C1024 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1025 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C1026 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1027 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1028 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1029 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1030 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.01fF
C1032 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.01fF
C1033 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1034 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C1035 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C1036 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1037 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1038 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C1039 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.01fF
C1040 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1041 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1042 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1043 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C1044 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1045 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C1046 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1047 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.02fF
C1048 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1049 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C1050 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1051 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C1052 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1053 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C1054 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1055 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C1056 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C1057 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C1058 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.93fF
C1059 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1060 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1061 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C1062 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C1063 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1064 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1065 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1066 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1067 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1068 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1069 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1070 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C1071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1072 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1073 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C1074 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1075 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C1076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C1077 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C1078 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# -0.00fF
C1079 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C1080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C1081 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1082 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.02fF
C1083 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1084 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1085 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.00fF
C1086 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C1087 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C1088 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C1089 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1090 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C1091 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1092 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C1093 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.02fF
C1094 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1095 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.01fF
C1096 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# -0.00fF
C1097 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C1098 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C1099 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C1100 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1101 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1102 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1103 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C1104 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1106 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1107 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1108 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C1109 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1110 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C1112 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C1113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C1114 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C1115 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C1116 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1117 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1118 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1119 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C1120 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C1121 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C1122 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1123 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1124 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1125 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1126 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1127 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1128 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1130 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# -0.00fF
C1131 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1132 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1133 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1134 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.01fF
C1135 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1136 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1137 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C1138 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1139 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C1140 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C1141 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1142 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C1143 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1144 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C1145 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.44fF
C1146 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1147 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C1148 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C1149 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C1150 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C1151 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1152 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.00fF
C1153 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C1155 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1156 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1157 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C1158 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C1159 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.01fF
C1160 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C1161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C1162 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1163 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1164 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1165 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C1166 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# -0.00fF
C1167 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1168 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1169 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1170 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C1171 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1172 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C1173 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1175 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C1176 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1177 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1178 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# -0.00fF
C1179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1180 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C1181 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1182 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1183 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C1184 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1185 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1186 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1187 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1188 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# -0.00fF
C1189 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1190 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C1191 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1192 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C1193 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1194 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# -0.00fF
C1195 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C1196 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C1197 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C1198 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C1199 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1200 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1201 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C1202 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1203 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# -0.00fF
C1204 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C1205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C1206 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1207 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1208 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C1209 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1210 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.02fF
C1211 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1212 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C1213 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C1214 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1215 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1216 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C1217 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C1218 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1220 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C1221 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1222 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C1223 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C1224 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1225 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1226 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1227 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C1228 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1229 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C1230 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1231 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1232 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C1233 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1234 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C1235 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C1236 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1237 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.02fF
C1238 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1239 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1240 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1241 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1242 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1243 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1244 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.02fF
C1245 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1246 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# -0.00fF
C1247 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C1248 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1249 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1250 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1251 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1252 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1253 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1254 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1255 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1256 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C1257 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C1258 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.01fF
C1259 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# -0.00fF
C1260 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C1261 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C1262 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.02fF
C1263 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C1264 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C1265 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C1266 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1267 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C1268 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# -0.00fF
C1269 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1270 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C1271 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1272 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1273 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C1274 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C1275 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# -0.00fF
C1276 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1277 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1278 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1279 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C1280 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C1281 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1282 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.01fF
C1283 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.02fF
C1284 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1285 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C1286 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1287 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C1288 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C1289 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1290 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1291 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.02fF
C1292 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1293 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1294 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1295 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C1296 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C1297 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.01fF
C1298 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C1299 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1300 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C1301 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C1302 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C1303 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# -0.00fF
C1304 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1305 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1306 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C1307 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.02fF
C1308 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1309 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C1310 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1311 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1312 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1313 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1314 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1315 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C1316 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C1317 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C1318 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C1319 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.02fF
C1320 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1321 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1322 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C1323 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1324 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C1325 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1326 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C1327 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C1328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1329 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1330 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C1331 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# -0.00fF
C1332 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1333 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C1334 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1335 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C1336 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1337 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1338 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1339 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C1340 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.02fF
C1341 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1342 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C1343 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1344 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C1345 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1346 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C1347 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1348 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# -0.00fF
C1349 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1350 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C1351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.00fF
C1352 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1353 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1354 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1355 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C1356 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C1357 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C1358 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.01fF
C1359 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1360 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C1361 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C1362 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C1363 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1364 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1365 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.01fF
C1366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C1367 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C1368 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1369 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# -0.00fF
C1370 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1371 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C1372 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C1373 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C1374 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1375 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1376 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C1378 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# -0.00fF
C1379 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1380 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C1381 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C1382 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1383 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C1384 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1385 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C1386 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# -0.00fF
C1388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1389 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C1390 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1391 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C1392 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.00fF
C1393 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.02fF
C1394 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C1395 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1396 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C1398 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C1399 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1400 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C1401 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1402 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1403 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.02fF
C1404 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.31fF
C1405 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1406 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.02fF
C1407 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1408 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.02fF
C1409 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C1410 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1411 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1413 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C1414 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1415 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1416 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.01fF
C1417 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1418 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C1419 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C1420 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1421 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C1422 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C1423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C1424 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C1425 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C1426 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C1427 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# -0.00fF
C1428 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# -0.00fF
C1429 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C1430 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C1431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C1432 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.01fF
C1433 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C1434 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1435 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C1436 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1437 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C1438 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.02fF
C1439 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1440 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1441 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.02fF
C1442 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1443 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C1444 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C1445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C1446 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C1447 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C1448 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.00fF
C1449 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1450 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C1451 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1452 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1453 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C1454 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# -0.00fF
C1455 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C1456 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1457 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C1458 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C1459 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C1460 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1461 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C1462 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.57fF
C1463 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C1464 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C1465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C1466 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C1467 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C1468 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C1469 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C1470 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1471 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1472 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C1473 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1474 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.01fF
C1475 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.42fF
C1476 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1477 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C1478 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1479 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C1480 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1481 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.01fF
C1482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C1483 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1484 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1485 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C1486 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1488 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1489 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1490 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1491 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1492 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1493 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1494 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1495 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.02fF
C1496 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1497 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1498 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1499 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C1500 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1501 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C1502 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C1503 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C1504 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C1505 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# -0.00fF
C1506 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C1507 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C1508 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.01fF
C1509 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1510 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1511 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1512 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C1513 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1515 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C1516 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.42fF
C1517 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1518 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1519 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C1520 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1521 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1522 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C1523 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1524 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C1525 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.27fF
C1526 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1527 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.01fF
C1528 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C1529 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.93fF
C1530 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1531 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C1532 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1533 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1534 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1535 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1536 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C1537 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C1538 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1540 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# -0.00fF
C1541 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.17fF
C1542 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C1543 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.01fF
C1544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1545 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1546 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1547 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1548 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1549 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C1550 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C1551 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1552 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.02fF
C1553 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C1554 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1555 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# -0.00fF
C1556 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1557 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1558 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C1559 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C1560 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1561 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1562 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C1563 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C1564 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C1565 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1566 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C1567 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1568 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1570 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.01fF
C1571 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C1572 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C1573 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C1574 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1575 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1576 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C1577 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1578 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1579 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1580 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# -0.00fF
C1581 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# -0.00fF
C1582 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1583 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C1584 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1585 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1586 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C1587 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C1588 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1589 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C1590 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1591 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C1593 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C1594 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C1595 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1596 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1597 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C1598 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1599 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1600 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C1601 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C1602 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1603 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1604 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C1605 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C1606 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1607 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C1608 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C1609 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C1610 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C1611 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.01fF
C1612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.02fF
C1613 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1614 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1615 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C1616 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1617 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.02fF
C1618 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C1619 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C1620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1621 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C1622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C1623 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# -0.00fF
C1624 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.02fF
C1625 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1626 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1627 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1628 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.01fF
C1629 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1630 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C1631 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1632 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1633 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# -0.00fF
C1634 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.01fF
C1635 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C1636 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.02fF
C1637 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C1638 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1639 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C1640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.02fF
C1642 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C1643 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C1644 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C1645 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1646 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1647 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1648 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C1649 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1650 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C1651 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C1652 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1653 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1654 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C1655 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1656 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C1657 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1658 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C1659 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C1660 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1661 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1662 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C1663 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1664 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1665 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C1666 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1667 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C1668 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1669 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C1670 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1671 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C1672 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1673 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1674 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C1675 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1676 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C1677 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1679 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1680 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C1682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C1683 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1684 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.01fF
C1685 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.00fF
C1686 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1687 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C1688 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C1689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.22fF
C1691 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C1692 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.02fF
C1693 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C1694 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# -0.00fF
C1695 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C1696 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1697 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1698 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1699 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1700 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.78fF
C1702 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C1703 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1704 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1705 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1706 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1707 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.02fF
C1708 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1709 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C1710 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C1711 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C1712 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C1713 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1714 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1715 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C1716 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1717 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1718 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C1719 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C1720 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1721 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C1722 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C1723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1724 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C1725 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1726 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.01fF
C1727 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1728 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1729 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1730 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1731 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1732 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1733 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# -0.00fF
C1734 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1735 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.02fF
C1736 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C1737 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1738 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C1739 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.01fF
C1740 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# -0.00fF
C1741 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C1742 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1743 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1744 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1745 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1746 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C1747 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1748 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1749 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1750 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# -0.00fF
C1751 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# -0.00fF
C1752 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1753 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C1754 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C1755 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1756 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C1757 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C1758 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C1759 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1760 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1761 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C1762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C1763 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1764 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1765 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C1766 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1767 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C1768 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C1769 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1770 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C1771 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1772 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# -0.00fF
C1773 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C1774 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1775 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C1776 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1777 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C1778 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1779 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.01fF
C1780 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C1781 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C1782 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1783 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1784 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C1785 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1786 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C1787 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1788 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C1789 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C1790 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C1791 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C1792 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C1793 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1794 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1795 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# -0.00fF
C1796 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C1797 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# -0.00fF
C1798 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1800 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# -0.00fF
C1801 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1802 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1803 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1804 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C1805 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1806 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C1807 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1808 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1809 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C1810 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C1811 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# -0.00fF
C1812 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C1813 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C1814 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C1815 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1816 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1817 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C1818 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C1819 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1820 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.00fF
C1821 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C1822 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C1823 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1824 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C1825 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1826 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.02fF
C1827 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1828 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.01fF
C1829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1830 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C1831 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1832 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C1833 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C1834 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1835 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1836 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C1837 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1838 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1839 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C1840 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C1841 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1842 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C1843 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C1844 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1845 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C1846 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.02fF
C1847 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C1848 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 1.18fF
C1849 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C1850 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C1851 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1852 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C1853 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1854 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1855 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1856 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1857 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.01fF
C1858 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C1859 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C1860 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1861 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1862 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C1863 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1864 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1865 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1866 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.02fF
C1867 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1868 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# -0.00fF
C1869 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.02fF
C1870 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1871 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1872 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C1873 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C1874 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C1875 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1876 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1877 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1878 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C1879 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C1880 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.02fF
C1881 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C1882 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1883 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1884 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C1885 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1886 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.02fF
C1887 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1888 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C1889 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C1890 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1891 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1892 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C1893 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1894 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1896 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C1897 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C1898 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1899 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C1900 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C1901 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1902 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1903 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1904 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C1905 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.00fF
C1906 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1907 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# 0.00fF
C1908 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1909 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1910 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1911 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1912 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.01fF
C1913 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.02fF
C1914 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1915 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1916 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C1917 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C1918 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1919 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.01fF
C1920 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C1921 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C1922 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1923 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C1924 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1925 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1926 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# -0.00fF
C1927 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1928 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C1929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.01fF
C1930 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1931 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C1932 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1933 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# -0.00fF
C1934 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C1935 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.01fF
C1936 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1937 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.02fF
C1938 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1939 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.01fF
C1940 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1941 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1942 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1943 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C1944 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C1945 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.02fF
C1946 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# -0.00fF
C1947 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C1948 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1949 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1950 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C1951 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.02fF
C1952 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.01fF
C1954 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1955 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1956 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1957 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C1958 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1959 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1960 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1961 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C1962 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1963 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1964 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# -0.00fF
C1965 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1966 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1967 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1968 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C1969 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1970 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1971 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C1972 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1973 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1974 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C1975 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1976 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C1977 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.01fF
C1978 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.02fF
C1979 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C1980 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1981 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1982 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1983 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1984 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1985 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# -0.00fF
C1986 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1987 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1988 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C1989 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1990 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C1991 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.02fF
C1992 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1994 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C1995 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C1996 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C1997 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1998 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C1999 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C2000 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2001 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C2002 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2003 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2004 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C2005 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.01fF
C2006 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C2007 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.01fF
C2008 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C2009 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2010 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C2011 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C2012 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2013 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# -0.00fF
C2014 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2016 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C2017 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C2018 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2019 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2020 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C2022 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.02fF
C2023 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C2024 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2025 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C2026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C2027 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2028 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C2029 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2030 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# -0.00fF
C2031 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C2032 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C2033 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2034 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C2035 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C2036 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.00fF
C2037 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C2038 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C2039 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# 0.02fF
C2040 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C2041 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C2042 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C2043 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2044 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C2045 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2046 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# -0.00fF
C2047 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2048 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C2049 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2050 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C2051 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C2052 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C2053 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C2054 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C2055 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2056 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C2057 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C2058 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2059 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C2060 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C2061 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C2062 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2063 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2064 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2065 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C2066 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2067 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C2068 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.02fF
C2069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C2070 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C2071 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2072 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.31fF
C2073 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C2074 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2075 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2076 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2077 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# -0.00fF
C2078 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2079 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2080 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2081 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2082 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.02fF
C2083 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2084 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2085 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C2086 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C2087 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C2088 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2089 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C2090 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2091 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C2092 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# -0.00fF
C2093 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C2095 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# -0.00fF
C2096 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C2097 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C2098 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C2099 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C2100 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C2101 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C2102 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2103 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.01fF
C2104 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2105 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C2106 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2107 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C2108 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C2109 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.42fF
C2110 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.02fF
C2111 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C2112 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C2113 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C2114 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2115 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.02fF
C2116 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C2117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.01fF
C2118 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2119 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C2120 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C2121 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C2122 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.02fF
C2123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C2124 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2125 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2126 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# -0.00fF
C2127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2128 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2129 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.00fF
C2130 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2131 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# -0.00fF
C2132 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2133 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C2134 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2135 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.02fF
C2136 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.01fF
C2137 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C2138 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C2139 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C2140 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2141 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C2142 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C2143 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2144 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C2145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.02fF
C2147 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2148 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C2149 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.57fF
C2150 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C2151 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C2152 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2153 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2154 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2155 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# -0.00fF
C2156 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2157 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2158 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2159 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2160 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.01fF
C2161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C2162 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2163 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2164 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2165 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C2166 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C2167 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2168 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C2169 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2170 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.01fF
C2171 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C2172 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.01fF
C2173 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2174 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# -0.00fF
C2175 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2176 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2177 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2178 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2179 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2180 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.01fF
C2181 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2182 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# -0.00fF
C2183 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2184 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2185 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2186 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2187 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# -0.00fF
C2188 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C2189 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# -0.00fF
C2190 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C2191 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C2192 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2193 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2194 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C2195 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C2196 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.02fF
C2197 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.02fF
C2198 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C2199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2200 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2201 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.48fF
C2202 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.02fF
C2203 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C2204 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C2206 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2207 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C2208 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2209 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C2210 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C2211 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.30fF
C2212 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C2213 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2214 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C2215 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2216 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C2217 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.01fF
C2218 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C2219 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.01fF
C2220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C2221 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2222 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2223 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2224 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C2225 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C2226 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2227 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.02fF
C2228 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C2229 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C2230 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C2231 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C2232 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2233 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C2234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C2235 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C2236 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C2237 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2238 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.02fF
C2239 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C2240 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C2241 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C2242 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C2243 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2244 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C2245 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C2246 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2247 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C2248 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2249 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2250 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2251 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.01fF
C2252 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C2253 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2254 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C2255 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C2256 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2257 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2258 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C2259 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C2260 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C2261 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# 0.01fF
C2262 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2263 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2264 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# -0.00fF
C2265 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2266 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C2267 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C2268 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2269 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C2270 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C2271 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C2272 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# -0.00fF
C2273 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2274 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2275 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.02fF
C2276 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# -0.00fF
C2277 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C2278 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2279 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2281 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2282 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.02fF
C2283 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C2284 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C2285 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2286 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C2287 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2288 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2289 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2290 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2291 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2292 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# -0.00fF
C2293 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C2294 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2295 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2296 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C2297 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C2298 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2299 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C2300 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2301 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# -0.00fF
C2302 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C2303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2304 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.01fF
C2305 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C2306 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C2307 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2308 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C2309 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C2310 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C2311 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2312 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C2313 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2314 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C2315 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2316 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2317 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 1.18fF
C2318 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2319 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2320 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.01fF
C2321 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2322 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C2323 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.01fF
C2324 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2325 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2326 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C2327 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C2329 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.01fF
C2330 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2331 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2332 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2333 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2334 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C2335 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2336 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2337 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2338 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2339 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C2340 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.02fF
C2341 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C2342 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.02fF
C2343 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.02fF
C2344 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C2345 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2346 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2347 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.02fF
C2348 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C2350 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2351 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C2352 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2353 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C2354 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C2355 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2356 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C2357 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2358 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2359 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# -0.00fF
C2360 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C2361 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C2362 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2363 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2364 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C2365 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C2366 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2367 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C2368 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2369 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.02fF
C2370 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2371 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.00fF
C2372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2373 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# -0.00fF
C2374 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2376 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C2377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C2378 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C2379 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C2380 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C2381 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C2382 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2383 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2384 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2385 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.02fF
C2386 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2388 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2389 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2390 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C2391 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C2392 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2393 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C2394 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2395 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2396 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2397 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2398 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C2399 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C2400 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.02fF
C2401 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2402 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C2403 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C2404 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C2405 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2406 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.44fF
C2407 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C2408 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2409 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C2410 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2411 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2412 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C2413 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C2414 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2415 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# -0.00fF
C2416 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C2417 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2418 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C2419 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C2420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C2421 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# -0.00fF
C2422 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.93fF
C2423 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2424 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2425 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C2426 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C2427 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2428 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.01fF
C2429 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C2430 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# -0.00fF
C2431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C2432 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C2433 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C2434 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2435 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2436 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C2437 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2438 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2439 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C2440 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C2441 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2442 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C2443 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2444 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2446 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C2447 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2448 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2449 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C2450 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2451 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2452 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.01fF
C2453 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2454 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.01fF
C2455 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C2456 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C2457 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C2458 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2459 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2460 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2461 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C2462 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2463 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C2464 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C2465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C2466 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C2467 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# -0.00fF
C2468 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C2469 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2470 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2471 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C2472 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C2473 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# -0.00fF
C2474 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.02fF
C2475 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C2476 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C2477 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C2478 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2479 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C2480 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2481 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C2482 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C2483 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2484 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C2485 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2486 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# -0.00fF
C2487 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C2488 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2489 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C2490 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2491 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C2492 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# -0.00fF
C2493 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2495 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C2496 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2497 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C2498 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2499 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C2500 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C2501 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C2502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2503 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C2504 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C2505 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2506 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C2507 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C2508 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C2509 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C2510 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2511 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2512 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2513 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2514 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2515 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.01fF
C2516 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C2517 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2518 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C2519 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2520 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2521 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2522 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C2523 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2524 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2525 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C2526 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C2527 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.01fF
C2528 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C2529 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2530 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C2531 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2532 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C2533 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2534 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C2535 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C2536 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2537 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C2538 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C2539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C2540 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C2541 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2542 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2543 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C2544 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C2545 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.02fF
C2546 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2547 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2548 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2549 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2550 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C2551 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2552 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C2553 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.02fF
C2554 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C2555 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2556 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2557 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2558 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C2560 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C2561 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2562 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C2563 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C2564 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2565 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C2566 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# -0.00fF
C2567 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2568 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C2569 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.02fF
C2570 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C2571 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C2572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C2573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.02fF
C2574 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C2575 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C2576 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C2577 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C2579 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C2580 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C2581 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C2582 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2583 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C2584 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C2585 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C2586 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C2587 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2588 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C2589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2590 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2591 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C2592 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C2593 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# -0.00fF
C2594 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C2595 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2596 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2597 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C2598 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C2599 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# -0.00fF
C2600 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C2601 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C2602 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C2603 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C2604 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# -0.00fF
C2605 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2606 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2607 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C2608 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2609 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2610 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C2611 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C2612 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2613 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C2615 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2616 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C2617 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2618 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# -0.00fF
C2619 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C2620 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C2622 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C2623 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C2625 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.00fF
C2626 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.01fF
C2627 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C2628 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C2629 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2630 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C2631 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C2632 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.02fF
C2633 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C2634 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C2635 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2636 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2637 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2638 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C2639 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C2640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C2641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2642 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2643 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C2644 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2645 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C2646 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.02fF
C2647 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.02fF
C2648 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2649 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C2650 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2651 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C2652 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2653 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C2654 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.02fF
C2655 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.02fF
C2656 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C2657 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2658 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.42fF
C2659 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2660 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C2661 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C2662 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2663 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# -0.00fF
C2664 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2665 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C2666 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2667 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2668 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.00fF
C2669 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C2671 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2672 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.02fF
C2673 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C2674 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2675 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C2676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2677 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C2678 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C2679 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2680 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C2681 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C2682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C2683 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# 0.00fF
C2684 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2686 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C2687 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C2688 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C2691 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C2692 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.02fF
C2693 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C2694 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2695 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C2696 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# -0.01fF
C2697 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C2698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C2699 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C2700 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C2701 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2702 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2703 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C2704 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C2705 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2706 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2707 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C2708 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2709 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C2710 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C2711 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2712 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C2713 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2714 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.27fF
C2715 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2716 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.02fF
C2717 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C2718 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.01fF
C2719 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C2720 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2721 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C2722 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2723 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C2724 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C2725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C2726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C2727 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C2728 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C2729 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.02fF
C2730 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C2731 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2732 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C2733 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C2734 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C2735 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C2736 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2738 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C2739 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C2740 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2741 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.01fF
C2742 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C2743 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2744 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C2745 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2746 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2747 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.02fF
C2748 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C2749 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2750 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2751 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.93fF
C2752 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C2753 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2754 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C2755 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2756 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.02fF
C2757 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2758 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C2759 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C2760 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2761 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.31fF
C2762 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.02fF
C2763 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.01fF
C2764 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2765 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C2766 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# -0.00fF
C2767 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2768 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C2769 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2770 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2771 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C2772 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2773 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C2774 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.02fF
C2775 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C2776 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2777 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C2778 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C2779 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2780 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# -0.00fF
C2781 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2782 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C2783 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C2784 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C2785 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2786 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2787 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C2788 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C2789 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.02fF
C2790 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.02fF
C2791 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C2792 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2793 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C2794 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C2795 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C2796 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.02fF
C2797 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2798 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.02fF
C2799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2800 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C2801 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C2802 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2803 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C2804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2805 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2806 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C2807 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2808 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C2809 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C2810 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C2811 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C2812 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# -0.00fF
C2813 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2814 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2815 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C2816 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C2817 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2818 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C2819 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C2820 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C2821 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2822 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2823 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2824 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.00fF
C2825 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.01fF
C2826 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# -0.00fF
C2827 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C2828 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.02fF
C2830 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2831 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C2832 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C2833 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C2834 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2835 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C2836 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2837 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2838 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2839 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2840 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C2841 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2842 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2843 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2844 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C2845 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2846 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2847 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C2848 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C2849 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2850 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2851 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.01fF
C2852 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2854 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2855 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C2856 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2857 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2858 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.01fF
C2859 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2860 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C2861 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2862 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C2863 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C2864 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.02fF
C2865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C2866 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2867 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C2868 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C2869 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C2870 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C2871 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C2872 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C2873 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C2874 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2875 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C2876 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C2877 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C2878 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.00fF
C2879 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2880 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.01fF
C2881 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C2882 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C2883 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C2884 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2885 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2886 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C2887 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C2888 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C2889 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C2890 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C2891 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2892 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2893 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C2894 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C2895 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2896 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.57fF
C2897 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C2898 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C2899 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C2900 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C2901 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C2902 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2903 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2904 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C2906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C2907 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2908 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2909 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2910 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C2911 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2912 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2913 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C2914 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.02fF
C2915 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2916 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C2917 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2918 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2919 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 1.18fF
C2920 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2921 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2922 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C2923 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2924 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2925 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C2926 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2927 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C2928 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C2929 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2930 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2931 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C2932 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.42fF
C2933 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C2934 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2935 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2936 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2937 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2938 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2939 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C2940 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2941 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2942 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2943 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C2944 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2945 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2946 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C2947 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C2948 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2949 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C2950 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.02fF
C2951 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2952 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C2953 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2954 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C2955 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C2956 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C2957 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C2958 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2959 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.02fF
C2960 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2961 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C2962 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2963 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C2964 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C2965 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2966 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2967 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C2968 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2969 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2970 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2971 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# -0.00fF
C2972 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C2973 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.01fF
C2974 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C2975 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2976 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2977 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C2978 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2979 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2980 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C2981 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.02fF
C2982 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C2983 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2984 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C2985 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2986 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2987 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2988 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.02fF
C2989 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2990 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C2991 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C2992 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.02fF
C2993 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C2994 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C2995 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C2996 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C2997 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.02fF
C2998 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2999 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3000 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3001 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C3002 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3003 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C3004 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C3005 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.02fF
C3006 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C3007 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.01fF
C3008 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C3009 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3010 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C3011 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C3012 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3013 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C3014 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3015 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C3016 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3017 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C3018 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.02fF
C3019 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3020 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# -0.00fF
C3021 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C3022 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3023 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3024 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3025 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3026 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C3027 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C3028 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C3029 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3030 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C3031 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C3032 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3033 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.01fF
C3034 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3035 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C3036 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3037 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3038 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C3039 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3040 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3041 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C3042 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C3043 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3044 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.02fF
C3045 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3046 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3047 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3048 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3049 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C3050 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.01fF
C3051 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# -0.00fF
C3052 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3053 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C3054 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3055 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C3056 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3057 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C3058 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# -0.00fF
C3059 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3060 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C3061 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3063 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3064 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C3065 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C3066 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3067 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3068 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3069 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C3070 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C3071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3072 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C3073 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# -0.00fF
C3074 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C3075 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.02fF
C3076 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# 0.02fF
C3077 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C3078 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# -0.00fF
C3079 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C3080 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C3081 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3082 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.02fF
C3083 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C3084 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3085 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C3086 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C3087 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.02fF
C3088 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.00fF
C3089 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C3090 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3091 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3092 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C3093 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C3094 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3095 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3096 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C3097 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3098 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# -0.00fF
C3099 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C3100 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.02fF
C3101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3102 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C3103 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C3104 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3105 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3106 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.02fF
C3107 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C3108 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C3109 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3110 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.01fF
C3111 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3112 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3113 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C3115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C3116 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C3118 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C3119 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3120 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3121 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.42fF
C3122 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C3123 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3124 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.02fF
C3125 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C3126 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3127 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3130 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3131 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3132 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3133 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3134 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C3135 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C3136 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.01fF
C3137 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.02fF
C3138 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3139 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C3141 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C3142 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.00fF
C3143 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.01fF
C3144 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# 0.00fF
C3145 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.02fF
C3146 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C3147 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3148 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3150 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.01fF
C3151 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3152 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C3153 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3154 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C3155 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C3156 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C3157 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C3158 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C3159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C3160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3162 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3163 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3164 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C3165 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3166 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.01fF
C3167 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3168 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C3169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C3170 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.02fF
C3171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# -0.00fF
C3172 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3173 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3174 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C3175 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C3176 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# -0.00fF
C3177 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C3178 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3179 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3183 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C3184 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3185 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3186 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C3187 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C3188 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3189 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C3190 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3191 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C3192 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C3193 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3194 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C3195 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C3196 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3197 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C3198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C3199 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3200 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C3201 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3202 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C3203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C3204 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3206 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# -0.00fF
C3207 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C3208 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C3209 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3210 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C3211 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C3212 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C3213 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C3214 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3215 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C3216 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3217 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3218 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C3219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C3220 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.01fF
C3221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3222 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C3223 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3224 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# -0.00fF
C3225 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C3226 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C3227 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C3228 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C3229 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3230 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3231 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C3232 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3233 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C3234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C3235 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C3236 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3237 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.02fF
C3238 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.01fF
C3239 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3240 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C3241 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3242 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3243 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C3244 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3245 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C3246 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3247 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3248 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C3249 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C3250 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# -0.00fF
C3251 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3252 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3253 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3254 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.01fF
C3255 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C3256 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3257 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3258 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.00fF
C3259 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3260 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.01fF
C3261 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3262 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3263 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3264 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C3265 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3266 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3267 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C3268 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3269 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C3270 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.02fF
C3271 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C3272 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C3273 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C3274 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.22fF
C3275 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C3276 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# 0.00fF
C3277 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3278 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C3279 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3280 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C3281 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C3282 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C3283 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C3284 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3285 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.01fF
C3286 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3287 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C3288 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3289 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.02fF
C3290 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3291 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C3292 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C3293 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3294 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C3295 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3296 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C3297 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.01fF
C3298 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C3299 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.01fF
C3300 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C3301 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3302 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3303 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3304 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3305 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3306 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3307 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C3308 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3309 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.02fF
C3310 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# -0.00fF
C3311 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.02fF
C3312 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3313 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# -0.00fF
C3314 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3315 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3316 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C3318 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3320 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C3321 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C3322 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3323 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C3324 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3325 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C3326 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C3327 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C3328 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3329 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C3330 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3331 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C3332 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3333 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C3334 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.02fF
C3335 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C3336 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C3337 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C3338 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3339 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C3340 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C3341 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3342 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3343 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C3344 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# 0.00fF
C3345 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.01fF
C3346 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C3347 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3348 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C3349 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C3350 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C3351 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C3352 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3353 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.01fF
C3354 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C3355 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3356 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3357 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C3358 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C3359 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3360 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3361 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3362 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# -0.00fF
C3363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C3364 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# -0.00fF
C3365 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C3366 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3367 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C3368 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C3369 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C3370 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# -0.00fF
C3371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3372 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3373 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.02fF
C3374 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C3375 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C3376 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3377 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3378 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C3379 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.93fF
C3380 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# -0.00fF
C3381 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3382 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3383 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.02fF
C3384 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C3385 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C3386 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# -0.00fF
C3387 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.44fF
C3389 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C3390 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C3391 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C3392 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C3393 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C3394 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C3395 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C3396 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.00fF
C3397 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.02fF
C3398 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C3399 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3400 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3401 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C3402 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C3405 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3406 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3407 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C3408 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# -0.00fF
C3409 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3410 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3411 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.48fF
C3413 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C3414 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3415 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C3416 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C3417 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3418 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C3419 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3420 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3421 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C3422 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.93fF
C3424 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C3426 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3427 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3428 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C3429 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3430 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C3431 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3432 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C3433 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C3434 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.02fF
C3435 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C3436 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C3437 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C3438 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C3440 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3441 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C3442 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# -0.00fF
C3443 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# -0.00fF
C3444 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C3445 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C3446 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C3447 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3448 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# -0.00fF
C3449 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C3450 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3451 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3452 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3453 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# -0.00fF
C3454 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C3455 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C3457 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3458 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C3459 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3460 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3461 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C3462 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C3463 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C3464 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.02fF
C3465 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3466 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.01fF
C3467 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C3468 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# 0.00fF
C3469 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3470 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3471 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C3472 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C3473 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3474 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3475 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C3476 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C3477 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C3478 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3479 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3480 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C3481 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.02fF
C3483 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C3484 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C3485 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3486 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3487 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3488 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C3489 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.02fF
C3490 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C3491 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3492 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3493 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.02fF
C3494 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C3495 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C3496 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.02fF
C3497 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3498 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C3499 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C3500 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C3501 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3502 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3503 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3504 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C3505 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# -0.00fF
C3506 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.42fF
C3507 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3508 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C3509 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.01fF
C3510 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3511 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C3512 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C3513 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3514 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C3515 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.01fF
C3516 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.02fF
C3517 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C3518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3519 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# -0.00fF
C3520 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C3521 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3522 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.02fF
C3523 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C3524 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3525 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3526 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C3527 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C3528 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3529 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3530 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C3531 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C3532 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C3533 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C3534 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C3535 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C3536 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C3537 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.02fF
C3538 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C3539 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C3540 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3541 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3542 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3543 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C3544 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C3545 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C3546 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C3547 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.00fF
C3548 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C3549 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C3550 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C3551 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3552 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C3553 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.02fF
C3554 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C3555 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C3556 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C3557 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C3558 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3559 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3560 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C3561 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3562 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3563 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C3564 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C3565 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# -0.00fF
C3566 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C3567 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C3568 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C3570 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3571 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.31fF
C3572 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.02fF
C3573 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.42fF
C3574 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3575 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C3576 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3577 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C3578 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3579 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3580 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.01fF
C3581 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3582 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C3583 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C3584 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C3585 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3586 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3587 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.02fF
C3588 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3589 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C3590 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C3591 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C3592 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3593 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C3594 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C3595 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C3596 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C3597 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.00fF
C3598 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3599 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3600 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C3601 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C3602 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3603 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C3604 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C3606 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3607 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3608 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3609 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C3610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C3611 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# -0.00fF
C3612 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C3613 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.02fF
C3614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3615 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C3616 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C3617 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C3618 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3619 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C3620 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.02fF
C3621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3622 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C3623 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3625 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3626 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C3627 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.02fF
C3628 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.27fF
C3629 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C3630 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3631 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C3632 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3633 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C3634 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C3635 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C3637 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.02fF
C3638 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3639 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C3640 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C3641 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.02fF
C3642 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.02fF
C3643 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C3644 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3645 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3646 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C3647 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C3648 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.01fF
C3649 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3650 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3651 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C3652 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3653 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3654 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3655 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3656 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3657 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C3658 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3659 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 1.18fF
C3660 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3661 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C3662 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3663 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3664 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3665 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C3666 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C3667 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3668 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C3669 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3670 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C3671 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3672 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3673 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C3674 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3675 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C3676 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3677 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3678 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C3679 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3680 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C3681 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C3682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C3683 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C3684 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.02fF
C3685 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C3686 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3687 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C3688 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C3689 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C3690 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3691 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# -0.00fF
C3692 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3693 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3694 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3695 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3696 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C3697 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C3698 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C3699 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C3700 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# -0.00fF
C3701 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3702 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3703 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C3704 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.02fF
C3705 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3706 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3708 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3709 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C3710 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C3711 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3712 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# -0.00fF
C3713 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3714 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C3715 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C3716 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3717 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C3718 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3719 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C3720 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C3721 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3722 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C3723 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C3724 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3725 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3726 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3727 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C3728 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C3729 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C3730 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3731 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# -0.00fF
C3732 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3733 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3734 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.02fF
C3735 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3736 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3737 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3738 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C3739 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3740 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C3741 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3742 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C3743 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C3744 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.02fF
C3745 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C3746 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C3747 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# -0.00fF
C3748 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# -0.00fF
C3749 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3750 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3751 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C3752 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C3753 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C3754 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C3755 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3756 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3757 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3758 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C3759 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C3760 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C3761 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3762 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C3763 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C3764 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3765 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C3766 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C3767 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3768 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3769 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3770 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C3771 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C3772 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3773 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3774 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# -0.00fF
C3775 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C3776 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.02fF
C3777 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3778 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3779 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C3780 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C3781 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C3782 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.02fF
C3783 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C3784 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C3785 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3786 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3787 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3788 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3789 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3790 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C3791 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3792 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3793 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3794 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C3795 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C3796 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.01fF
C3797 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3798 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.27fF
C3799 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C3800 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.02fF
C3801 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C3802 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3803 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C3805 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C3806 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3807 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.02fF
C3808 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3809 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C3810 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3811 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3812 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C3813 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C3814 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C3815 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3816 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C3817 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C3818 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3819 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3820 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3821 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C3822 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.19fF
C3823 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.02fF
C3824 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3825 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3826 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3827 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.02fF
C3828 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C3830 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3831 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3832 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.02fF
C3833 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C3834 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C3835 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C3836 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3837 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3838 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3839 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3840 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C3841 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3842 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C3843 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3844 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# 0.01fF
C3845 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C3846 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3847 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C3848 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C3849 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C3850 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.00fF
C3851 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# -0.00fF
C3852 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C3853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C3854 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C3855 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C3856 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C3857 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3858 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.02fF
C3859 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3860 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# -0.00fF
C3861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3862 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C3863 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C3864 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3865 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C3866 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3867 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# -0.00fF
C3868 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.01fF
C3869 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C3870 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C3871 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.02fF
C3872 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C3873 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.02fF
C3874 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3875 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.02fF
C3876 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C3877 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3878 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C3879 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C3880 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C3881 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3882 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3883 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.02fF
C3884 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C3885 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.02fF
C3886 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C3887 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C3888 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.02fF
C3889 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C3890 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3891 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C3892 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.01fF
C3893 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3894 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3895 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3896 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3897 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3898 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# -0.00fF
C3899 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3900 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3901 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.02fF
C3902 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# -0.00fF
C3903 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3904 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C3905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.02fF
C3906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# -0.00fF
C3907 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C3908 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3909 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3910 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C3911 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3912 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3913 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3914 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3915 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C3916 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C3917 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C3918 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C3919 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C3920 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C3921 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3922 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.01fF
C3923 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C3924 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3925 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C3926 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.02fF
C3927 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3928 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3929 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C3930 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C3931 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3932 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C3933 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3934 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C3935 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C3936 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3937 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C3938 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C3939 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3940 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3941 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.01fF
C3942 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# -0.00fF
C3943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C3944 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3945 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3946 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C3947 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C3948 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3949 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3950 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# -0.00fF
C3951 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3952 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C3953 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C3954 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C3955 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3956 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C3957 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3958 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C3959 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3960 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C3961 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C3962 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C3963 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3964 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C3965 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C3966 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C3967 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3968 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3969 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C3970 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C3971 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3972 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3973 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3974 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3975 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3976 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C3977 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3978 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3979 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3980 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3981 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C3982 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C3983 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C3984 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3985 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.00fF
C3986 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3987 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C3988 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3989 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C3990 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.02fF
C3991 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C3992 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C3993 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C3994 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C3995 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3996 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C3997 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C3998 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C3999 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C4000 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C4001 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4002 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.01fF
C4003 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C4004 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4006 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# -0.00fF
C4007 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4008 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C4009 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4010 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.01fF
C4011 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4012 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4013 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C4014 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.02fF
C4015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C4016 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C4017 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C4018 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4019 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4020 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.00fF
C4021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# -0.00fF
C4022 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C4023 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.02fF
C4024 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C4025 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C4026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4027 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C4028 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C4029 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4030 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C4032 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C4033 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C4034 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.01fF
C4035 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# -0.00fF
C4036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C4037 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4038 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C4039 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4040 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C4041 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C4042 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.01fF
C4043 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4044 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C4045 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4046 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.02fF
C4047 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C4048 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C4049 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4050 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C4051 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.31fF
C4052 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C4053 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C4054 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C4055 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.01fF
C4056 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C4057 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C4058 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C4059 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4060 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.02fF
C4061 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C4062 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4063 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C4064 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C4065 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4066 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# -0.00fF
C4067 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4068 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C4069 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.57fF
C4070 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4071 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.01fF
C4072 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.00fF
C4073 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4074 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4075 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C4076 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4077 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C4078 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C4079 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C4080 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# -0.00fF
C4081 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4082 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4083 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4084 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4085 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C4086 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C4087 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.27fF
C4088 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C4089 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4090 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4091 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C4092 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C4093 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C4094 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4095 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4096 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C4097 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4098 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.02fF
C4099 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C4100 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4101 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C4102 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4103 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C4104 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C4105 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4106 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C4107 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4108 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.02fF
C4109 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.02fF
C4110 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4111 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C4112 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.02fF
C4113 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4114 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C4115 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4118 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C4119 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.02fF
C4120 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.02fF
C4121 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C4122 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C4123 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.02fF
C4124 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4125 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C4126 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C4127 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C4128 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C4129 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4130 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4131 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4132 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C4133 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4134 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C4135 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C4136 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C4137 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4138 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C4139 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4140 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4141 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.02fF
C4142 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C4143 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4144 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4145 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C4146 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4147 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4148 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C4149 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4150 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.01fF
C4151 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.01fF
C4152 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4153 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# -0.00fF
C4154 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C4155 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4156 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C4157 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.01fF
C4158 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C4159 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# -0.00fF
C4161 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.02fF
C4162 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.02fF
C4163 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C4164 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C4165 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4166 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C4167 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4168 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C4169 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4170 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.02fF
C4171 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4172 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C4173 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4174 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C4175 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C4176 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C4177 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4178 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C4179 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C4180 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C4181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C4182 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C4183 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4184 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C4185 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4186 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C4187 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C4188 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4189 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4190 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C4191 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.02fF
C4192 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C4193 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# -0.00fF
C4194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4195 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C4196 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C4197 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C4198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.02fF
C4199 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C4200 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4201 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C4202 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C4203 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C4205 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4206 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.27fF
C4207 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4208 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C4209 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C4210 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C4211 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C4212 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4213 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4214 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.02fF
C4215 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C4216 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4217 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# -0.00fF
C4218 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C4219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C4220 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C4221 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4222 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.19fF
C4223 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4224 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C4225 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4226 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C4227 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.02fF
C4228 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4229 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4230 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C4231 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 1.18fF
C4232 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C4233 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4234 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.02fF
C4235 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4236 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C4237 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4238 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C4239 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C4240 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C4241 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4242 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4243 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.02fF
C4244 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4245 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C4246 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# -0.00fF
C4247 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4248 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4249 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.42fF
C4250 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4251 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C4252 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C4253 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C4254 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C4255 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.01fF
C4256 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C4257 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.02fF
C4258 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C4259 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.02fF
C4260 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C4261 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C4262 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.57fF
C4263 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C4264 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C4265 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4266 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.01fF
C4268 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C4269 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C4270 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C4271 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4272 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.22fF
C4273 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C4274 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# -0.00fF
C4275 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4276 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C4277 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C4278 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C4279 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C4280 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4281 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4283 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4284 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C4285 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4286 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C4287 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C4288 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C4289 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4290 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4291 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4292 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4293 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# -0.00fF
C4294 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4295 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4296 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4297 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4298 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C4299 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C4300 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4301 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C4302 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.02fF
C4303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4304 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C4305 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C4306 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4307 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C4308 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C4309 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C4310 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.42fF
C4311 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C4312 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4313 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C4314 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C4315 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4316 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4317 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C4318 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C4319 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4320 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4321 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4322 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4323 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C4324 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C4325 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C4326 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4327 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C4328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4329 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.00fF
C4330 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4331 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4332 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C4333 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4334 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4335 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C4336 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C4337 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4338 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C4339 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C4340 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.02fF
C4341 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C4342 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C4343 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4344 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C4345 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4346 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C4347 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4348 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C4349 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4350 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# -0.00fF
C4351 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4352 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C4353 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# -0.00fF
C4354 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4355 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4356 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C4357 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C4358 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.02fF
C4359 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4360 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C4361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C4362 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4363 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C4364 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C4365 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4366 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.01fF
C4367 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C4368 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C4369 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C4372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C4373 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C4374 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.02fF
C4375 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C4376 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4378 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4379 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4380 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4381 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C4382 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C4383 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C4384 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C4385 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C4386 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4387 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C4388 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.02fF
C4389 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4390 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C4391 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C4392 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C4393 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4394 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4395 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C4396 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C4397 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C4398 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.01fF
C4399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C4400 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4401 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.01fF
C4402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.02fF
C4403 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4404 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C4405 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C4406 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C4407 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.02fF
C4408 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4409 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C4410 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C4411 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C4412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C4413 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# -0.00fF
C4414 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C4415 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.02fF
C4416 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4417 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C4418 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# 0.00fF
C4419 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4420 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4421 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4422 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.57fF
C4423 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4424 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4425 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.02fF
C4426 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# -0.00fF
C4427 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C4428 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4429 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.31fF
C4430 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C4431 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C4432 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C4433 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C4434 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C4435 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C4436 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C4437 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C4438 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C4439 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.27fF
C4440 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4441 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C4442 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C4443 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.01fF
C4444 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# -0.00fF
C4445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4446 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4447 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C4448 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4449 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4450 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C4451 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4452 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C4453 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C4454 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4455 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4456 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C4457 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C4458 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4459 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C4460 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C4461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C4462 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4463 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C4464 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C4465 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.01fF
C4466 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4467 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C4468 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4469 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C4470 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C4471 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4472 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# 0.02fF
C4473 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4474 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4475 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4476 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.02fF
C4477 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C4478 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4479 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4480 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C4481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4482 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.02fF
C4483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C4484 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4485 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C4486 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4487 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C4488 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4489 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C4490 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C4491 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4492 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C4493 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C4494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C4495 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C4496 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C4497 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4498 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4499 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.01fF
C4500 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C4501 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# -0.00fF
C4502 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4503 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4504 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C4505 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4506 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C4507 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.02fF
C4508 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C4509 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C4510 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C4511 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C4512 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4513 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C4514 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4515 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C4516 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4517 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C4518 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C4519 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4520 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4521 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C4522 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C4523 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4524 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4525 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.02fF
C4526 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C4527 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4528 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C4529 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4530 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4531 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4532 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C4533 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4534 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4535 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C4536 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C4537 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C4538 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C4539 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4540 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4541 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C4542 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# -0.00fF
C4543 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C4544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4545 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4546 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C4547 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4548 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C4549 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4550 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4551 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C4552 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4553 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4554 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4555 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4556 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C4557 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4558 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C4559 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C4560 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C4561 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C4562 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C4563 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C4564 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4565 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C4566 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4567 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C4568 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4569 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C4570 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C4571 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.02fF
C4572 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.01fF
C4573 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4574 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C4575 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 1.18fF
C4576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4577 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C4578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C4579 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C4580 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.02fF
C4581 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4582 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C4583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4584 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C4585 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4586 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C4587 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C4588 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4589 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4590 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C4591 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4592 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.02fF
C4593 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4594 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C4595 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C4597 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.01fF
C4598 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C4599 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4600 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# -0.00fF
C4601 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C4602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C4603 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C4604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C4605 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C4606 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C4607 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C4608 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C4609 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C4610 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.01fF
C4611 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C4612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4613 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4614 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C4615 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4616 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C4617 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C4618 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4619 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C4620 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C4621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C4622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C4623 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C4624 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C4625 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C4626 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C4627 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4628 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4629 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4630 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C4631 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C4632 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C4633 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C4634 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# -0.00fF
C4635 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4636 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# 0.00fF
C4637 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4638 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C4639 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C4640 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C4641 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C4642 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4643 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C4644 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C4645 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.01fF
C4646 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C4647 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4648 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C4649 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4650 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C4651 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C4652 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4653 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C4654 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C4655 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4656 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4657 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C4658 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4659 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C4660 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C4661 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C4662 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C4663 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C4664 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C4665 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# -0.00fF
C4666 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4667 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4668 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C4669 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C4670 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C4671 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C4672 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C4673 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C4674 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4675 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C4676 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4677 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4678 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C4679 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C4680 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4681 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.02fF
C4682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C4683 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4684 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C4685 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4686 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4687 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C4688 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4689 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C4691 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4692 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C4693 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4694 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C4695 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C4696 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C4697 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C4698 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.02fF
C4699 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C4700 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# -0.00fF
C4701 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4702 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.02fF
C4703 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4704 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4705 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4706 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C4707 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C4708 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C4709 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4710 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# -0.00fF
C4711 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C4712 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4713 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4714 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C4715 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4716 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C4717 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4718 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4719 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# -0.00fF
C4720 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4721 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C4722 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C4723 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C4724 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C4725 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C4726 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C4727 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C4728 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4729 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C4730 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C4731 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C4732 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4733 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4734 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C4735 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4736 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C4737 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C4738 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4739 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C4740 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# 0.00fF
C4741 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C4742 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C4743 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4744 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C4745 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C4746 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4747 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4748 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C4749 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C4750 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4751 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C4752 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C4753 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4754 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C4755 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# -0.00fF
C4756 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C4757 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.02fF
C4758 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C4759 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4760 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4761 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4762 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C4763 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4764 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C4765 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4766 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4767 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C4768 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C4769 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4770 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4771 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4772 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C4773 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4774 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4775 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4776 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C4777 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C4778 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C4779 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4780 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.01fF
C4781 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4782 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.48fF
C4783 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4784 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4785 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C4786 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C4787 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C4788 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.02fF
C4789 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4790 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C4791 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C4792 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4793 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C4794 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C4795 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4796 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C4797 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4798 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C4799 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C4800 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4801 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4802 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C4803 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.01fF
C4804 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C4805 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4806 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C4807 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C4808 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4809 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4810 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4811 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4812 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C4813 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C4814 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C4815 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.00fF
C4816 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C4817 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4818 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.01fF
C4819 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C4820 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C4821 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C4822 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.93fF
C4823 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C4824 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C4825 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C4826 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C4827 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C4828 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4829 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C4830 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C4831 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C4832 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C4833 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C4834 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4835 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4836 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4837 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C4838 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.00fF
C4839 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# -0.00fF
C4840 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C4841 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C4842 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# -0.00fF
C4843 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# -0.00fF
C4844 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.93fF
C4845 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4846 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4847 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C4848 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C4849 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C4850 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C4851 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.02fF
C4852 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C4853 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4854 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C4855 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C4856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# VSUBS 1.08fF
C4857 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# VSUBS 1.03fF
C4858 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# VSUBS 0.11fF
C4859 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# VSUBS 0.17fF
C4860 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# VSUBS 0.10fF
C4861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# VSUBS 0.09fF
C4862 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# VSUBS 0.11fF
C4863 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# VSUBS 0.11fF
C4864 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# VSUBS 0.12fF
C4865 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# VSUBS 0.11fF
C4866 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# VSUBS 0.12fF
C4867 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# VSUBS 0.12fF
C4868 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# VSUBS 0.12fF
C4869 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# VSUBS 0.12fF
C4870 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# VSUBS 0.12fF
C4871 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# VSUBS 0.12fF
C4872 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# VSUBS 0.12fF
C4873 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# VSUBS 0.12fF
C4874 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# VSUBS 0.12fF
C4875 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# VSUBS 0.12fF
C4876 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# VSUBS 0.12fF
C4877 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# VSUBS 0.12fF
C4878 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# VSUBS 0.12fF
C4879 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# VSUBS 0.12fF
C4880 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# VSUBS 0.12fF
C4881 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# VSUBS 0.12fF
C4882 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# VSUBS 0.12fF
C4883 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# VSUBS 0.12fF
C4884 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# VSUBS 0.12fF
C4885 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# VSUBS 0.12fF
C4886 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# VSUBS 0.12fF
C4887 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# VSUBS 0.12fF
C4888 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# VSUBS 0.12fF
C4889 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# VSUBS 0.12fF
C4890 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# VSUBS 0.12fF
C4891 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# VSUBS 0.12fF
C4892 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# VSUBS 0.12fF
C4893 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# VSUBS 0.12fF
C4894 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# VSUBS 0.12fF
C4895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# VSUBS 0.12fF
C4896 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# VSUBS 0.12fF
C4897 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# VSUBS 0.12fF
C4898 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# VSUBS 0.20fF
C4899 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# VSUBS 0.13fF
C4900 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# VSUBS 1.08fF
C4901 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# VSUBS 1.03fF
C4902 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# VSUBS 0.11fF
C4903 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# VSUBS 0.17fF
C4904 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# VSUBS 0.10fF
C4905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# VSUBS 0.09fF
C4906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# VSUBS 0.11fF
C4907 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# VSUBS 0.11fF
C4908 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# VSUBS 0.12fF
C4909 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# VSUBS 0.11fF
C4910 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# VSUBS 0.12fF
C4911 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# VSUBS 0.12fF
C4912 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# VSUBS 0.12fF
C4913 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# VSUBS 0.12fF
C4914 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# VSUBS 0.12fF
C4915 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# VSUBS 0.12fF
C4916 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# VSUBS 0.12fF
C4917 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# VSUBS 0.12fF
C4918 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# VSUBS 0.12fF
C4919 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# VSUBS 0.12fF
C4920 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# VSUBS 0.12fF
C4921 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# VSUBS 0.12fF
C4922 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# VSUBS 0.12fF
C4923 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# VSUBS 0.12fF
C4924 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# VSUBS 0.12fF
C4925 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# VSUBS 0.12fF
C4926 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# VSUBS 0.12fF
C4927 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# VSUBS 0.12fF
C4928 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# VSUBS 0.12fF
C4929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# VSUBS 0.12fF
C4930 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# VSUBS 0.12fF
C4931 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# VSUBS 0.12fF
C4932 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# VSUBS 0.12fF
C4933 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# VSUBS 0.12fF
C4934 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# VSUBS 0.12fF
C4935 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# VSUBS 0.12fF
C4936 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# VSUBS 0.12fF
C4937 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# VSUBS 0.12fF
C4938 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# VSUBS 0.12fF
C4939 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# VSUBS 0.12fF
C4940 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# VSUBS 0.12fF
C4941 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# VSUBS 0.12fF
C4942 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# VSUBS 0.20fF
C4943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# VSUBS 0.13fF
C4944 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# VSUBS 1.08fF
C4945 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# VSUBS 1.03fF
C4946 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# VSUBS 0.11fF
C4947 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# VSUBS 0.17fF
C4948 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# VSUBS 0.10fF
C4949 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# VSUBS 0.09fF
C4950 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# VSUBS 0.11fF
C4951 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# VSUBS 0.11fF
C4952 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# VSUBS 0.12fF
C4953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# VSUBS 0.11fF
C4954 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# VSUBS 0.12fF
C4955 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# VSUBS 0.12fF
C4956 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# VSUBS 0.12fF
C4957 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# VSUBS 0.12fF
C4958 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# VSUBS 0.12fF
C4959 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# VSUBS 0.12fF
C4960 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# VSUBS 0.12fF
C4961 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# VSUBS 0.12fF
C4962 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# VSUBS 0.12fF
C4963 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# VSUBS 0.12fF
C4964 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# VSUBS 0.12fF
C4965 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# VSUBS 0.12fF
C4966 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# VSUBS 0.12fF
C4967 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# VSUBS 0.12fF
C4968 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# VSUBS 0.12fF
C4969 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# VSUBS 0.12fF
C4970 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# VSUBS 0.12fF
C4971 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# VSUBS 0.12fF
C4972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# VSUBS 0.12fF
C4973 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# VSUBS 0.12fF
C4974 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# VSUBS 0.12fF
C4975 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# VSUBS 0.12fF
C4976 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# VSUBS 0.12fF
C4977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# VSUBS 0.12fF
C4978 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# VSUBS 0.12fF
C4979 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# VSUBS 0.12fF
C4980 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# VSUBS 0.12fF
C4981 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# VSUBS 0.12fF
C4982 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# VSUBS 0.12fF
C4983 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# VSUBS 0.12fF
C4984 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# VSUBS 0.12fF
C4985 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# VSUBS 0.12fF
C4986 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS 0.20fF
C4987 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# VSUBS 0.13fF
C4988 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# VSUBS 1.08fF
C4989 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# VSUBS 1.03fF
C4990 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# VSUBS 0.11fF
C4991 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# VSUBS 0.17fF
C4992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# VSUBS 0.10fF
C4993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# VSUBS 0.09fF
C4994 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# VSUBS 0.11fF
C4995 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# VSUBS 0.11fF
C4996 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# VSUBS 0.12fF
C4997 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# VSUBS 0.11fF
C4998 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# VSUBS 0.12fF
C4999 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# VSUBS 0.12fF
C5000 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# VSUBS 0.12fF
C5001 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# VSUBS 0.12fF
C5002 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# VSUBS 0.12fF
C5003 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# VSUBS 0.12fF
C5004 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# VSUBS 0.12fF
C5005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# VSUBS 0.12fF
C5006 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# VSUBS 0.12fF
C5007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# VSUBS 0.12fF
C5008 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# VSUBS 0.12fF
C5009 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# VSUBS 0.12fF
C5010 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# VSUBS 0.12fF
C5011 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# VSUBS 0.12fF
C5012 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# VSUBS 0.12fF
C5013 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# VSUBS 0.12fF
C5014 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# VSUBS 0.12fF
C5015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# VSUBS 0.12fF
C5016 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# VSUBS 0.12fF
C5017 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# VSUBS 0.12fF
C5018 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# VSUBS 0.12fF
C5019 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# VSUBS 0.12fF
C5020 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# VSUBS 0.12fF
C5021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# VSUBS 0.12fF
C5022 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# VSUBS 0.12fF
C5023 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# VSUBS 0.12fF
C5024 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# VSUBS 0.12fF
C5025 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# VSUBS 0.12fF
C5026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# VSUBS 0.12fF
C5027 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# VSUBS 0.12fF
C5028 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# VSUBS 0.12fF
C5029 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# VSUBS 0.12fF
C5030 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# VSUBS 0.20fF
C5031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# VSUBS 0.13fF
C5032 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# VSUBS 1.08fF
C5033 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# VSUBS 1.03fF
C5034 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# VSUBS 0.11fF
C5035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# VSUBS 0.17fF
C5036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# VSUBS 0.10fF
C5037 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# VSUBS 0.09fF
C5038 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# VSUBS 0.11fF
C5039 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# VSUBS 0.11fF
C5040 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# VSUBS 0.12fF
C5041 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# VSUBS 0.11fF
C5042 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# VSUBS 0.12fF
C5043 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# VSUBS 0.12fF
C5044 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# VSUBS 0.12fF
C5045 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# VSUBS 0.12fF
C5046 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# VSUBS 0.12fF
C5047 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# VSUBS 0.12fF
C5048 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# VSUBS 0.12fF
C5049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# VSUBS 0.12fF
C5050 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# VSUBS 0.12fF
C5051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# VSUBS 0.12fF
C5052 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# VSUBS 0.12fF
C5053 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# VSUBS 0.12fF
C5054 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# VSUBS 0.12fF
C5055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# VSUBS 0.12fF
C5056 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# VSUBS 0.12fF
C5057 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# VSUBS 0.12fF
C5058 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# VSUBS 0.12fF
C5059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# VSUBS 0.12fF
C5060 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# VSUBS 0.12fF
C5061 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# VSUBS 0.12fF
C5062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# VSUBS 0.12fF
C5063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# VSUBS 0.12fF
C5064 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# VSUBS 0.12fF
C5065 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# VSUBS 0.12fF
C5066 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# VSUBS 0.12fF
C5067 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# VSUBS 0.12fF
C5068 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# VSUBS 0.12fF
C5069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# VSUBS 0.12fF
C5070 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# VSUBS 0.12fF
C5071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# VSUBS 0.12fF
C5072 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# VSUBS 0.12fF
C5073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# VSUBS 0.12fF
C5074 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# VSUBS 0.20fF
C5075 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# VSUBS 0.13fF
C5076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# VSUBS 1.08fF
C5077 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# VSUBS 1.03fF
C5078 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# VSUBS 0.11fF
C5079 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# VSUBS 0.17fF
C5080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# VSUBS 0.10fF
C5081 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# VSUBS 0.09fF
C5082 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# VSUBS 0.11fF
C5083 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# VSUBS 0.11fF
C5084 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# VSUBS 0.12fF
C5085 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# VSUBS 0.11fF
C5086 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# VSUBS 0.12fF
C5087 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# VSUBS 0.12fF
C5088 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# VSUBS 0.12fF
C5089 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# VSUBS 0.12fF
C5090 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# VSUBS 0.12fF
C5091 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# VSUBS 0.12fF
C5092 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# VSUBS 0.12fF
C5093 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# VSUBS 0.12fF
C5094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# VSUBS 0.12fF
C5095 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# VSUBS 0.12fF
C5096 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# VSUBS 0.12fF
C5097 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# VSUBS 0.12fF
C5098 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# VSUBS 0.12fF
C5099 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# VSUBS 0.12fF
C5100 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# VSUBS 0.12fF
C5101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# VSUBS 0.12fF
C5102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# VSUBS 0.12fF
C5103 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# VSUBS 0.12fF
C5104 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# VSUBS 0.12fF
C5105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# VSUBS 0.12fF
C5106 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# VSUBS 0.12fF
C5107 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# VSUBS 0.12fF
C5108 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# VSUBS 0.12fF
C5109 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# VSUBS 0.12fF
C5110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# VSUBS 0.12fF
C5111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# VSUBS 0.12fF
C5112 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# VSUBS 0.12fF
C5113 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# VSUBS 0.12fF
C5114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# VSUBS 0.12fF
C5115 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# VSUBS 0.12fF
C5116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# VSUBS 0.12fF
C5117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# VSUBS 0.12fF
C5118 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# VSUBS 0.20fF
C5119 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# VSUBS 0.13fF
C5120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# VSUBS 1.08fF
C5121 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# VSUBS 1.03fF
C5122 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# VSUBS 0.11fF
C5123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# VSUBS 0.17fF
C5124 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# VSUBS 0.10fF
C5125 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# VSUBS 0.09fF
C5126 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# VSUBS 0.11fF
C5127 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# VSUBS 0.11fF
C5128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# VSUBS 0.12fF
C5129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# VSUBS 0.11fF
C5130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# VSUBS 0.12fF
C5131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# VSUBS 0.12fF
C5132 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# VSUBS 0.12fF
C5133 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# VSUBS 0.12fF
C5134 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# VSUBS 0.12fF
C5135 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# VSUBS 0.12fF
C5136 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# VSUBS 0.12fF
C5137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# VSUBS 0.12fF
C5138 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# VSUBS 0.12fF
C5139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# VSUBS 0.12fF
C5140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# VSUBS 0.12fF
C5141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# VSUBS 0.12fF
C5142 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# VSUBS 0.12fF
C5143 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# VSUBS 0.12fF
C5144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# VSUBS 0.12fF
C5145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# VSUBS 0.12fF
C5146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# VSUBS 0.12fF
C5147 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# VSUBS 0.12fF
C5148 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# VSUBS 0.12fF
C5149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# VSUBS 0.12fF
C5150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# VSUBS 0.12fF
C5151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# VSUBS 0.12fF
C5152 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# VSUBS 0.12fF
C5153 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# VSUBS 0.12fF
C5154 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# VSUBS 0.12fF
C5155 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# VSUBS 0.12fF
C5156 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# VSUBS 0.12fF
C5157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# VSUBS 0.12fF
C5158 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# VSUBS 0.12fF
C5159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# VSUBS 0.12fF
C5160 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# VSUBS 0.12fF
C5161 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# VSUBS 0.12fF
C5162 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# VSUBS 0.20fF
C5163 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# VSUBS 0.13fF
C5164 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# VSUBS 1.08fF
C5165 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# VSUBS 1.03fF
C5166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# VSUBS 0.11fF
C5167 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# VSUBS 0.17fF
C5168 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# VSUBS 0.10fF
C5169 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# VSUBS 0.09fF
C5170 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# VSUBS 0.11fF
C5171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# VSUBS 0.11fF
C5172 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# VSUBS 0.12fF
C5173 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# VSUBS 0.11fF
C5174 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# VSUBS 0.12fF
C5175 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# VSUBS 0.12fF
C5176 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# VSUBS 0.12fF
C5177 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# VSUBS 0.12fF
C5178 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# VSUBS 0.12fF
C5179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# VSUBS 0.12fF
C5180 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# VSUBS 0.12fF
C5181 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# VSUBS 0.12fF
C5182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# VSUBS 0.12fF
C5183 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# VSUBS 0.12fF
C5184 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# VSUBS 0.12fF
C5185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# VSUBS 0.12fF
C5186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# VSUBS 0.12fF
C5187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# VSUBS 0.12fF
C5188 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# VSUBS 0.12fF
C5189 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# VSUBS 0.12fF
C5190 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# VSUBS 0.12fF
C5191 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# VSUBS 0.12fF
C5192 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# VSUBS 0.12fF
C5193 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# VSUBS 0.12fF
C5194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# VSUBS 0.12fF
C5195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# VSUBS 0.12fF
C5196 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# VSUBS 0.12fF
C5197 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# VSUBS 0.12fF
C5198 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# VSUBS 0.12fF
C5199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# VSUBS 0.12fF
C5200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# VSUBS 0.12fF
C5201 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# VSUBS 0.12fF
C5202 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# VSUBS 0.12fF
C5203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# VSUBS 0.12fF
C5204 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# VSUBS 0.12fF
C5205 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# VSUBS 0.12fF
C5206 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# VSUBS 0.20fF
C5207 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# VSUBS 0.13fF
.ends

.subckt comparator_v2 clk outp VSS sky130_fd_sc_hd__buf_2_1/a_27_47# outn sky130_fd_sc_hd__buf_2_0/X
+ sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_1/X
+ VDD li_n2324_818# li_940_3458# li_940_818# ip sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ in sky130_fd_sc_hd__buf_2_1/A
Xlatch_pmos_pair_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VDD VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD latch_pmos_pair
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__buf_2_1/X outp VSS VDD outn VSS VDD sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__buf_2_0/X outn VSS VDD outp VSS VDD sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_pr__pfet_01v8_VCG74W_1 li_940_3458# li_940_3458# li_940_3458# clk VDD VDD
+ clk clk li_940_3458# li_940_3458# li_940_3458# clk VDD VDD clk clk VDD li_940_3458#
+ clk clk VDD clk clk clk VDD VDD clk clk li_940_3458# li_940_3458# clk VDD clk clk
+ VSS sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk VDD sky130_fd_sc_hd__buf_2_1/A clk
+ clk VDD clk clk clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ clk VDD clk clk VSS sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_sc_hd__buf_2_0 sky130_fd_sc_hd__buf_2_0/A VSS VDD sky130_fd_sc_hd__buf_2_0/X
+ VSS VDD sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_1 sky130_fd_sc_hd__buf_2_1/A VSS VDD sky130_fd_sc_hd__buf_2_1/X
+ VSS VDD sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_0 clk sky130_fd_sc_hd__buf_2_0/A clk VDD VDD clk sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A clk sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A clk clk VDD VDD clk clk clk sky130_fd_sc_hd__buf_2_0/A
+ clk clk clk clk VSS precharge_pmos
Xcurrent_tail_0 li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# VSS VSS VSS
+ li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS VSS VSS li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS li_n2324_818# li_n2324_818# VSS VSS VSS clk li_n2324_818# VSS current_tail
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_1 clk li_940_818# clk VDD VDD clk li_940_818# li_940_818# li_940_818#
+ clk li_940_818# VDD VDD clk VDD VDD clk clk li_940_818# VDD li_940_818# li_940_818#
+ clk clk VDD VDD clk clk clk li_940_818# clk clk clk clk VSS precharge_pmos
Xlatch_nmos_pair_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A latch_nmos_pair
Xinput_diff_pair_0 ip ip ip in in VSS ip in in in in VSS li_940_3458# ip ip ip in
+ ip li_n2324_818# ip ip in ip ip ip in in in ip ip ip in ip in ip in ip in in ip
+ ip VSS ip ip in ip li_n2324_818# ip ip in in in ip ip ip in in in li_940_3458# in
+ in ip ip in ip in ip ip ip VSS ip in ip ip ip in in in ip ip in in ip in VSS ip
+ in in in in in ip in li_940_818# ip ip in ip ip li_n2324_818# in in ip ip ip in
+ ip ip ip ip in in in in in in VSS ip in in ip ip ip ip ip in in ip ip in in ip li_940_818#
+ ip ip in li_n2324_818# in in in VSS ip in in ip ip ip in ip ip ip in in ip in ip
+ in ip ip ip in in in in in VSS in ip li_n2324_818# ip ip in ip ip in ip ip in ip
+ ip li_940_3458# in in ip ip ip in in in ip ip in ip ip in in in VSS ip in VSS VSS
+ in in ip ip in in ip ip ip in in ip ip li_940_3458# in ip in ip ip in li_n2324_818#
+ ip in in in in in in ip ip in in ip ip ip ip VSS ip ip ip in in in in ip ip in ip
+ ip ip in in ip ip in in ip in in li_n2324_818# in in in in ip in in ip in ip li_940_818#
+ VSS ip ip ip ip in in ip ip VSS in in in ip in in ip ip ip in in ip in in VSS in
+ in li_n2324_818# ip in in in ip ip ip ip in in ip ip li_940_818# in ip ip in in
+ in ip in ip in ip ip ip in in in ip ip ip ip in in in ip ip in in in in ip VSS VSS
+ in in ip ip in in in input_diff_pair
C0 VDD li_940_818# 2.07fF
C1 clk sky130_fd_sc_hd__buf_2_0/A 3.33fF
C2 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_0/A 0.06fF
C3 outp VSS 0.44fF
C4 outn VSS 0.57fF
C5 sky130_fd_sc_hd__buf_2_0/X VDD 0.20fF
C6 VSS sky130_fd_sc_hd__buf_2_0/A 2.10fF
C7 sky130_fd_sc_hd__buf_2_1/A outp 0.05fF
C8 clk VDD 14.97fF
C9 sky130_fd_sc_hd__buf_2_1/A outn 0.03fF
C10 sky130_fd_sc_hd__buf_2_1/X VDD 0.24fF
C11 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A 76.00fF
C12 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_0/a_27_47# 0.11fF
C13 li_940_818# li_940_3458# 4.44fF
C14 li_n2324_818# in 49.83fF
C15 outn outp 1.34fF
C16 VSS VDD 0.85fF
C17 outp sky130_fd_sc_hd__buf_2_0/A 0.04fF
C18 outn sky130_fd_sc_hd__buf_2_0/A 0.05fF
C19 sky130_fd_sc_hd__buf_2_1/A VDD 26.42fF
C20 clk li_940_3458# 2.09fF
C21 VSS sky130_fd_sc_hd__buf_2_0/a_27_47# 0.03fF
C22 outp VDD 0.83fF
C23 li_940_818# ip 35.81fF
C24 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/a_27_47# 0.02fF
C25 outn VDD 0.93fF
C26 VSS li_940_3458# 1.22fF
C27 VDD sky130_fd_sc_hd__buf_2_0/A 30.94fF
C28 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.03fF
C29 sky130_fd_sc_hd__buf_2_1/A li_940_3458# 9.09fF
C30 outp sky130_fd_sc_hd__buf_2_0/a_27_47# 0.04fF
C31 outn sky130_fd_sc_hd__buf_2_0/a_27_47# 0.02fF
C32 clk ip 0.62fF
C33 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.01fF
C34 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.02fF
C35 sky130_fd_sc_hd__buf_2_0/A li_940_3458# 18.81fF
C36 VSS ip 2.78fF
C37 sky130_fd_sc_hd__buf_2_0/a_27_47# VDD 0.07fF
C38 sky130_fd_sc_hd__buf_2_1/A ip 1.73fF
C39 li_n2324_818# li_940_818# 2.99fF
C40 VDD li_940_3458# 2.18fF
C41 in li_940_818# 12.98fF
C42 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_0/X 0.03fF
C43 sky130_fd_sc_hd__buf_2_0/A ip 2.05fF
C44 li_n2324_818# clk 6.63fF
C45 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.01fF
C46 clk in 0.47fF
C47 li_n2324_818# VSS 3.07fF
C48 VDD ip 0.03fF
C49 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.24fF
C50 VSS in 1.52fF
C51 sky130_fd_sc_hd__buf_2_1/A li_n2324_818# 0.95fF
C52 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.00fF
C53 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.11fF
C54 sky130_fd_sc_hd__buf_2_1/A in 0.67fF
C55 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_0/X 0.01fF
C56 sky130_fd_sc_hd__nand2_4_1/a_27_47# outp 0.09fF
C57 sky130_fd_sc_hd__buf_2_1/a_27_47# VSS 0.04fF
C58 ip li_940_3458# 13.70fF
C59 sky130_fd_sc_hd__nand2_4_1/a_27_47# outn 0.06fF
C60 li_n2324_818# sky130_fd_sc_hd__buf_2_0/A 1.31fF
C61 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.00fF
C62 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.05fF
C63 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.03fF
C64 in sky130_fd_sc_hd__buf_2_0/A 1.07fF
C65 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.28fF
C66 sky130_fd_sc_hd__buf_2_1/a_27_47# outp 0.02fF
C67 sky130_fd_sc_hd__buf_2_1/a_27_47# outn 0.04fF
C68 li_n2324_818# VDD 0.09fF
C69 sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.02fF
C70 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.00fF
C71 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.02fF
C72 in VDD 0.01fF
C73 sky130_fd_sc_hd__nand2_4_0/a_27_47# outp 0.08fF
C74 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_0/a_27_47# 0.02fF
C75 sky130_fd_sc_hd__nand2_4_0/a_27_47# outn 0.18fF
C76 clk li_940_818# 4.02fF
C77 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.00fF
C78 sky130_fd_sc_hd__buf_2_1/a_27_47# VDD 0.09fF
C79 li_n2324_818# li_940_3458# 4.64fF
C80 in li_940_3458# 37.79fF
C81 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_0/X 0.11fF
C82 VSS li_940_818# 0.96fF
C83 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_0/a_27_47# 0.06fF
C84 sky130_fd_sc_hd__nand2_4_0/a_27_47# VDD 0.01fF
C85 sky130_fd_sc_hd__buf_2_1/A li_940_818# 21.09fF
C86 sky130_fd_sc_hd__buf_2_0/X VSS 0.04fF
C87 VSS clk 1.71fF
C88 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/X 0.04fF
C89 sky130_fd_sc_hd__buf_2_1/X VSS 0.05fF
C90 li_n2324_818# ip 48.05fF
C91 in ip 30.51fF
C92 li_940_818# sky130_fd_sc_hd__buf_2_0/A 9.11fF
C93 sky130_fd_sc_hd__buf_2_1/A clk 3.03fF
C94 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_1/A 0.09fF
C95 sky130_fd_sc_hd__buf_2_0/X outp 0.20fF
C96 sky130_fd_sc_hd__buf_2_0/X outn 0.03fF
C97 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_0/A 0.10fF
C98 sky130_fd_sc_hd__buf_2_1/A VSS 1.57fF
C99 sky130_fd_sc_hd__buf_2_1/X outp 0.03fF
C100 sky130_fd_sc_hd__buf_2_1/X outn 0.23fF
C101 li_940_3458# 0 -1568.83fF
C102 li_940_818# 0 -2217.21fF
C103 outn 0 21.70fF
C104 in 0 -297.33fF
C105 li_n2324_818# 0 -3691.32fF
C106 ip 0 -420.77fF
C107 VSS 0 -39.09fF
C108 sky130_fd_sc_hd__buf_2_0/A 0 -9.07fF
C109 sky130_fd_sc_hd__buf_2_1/A 0 -133.79fF
C110 VDD 0 -358.52fF
C111 clk 0 100.72fF
C112 sky130_fd_sc_hd__buf_2_1/a_27_47# 0 0.15fF
C113 sky130_fd_sc_hd__buf_2_0/a_27_47# 0 0.15fF
C114 outp 0 26.34fF
C115 sky130_fd_sc_hd__buf_2_0/X 0 43.25fF
C116 sky130_fd_sc_hd__nand2_4_1/a_27_47# 0 0.06fF
C117 sky130_fd_sc_hd__buf_2_1/X 0 23.78fF
C118 sky130_fd_sc_hd__nand2_4_0/a_27_47# 0 0.06fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CFEPS5 a_n275_n238# a_n129_n152# a_n173_n64#
X0 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=8.32e+11p pd=7.76e+06u as=0p ps=0u w=650000u l=150000u
X1 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 a_n129_n152# a_n173_n64# 0.38fF
C1 a_n173_n64# a_n275_n238# 0.40fF
C2 a_n129_n152# a_n275_n238# 0.60fF
.ends

.subckt analog_top_v2 ip in rst_n i_bias_1 i_bias_2 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1
+ debug op a_probe_0 a_probe_1 a_probe_2 a_probe_3 clk d_probe_0 d_probe_1 d_probe_2
+ d_probe_3 d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1
+ VDD VSS
Xesd_cell_5 i_bias_2 VDD VSS esd_cell_flat
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_2 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_18 sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_29 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_12_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_31 clock_v2_0/p2d VDD transmission_gate_31/nmos_tgate_0/w_n646_n262#
+ onebit_dac_1/out transmission_gate_31/out clock_v2_0/p2d_b VSS transmission_gate
Xtransmission_gate_20 clock_v2_0/p1d VDD transmission_gate_20/nmos_tgate_0/w_n646_n262#
+ a_mux2_en_0/in1 transmission_gate_21/in clock_v2_0/p1d_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_70 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_19 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_6 in VDD VSS esd_cell_flat
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_3 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__decap_12_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_32 clock_v2_0/p2d VDD transmission_gate_32/nmos_tgate_0/w_n646_n262#
+ onebit_dac_0/out transmission_gate_32/out clock_v2_0/p2d_b VSS transmission_gate
Xtransmission_gate_21 clock_v2_0/p2d VDD transmission_gate_21/nmos_tgate_0/w_n646_n262#
+ transmission_gate_21/in transmission_gate_21/out clock_v2_0/p2d_b VSS transmission_gate
Xtransmission_gate_10 clock_v2_0/p1d VDD transmission_gate_10/nmos_tgate_0/w_n646_n262#
+ ip transmission_gate_32/out clock_v2_0/p1d_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_60 sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_71 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_4 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xesd_cell_7 ip VDD VSS esd_cell_flat
Xsky130_fd_sc_hd__decap_12_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_22 ota_v2_0/p2 VDD transmission_gate_22/nmos_tgate_0/w_n646_n262#
+ transmission_gate_23/in ota_v2_0/ip ota_v2_0/p2_b VSS transmission_gate
Xtransmission_gate_11 clock_v2_0/p1d VDD transmission_gate_11/nmos_tgate_0/w_n646_n262#
+ in transmission_gate_31/out clock_v2_0/p1d_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_50 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_61 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_5 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_23 ota_v2_0/p1 VDD transmission_gate_23/nmos_tgate_0/w_n646_n262#
+ transmission_gate_23/in ota_v2_0/cm ota_v2_0/p1_b VSS transmission_gate
Xtransmission_gate_12 clock_v2_0/Bd VDD transmission_gate_12/nmos_tgate_0/w_n646_n262#
+ ota_w_test_v2_0/on a_mux2_en_0/in0 clock_v2_0/Bd_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_40 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_51 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_62 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_16_0 rst_n VSS VDD transmission_gate_7/en VSS VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__decap_12_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_6 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_24 ota_v2_0/p1 VDD transmission_gate_24/nmos_tgate_0/w_n646_n262#
+ transmission_gate_25/in ota_v2_0/cm ota_v2_0/p1_b VSS transmission_gate
Xtransmission_gate_13 clock_v2_0/Ad VDD transmission_gate_13/nmos_tgate_0/w_n646_n262#
+ ota_w_test_v2_0/on a_mux2_en_0/in1 clock_v2_0/Ad_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_30 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_41 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_52 transmission_gate_23/in transmission_gate_21/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_63 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_16_1 sky130_fd_sc_hd__clkinv_4_0/Y VSS VDD d_probe_1 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xota_v2_0 ota_v2_0/ip ota_v2_0/in ota_v2_0/op i_bias_2 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580#
+ ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_v2_0/sc_cmfb_0/transmission_gate_3/out
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_v2_0/sc_cmfb_0/transmission_gate_8/in
+ ota_v2_0/ota_v2_without_cmfb_0/li_11121_570# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480#
+ ota_v2_0/ota_v2_without_cmfb_0/li_8434_570# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580#
+ ota_v2_0/on ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# ota_v2_0/sc_cmfb_0/transmission_gate_6/in
+ ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580#
+ ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/sc_cmfb_0/bias_a VDD ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480#
+ ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# ota_v2_0/ota_v2_without_cmfb_0/bias_b
+ ota_v2_0/p1_b ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480#
+ ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/sc_cmfb_0/transmission_gate_9/in
+ ota_v2_0/sc_cmfb_0/cmc ota_v2_0/ota_v2_without_cmfb_0/m1_18877_3928# ota_v2_0/sc_cmfb_0/transmission_gate_4/out
+ ota_v2_0/cm ota_v2_0/p2_b ota_v2_0/p2 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399#
+ ota_v2_0/p1 ota_v2_0/ota_v2_without_cmfb_0/bias_d ota_v2_0/ota_v2_without_cmfb_0/m1_15613_3568#
+ VSS ota_v2
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_7 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_25 ota_v2_0/p2 VDD transmission_gate_25/nmos_tgate_0/w_n646_n262#
+ transmission_gate_25/in ota_v2_0/in ota_v2_0/p2_b VSS transmission_gate
Xtransmission_gate_14 clock_v2_0/Ad VDD transmission_gate_14/nmos_tgate_0/w_n646_n262#
+ ota_w_test_v2_0/op a_mux2_en_0/in0 clock_v2_0/Ad_b VSS transmission_gate
Xsky130_fd_sc_hd__clkinv_16_2 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD d_probe_2 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_20 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_31 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_42 transmission_gate_25/in transmission_gate_21/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_53 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_64 sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__mux4_1_0/X VSS VDD sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__clkinv_4_0/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_8 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_26 transmission_gate_7/en VDD transmission_gate_26/nmos_tgate_0/w_n646_n262#
+ ota_v2_0/cm ota_v2_0/in rst_n VSS transmission_gate
Xtransmission_gate_15 clock_v2_0/Bd VDD transmission_gate_15/nmos_tgate_0/w_n646_n262#
+ ota_w_test_v2_0/op a_mux2_en_0/in1 clock_v2_0/Bd_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_10 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_21 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_32 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_43 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_54 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_65 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_16_3 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD d_probe_3 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_9 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__mux4_1_1/X VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__clkinv_4_1/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_27 transmission_gate_7/en VDD transmission_gate_27/nmos_tgate_0/w_n646_n262#
+ ota_v2_0/cm ota_v2_0/ip rst_n VSS transmission_gate
Xtransmission_gate_16 transmission_gate_7/en VDD transmission_gate_16/nmos_tgate_0/w_n646_n262#
+ a_mux2_en_0/in1 a_mux2_en_0/in0 rst_n VSS transmission_gate
Xsky130_fd_sc_hd__clkinv_16_4 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD d_probe_0 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_11 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_22 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_33 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_44 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_55 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_66 sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__mux4_1_2/X VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__clkinv_4_2/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_28 transmission_gate_7/en VDD transmission_gate_28/nmos_tgate_0/w_n646_n262#
+ ota_v2_0/on ota_v2_0/op rst_n VSS transmission_gate
Xtransmission_gate_17 clock_v2_0/p2d VDD transmission_gate_17/nmos_tgate_0/w_n646_n262#
+ onebit_dac_0/out transmission_gate_30/out clock_v2_0/p2d_b VSS transmission_gate
Xonebit_dac_0 op VDD VDD onebit_dac_1/v_b VSS onebit_dac_0/out VSS onebit_dac
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_12 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_23 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_34 transmission_gate_25/in transmission_gate_30/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_45 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_56 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_67 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__mux4_1_3/X VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__clkinv_4_3/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_29 clock_v2_0/p1d VDD transmission_gate_29/nmos_tgate_0/w_n646_n262#
+ in transmission_gate_29/out clock_v2_0/p1d_b VSS transmission_gate
Xtransmission_gate_18 clock_v2_0/p2d VDD transmission_gate_18/nmos_tgate_0/w_n646_n262#
+ onebit_dac_1/out transmission_gate_29/out clock_v2_0/p2d_b VSS transmission_gate
Xa_mux2_en_0 debug a_mux2_en_0/in0 a_mux2_en_0/in1 a_probe_0 a_mux2_en_0/transmission_gate_1/en_b
+ a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in a_mux2_en_0/switch_5t_mux2_1/en
+ VDD a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in a_mux2_en_0/switch_5t_mux2_1/in
+ VSS a_mod_grp_ctrl_0 a_mux2_en_0/switch_5t_mux2_0/in a_mux2_en
Xonebit_dac_1 op VDD VSS onebit_dac_1/v_b VDD onebit_dac_1/out VSS onebit_dac
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_13 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_24 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_35 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_46 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_57 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_68 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_1 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xota_w_test_v2_0 ota_w_test_v2_0/ip ota_w_test_v2_0/in ota_w_test_v2_0/op ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651#
+ ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8434_570#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# a_mux4_en_0/in1 ota_w_test_v2_0/on
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# a_mux4_en_1/in0 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in
+ VDD ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# a_mux4_en_0/in2
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# ota_v2_0/p1_b ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# i_bias_1 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in
+ ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_18877_3928# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out
+ VSS a_mux4_en_0/in0 ota_v2_0/p2_b ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570#
+ ota_v2_0/p2 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# a_mux4_en_1/in1
+ ota_v2_0/p1 a_mux4_en_1/in2 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_15613_3568#
+ ota_w_test_v2
Xtransmission_gate_19 clock_v2_0/p1d VDD transmission_gate_19/nmos_tgate_0/w_n646_n262#
+ a_mux2_en_0/in0 transmission_gate_21/out clock_v2_0/p1d_b VSS transmission_gate
Xa_mux2_en_1 debug ota_v2_0/op ota_v2_0/on a_probe_1 a_mux2_en_1/transmission_gate_1/en_b
+ a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in a_mux2_en_1/switch_5t_mux2_1/en
+ VDD a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in a_mux2_en_1/switch_5t_mux2_1/in
+ VSS a_mod_grp_ctrl_0 a_mux2_en_1/switch_5t_mux2_0/in a_mux2_en
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_14 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_25 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_36 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_47 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_58 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_69 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__mux4_1_0 ota_v2_0/p2 clock_v2_0/B ota_v2_0/p2_b clock_v2_0/B_b d_clk_grp_1_ctrl_0
+ d_clk_grp_1_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_27_413#
+ sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__mux4_1_0/a_834_97#
+ sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_193_413#
+ sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__pfet_01v8_hvt_XAYTAL_0 onebit_dac_1/v_b VDD VDD VSS sky130_fd_pr__pfet_01v8_hvt_XAYTAL
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_2 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_15 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_26 transmission_gate_25/in transmission_gate_21/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_37 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_48 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_59 sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_3 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__mux4_1_1 clock_v2_0/p1d clock_v2_0/Ad clock_v2_0/p1d_b clock_v2_0/Ad_b
+ d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__mux4_1_1/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_1/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_27_413#
+ sky130_fd_sc_hd__mux4_1_1/a_923_363# sky130_fd_sc_hd__mux4_1_1/a_193_47# sky130_fd_sc_hd__mux4_1_1/a_834_97#
+ sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_193_413#
+ sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_16 sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_27 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_38 transmission_gate_23/in transmission_gate_29/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_49 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__mux4_1_2 clock_v2_0/p2d clock_v2_0/Bd clock_v2_0/p2d_b clock_v2_0/Bd_b
+ d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_27_413#
+ sky130_fd_sc_hd__mux4_1_2/a_923_363# sky130_fd_sc_hd__mux4_1_2/a_193_47# sky130_fd_sc_hd__mux4_1_2/a_834_97#
+ sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_193_413#
+ sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_4 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_0 clock_v2_0/A VDD transmission_gate_0/nmos_tgate_0/w_n646_n262#
+ transmission_gate_2/in ota_w_test_v2_0/in clock_v2_0/A_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_17 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_28 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_39 ota_v2_0/on ota_v2_0/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_5 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__mux4_1_3 ota_v2_0/p1 clock_v2_0/A ota_v2_0/p1_b clock_v2_0/A_b d_clk_grp_1_ctrl_0
+ d_clk_grp_1_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_27_413#
+ sky130_fd_sc_hd__mux4_1_3/a_923_363# sky130_fd_sc_hd__mux4_1_3/a_193_47# sky130_fd_sc_hd__mux4_1_3/a_834_97#
+ sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_193_413#
+ sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_18 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_29 transmission_gate_23/in transmission_gate_21/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_1 clock_v2_0/B VDD transmission_gate_1/nmos_tgate_0/w_n646_n262#
+ transmission_gate_3/in ota_w_test_v2_0/in clock_v2_0/B_b VSS transmission_gate
Xclock_v2_0 clk clock_v2_0/p2d_b clock_v2_0/p2d ota_v2_0/p2_b ota_v2_0/p2 clock_v2_0/p1d_b
+ clock_v2_0/p1d ota_v2_0/p1_b ota_v2_0/p1 clock_v2_0/Ad_b clock_v2_0/Ad clock_v2_0/A_b
+ clock_v2_0/A clock_v2_0/Bd_b clock_v2_0/Bd clock_v2_0/B_b clock_v2_0/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/A
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_439_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_218_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_218_374#
+ clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B
+ clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
+ clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_592_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_535_374# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A clock_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A
+ VSS VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y
+ clock_v2
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_6 sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_2 clock_v2_0/B VDD transmission_gate_2/nmos_tgate_0/w_n646_n262#
+ transmission_gate_2/in ota_w_test_v2_0/ip clock_v2_0/B_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_19 ota_v2_0/op ota_v2_0/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_7 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_3 clock_v2_0/A VDD transmission_gate_3/nmos_tgate_0/w_n646_n262#
+ transmission_gate_3/in ota_w_test_v2_0/ip clock_v2_0/A_b VSS transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_8 transmission_gate_8/in transmission_gate_32/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_9 transmission_gate_8/in transmission_gate_32/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_4 ota_v2_0/p2 VDD transmission_gate_4/nmos_tgate_0/w_n646_n262#
+ transmission_gate_8/in transmission_gate_2/in ota_v2_0/p2_b VSS transmission_gate
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_5 ota_v2_0/p2 VDD transmission_gate_5/nmos_tgate_0/w_n646_n262#
+ transmission_gate_9/in transmission_gate_3/in ota_v2_0/p2_b VSS transmission_gate
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_6 transmission_gate_7/en VDD transmission_gate_6/nmos_tgate_0/w_n646_n262#
+ a_mux4_en_0/in0 transmission_gate_2/in rst_n VSS transmission_gate
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_7 transmission_gate_7/en VDD transmission_gate_7/nmos_tgate_0/w_n646_n262#
+ a_mux4_en_0/in0 transmission_gate_3/in rst_n VSS transmission_gate
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_8 ota_v2_0/p1 VDD transmission_gate_8/nmos_tgate_0/w_n646_n262#
+ transmission_gate_8/in a_mux4_en_0/in0 ota_v2_0/p1_b VSS transmission_gate
Xsky130_fd_sc_hd__decap_12_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xtransmission_gate_9 ota_v2_0/p1 VDD transmission_gate_9/nmos_tgate_0/w_n646_n262#
+ transmission_gate_9/in a_mux4_en_0/in0 ota_v2_0/p1_b VSS transmission_gate
Xsky130_fd_sc_hd__decap_12_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xa_mux4_en_0 debug a_mux4_en_0/in0 a_mux4_en_0/in1 a_mux4_en_0/in2 a_mux4_en_0/in3
+ a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y a_mux4_en_0/switch_5t_mux4_1/en a_mux4_en_0/sky130_fd_sc_hd__nand2_1_2/a_113_47#
+ a_mux4_en_0/switch_5t_mux4_1/in a_mux4_en_0/switch_5t_mux4_1/en_b a_mux4_en_0/switch_5t_mux4_0/a_300_216#
+ a_mux4_en_0/switch_5t_mux4_3/en a_mux4_en_0/switch_5t_mux4_0/en a_mux4_en_0/sky130_fd_sc_hd__nand2_1_3/a_113_47#
+ a_mux4_en_0/switch_5t_mux4_1/a_300_216# a_mux4_en_0/switch_5t_mux4_2/a_300_216#
+ a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y a_mux4_en_0/switch_5t_mux4_3/a_300_216# a_mux4_en_0/transmission_gate_3/en_b
+ a_mux4_en_0/sky130_fd_sc_hd__nand2_1_0/a_113_47# a_mux4_en_0/switch_5t_mux4_2/en_b
+ a_mux4_en_0/switch_5t_mux4_3/in a_mux4_en_0/switch_5t_mux4_2/en a_probe_2 a_mux4_en_0/switch_5t_mux4_0/en_b
+ a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_0/in VDD a_mod_grp_ctrl_1 a_mux4_en_0/switch_5t_mux4_2/in
+ a_mux4_en_0/switch_5t_mux4_3/en_b VSS a_mux4_en_0/sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ a_mux4_en
Xa_mux4_en_1 debug a_mux4_en_1/in0 a_mux4_en_1/in1 a_mux4_en_1/in2 a_mux4_en_1/in3
+ a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y a_mux4_en_1/switch_5t_mux4_1/en a_mux4_en_1/sky130_fd_sc_hd__nand2_1_2/a_113_47#
+ a_mux4_en_1/switch_5t_mux4_1/in a_mux4_en_1/switch_5t_mux4_1/en_b a_mux4_en_1/switch_5t_mux4_0/a_300_216#
+ a_mux4_en_1/switch_5t_mux4_3/en a_mux4_en_1/switch_5t_mux4_0/en a_mux4_en_1/sky130_fd_sc_hd__nand2_1_3/a_113_47#
+ a_mux4_en_1/switch_5t_mux4_1/a_300_216# a_mux4_en_1/switch_5t_mux4_2/a_300_216#
+ a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y a_mux4_en_1/switch_5t_mux4_3/a_300_216# a_mux4_en_1/transmission_gate_3/en_b
+ a_mux4_en_1/sky130_fd_sc_hd__nand2_1_0/a_113_47# a_mux4_en_1/switch_5t_mux4_2/en_b
+ a_mux4_en_1/switch_5t_mux4_3/in a_mux4_en_1/switch_5t_mux4_2/en a_probe_3 a_mux4_en_1/switch_5t_mux4_0/en_b
+ a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_0/in VDD a_mod_grp_ctrl_1 a_mux4_en_1/switch_5t_mux4_2/in
+ a_mux4_en_1/switch_5t_mux4_3/en_b VSS a_mux4_en_1/sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ a_mux4_en
Xsky130_fd_sc_hd__decap_12_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_40 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_30 sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_41 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_20 sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_31 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_42 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_10 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_21 sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_32 transmission_gate_9/in transmission_gate_31/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_43 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_11 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_22 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_33 transmission_gate_9/in transmission_gate_31/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_44 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_12 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_23 sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_34 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_TABSMU_0 ota_v2_0/on VSS VSS sky130_fd_pr__cap_mim_m3_1_TABSMU
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_45 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xcomparator_v2_0 ota_v2_0/p1_b op VSS comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47#
+ onebit_dac_1/v_b comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X
+ VDD comparator_v2_0/li_n2324_818# comparator_v2_0/li_940_3458# comparator_v2_0/li_940_818#
+ ota_v2_0/op comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ ota_v2_0/on comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A comparator_v2
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_13 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_24 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_35 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_46 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_0 a_probe_2 VDD VSS esd_cell_flat
Xsky130_fd_pr__cap_mim_m3_1_TABSMU_1 ota_v2_0/op VSS VSS sky130_fd_pr__cap_mim_m3_1_TABSMU
Xesd_cell_1 a_probe_3 VDD VSS esd_cell_flat
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_14 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_25 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_36 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_47 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_15 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_26 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_37 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__nfet_01v8_CFEPS5_0 VSS onebit_dac_1/v_b VSS sky130_fd_pr__nfet_01v8_CFEPS5
Xesd_cell_2 a_probe_0 VDD VSS esd_cell_flat
Xesd_cell_3 a_probe_1 VDD VSS esd_cell_flat
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_0 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_16 transmission_gate_2/in a_mux2_en_0/in0 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_27 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_38 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_17 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_28 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_39 transmission_gate_3/in a_mux2_en_0/in1 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_4 i_bias_1 VDD VSS esd_cell_flat
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_30 clock_v2_0/p1d VDD transmission_gate_30/nmos_tgate_0/w_n646_n262#
+ ip transmission_gate_30/out clock_v2_0/p1d_b VSS transmission_gate
C0 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p1 -0.00fF
C1 onebit_dac_1/out a_mux4_en_1/in0 0.18fF
C2 clock_v2_0/p2d_b clock_v2_0/A 0.79fF
C3 clock_v2_0/p1d_b clock_v2_0/Bd_b 1.03fF
C4 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.03fF
C5 ota_v2_0/ip transmission_gate_7/en 0.18fF
C6 comparator_v2_0/li_940_818# ota_v2_0/p1_b 1.53fF
C7 a_mux4_en_1/in2 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# -0.00fF
C8 ota_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.00fF
C9 a_mux4_en_1/switch_5t_mux4_3/en a_mux4_en_1/switch_5t_mux4_3/in 0.00fF
C10 sky130_fd_sc_hd__mux4_1_1/a_668_97# clock_v2_0/Ad_b 0.00fF
C11 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_w_test_v2_0/ip -0.00fF
C12 debug a_mux4_en_0/switch_5t_mux4_3/en 0.11fF
C13 clock_v2_0/p2d clock_v2_0/Bd_b 1.17fF
C14 a_mod_grp_ctrl_0 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C15 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C16 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.00fF
C17 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.07fF
C18 ota_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/p1_b 0.00fF
C19 transmission_gate_31/out ip 0.03fF
C20 a_mux4_en_1/in2 a_mux4_en_1/switch_5t_mux4_3/in 0.00fF
C21 ota_v2_0/p1 clock_v2_0/A 1.80fF
C22 ota_w_test_v2_0/on ota_v2_0/p2_b -0.01fF
C23 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.00fF
C24 sky130_fd_sc_hd__mux4_1_3/a_757_363# clock_v2_0/B_b 0.00fF
C25 a_mux2_en_0/in0 ota_v2_0/p1_b 0.05fF
C26 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.00fF
C27 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/Bd_b 0.07fF
C28 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210# ota_v2_0/on 0.03fF
C29 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# -0.04fF
C30 ota_v2_0/op VDD 24.55fF
C31 clock_v2_0/Ad clock_v2_0/Bd_b 1.54fF
C32 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# 0.02fF
C33 ota_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/p2_b 0.00fF
C34 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C35 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.01fF
C36 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p2 0.01fF
C37 clock_v2_0/p1d_b VDD 9.58fF
C38 a_mux4_en_0/in0 transmission_gate_7/en 1.73fF
C39 a_mux4_en_1/in0 ota_v2_0/p1_b 0.00fF
C40 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.01fF
C41 sky130_fd_sc_hd__mux4_1_1/a_193_47# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.01fF
C42 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/op 1.31fF
C43 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# 0.09fF
C44 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# VDD 1.90fF
C45 clock_v2_0/p2d VDD 8.73fF
C46 clock_v2_0/B clock_v2_0/p1d 1.00fF
C47 clock_v2_0/Bd clock_v2_0/p1d 0.82fF
C48 sky130_fd_sc_hd__mux4_1_0/X VDD 1.01fF
C49 sky130_fd_sc_hd__mux4_1_2/a_247_21# clock_v2_0/Bd_b 0.12fF
C50 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.00fF
C51 sky130_fd_sc_hd__mux4_1_3/a_834_97# clock_v2_0/B_b 0.00fF
C52 sky130_fd_sc_hd__clkinv_4_3/Y VDD 0.63fF
C53 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# ota_v2_0/ip 0.11fF
C54 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/m3_n1030_n980# transmission_gate_2/in 0.17fF
C55 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VDD 0.03fF
C56 sky130_fd_sc_hd__mux4_1_0/a_27_47# clock_v2_0/A 0.00fF
C57 d_clk_grp_2_ctrl_1 clock_v2_0/Bd 0.01fF
C58 a_mux4_en_0/in2 ota_w_test_v2_0/ip 0.26fF
C59 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/c1_n260_n210# 0.03fF
C60 transmission_gate_8/in transmission_gate_2/in 2.48fF
C61 sky130_fd_sc_hd__mux4_1_2/a_1478_413# clock_v2_0/Bd_b 0.00fF
C62 a_mux4_en_1/in1 a_mux4_en_1/switch_5t_mux4_0/in -0.00fF
C63 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.02fF
C64 sky130_fd_sc_hd__mux4_1_2/a_277_47# VDD 0.12fF
C65 ota_w_test_v2_0/on ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out -0.01fF
C66 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in 0.00fF
C67 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.00fF
C68 VDD clock_v2_0/Ad 2.18fF
C69 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/m3_n1030_n980# 0.12fF
C70 debug a_mux4_en_1/switch_5t_mux4_2/a_300_216# 0.13fF
C71 d_probe_3 d_clk_grp_2_ctrl_1 1.14fF
C72 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/p1d 0.00fF
C73 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980# 0.09fF
C74 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.00fF
C75 transmission_gate_30/out ota_v2_0/op 0.01fF
C76 d_clk_grp_2_ctrl_0 clock_v2_0/p1d 0.00fF
C77 sky130_fd_sc_hd__mux4_1_2/a_247_21# VDD 0.07fF
C78 ota_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/p2_b 0.01fF
C79 onebit_dac_0/out clock_v2_0/p2d_b 0.99fF
C80 onebit_dac_1/out VDD 1.16fF
C81 rst_n clock_v2_0/p2d_b 0.57fF
C82 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.08fF
C83 transmission_gate_30/out clock_v2_0/p1d_b 0.33fF
C84 ota_v2_0/p1_b clock_v2_0/Bd_b 1.44fF
C85 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 2.73fF
C86 sky130_fd_sc_hd__mux4_1_1/a_277_47# ota_v2_0/p2_b 0.00fF
C87 sky130_fd_sc_hd__mux4_1_2/a_1478_413# VDD 0.14fF
C88 transmission_gate_2/in clock_v2_0/A 0.49fF
C89 transmission_gate_30/out clock_v2_0/p2d 0.14fF
C90 a_mod_grp_ctrl_0 a_mux2_en_1/switch_5t_mux2_1/in -0.00fF
C91 a_mux2_en_0/in0 ota_v2_0/p2_b 0.05fF
C92 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/c1_n930_n880# 0.07fF
C93 rst_n ota_v2_0/p1 0.76fF
C94 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in -0.00fF
C95 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.00fF
C96 transmission_gate_29/out onebit_dac_0/out 0.03fF
C97 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y -0.00fF
C98 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y VDD 0.14fF
C99 a_mux4_en_0/in0 transmission_gate_3/in 0.36fF
C100 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/c1_n260_n210# -0.07fF
C101 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C102 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.12fF
C103 a_mux4_en_1/in0 ota_v2_0/p2_b 0.00fF
C104 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# ota_v2_0/ip 0.03fF
C105 a_mux4_en_1/switch_5t_mux4_1/in a_mux4_en_1/switch_5t_mux4_0/in -0.00fF
C106 a_mux2_en_0/switch_5t_mux2_1/en VDD 0.24fF
C107 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C108 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C109 i_bias_2 ota_v2_0/sc_cmfb_0/bias_a 0.01fF
C110 VDD ota_v2_0/p1_b 17.95fF
C111 ota_w_test_v2_0/on ota_w_test_v2_0/ip 0.42fF
C112 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# -0.00fF
C113 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C114 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C115 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y -0.00fF
C116 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.35fF
C117 onebit_dac_1/out transmission_gate_30/out 0.03fF
C118 a_mux2_en_1/switch_5t_mux2_1/en VDD 0.24fF
C119 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X -0.00fF
C120 sky130_fd_sc_hd__mux4_1_0/a_247_21# ota_v2_0/p2_b 0.08fF
C121 ota_v2_0/p2 transmission_gate_9/in 0.59fF
C122 a_mux4_en_1/switch_5t_mux4_1/in a_mux4_en_1/switch_5t_mux4_1/en -0.00fF
C123 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_1/en_b 0.14fF
C124 clock_v2_0/Bd clock_v2_0/A 0.47fF
C125 clock_v2_0/B clock_v2_0/A 0.92fF
C126 onebit_dac_1/v_b op 2.11fF
C127 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A -0.00fF
C128 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.03fF
C129 sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/m3_n1030_n980# 0.09fF
C130 a_mux2_en_0/switch_5t_mux2_1/in a_mux2_en_0/in0 0.05fF
C131 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/Bd_b 0.00fF
C132 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# ota_v2_0/op 0.31fF
C133 ota_v2_0/p2 ota_w_test_v2_0/op 0.00fF
C134 ota_v2_0/cm ota_v2_0/p2 0.10fF
C135 transmission_gate_7/en clock_v2_0/Ad_b 0.33fF
C136 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# -0.09fF
C137 comparator_v2_0/li_n2324_818# ota_v2_0/op 0.01fF
C138 ota_v2_0/p2_b clock_v2_0/Bd_b 0.91fF
C139 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C140 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X -0.01fF
C141 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# -0.00fF
C142 a_mux4_en_0/switch_5t_mux4_0/in a_mux4_en_0/switch_5t_mux4_0/en_b -0.00fF
C143 a_mux4_en_0/switch_5t_mux4_3/en a_mux4_en_0/switch_5t_mux4_3/a_300_216# -0.00fF
C144 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A -0.00fF
C145 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# 0.03fF
C146 ota_v2_0/in ota_v2_0/ip 2.02fF
C147 a_mux4_en_0/switch_5t_mux4_1/en VDD 0.12fF
C148 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_193_47# -0.00fF
C149 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# transmission_gate_3/in 1.64fF
C150 clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y VDD 0.13fF
C151 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.13fF
C152 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.09fF
C153 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# -0.01fF
C154 clock_v2_0/p1d_b clock_v2_0/p1d 27.04fF
C155 sky130_fd_sc_hd__mux4_1_0/a_668_97# VDD 0.01fF
C156 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.00fF
C157 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# ota_v2_0/ip 0.03fF
C158 sky130_fd_sc_hd__mux4_1_3/a_27_413# ota_v2_0/p1 -0.00fF
C159 rst_n transmission_gate_2/in 0.12fF
C160 a_mux2_en_0/in1 a_mux2_en_0/switch_5t_mux2_0/in 0.04fF
C161 debug ota_v2_0/op -0.00fF
C162 clock_v2_0/p1d_b d_clk_grp_2_ctrl_1 0.13fF
C163 sky130_fd_sc_hd__mux4_1_1/a_834_97# VDD 0.01fF
C164 clock_v2_0/p2d clock_v2_0/p1d 1.04fF
C165 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# 0.03fF
C166 a_mux4_en_0/in2 a_mux4_en_0/in3 0.00fF
C167 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C168 transmission_gate_31/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# -0.27fF
C169 sky130_fd_sc_hd__mux4_1_3/a_277_47# clock_v2_0/A 0.00fF
C170 clock_v2_0/p2d d_clk_grp_2_ctrl_1 0.02fF
C171 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.09fF
C172 a_mux4_en_0/switch_5t_mux4_2/in VDD 0.60fF
C173 a_mux2_en_0/switch_5t_mux2_1/en a_mod_grp_ctrl_1 3.61fF
C174 transmission_gate_23/in ota_v2_0/p2 0.57fF
C175 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.09fF
C176 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# 0.09fF
C177 ota_v2_0/p2_b VDD 16.24fF
C178 transmission_gate_25/in VDD 0.77fF
C179 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C180 a_mux4_en_1/in1 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C181 a_mux2_en_1/switch_5t_mux2_0/in ota_v2_0/on 0.04fF
C182 clock_v2_0/Ad clock_v2_0/p1d 1.95fF
C183 sky130_fd_sc_hd__mux4_1_2/a_277_47# d_clk_grp_2_ctrl_1 0.15fF
C184 sky130_fd_sc_hd__clkinv_4_1/Y d_probe_3 0.06fF
C185 a_mux2_en_1/switch_5t_mux2_1/en a_mod_grp_ctrl_1 0.32fF
C186 a_mux2_en_0/in0 ota_w_test_v2_0/ip 0.56fF
C187 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C188 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_v2_0/sc_cmfb_0/cmc -0.00fF
C189 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__clkinv_4_0/Y 0.00fF
C190 d_clk_grp_2_ctrl_1 clock_v2_0/Ad 0.01fF
C191 ota_v2_0/in ota_v2_0/ota_v2_without_cmfb_0/m1_18877_3928# 0.00fF
C192 ota_v2_0/ota_v2_without_cmfb_0/bias_d VDD 2.73fF
C193 a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in VDD 0.59fF
C194 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C195 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C196 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/p2 0.00fF
C197 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# -0.01fF
C198 a_mux4_en_1/switch_5t_mux4_3/en_b a_mux4_en_1/switch_5t_mux4_2/en -0.00fF
C199 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VDD -0.00fF
C200 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.00fF
C201 a_mux4_en_0/switch_5t_mux4_0/en a_mod_grp_ctrl_0 0.29fF
C202 rst_n clock_v2_0/B 0.33fF
C203 rst_n clock_v2_0/Bd 0.28fF
C204 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# -0.12fF
C205 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C206 d_clk_grp_1_ctrl_0 VDD 6.43fF
C207 sky130_fd_sc_hd__mux4_1_2/a_247_21# d_clk_grp_2_ctrl_1 0.01fF
C208 a_mux4_en_1/switch_5t_mux4_2/en a_mux4_en_1/switch_5t_mux4_2/en_b -0.00fF
C209 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# ota_v2_0/ip 0.12fF
C210 VDD comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A 3.93fF
C211 ota_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/p1 0.07fF
C212 a_mux4_en_0/switch_5t_mux4_1/en a_mod_grp_ctrl_1 0.08fF
C213 a_mux2_en_0/switch_5t_mux2_1/in VDD 0.44fF
C214 sky130_fd_sc_hd__mux4_1_2/a_1478_413# d_clk_grp_2_ctrl_1 0.00fF
C215 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.13fF
C216 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out VDD 2.54fF
C217 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.00fF
C218 sky130_fd_sc_hd__mux4_1_0/a_277_47# clock_v2_0/B_b 0.06fF
C219 sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.02fF
C220 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# 0.09fF
C221 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C222 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.01fF
C223 transmission_gate_30/out transmission_gate_25/in 0.24fF
C224 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# 0.14fF
C225 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.03fF
C226 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.00fF
C227 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# ota_v2_0/op 0.03fF
C228 comparator_v2_0/li_n2324_818# ota_v2_0/p1_b 0.87fF
C229 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VDD 0.09fF
C230 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.06fF
C231 a_mux4_en_1/in1 a_mux4_en_0/in0 0.62fF
C232 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C233 sky130_fd_sc_hd__mux4_1_2/X clock_v2_0/p2d_b 0.00fF
C234 sky130_fd_sc_hd__mux4_1_0/a_923_363# VDD 0.01fF
C235 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/Bd 0.00fF
C236 sky130_fd_sc_hd__clkinv_4_2/Y VDD 1.22fF
C237 a_mux2_en_0/in1 ota_w_test_v2_0/op 0.93fF
C238 a_mux4_en_1/in2 in 1.21fF
C239 ota_v2_0/p1_b clock_v2_0/p1d 18.64fF
C240 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# clock_v2_0/p1d_b 0.02fF
C241 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# 0.12fF
C242 a_mux4_en_0/switch_5t_mux4_2/in a_mod_grp_ctrl_1 -0.00fF
C243 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C244 a_mux4_en_0/switch_5t_mux4_0/en_b a_mux4_en_0/switch_5t_mux4_1/en_b 0.00fF
C245 clock_v2_0/p1d_b clock_v2_0/A 0.85fF
C246 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C247 sky130_fd_sc_hd__mux4_1_1/a_668_97# clock_v2_0/Bd_b 0.00fF
C248 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D clk 0.00fF
C249 a_mod_grp_ctrl_0 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y 0.01fF
C250 debug a_mux2_en_0/switch_5t_mux2_1/en 5.25fF
C251 clock_v2_0/p2d clock_v2_0/A 0.76fF
C252 a_mux2_en_0/in1 in 0.30fF
C253 i_bias_1 ip 0.17fF
C254 sky130_fd_sc_hd__mux4_1_0/a_834_97# ota_v2_0/p1_b 0.00fF
C255 d_probe_0 sky130_fd_sc_hd__clkinv_4_0/Y 0.08fF
C256 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.02fF
C257 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C258 VDD a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.14fF
C259 a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in a_mod_grp_ctrl_1 0.14fF
C260 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C261 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.01fF
C262 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/p2d_b 0.04fF
C263 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y -0.00fF
C264 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y VDD 1.63fF
C265 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/c1_n260_n210# ota_v2_0/op 0.06fF
C266 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# 0.09fF
C267 a_mux2_en_1/switch_5t_mux2_1/en debug 0.42fF
C268 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.00fF
C269 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_w_test_v2_0/in 0.06fF
C270 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C271 sky130_fd_sc_hd__mux4_1_0/a_1290_413# clock_v2_0/B 0.00fF
C272 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.00fF
C273 clock_v2_0/Ad clock_v2_0/A 8.16fF
C274 sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980# transmission_gate_3/in 0.17fF
C275 transmission_gate_31/out transmission_gate_32/out 0.62fF
C276 a_mux2_en_0/in0 a_mux2_en_0/transmission_gate_1/en_b 0.00fF
C277 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_2/en 0.13fF
C278 sky130_fd_sc_hd__mux4_1_3/a_27_413# clock_v2_0/B 0.00fF
C279 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# a_mux4_en_0/in2 0.07fF
C280 VDD clk 5.10fF
C281 sky130_fd_sc_hd__mux4_1_1/a_668_97# VDD 0.01fF
C282 ota_w_test_v2_0/ip VDD 2.20fF
C283 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out VDD 1.89fF
C284 sky130_fd_sc_hd__mux4_1_3/a_750_97# VDD 0.07fF
C285 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47# clock_v2_0/Bd_b -0.00fF
C286 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/c1_n930_n880# -0.01fF
C287 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# 0.09fF
C288 ota_v2_0/cm ota_v2_0/on 0.31fF
C289 a_mux4_en_0/in0 ip 0.25fF
C290 transmission_gate_8/in ota_v2_0/p1_b 0.43fF
C291 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# -0.12fF
C292 transmission_gate_32/out ip 0.06fF
C293 debug a_mux4_en_0/switch_5t_mux4_1/en 0.12fF
C294 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VDD 0.00fF
C295 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B -0.00fF
C296 ota_v2_0/in transmission_gate_21/in 0.43fF
C297 i_bias_2 a_mod_grp_ctrl_0 0.17fF
C298 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C299 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# -0.06fF
C300 sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C301 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# ota_v2_0/in 0.23fF
C302 ota_v2_0/p2_b clock_v2_0/p1d 2.90fF
C303 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p1_b -0.00fF
C304 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C305 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C306 clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y VDD -0.00fF
C307 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_247_21# -0.00fF
C308 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C309 onebit_dac_0/out ota_v2_0/op 0.16fF
C310 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C311 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C312 a_mux4_en_0/in2 ota_w_test_v2_0/in 0.24fF
C313 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/c1_n930_n880# 0.07fF
C314 rst_n ota_v2_0/op 0.16fF
C315 debug a_mux4_en_0/switch_5t_mux4_2/in 0.67fF
C316 ota_v2_0/p2_b sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.01fF
C317 transmission_gate_23/in ota_v2_0/on 0.27fF
C318 clock_v2_0/p1d_b rst_n 0.61fF
C319 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C320 clock_v2_0/A ota_v2_0/p1_b 1.55fF
C321 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C322 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in ota_w_test_v2_0/op 0.00fF
C323 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y a_mod_grp_ctrl_1 0.00fF
C324 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C325 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# 0.07fF
C326 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/c1_n930_n880# -0.01fF
C327 a_mux2_en_0/in0 transmission_gate_7/en 0.13fF
C328 clock_v2_0/p2d onebit_dac_0/out 1.23fF
C329 clock_v2_0/p2d rst_n 0.57fF
C330 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VDD 0.80fF
C331 a_mod_grp_ctrl_0 a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in -0.00fF
C332 a_mux4_en_1/in2 a_mux4_en_1/transmission_gate_3/en_b 0.03fF
C333 debug a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in 0.14fF
C334 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C335 sky130_fd_sc_hd__mux4_1_2/a_668_97# clock_v2_0/Ad_b 0.00fF
C336 clock_v2_0/p2d_b sky130_fd_sc_hd__mux4_1_2/a_1290_413# -0.00fF
C337 a_mux2_en_1/switch_5t_mux2_1/in VDD 0.44fF
C338 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C339 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# VDD 0.31fF
C340 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.00fF
C341 sky130_fd_sc_hd__mux4_1_3/a_668_97# clock_v2_0/B_b 0.00fF
C342 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/on 0.00fF
C343 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# -0.12fF
C344 a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in a_mod_grp_ctrl_0 0.01fF
C345 rst_n clock_v2_0/Ad 0.28fF
C346 transmission_gate_8/in ota_v2_0/p2_b 0.44fF
C347 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/c1_n260_n210# 0.03fF
C348 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980# -0.05fF
C349 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# -0.01fF
C350 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/c1_n930_n880# 0.07fF
C351 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C352 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.04fF
C353 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C354 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# 0.00fF
C355 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VDD 0.57fF
C356 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# -0.00fF
C357 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# -0.01fF
C358 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# transmission_gate_21/in 0.03fF
C359 debug a_mux2_en_0/switch_5t_mux2_1/in -0.00fF
C360 a_mux4_en_1/switch_5t_mux4_3/en a_mux4_en_1/switch_5t_mux4_2/en 0.00fF
C361 clock_v2_0/A_b clock_v2_0/p2d_b 0.70fF
C362 clock_v2_0/p2d_b clock_v2_0/B_b 0.78fF
C363 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A -0.00fF
C364 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.00fF
C365 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A ota_v2_0/p1_b -0.00fF
C366 onebit_dac_1/out onebit_dac_0/out 6.34fF
C367 a_mux2_en_0/transmission_gate_1/en_b VDD 0.21fF
C368 sky130_fd_sc_hd__mux4_1_0/a_750_97# clock_v2_0/Ad_b 0.00fF
C369 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.03fF
C370 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.09fF
C371 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210# 0.03fF
C372 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p2_b 0.01fF
C373 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.00fF
C374 sky130_fd_sc_hd__mux4_1_3/a_193_413# VDD 0.02fF
C375 a_mux4_en_1/switch_5t_mux4_1/en_b VDD 0.94fF
C376 ota_v2_0/p1 clock_v2_0/B_b 0.96fF
C377 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VDD 0.08fF
C378 clock_v2_0/A_b ota_v2_0/p1 1.01fF
C379 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.00fF
C380 a_mux4_en_0/in2 a_mux4_en_1/in1 0.43fF
C381 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# -0.00fF
C382 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y 0.13fF
C383 clock_v2_0/p2d_b ota_v2_0/p2 5.67fF
C384 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/Ad 0.01fF
C385 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/switch_5t_mux4_2/en_b -0.00fF
C386 transmission_gate_7/en clock_v2_0/Bd_b 0.29fF
C387 ota_v2_0/p2_b clock_v2_0/A 1.12fF
C388 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/Bd 0.01fF
C389 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# 0.13fF
C390 a_mux2_en_0/in0 transmission_gate_3/in 0.35fF
C391 a_mux4_en_0/switch_5t_mux4_0/en_b a_mux4_en_0/switch_5t_mux4_0/a_300_216# -0.00fF
C392 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.01fF
C393 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VDD 0.11fF
C394 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/X 0.02fF
C395 sky130_fd_sc_hd__mux4_1_0/a_757_363# clock_v2_0/B_b 0.01fF
C396 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C397 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/X 0.00fF
C398 sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/c1_n260_n210# clock_v2_0/p1d_b 0.02fF
C399 a_mux4_en_1/in1 a_mux4_en_0/in1 1.08fF
C400 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# -0.00fF
C401 ota_v2_0/p1 ota_v2_0/p2 6.27fF
C402 a_mux4_en_0/in3 VDD 0.31fF
C403 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VDD -0.00fF
C404 a_mux4_en_1/in2 a_mux4_en_0/switch_5t_mux4_3/in 0.08fF
C405 rst_n ota_v2_0/p1_b 0.83fF
C406 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# -0.21fF
C407 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_w_test_v2_0/ip -0.54fF
C408 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# 0.11fF
C409 sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# 0.03fF
C410 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C411 clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C412 transmission_gate_7/en VDD 5.09fF
C413 a_mux4_en_0/in0 a_mux4_en_0/switch_5t_mux4_1/in -0.00fF
C414 a_mux4_en_1/switch_5t_mux4_1/in a_mod_grp_ctrl_0 0.00fF
C415 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.01fF
C416 sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C417 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.00fF
C418 a_probe_1 a_mod_grp_ctrl_0 0.20fF
C419 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.00fF
C420 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# 0.09fF
C421 ota_v2_0/p2 sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.05fF
C422 a_mux4_en_0/in2 ip 0.25fF
C423 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.00fF
C424 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# 0.07fF
C425 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.13fF
C426 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.12fF
C427 a_mux4_en_0/switch_5t_mux4_1/a_300_216# a_mux4_en_0/switch_5t_mux4_1/en_b -0.00fF
C428 a_mux4_en_1/switch_5t_mux4_2/a_300_216# a_mux4_en_1/switch_5t_mux4_2/en_b -0.00fF
C429 a_mux4_en_1/switch_5t_mux4_1/en_b a_mod_grp_ctrl_1 0.08fF
C430 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C431 a_mux4_en_0/switch_5t_mux4_3/en_b a_mux4_en_0/switch_5t_mux4_3/in -0.00fF
C432 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A -0.01fF
C433 transmission_gate_2/in clock_v2_0/B_b 0.43fF
C434 clock_v2_0/A_b transmission_gate_2/in 0.42fF
C435 a_mux4_en_0/in1 ip 0.40fF
C436 transmission_gate_21/out ota_v2_0/p2 0.06fF
C437 a_mux2_en_0/in0 ota_w_test_v2_0/in 0.23fF
C438 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.09fF
C439 transmission_gate_31/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980# 1.14fF
C440 ota_v2_0/p1 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in 0.01fF
C441 a_mux4_en_0/switch_5t_mux4_0/en VDD 0.01fF
C442 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X -0.00fF
C443 ota_v2_0/p2_b sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C444 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# 0.03fF
C445 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/ip 0.00fF
C446 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A 0.02fF
C447 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/X 0.01fF
C448 sky130_fd_sc_hd__mux4_1_2/a_1290_413# clock_v2_0/Bd 0.00fF
C449 d_probe_3 d_probe_2 1.23fF
C450 ota_v2_0/cm transmission_gate_23/in 0.12fF
C451 ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_v2_0/on 0.00fF
C452 rst_n ota_v2_0/p2_b 1.02fF
C453 ota_v2_0/p2 transmission_gate_2/in 0.12fF
C454 a_mux4_en_0/switch_5t_mux4_2/en_b a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C455 sky130_fd_sc_hd__mux4_1_3/a_27_413# ota_v2_0/p1_b 0.02fF
C456 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# 0.03fF
C457 clock_v2_0/p2d sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# 0.09fF
C458 VDD transmission_gate_3/in 3.15fF
C459 debug a_mux2_en_1/switch_5t_mux2_1/in -0.00fF
C460 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.11fF
C461 ota_v2_0/sc_cmfb_0/transmission_gate_7/in VDD 0.67fF
C462 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_3/a_113_47# a_mux4_en_0/switch_5t_mux4_0/en_b -0.00fF
C463 transmission_gate_25/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# 0.49fF
C464 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in -0.00fF
C465 clock_v2_0/A_b clock_v2_0/B 1.20fF
C466 clock_v2_0/A_b clock_v2_0/Bd 0.42fF
C467 clock_v2_0/Bd clock_v2_0/B_b 18.03fF
C468 clock_v2_0/B clock_v2_0/B_b 19.88fF
C469 ota_v2_0/cm ota_v2_0/sc_cmfb_0/cmc 0.00fF
C470 ota_w_test_v2_0/ip clock_v2_0/A 0.18fF
C471 a_mux4_en_0/in3 a_mux4_en_0/transmission_gate_3/en_b 0.03fF
C472 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VDD -0.00fF
C473 sky130_fd_sc_hd__mux4_1_3/a_750_97# clock_v2_0/A 0.00fF
C474 sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__mux4_1_1/a_27_47# -0.00fF
C475 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.21fF
C476 a_mux2_en_0/in1 ota_v2_0/p1 0.07fF
C477 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# transmission_gate_21/out 0.03fF
C478 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.03fF
C479 transmission_gate_30/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.53fF
C480 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# 0.04fF
C481 sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/c1_n260_n210# ota_v2_0/op 0.03fF
C482 a_mux4_en_1/switch_5t_mux4_0/in a_mod_grp_ctrl_0 0.00fF
C483 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y VDD 0.13fF
C484 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21# clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C485 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# -0.00fF
C486 sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/c1_n260_n210# ota_v2_0/op 0.06fF
C487 ota_v2_0/p2 ota_v2_0/sc_cmfb_0/transmission_gate_4/out 0.00fF
C488 debug a_mux2_en_0/transmission_gate_1/en_b -0.00fF
C489 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/X 0.01fF
C490 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# -0.12fF
C491 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.03fF
C492 a_mux2_en_1/transmission_gate_1/en_b VDD 0.21fF
C493 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/c1_n260_n210# 0.02fF
C494 ota_v2_0/p2 clock_v2_0/Bd 0.86fF
C495 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# 0.09fF
C496 ota_v2_0/p2 clock_v2_0/B 3.21fF
C497 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.01fF
C498 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.02fF
C499 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_592_47# clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C500 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/p2d_b 0.15fF
C501 a_mux4_en_0/switch_5t_mux4_0/en a_mod_grp_ctrl_1 0.20fF
C502 debug a_mux4_en_1/switch_5t_mux4_1/en_b 0.16fF
C503 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in a_mod_grp_ctrl_0 -0.00fF
C504 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_1/en 0.19fF
C505 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/m3_n1030_n980# 0.09fF
C506 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.06fF
C507 sky130_fd_sc_hd__mux4_1_1/a_193_47# clock_v2_0/p1d 0.02fF
C508 ota_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/p1_b 0.00fF
C509 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C510 clock_v2_0/p2d_b ota_v2_0/on 0.07fF
C511 a_mux4_en_0/switch_5t_mux4_2/en VDD 0.15fF
C512 sky130_fd_sc_hd__mux4_1_0/a_1290_413# ota_v2_0/p2_b -0.00fF
C513 transmission_gate_30/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.03fF
C514 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/Ad 0.00fF
C515 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0.01fF
C516 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.06fF
C517 sky130_fd_sc_hd__mux4_1_3/a_277_47# clock_v2_0/B_b 0.00fF
C518 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# ota_v2_0/ip 0.03fF
C519 a_mux4_en_1/in1 a_mux4_en_1/in0 0.59fF
C520 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# -0.12fF
C521 sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/m3_n1030_n980# -0.06fF
C522 debug a_mux4_en_0/in3 0.03fF
C523 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# ota_v2_0/on 0.03fF
C524 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# ota_v2_0/ip 0.23fF
C525 ota_v2_0/p1 ota_v2_0/on 0.23fF
C526 ota_w_test_v2_0/in VDD 0.64fF
C527 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_1/in 0.00fF
C528 transmission_gate_7/en clock_v2_0/p1d 0.59fF
C529 sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C530 transmission_gate_29/out ota_v2_0/on 0.04fF
C531 i_bias_2 VDD 4.19fF
C532 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/c1_n930_n880# 0.07fF
C533 onebit_dac_1/v_b comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# -0.00fF
C534 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# 0.03fF
C535 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.02fF
C536 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# 3.46fF
C537 sky130_fd_sc_hd__mux4_1_0/a_27_413# clock_v2_0/B 0.01fF
C538 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# 0.04fF
C539 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# -0.14fF
C540 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C541 op comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# -0.00fF
C542 ota_v2_0/in VDD 1.65fF
C543 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# ota_v2_0/op 0.12fF
C544 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y a_mod_grp_ctrl_1 0.02fF
C545 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/X 0.01fF
C546 sky130_fd_sc_hd__mux4_1_3/a_27_413# d_clk_grp_1_ctrl_0 0.00fF
C547 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C548 sky130_fd_sc_hd__mux4_1_1/X clock_v2_0/Ad_b 0.00fF
C549 a_mux2_en_0/in0 ip 0.70fF
C550 sky130_fd_sc_hd__mux4_1_2/a_668_97# clock_v2_0/Bd_b 0.00fF
C551 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# 0.04fF
C552 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/p1 0.05fF
C553 ota_v2_0/in ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# 0.11fF
C554 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210# -0.04fF
C555 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p1 0.00fF
C556 a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in VDD 0.60fF
C557 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# transmission_gate_9/in 1.53fF
C558 op VDD 27.49fF
C559 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__clkinv_4_0/Y 0.16fF
C560 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/c1_n930_n880# -0.01fF
C561 a_mux4_en_0/switch_5t_mux4_3/en_b a_mux4_en_0/switch_5t_mux4_3/en 0.00fF
C562 a_mux4_en_1/in0 ip 0.19fF
C563 sky130_fd_sc_hd__clkinv_4_0/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.22fF
C564 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.02fF
C565 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.00fF
C566 sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980# -0.01fF
C567 a_mux4_en_0/switch_5t_mux4_2/en a_mod_grp_ctrl_1 0.08fF
C568 debug a_mux4_en_0/switch_5t_mux4_0/en 0.13fF
C569 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# -0.26fF
C570 a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in VDD 0.58fF
C571 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# -0.00fF
C572 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C573 clock_v2_0/A_b clock_v2_0/p1d_b 0.76fF
C574 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.01fF
C575 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.04fF
C576 clock_v2_0/p1d_b clock_v2_0/B_b 0.96fF
C577 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# -0.00fF
C578 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VDD -0.00fF
C579 a_mux2_en_0/in1 clock_v2_0/Bd 0.11fF
C580 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651# 0.00fF
C581 transmission_gate_30/out ota_v2_0/in 1.37fF
C582 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# transmission_gate_3/in 0.13fF
C583 sky130_fd_sc_hd__mux4_1_2/a_668_97# VDD 0.01fF
C584 clock_v2_0/p2d clock_v2_0/B_b 0.75fF
C585 i_bias_2 a_mod_grp_ctrl_1 0.13fF
C586 clock_v2_0/A_b clock_v2_0/p2d 0.68fF
C587 a_mux4_en_1/in1 VDD 5.81fF
C588 sky130_fd_sc_hd__mux4_1_0/X clock_v2_0/B_b 0.00fF
C589 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/c1_n260_n210# 0.03fF
C590 a_mux4_en_1/in1 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.02fF
C591 clock_v2_0/p2d_b sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.09fF
C592 ota_v2_0/p2 ota_v2_0/op 0.05fF
C593 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/ota_v2_without_cmfb_0/bias_b 0.06fF
C594 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C595 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.02fF
C596 sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/c1_n260_n210# ota_v2_0/op 0.03fF
C597 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# 0.09fF
C598 ota_v2_0/ip transmission_gate_21/in 1.55fF
C599 transmission_gate_7/en clock_v2_0/A 0.30fF
C600 clock_v2_0/p1d_b ota_v2_0/p2 0.92fF
C601 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# VDD 0.26fF
C602 clock_v2_0/B_b clock_v2_0/Ad 0.93fF
C603 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C604 clock_v2_0/A_b clock_v2_0/Ad 17.92fF
C605 clock_v2_0/p2d ota_v2_0/p2 8.55fF
C606 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.01fF
C607 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.01fF
C608 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# -0.00fF
C609 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD 0.06fF
C610 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210# 0.03fF
C611 sky130_fd_sc_hd__mux4_1_0/a_750_97# VDD 0.16fF
C612 sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# 0.03fF
C613 debug a_mux2_en_1/transmission_gate_1/en_b -0.00fF
C614 sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C615 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/Bd 0.00fF
C616 a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in a_mod_grp_ctrl_1 0.23fF
C617 sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# 0.03fF
C618 a_mod_grp_ctrl_0 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.01fF
C619 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/Ad_b 0.14fF
C620 ota_v2_0/p2 clock_v2_0/Ad 0.93fF
C621 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.01fF
C622 a_mux4_en_0/in0 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# 0.00fF
C623 transmission_gate_31/out VDD 0.82fF
C624 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.09fF
C625 transmission_gate_2/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/m3_n1030_n980# 1.65fF
C626 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# 0.03fF
C627 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.00fF
C628 sky130_fd_sc_hd__mux4_1_2/a_193_413# VDD 0.06fF
C629 a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in a_mod_grp_ctrl_1 0.14fF
C630 VDD ip 5.17fF
C631 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C632 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_w_test_v2_0/in 0.04fF
C633 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651# a_mux4_en_0/in1 -0.00fF
C634 debug a_mux4_en_0/switch_5t_mux4_2/en 0.12fF
C635 a_mux4_en_1/switch_5t_mux4_1/in VDD 1.35fF
C636 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.01fF
C637 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# 0.03fF
C638 ota_v2_0/cm clock_v2_0/p2d_b 0.07fF
C639 ota_v2_0/p1 transmission_gate_9/in 0.65fF
C640 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# -0.14fF
C641 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.02fF
C642 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210# ota_v2_0/op 0.03fF
C643 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_15613_3568# VDD 0.01fF
C644 a_probe_1 VDD 4.63fF
C645 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C646 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/sky130_fd_sc_hd__nand2_1_3/a_113_47# -0.00fF
C647 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C648 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210# 0.02fF
C649 clock_v2_0/B_b ota_v2_0/p1_b 1.14fF
C650 clock_v2_0/A_b ota_v2_0/p1_b 3.79fF
C651 debug i_bias_2 0.15fF
C652 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C653 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__clkinv_4_2/Y 0.17fF
C654 clock_v2_0/A transmission_gate_3/in 0.57fF
C655 ota_v2_0/p1 ota_w_test_v2_0/op -0.04fF
C656 ota_v2_0/cm ota_v2_0/p1 0.24fF
C657 a_mux4_en_0/in2 a_mux4_en_0/in0 0.73fF
C658 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A -0.00fF
C659 sky130_fd_sc_hd__mux4_1_0/a_27_413# clock_v2_0/Ad 0.00fF
C660 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00fF
C661 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C662 rst_n transmission_gate_7/en 18.57fF
C663 in transmission_gate_29/out 0.05fF
C664 ota_v2_0/p2 ota_v2_0/p1_b 14.84fF
C665 sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# -0.04fF
C666 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# VDD 0.58fF
C667 transmission_gate_30/out ip 0.01fF
C668 sky130_fd_sc_hd__mux4_1_3/a_27_47# VDD 0.00fF
C669 a_mux4_en_0/in0 a_mux4_en_0/in1 0.76fF
C670 sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/c1_n930_n880# -0.06fF
C671 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.00fF
C672 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C673 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.09fF
C674 debug a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in 0.40fF
C675 transmission_gate_23/in ota_v2_0/p1 0.70fF
C676 a_mux2_en_0/in1 clock_v2_0/p1d_b 0.47fF
C677 transmission_gate_29/out transmission_gate_23/in 0.23fF
C678 sky130_fd_sc_hd__mux4_1_1/a_247_21# clock_v2_0/Ad_b 0.12fF
C679 sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.01fF
C680 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# -0.01fF
C681 a_mux4_en_1/in1 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# 0.01fF
C682 a_mux4_en_1/switch_5t_mux4_1/in a_mod_grp_ctrl_1 0.00fF
C683 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C684 sky130_fd_sc_hd__mux4_1_0/a_668_97# clock_v2_0/B_b 0.00fF
C685 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C686 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# -0.06fF
C687 a_mux4_en_0/switch_5t_mux4_2/en_b a_mux4_en_0/switch_5t_mux4_2/en -0.00fF
C688 debug a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in 0.14fF
C689 d_clk_grp_1_ctrl_0 d_probe_2 1.19fF
C690 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# transmission_gate_3/in 0.17fF
C691 a_probe_1 a_mod_grp_ctrl_1 0.31fF
C692 transmission_gate_2/in transmission_gate_9/in 0.29fF
C693 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C694 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD 0.01fF
C695 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/B_b 0.00fF
C696 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# 0.12fF
C697 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/sc_cmfb_0/bias_a 0.00fF
C698 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/p1 -0.03fF
C699 clock_v2_0/A_b ota_v2_0/p2_b 1.18fF
C700 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD 0.00fF
C701 ota_v2_0/p2_b clock_v2_0/B_b 3.41fF
C702 ota_v2_0/ota_v2_without_cmfb_0/bias_b VDD 7.93fF
C703 a_mux4_en_1/switch_5t_mux4_0/in VDD 1.02fF
C704 onebit_dac_1/out a_mux4_en_1/in2 0.10fF
C705 ota_w_test_v2_0/in clock_v2_0/A 0.19fF
C706 a_mux2_en_0/in1 clock_v2_0/Ad 0.27fF
C707 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_v2_0/sc_cmfb_0/transmission_gate_6/in -0.00fF
C708 debug a_mux4_en_1/in1 0.03fF
C709 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y -0.00fF
C710 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A VDD 0.47fF
C711 a_probe_0 a_mod_grp_ctrl_0 0.20fF
C712 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/X 0.01fF
C713 d_clk_grp_1_ctrl_1 d_probe_1 1.18fF
C714 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_3/X 0.07fF
C715 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.12fF
C716 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/p1_b 0.00fF
C717 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A -0.00fF
C718 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C719 ota_v2_0/op ota_v2_0/on 3.50fF
C720 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__clkinv_4_3/Y 0.10fF
C721 rst_n transmission_gate_3/in 1.13fF
C722 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# 0.09fF
C723 ota_v2_0/sc_cmfb_0/transmission_gate_6/in VDD 3.23fF
C724 onebit_dac_1/out a_mux2_en_0/in1 0.36fF
C725 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/c1_n930_n880# 0.07fF
C726 a_mux4_en_1/switch_5t_mux4_1/en VDD 0.12fF
C727 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in VDD 0.60fF
C728 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VDD 0.00fF
C729 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_750_97# -0.00fF
C730 sky130_fd_sc_hd__clkinv_4_2/Y d_probe_2 0.09fF
C731 ota_v2_0/p2_b ota_v2_0/p2 33.03fF
C732 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_3/a_277_47# -0.00fF
C733 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# 0.03fF
C734 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/c1_n930_n880# 0.07fF
C735 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# 0.04fF
C736 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.08fF
C737 sky130_fd_sc_hd__mux4_1_0/a_750_97# d_clk_grp_2_ctrl_1 0.00fF
C738 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C739 ota_v2_0/p2 transmission_gate_25/in 0.57fF
C740 clock_v2_0/p2d ota_v2_0/on 0.49fF
C741 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VDD -0.01fF
C742 clock_v2_0/A_b d_clk_grp_1_ctrl_0 0.07fF
C743 d_clk_grp_1_ctrl_0 clock_v2_0/B_b 0.14fF
C744 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# transmission_gate_23/in 0.01fF
C745 transmission_gate_31/out clock_v2_0/p1d 0.14fF
C746 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.03fF
C747 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# 0.03fF
C748 sky130_fd_sc_hd__mux4_1_2/a_193_413# clock_v2_0/p1d 0.00fF
C749 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.00fF
C750 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S 0.21fF
C751 ip clock_v2_0/p1d 1.49fF
C752 a_mux4_en_0/switch_5t_mux4_1/in VDD 0.93fF
C753 ota_w_test_v2_0/op clock_v2_0/Bd 0.52fF
C754 d_clk_grp_1_ctrl_0 ota_v2_0/p2 0.03fF
C755 a_mux2_en_0/in1 ota_v2_0/p1_b 0.05fF
C756 a_mux4_en_0/in2 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# 0.08fF
C757 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# transmission_gate_3/in 0.13fF
C758 sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.02fF
C759 debug a_mux4_en_1/switch_5t_mux4_1/in 0.18fF
C760 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# -0.01fF
C761 transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/c1_n930_n880# -0.84fF
C762 onebit_dac_1/out ota_v2_0/on 0.16fF
C763 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.07fF
C764 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C765 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# ota_v2_0/ip 0.03fF
C766 sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C767 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/p2 -0.00fF
C768 a_mux4_en_1/switch_5t_mux4_0/in a_mod_grp_ctrl_1 0.00fF
C769 debug a_probe_1 0.31fF
C770 ota_v2_0/p2_b sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.04fF
C771 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A -0.01fF
C772 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C773 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.02fF
C774 ota_v2_0/p2_b ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in 0.00fF
C775 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# 0.07fF
C776 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_247_21# -0.01fF
C777 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.26fF
C778 sky130_fd_sc_hd__mux4_1_3/X ota_v2_0/p1_b 0.00fF
C779 i_bias_2 onebit_dac_0/out 0.17fF
C780 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.03fF
C781 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# ota_v2_0/in 0.03fF
C782 a_mux4_en_1/switch_5t_mux4_1/en a_mod_grp_ctrl_1 0.08fF
C783 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.00fF
C784 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in a_mod_grp_ctrl_1 0.16fF
C785 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.00fF
C786 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# 0.11fF
C787 a_mux2_en_0/in0 a_mux4_en_0/in0 0.18fF
C788 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.09fF
C789 transmission_gate_32/out a_mux2_en_0/in0 -1.11fF
C790 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# -0.00fF
C791 sky130_fd_sc_hd__mux4_1_1/a_668_97# clock_v2_0/B_b 0.00fF
C792 sky130_fd_sc_hd__mux4_1_1/X VDD 1.03fF
C793 ota_v2_0/on ota_v2_0/p1_b 0.18fF
C794 onebit_dac_1/v_b VDD 3.36fF
C795 a_mux4_en_1/in2 a_mux4_en_0/switch_5t_mux4_2/in 0.08fF
C796 clock_v2_0/A_b ota_w_test_v2_0/ip 0.26fF
C797 clock_v2_0/B_b ota_w_test_v2_0/ip 0.16fF
C798 ota_v2_0/in rst_n 0.09fF
C799 a_mux4_en_0/in0 a_mux4_en_1/in0 0.01fF
C800 sky130_fd_sc_hd__mux4_1_3/a_750_97# clock_v2_0/B_b 0.00fF
C801 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.12fF
C802 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C803 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# -0.21fF
C804 a_mux4_en_1/in1 a_mux4_en_1/switch_5t_mux4_2/in -0.00fF
C805 a_mux4_en_0/switch_5t_mux4_1/in a_mod_grp_ctrl_1 0.00fF
C806 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.02fF
C807 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C808 a_mux4_en_0/in2 a_mux4_en_0/in1 0.11fF
C809 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# 0.13fF
C810 ota_v2_0/ota_v2_without_cmfb_0/m1_15613_3568# VDD 0.01fF
C811 a_mux2_en_0/in1 ota_v2_0/p2_b 0.05fF
C812 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y -0.00fF
C813 ota_w_test_v2_0/on clock_v2_0/Ad_b 0.07fF
C814 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/c1_n260_n210# 0.03fF
C815 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C816 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# 0.12fF
C817 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# -0.00fF
C818 sky130_fd_sc_hd__mux4_1_1/a_1290_413# clock_v2_0/p1d_b -0.00fF
C819 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/c1_n260_n210# ota_v2_0/on 0.06fF
C820 ota_v2_0/sc_cmfb_0/bias_a VDD 7.94fF
C821 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C822 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# 0.12fF
C823 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651# VDD 0.30fF
C824 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/p1_b 0.00fF
C825 a_mux4_en_0/transmission_gate_3/en_b a_mux4_en_0/switch_5t_mux4_1/in 0.00fF
C826 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.04fF
C827 sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.03fF
C828 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p1_b -0.02fF
C829 a_mux4_en_1/switch_5t_mux4_1/en_b a_mux4_en_1/switch_5t_mux4_2/en_b 0.00fF
C830 debug a_mux4_en_1/switch_5t_mux4_0/in 0.18fF
C831 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/Bd_b 0.00fF
C832 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/sc_cmfb_0/bias_a -0.00fF
C833 ota_v2_0/ip VDD 1.01fF
C834 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VDD 0.09fF
C835 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/switch_5t_mux4_3/en_b -0.00fF
C836 sky130_fd_sc_hd__mux4_1_3/a_757_363# ota_v2_0/p1_b 0.06fF
C837 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C838 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# VDD 0.03fF
C839 sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980# 0.17fF
C840 i_bias_1 VDD 4.25fF
C841 a_mux4_en_1/in1 onebit_dac_0/out 0.14fF
C842 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C843 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# 0.03fF
C844 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y VDD 0.13fF
C845 sky130_fd_sc_hd__mux4_1_1/a_1290_413# clock_v2_0/Ad 0.00fF
C846 sky130_fd_sc_hd__mux4_1_0/a_277_47# clock_v2_0/B -0.00fF
C847 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C848 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C849 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.03fF
C850 ota_v2_0/cm ota_v2_0/op 0.31fF
C851 debug a_mux4_en_1/switch_5t_mux4_1/en 0.12fF
C852 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/ip 0.00fF
C853 a_mux2_en_1/switch_5t_mux2_1/en a_mux2_en_1/switch_5t_mux2_0/in -0.02fF
C854 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in debug 0.15fF
C855 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD 0.06fF
C856 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.02fF
C857 ota_w_test_v2_0/on a_mux4_en_0/in2 0.56fF
C858 ota_v2_0/p2_b ota_v2_0/on 0.08fF
C859 transmission_gate_31/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# 0.41fF
C860 a_mux4_en_1/switch_5t_mux4_1/in a_mux4_en_1/switch_5t_mux4_2/in -0.00fF
C861 a_mux2_en_0/switch_5t_mux2_0/in a_mux2_en_0/switch_5t_mux2_1/en -0.02fF
C862 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C863 sky130_fd_sc_hd__mux4_1_3/a_27_47# clock_v2_0/A -0.00fF
C864 sky130_fd_sc_hd__mux4_1_3/a_834_97# ota_v2_0/p1_b 0.01fF
C865 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C866 ota_v2_0/cm clock_v2_0/p2d 0.07fF
C867 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/X 0.00fF
C868 sky130_fd_sc_hd__mux4_1_1/a_750_97# VDD 0.17fF
C869 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.25fF
C870 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0.00fF
C871 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# -0.14fF
C872 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# 0.03fF
C873 a_mux4_en_0/switch_5t_mux4_3/en a_mux4_en_0/switch_5t_mux4_3/in 0.00fF
C874 ota_v2_0/p1 clock_v2_0/p2d_b 2.42fF
C875 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A 0.38fF
C876 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210# -0.07fF
C877 transmission_gate_32/out VDD 1.44fF
C878 a_mux4_en_0/in0 VDD 8.05fF
C879 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.00fF
C880 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210# 0.03fF
C881 transmission_gate_29/out clock_v2_0/p2d_b 0.30fF
C882 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# a_mux4_en_0/in0 0.03fF
C883 in clock_v2_0/p1d_b 1.02fF
C884 m5_41088_30705# transmission_gate_9/in 0.19fF
C885 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X -0.00fF
C886 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/c1_n260_n210# ota_v2_0/op 0.06fF
C887 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/c1_n930_n880# 0.07fF
C888 debug a_mux4_en_0/switch_5t_mux4_1/in 0.67fF
C889 in clock_v2_0/p2d 0.18fF
C890 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# 0.13fF
C891 transmission_gate_30/out ota_v2_0/ip 0.03fF
C892 transmission_gate_31/out onebit_dac_0/out 0.09fF
C893 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/Ad_b 0.07fF
C894 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C895 ota_w_test_v2_0/op clock_v2_0/Ad 0.50fF
C896 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# 0.14fF
C897 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.01fF
C898 a_mux2_en_0/in0 clock_v2_0/Ad_b 0.23fF
C899 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/p2_b 0.00fF
C900 onebit_dac_0/out ip 0.17fF
C901 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.05fF
C902 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/switch_5t_mux4_1/en_b 0.00fF
C903 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.01fF
C904 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p2_b 0.01fF
C905 sky130_fd_sc_hd__mux4_1_1/a_27_47# VDD 0.01fF
C906 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# 0.03fF
C907 a_mux4_en_1/in0 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# -0.00fF
C908 a_mux4_en_1/switch_5t_mux4_2/a_300_216# a_mux4_en_1/switch_5t_mux4_2/en -0.00fF
C909 ota_v2_0/p2_b sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.00fF
C910 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/op 0.38fF
C911 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y a_mod_grp_ctrl_1 0.02fF
C912 sky130_fd_sc_hd__mux4_1_3/a_193_413# ota_v2_0/p2 0.00fF
C913 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# 0.07fF
C914 a_mux2_en_0/in1 ota_w_test_v2_0/ip 0.47fF
C915 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.00fF
C916 sky130_fd_sc_hd__mux4_1_0/a_193_413# VDD 0.05fF
C917 sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.00fF
C918 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.03fF
C919 onebit_dac_1/out in 0.17fF
C920 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clk 0.02fF
C921 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210# 0.03fF
C922 sky130_fd_sc_hd__mux4_1_3/a_247_21# ota_v2_0/p1_b 0.04fF
C923 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y VDD 0.21fF
C924 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C925 ota_v2_0/p1_b transmission_gate_9/in 0.50fF
C926 transmission_gate_21/out clock_v2_0/p2d_b 0.16fF
C927 sky130_fd_sc_hd__mux4_1_1/X d_clk_grp_2_ctrl_1 0.00fF
C928 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.12fF
C929 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C930 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A -0.00fF
C931 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.01fF
C932 sky130_fd_sc_hd__mux4_1_1/a_27_413# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C933 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VDD 0.08fF
C934 sky130_fd_sc_hd__mux4_1_3/a_834_97# ota_v2_0/p2_b 0.00fF
C935 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/m3_n1030_n980# transmission_gate_3/in 0.17fF
C936 clock_v2_0/A_b transmission_gate_7/en 0.28fF
C937 transmission_gate_7/en clock_v2_0/B_b 0.29fF
C938 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y -0.00fF
C939 sky130_fd_sc_hd__mux4_1_3/a_1478_413# ota_v2_0/p1 -0.00fF
C940 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/c1_n260_n210# 0.03fF
C941 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_757_363# -0.00fF
C942 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.03fF
C943 ota_v2_0/p1 transmission_gate_21/out 0.07fF
C944 ota_w_test_v2_0/op ota_v2_0/p1_b 0.01fF
C945 ota_v2_0/cm ota_v2_0/p1_b 0.30fF
C946 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.01fF
C947 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C948 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# 0.13fF
C949 clock_v2_0/Ad_b clock_v2_0/Bd_b 6.24fF
C950 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# ota_v2_0/op 0.03fF
C951 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_w_test_v2_0/op -0.00fF
C952 a_mux4_en_0/in2 a_mux4_en_1/in0 0.35fF
C953 a_mux4_en_0/switch_5t_mux4_1/en a_mux4_en_0/switch_5t_mux4_0/en_b -0.00fF
C954 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/a_923_363# 0.02fF
C955 sky130_fd_sc_hd__mux4_1_1/a_247_21# VDD 0.06fF
C956 sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C957 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# ota_v2_0/ip 0.14fF
C958 a_probe_0 VDD 4.64fF
C959 ota_v2_0/p2 transmission_gate_7/en 0.72fF
C960 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C961 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# clock_v2_0/p1d_b 0.02fF
C962 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C963 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C964 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.06fF
C965 a_mux4_en_1/in0 a_mux4_en_0/in1 0.25fF
C966 a_mux4_en_0/in0 a_mux4_en_0/transmission_gate_3/en_b 0.03fF
C967 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_18877_3928# ota_w_test_v2_0/in 0.00fF
C968 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C969 clock_v2_0/p2d sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/c1_n930_n880# 0.09fF
C970 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VDD 0.05fF
C971 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C972 d_probe_1 VDD 6.81fF
C973 transmission_gate_23/in ota_v2_0/p1_b 0.25fF
C974 VDD clock_v2_0/Ad_b 3.09fF
C975 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# VDD 2.04fF
C976 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VDD 0.31fF
C977 d_clk_grp_1_ctrl_1 VDD 6.38fF
C978 clock_v2_0/p2d_b sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.01fF
C979 sky130_fd_sc_hd__mux4_1_1/a_193_413# VDD 0.05fF
C980 transmission_gate_21/in VDD 1.04fF
C981 clock_v2_0/p2d_b clock_v2_0/B 0.87fF
C982 clock_v2_0/p2d_b clock_v2_0/Bd 1.82fF
C983 ota_v2_0/p2_b transmission_gate_9/in 0.42fF
C984 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.02fF
C985 ota_v2_0/p1 ota_v2_0/sc_cmfb_0/transmission_gate_4/out 0.06fF
C986 clock_v2_0/A_b transmission_gate_3/in 0.42fF
C987 clock_v2_0/B_b transmission_gate_3/in 0.50fF
C988 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210# ota_v2_0/on 0.03fF
C989 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/p1d 0.00fF
C990 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# transmission_gate_21/out 0.38fF
C991 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# 0.04fF
C992 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# 0.09fF
C993 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/p1_b -0.02fF
C994 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VDD 0.55fF
C995 ota_v2_0/p1 clock_v2_0/Bd 1.34fF
C996 ota_v2_0/p1 clock_v2_0/B 1.13fF
C997 ota_w_test_v2_0/on a_mux2_en_0/in0 1.02fF
C998 transmission_gate_32/out clock_v2_0/p1d 0.15fF
C999 a_mod_grp_ctrl_0 VDD 11.70fF
C1000 sky130_fd_sc_hd__mux4_1_1/a_750_97# d_clk_grp_2_ctrl_1 0.09fF
C1001 ota_v2_0/p2_b ota_w_test_v2_0/op -0.05fF
C1002 ota_v2_0/cm ota_v2_0/p2_b 0.07fF
C1003 comparator_v2_0/li_940_818# comparator_v2_0/li_940_3458# -0.00fF
C1004 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_750_97# -0.00fF
C1005 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C1006 ota_v2_0/cm transmission_gate_25/in 0.08fF
C1007 transmission_gate_31/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/c1_n930_n880# -0.36fF
C1008 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VDD -0.00fF
C1009 sky130_fd_sc_hd__mux4_1_2/a_923_363# VDD 0.01fF
C1010 ota_v2_0/p2 transmission_gate_3/in 0.10fF
C1011 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VDD 0.57fF
C1012 debug a_mux4_en_0/in0 0.03fF
C1013 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C1014 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.04fF
C1015 d_clk_grp_2_ctrl_0 clock_v2_0/p2d_b 0.18fF
C1016 ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p2 0.04fF
C1017 a_mux4_en_1/in2 a_mux4_en_0/in3 0.11fF
C1018 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C1019 a_probe_0 a_mod_grp_ctrl_1 0.31fF
C1020 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_v2_0/on 0.01fF
C1021 a_mux4_en_0/in2 VDD 10.00fF
C1022 a_mux4_en_0/switch_5t_mux4_0/en a_mux4_en_0/switch_5t_mux4_0/in -0.03fF
C1023 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# -0.12fF
C1024 a_mux4_en_0/switch_5t_mux4_2/en a_mux4_en_0/switch_5t_mux4_2/a_300_216# -0.00fF
C1025 sky130_fd_sc_hd__mux4_1_3/a_1290_413# VDD 0.05fF
C1026 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/p1d 0.10fF
C1027 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# -0.01fF
C1028 ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_v2_0/op 0.01fF
C1029 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.21fF
C1030 sky130_fd_sc_hd__mux4_1_0/a_27_47# clock_v2_0/B 0.01fF
C1031 a_mux4_en_0/in1 VDD 6.81fF
C1032 d_probe_0 sky130_fd_sc_hd__clkinv_4_3/Y 1.85fF
C1033 sky130_fd_sc_hd__mux4_1_0/a_193_413# clock_v2_0/p1d 0.00fF
C1034 transmission_gate_23/in ota_v2_0/p2_b 0.31fF
C1035 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# a_mux4_en_0/in1 0.02fF
C1036 a_mux4_en_0/switch_5t_mux4_2/en_b a_mux4_en_0/sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C1037 sky130_fd_sc_hd__mux4_1_0/a_277_47# ota_v2_0/p1_b 0.00fF
C1038 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# 0.29fF
C1039 transmission_gate_23/in transmission_gate_25/in 0.49fF
C1040 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_3/a_277_47# -0.00fF
C1041 sky130_fd_sc_hd__mux4_1_1/a_1478_413# VDD 0.13fF
C1042 transmission_gate_8/in a_mux4_en_0/in0 0.03fF
C1043 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_1/X 0.17fF
C1044 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# ota_v2_0/on 0.03fF
C1045 transmission_gate_8/in transmission_gate_32/out 0.07fF
C1046 sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C1047 a_mux2_en_0/in1 transmission_gate_7/en 0.62fF
C1048 transmission_gate_2/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980# 0.17fF
C1049 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VDD 0.00fF
C1050 ota_w_test_v2_0/on clock_v2_0/Bd_b 0.49fF
C1051 ota_w_test_v2_0/in clock_v2_0/B_b 0.18fF
C1052 clock_v2_0/A_b ota_w_test_v2_0/in 0.24fF
C1053 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# ota_v2_0/in 0.27fF
C1054 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# 0.03fF
C1055 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X -0.00fF
C1056 a_mux4_en_0/switch_5t_mux4_0/en_b a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C1057 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X VDD 0.11fF
C1058 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.09fF
C1059 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# 0.13fF
C1060 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1 9.83fF
C1061 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C1062 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C1063 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980# transmission_gate_2/in 0.17fF
C1064 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# -0.21fF
C1065 transmission_gate_2/in clock_v2_0/B 0.52fF
C1066 sky130_fd_sc_hd__mux4_1_1/a_247_21# clock_v2_0/p1d 0.01fF
C1067 transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980# 1.59fF
C1068 onebit_dac_0/out onebit_dac_1/v_b 0.32fF
C1069 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C1070 sky130_fd_sc_hd__mux4_1_1/a_247_21# d_clk_grp_2_ctrl_1 0.01fF
C1071 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/c1_n260_n210# 0.03fF
C1072 ota_w_test_v2_0/on VDD 3.99fF
C1073 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980# 0.17fF
C1074 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C1075 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.01fF
C1076 clock_v2_0/p2d_b ota_v2_0/op 0.43fF
C1077 a_mod_grp_ctrl_0 a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C1078 debug a_probe_0 0.31fF
C1079 transmission_gate_7/en ota_v2_0/on -0.16fF
C1080 sky130_fd_sc_hd__mux4_1_1/a_757_363# clock_v2_0/Ad_b 0.01fF
C1081 ota_v2_0/in ota_v2_0/p2 0.10fF
C1082 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# 0.03fF
C1083 clock_v2_0/p1d_b clock_v2_0/p2d_b 10.67fF
C1084 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# 0.05fF
C1085 ota_v2_0/sc_cmfb_0/transmission_gate_8/in VDD 0.88fF
C1086 ota_w_test_v2_0/op ota_w_test_v2_0/ip 0.09fF
C1087 clock_v2_0/Ad_b clock_v2_0/p1d 1.12fF
C1088 ota_w_test_v2_0/op ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out 0.00fF
C1089 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.10fF
C1090 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/m3_n1030_n980# 0.09fF
C1091 sky130_fd_sc_hd__mux4_1_0/a_277_47# ota_v2_0/p2_b 0.05fF
C1092 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.01fF
C1093 ota_v2_0/p1 ota_v2_0/op 0.05fF
C1094 clock_v2_0/p2d clock_v2_0/p2d_b 27.11fF
C1095 d_clk_grp_2_ctrl_1 clock_v2_0/Ad_b 0.02fF
C1096 transmission_gate_21/in clock_v2_0/p1d 0.18fF
C1097 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# 0.07fF
C1098 a_mux2_en_0/in1 transmission_gate_3/in -11.45fF
C1099 transmission_gate_29/out ota_v2_0/op 0.20fF
C1100 clock_v2_0/B clock_v2_0/Bd 8.12fF
C1101 d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_1 0.01fF
C1102 a_mux4_en_0/in2 a_mux4_en_0/transmission_gate_3/en_b 0.03fF
C1103 comparator_v2_0/li_940_3458# VDD 1.47fF
C1104 a_mux4_en_1/switch_5t_mux4_1/a_300_216# a_mux4_en_1/switch_5t_mux4_1/en_b -0.00fF
C1105 clock_v2_0/p1d_b ota_v2_0/p1 5.38fF
C1106 ota_v2_0/ota_v2_without_cmfb_0/bias_c VDD 4.53fF
C1107 transmission_gate_29/out clock_v2_0/p1d_b 0.16fF
C1108 clock_v2_0/p2d ota_v2_0/p1 1.61fF
C1109 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/p2d_b 0.05fF
C1110 ota_w_test_v2_0/on m2_72825_34855# 0.25fF
C1111 onebit_dac_0/out i_bias_1 0.15fF
C1112 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/Bd_b 0.00fF
C1113 rst_n ota_v2_0/ip 0.24fF
C1114 clock_v2_0/p2d_b clock_v2_0/Ad 0.93fF
C1115 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C1116 clock_v2_0/p2d transmission_gate_29/out 0.14fF
C1117 a_mux4_en_0/in1 a_mux4_en_0/transmission_gate_3/en_b 0.03fF
C1118 a_mux2_en_0/in0 clock_v2_0/Bd_b 0.21fF
C1119 clock_v2_0/p2d sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/c1_n930_n880# 0.09fF
C1120 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A -0.00fF
C1121 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/Bd 0.01fF
C1122 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C1123 clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y VDD 0.13fF
C1124 sky130_fd_sc_hd__mux4_1_0/a_277_47# d_clk_grp_1_ctrl_0 0.07fF
C1125 comparator_v2_0/li_940_818# VDD 4.95fF
C1126 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210# 0.03fF
C1127 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C1128 d_clk_grp_2_ctrl_0 clock_v2_0/Bd 0.01fF
C1129 debug a_mod_grp_ctrl_0 7.42fF
C1130 a_mux4_en_0/switch_5t_mux4_1/en a_mux4_en_0/switch_5t_mux4_1/a_300_216# -0.00fF
C1131 ota_v2_0/p1 clock_v2_0/Ad 3.02fF
C1132 clock_v2_0/p2d_b sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.08fF
C1133 onebit_dac_1/out clock_v2_0/p2d_b 0.85fF
C1134 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C1135 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# ota_v2_0/in 0.11fF
C1136 ota_v2_0/sc_cmfb_0/transmission_gate_9/in VDD 0.58fF
C1137 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C1138 sky130_fd_sc_hd__mux4_1_2/a_1478_413# clock_v2_0/p2d_b -0.00fF
C1139 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1140 sky130_fd_sc_hd__mux4_1_0/a_750_97# clock_v2_0/B_b 0.13fF
C1141 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980# VDD 0.25fF
C1142 ota_v2_0/cm ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# -0.00fF
C1143 sky130_fd_sc_hd__mux4_1_1/a_277_47# VDD 0.11fF
C1144 transmission_gate_21/out ota_v2_0/op -0.00fF
C1145 transmission_gate_32/out onebit_dac_0/out 0.02fF
C1146 onebit_dac_0/out a_mux4_en_0/in0 0.22fF
C1147 a_mux4_en_0/in2 debug 0.03fF
C1148 rst_n a_mux4_en_0/in0 0.97fF
C1149 ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/on 0.05fF
C1150 a_mux2_en_0/in0 VDD 14.74fF
C1151 onebit_dac_1/out transmission_gate_29/out -0.18fF
C1152 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.01fF
C1153 clock_v2_0/p1d_b transmission_gate_21/out 0.20fF
C1154 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C1155 sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/c1_n930_n880# -0.01fF
C1156 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210# transmission_gate_23/in 0.01fF
C1157 a_mux2_en_0/in1 ota_w_test_v2_0/in 0.62fF
C1158 clock_v2_0/p2d transmission_gate_21/out 0.13fF
C1159 debug a_mux4_en_0/in1 0.03fF
C1160 a_mux4_en_1/in0 VDD 6.36fF
C1161 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_3/a_300_216# 1.43fF
C1162 sky130_fd_sc_hd__mux4_1_0/a_750_97# ota_v2_0/p2 0.00fF
C1163 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C1164 clock_v2_0/p2d_b ota_v2_0/p1_b 1.99fF
C1165 sky130_fd_sc_hd__mux4_1_1/a_1478_413# d_clk_grp_2_ctrl_1 0.00fF
C1166 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/c1_n930_n880# 0.07fF
C1167 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/switch_5t_mux4_3/in -0.00fF
C1168 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47# -0.00fF
C1169 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_3/a_247_21# -0.00fF
C1170 ota_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# -0.00fF
C1171 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/switch_5t_mux4_1/in 0.00fF
C1172 d_clk_grp_1_ctrl_1 clock_v2_0/A 0.01fF
C1173 clock_v2_0/A clock_v2_0/Ad_b 4.82fF
C1174 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# -0.02fF
C1175 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# 0.03fF
C1176 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# 0.07fF
C1177 a_mux4_en_0/switch_5t_mux4_3/en_b a_mux4_en_0/switch_5t_mux4_2/en -0.00fF
C1178 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y -0.00fF
C1179 ota_v2_0/p1 ota_v2_0/p1_b 35.51fF
C1180 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_1/a_113_47# a_mux4_en_1/switch_5t_mux4_2/en_b 0.00fF
C1181 sky130_fd_sc_hd__mux4_1_0/a_247_21# VDD 0.06fF
C1182 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.02fF
C1183 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# 0.07fF
C1184 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_218_374# 0.01fF
C1185 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# ota_v2_0/on 0.06fF
C1186 transmission_gate_30/out a_mux2_en_0/in0 0.06fF
C1187 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD 0.00fF
C1188 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.21fF
C1189 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_2/en_b 0.41fF
C1190 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.03fF
C1191 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/c1_n260_n210# ota_v2_0/on 0.03fF
C1192 ota_v2_0/sc_cmfb_0/transmission_gate_4/out ota_v2_0/op 0.00fF
C1193 clock_v2_0/p2d sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# 0.09fF
C1194 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.01fF
C1195 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/c1_n260_n210# -0.14fF
C1196 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# 0.07fF
C1197 sky130_fd_sc_hd__mux4_1_0/a_757_363# ota_v2_0/p1_b 0.00fF
C1198 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# 0.03fF
C1199 ota_v2_0/cm ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.03fF
C1200 VDD clock_v2_0/Bd_b 2.95fF
C1201 a_mux4_en_1/in1 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# 0.04fF
C1202 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y -0.00fF
C1203 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C1204 comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.33fF
C1205 clock_v2_0/p1d_b clock_v2_0/Bd 2.90fF
C1206 clock_v2_0/p1d_b clock_v2_0/B 0.93fF
C1207 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD 0.08fF
C1208 a_mux4_en_1/in2 a_mux4_en_1/in1 0.55fF
C1209 sky130_fd_sc_hd__clkinv_4_1/Y d_probe_1 0.06fF
C1210 comparator_v2_0/li_n2324_818# comparator_v2_0/li_940_3458# -0.00fF
C1211 clock_v2_0/p2d clock_v2_0/B 0.84fF
C1212 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.00fF
C1213 clock_v2_0/p2d clock_v2_0/Bd 2.52fF
C1214 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/p2d_b 0.00fF
C1215 sky130_fd_sc_hd__mux4_1_3/a_1290_413# clock_v2_0/A 0.00fF
C1216 sky130_fd_sc_hd__mux4_1_2/a_193_47# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.01fF
C1217 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_1/X 0.07fF
C1218 in a_mux4_en_0/in3 0.03fF
C1219 sky130_fd_sc_hd__mux4_1_3/a_1478_413# ota_v2_0/p1_b -0.00fF
C1220 ota_v2_0/cm transmission_gate_7/en 1.22fF
C1221 ota_v2_0/p2_b clock_v2_0/p2d_b 9.21fF
C1222 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.08fF
C1223 ota_v2_0/in ota_v2_0/on -0.00fF
C1224 transmission_gate_21/out ota_v2_0/p1_b 0.05fF
C1225 ota_v2_0/p2 sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.00fF
C1226 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_2/in 0.00fF
C1227 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/Bd 0.00fF
C1228 a_mux4_en_0/switch_5t_mux4_0/en a_mux4_en_0/switch_5t_mux4_0/en_b -0.01fF
C1229 clock_v2_0/Bd clock_v2_0/Ad 0.83fF
C1230 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VDD 0.11fF
C1231 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X -0.00fF
C1232 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C1233 clock_v2_0/B clock_v2_0/Ad 0.85fF
C1234 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# ota_v2_0/on 0.01fF
C1235 comparator_v2_0/li_940_818# comparator_v2_0/li_n2324_818# -0.00fF
C1236 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.00fF
C1237 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.05fF
C1238 d_clk_grp_2_ctrl_0 clock_v2_0/p1d_b 0.13fF
C1239 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# 0.09fF
C1240 ota_v2_0/p1 ota_v2_0/p2_b 4.20fF
C1241 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# 0.07fF
C1242 a_mux4_en_0/switch_5t_mux4_0/en a_mux4_en_0/switch_5t_mux4_0/a_300_216# -0.00fF
C1243 rst_n clock_v2_0/Ad_b 0.33fF
C1244 ota_v2_0/p1 transmission_gate_25/in 0.67fF
C1245 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# VDD 3.53fF
C1246 d_clk_grp_2_ctrl_0 clock_v2_0/p2d 0.03fF
C1247 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/switch_5t_mux4_0/in -0.00fF
C1248 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.01fF
C1249 sky130_fd_sc_hd__mux4_1_2/a_247_21# clock_v2_0/Bd 0.01fF
C1250 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.12fF
C1251 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00fF
C1252 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.02fF
C1253 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD 0.00fF
C1254 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B VDD 0.00fF
C1255 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/Ad 0.00fF
C1256 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_3/a_300_216# 1.71fF
C1257 sky130_fd_sc_hd__mux4_1_0/a_757_363# ota_v2_0/p2_b 0.10fF
C1258 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.07fF
C1259 ota_w_test_v2_0/on ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in -0.01fF
C1260 a_mux4_en_1/in2 ip 0.53fF
C1261 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# 0.03fF
C1262 a_mux4_en_1/in2 a_mux4_en_1/switch_5t_mux4_1/in 0.08fF
C1263 d_clk_grp_2_ctrl_0 clock_v2_0/Ad 0.00fF
C1264 transmission_gate_31/out a_mux2_en_0/in1 0.40fF
C1265 transmission_gate_3/in transmission_gate_9/in 2.35fF
C1266 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/switch_5t_mux4_1/en -0.00fF
C1267 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C1268 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C1269 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# 0.11fF
C1270 d_clk_grp_1_ctrl_0 ota_v2_0/p1 0.00fF
C1271 a_mux2_en_0/in0 clock_v2_0/p1d 0.76fF
C1272 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# 0.12fF
C1273 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_0/a_300_216# 0.26fF
C1274 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.01fF
C1275 sky130_fd_sc_hd__mux4_1_1/a_277_47# d_clk_grp_2_ctrl_1 0.12fF
C1276 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.00fF
C1277 transmission_gate_30/out VDD 0.61fF
C1278 a_mux2_en_0/in1 ip 0.33fF
C1279 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VDD 0.00fF
C1280 ota_v2_0/sc_cmfb_0/transmission_gate_4/out ota_v2_0/p1_b 0.01fF
C1281 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.20fF
C1282 ota_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p2 0.02fF
C1283 ota_v2_0/p1 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out 0.03fF
C1284 debug a_mux2_en_0/in0 -0.00fF
C1285 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C1286 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C1287 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# clock_v2_0/p1d_b 0.02fF
C1288 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_193_413# 0.01fF
C1289 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.01fF
C1290 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# 0.07fF
C1291 a_mux4_en_0/in2 onebit_dac_0/out 0.23fF
C1292 clock_v2_0/Bd ota_v2_0/p1_b 0.92fF
C1293 clock_v2_0/B ota_v2_0/p1_b 1.26fF
C1294 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VDD 0.07fF
C1295 sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# 0.01fF
C1296 transmission_gate_21/out ota_v2_0/p2_b 0.05fF
C1297 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VDD 0.00fF
C1298 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C1299 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980# 0.09fF
C1300 debug a_mux4_en_1/in0 0.03fF
C1301 m1_86360_35183# ota_v2_0/on 0.12fF
C1302 transmission_gate_21/out transmission_gate_25/in 0.10fF
C1303 VDD a_mod_grp_ctrl_1 11.29fF
C1304 onebit_dac_0/out a_mux4_en_0/in1 0.17fF
C1305 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# -0.00fF
C1306 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C1307 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.03fF
C1308 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C1309 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# transmission_gate_32/out -1.21fF
C1310 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.09fF
C1311 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X -0.00fF
C1312 ota_v2_0/p2_b transmission_gate_2/in 0.22fF
C1313 sky130_fd_sc_hd__clkinv_4_0/Y sky130_fd_sc_hd__mux4_1_1/X 0.01fF
C1314 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_1478_413# -0.00fF
C1315 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210# ota_v2_0/on -0.06fF
C1316 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y VDD 0.13fF
C1317 clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y VDD 0.12fF
C1318 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.01fF
C1319 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_193_47# 0.01fF
C1320 sky130_fd_sc_hd__mux4_1_1/a_757_363# clock_v2_0/Bd_b 0.00fF
C1321 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# -0.00fF
C1322 a_mux4_en_0/transmission_gate_3/en_b VDD 0.73fF
C1323 clock_v2_0/Bd_b clock_v2_0/p1d 0.81fF
C1324 clock_v2_0/p2d ota_v2_0/op 0.23fF
C1325 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# -0.02fF
C1326 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# 0.00fF
C1327 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# -0.00fF
C1328 clock_v2_0/p2d clock_v2_0/p1d_b 2.11fF
C1329 d_clk_grp_2_ctrl_1 clock_v2_0/Bd_b 0.02fF
C1330 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0.16fF
C1331 sky130_fd_sc_hd__mux4_1_3/a_277_47# ota_v2_0/p1_b 0.04fF
C1332 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.01fF
C1333 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# -0.00fF
C1334 a_mux4_en_0/switch_5t_mux4_0/in a_mux4_en_0/switch_5t_mux4_1/in 0.00fF
C1335 a_mux4_en_1/switch_5t_mux4_0/en a_mux4_en_1/switch_5t_mux4_0/in -0.03fF
C1336 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.00fF
C1337 ota_v2_0/p1 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out 0.02fF
C1338 ota_v2_0/p2_b ota_v2_0/sc_cmfb_0/transmission_gate_4/out 0.01fF
C1339 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_3/a_750_97# -0.00fF
C1340 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# 0.04fF
C1341 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.00fF
C1342 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C1343 comparator_v2_0/li_n2324_818# VDD 2.80fF
C1344 a_mux4_en_1/in2 a_mux4_en_1/switch_5t_mux4_0/in 0.08fF
C1345 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C1346 sky130_fd_sc_hd__mux4_1_2/a_27_413# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.01fF
C1347 ota_v2_0/p2_b clock_v2_0/Bd 0.82fF
C1348 ota_v2_0/p2_b clock_v2_0/B 2.41fF
C1349 clock_v2_0/p1d_b clock_v2_0/Ad 1.65fF
C1350 sky130_fd_sc_hd__mux4_1_1/a_757_363# VDD 0.06fF
C1351 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# 0.03fF
C1352 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_277_47# -0.00fF
C1353 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11122_5650# VDD 0.28fF
C1354 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/c1_n260_n210# 0.03fF
C1355 clock_v2_0/p2d clock_v2_0/Ad 1.04fF
C1356 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A -0.00fF
C1357 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.03fF
C1358 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C1359 VDD clock_v2_0/p1d 36.15fF
C1360 a_mux4_en_1/switch_5t_mux4_0/en a_mux4_en_1/switch_5t_mux4_1/en -0.00fF
C1361 onebit_dac_1/out ota_v2_0/op 0.42fF
C1362 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C1363 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.00fF
C1364 d_clk_grp_2_ctrl_1 VDD 6.60fF
C1365 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# ota_v2_0/on 0.03fF
C1366 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# ota_v2_0/ip 0.03fF
C1367 ota_v2_0/cm ota_v2_0/in 0.26fF
C1368 sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/c1_n260_n210# -0.07fF
C1369 sky130_fd_sc_hd__mux4_1_0/a_834_97# VDD 0.01fF
C1370 debug VDD 8.90fF
C1371 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C1372 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1373 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.00fF
C1374 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.01fF
C1375 sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# 0.12fF
C1376 onebit_dac_1/out clock_v2_0/p2d 1.27fF
C1377 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# -0.06fF
C1378 d_clk_grp_1_ctrl_0 clock_v2_0/B 0.01fF
C1379 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0.00fF
C1380 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C1381 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.03fF
C1382 a_mux4_en_0/transmission_gate_3/en_b a_mod_grp_ctrl_1 0.00fF
C1383 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C1384 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/p2 0.01fF
C1385 a_mux4_en_1/in2 a_mux4_en_0/switch_5t_mux4_1/in 0.08fF
C1386 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C1387 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.01fF
C1388 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# 0.13fF
C1389 ota_v2_0/op ota_v2_0/p1_b 0.07fF
C1390 sky130_fd_sc_hd__mux4_1_3/a_923_363# sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.00fF
C1391 ota_v2_0/p2_b sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C1392 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0.01fF
C1393 transmission_gate_30/out clock_v2_0/p1d 0.14fF
C1394 clock_v2_0/p1d_b ota_v2_0/p1_b 8.83fF
C1395 transmission_gate_8/in VDD 0.12fF
C1396 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/c1_n930_n880# 0.07fF
C1397 VDD a_mux4_en_1/switch_5t_mux4_3/a_300_216# 0.23fF
C1398 clock_v2_0/A clock_v2_0/Bd_b 0.52fF
C1399 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD 0.07fF
C1400 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C1401 ota_v2_0/ip ota_v2_0/p2 0.10fF
C1402 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# 0.28fF
C1403 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/c1_n930_n880# 0.07fF
C1404 clock_v2_0/p2d ota_v2_0/p1_b 0.95fF
C1405 d_clk_grp_2_ctrl_0 d_clk_grp_1_ctrl_0 0.01fF
C1406 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.11fF
C1407 transmission_gate_2/in ota_w_test_v2_0/ip 0.00fF
C1408 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# -0.01fF
C1409 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C1410 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C1411 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X -0.00fF
C1412 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_535_374# 0.00fF
C1413 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# a_mux4_en_1/in0 0.00fF
C1414 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in VDD 1.03fF
C1415 a_mux2_en_0/in0 onebit_dac_0/out 0.31fF
C1416 ota_v2_0/in ota_v2_0/sc_cmfb_0/cmc 0.31fF
C1417 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210# -0.07fF
C1418 clock_v2_0/Ad ota_v2_0/p1_b 1.00fF
C1419 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C1420 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.02fF
C1421 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.00fF
C1422 d_probe_3 sky130_fd_sc_hd__clkinv_4_2/Y 2.12fF
C1423 rst_n a_mux2_en_0/in0 0.13fF
C1424 in a_mux4_en_1/in1 0.20fF
C1425 a_mod_grp_ctrl_0 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_2/a_113_47# -0.00fF
C1426 a_mod_grp_ctrl_0 a_probe_3 2.56fF
C1427 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# VDD 0.60fF
C1428 debug a_mod_grp_ctrl_1 8.05fF
C1429 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# 0.07fF
C1430 a_mux4_en_0/switch_5t_mux4_1/in a_mux4_en_0/switch_5t_mux4_1/en_b -0.00fF
C1431 a_mux4_en_0/switch_5t_mux4_2/en_b VDD 1.01fF
C1432 onebit_dac_0/out a_mux4_en_1/in0 0.18fF
C1433 VDD clock_v2_0/A 2.31fF
C1434 transmission_gate_31/out transmission_gate_9/in 0.32fF
C1435 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B VDD -0.00fF
C1436 a_mux4_en_0/in0 ota_v2_0/p2 0.09fF
C1437 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD 0.00fF
C1438 sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C1439 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# transmission_gate_3/in 0.12fF
C1440 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/m3_n1030_n980# 0.17fF
C1441 clock_v2_0/B ota_w_test_v2_0/ip 0.11fF
C1442 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD 0.00fF
C1443 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/p1d_b 0.01fF
C1444 ota_v2_0/p2_b ota_v2_0/op 0.07fF
C1445 clock_v2_0/p2d_b transmission_gate_7/en 0.58fF
C1446 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD -0.00fF
C1447 debug a_mux4_en_0/transmission_gate_3/en_b -0.01fF
C1448 transmission_gate_25/in ota_v2_0/op 0.58fF
C1449 clock_v2_0/p1d_b ota_v2_0/p2_b 0.99fF
C1450 a_mux4_en_1/switch_5t_mux4_3/a_300_216# a_mod_grp_ctrl_1 0.04fF
C1451 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C1452 ota_v2_0/p2 sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C1453 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# -0.00fF
C1454 transmission_gate_31/out in 0.01fF
C1455 clock_v2_0/p1d_b transmission_gate_25/in 1.90fF
C1456 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C1457 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# VDD 0.06fF
C1458 clock_v2_0/p2d ota_v2_0/p2_b 18.47fF
C1459 ota_v2_0/p1 transmission_gate_7/en 0.76fF
C1460 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X -0.00fF
C1461 sky130_fd_sc_hd__mux4_1_0/X ota_v2_0/p2_b 0.00fF
C1462 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A VDD 13.63fF
C1463 a_mux4_en_1/switch_5t_mux4_2/in VDD 0.77fF
C1464 a_mux4_en_1/switch_5t_mux4_3/en_b a_mod_grp_ctrl_0 1.01fF
C1465 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C1466 d_probe_1 d_probe_2 0.10fF
C1467 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/c1_n260_n210# ota_v2_0/on 0.01fF
C1468 in ip 2.22fF
C1469 rst_n clock_v2_0/Bd_b 0.29fF
C1470 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.01fF
C1471 sky130_fd_sc_hd__clkinv_4_1/Y VDD 0.99fF
C1472 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0.09fF
C1473 a_mux4_en_1/switch_5t_mux4_1/a_300_216# a_mux4_en_1/switch_5t_mux4_1/en -0.00fF
C1474 d_clk_grp_1_ctrl_1 d_probe_2 0.10fF
C1475 d_clk_grp_2_ctrl_1 clock_v2_0/p1d 0.01fF
C1476 a_mux4_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0.19fF
C1477 ota_v2_0/p2_b clock_v2_0/Ad 1.13fF
C1478 a_mux4_en_1/in2 i_bias_1 1.54fF
C1479 a_mux4_en_1/in3 VDD 0.27fF
C1480 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_2/en_b 0.28fF
C1481 sky130_fd_sc_hd__clkinv_4_0/Y d_probe_1 1.70fF
C1482 d_clk_grp_1_ctrl_0 clock_v2_0/p1d_b 0.04fF
C1483 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X -0.00fF
C1484 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# -0.00fF
C1485 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C1486 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.00fF
C1487 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C1488 a_mux4_en_0/switch_5t_mux4_2/en_b a_mod_grp_ctrl_1 0.08fF
C1489 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VDD 0.14fF
C1490 a_mux4_en_0/switch_5t_mux4_3/a_300_216# VDD 0.23fF
C1491 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C1492 onebit_dac_1/v_b ota_v2_0/on 0.00fF
C1493 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# 0.13fF
C1494 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# ota_v2_0/ip 0.13fF
C1495 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# -0.09fF
C1496 a_mux4_en_0/in0 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# -0.00fF
C1497 onebit_dac_0/out VDD 1.26fF
C1498 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.01fF
C1499 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# -0.00fF
C1500 rst_n VDD 10.15fF
C1501 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# 0.04fF
C1502 a_mux4_en_1/switch_5t_mux4_0/a_300_216# VDD 0.22fF
C1503 a_mux4_en_1/in2 a_mux4_en_0/in0 0.58fF
C1504 a_mux4_en_1/in1 a_mux4_en_1/transmission_gate_3/en_b 0.03fF
C1505 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD -0.00fF
C1506 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A VDD 1.26fF
C1507 clock_v2_0/A_b d_clk_grp_1_ctrl_1 0.02fF
C1508 d_clk_grp_1_ctrl_1 clock_v2_0/B_b 0.02fF
C1509 clock_v2_0/A_b clock_v2_0/Ad_b 8.17fF
C1510 clock_v2_0/B_b clock_v2_0/Ad_b 0.94fF
C1511 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# 0.03fF
C1512 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# transmission_gate_29/out 0.53fF
C1513 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# transmission_gate_3/in 0.13fF
C1514 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# ota_v2_0/on 0.06fF
C1515 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/on -0.00fF
C1516 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VDD 0.00fF
C1517 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# 0.12fF
C1518 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980# 0.12fF
C1519 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_2/a_300_216# 0.60fF
C1520 a_mux2_en_0/in1 a_mux4_en_0/in0 0.22fF
C1521 ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p1 0.01fF
C1522 a_mux4_en_1/switch_5t_mux4_2/in a_mod_grp_ctrl_1 -0.00fF
C1523 debug a_mux4_en_1/switch_5t_mux4_3/a_300_216# 0.33fF
C1524 ota_v2_0/p2 clock_v2_0/Ad_b 1.05fF
C1525 transmission_gate_7/en transmission_gate_2/in 0.13fF
C1526 ota_v2_0/p2_b ota_v2_0/p1_b 6.65fF
C1527 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y -0.00fF
C1528 d_clk_grp_1_ctrl_1 ota_v2_0/p2 0.02fF
C1529 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.03fF
C1530 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C1531 sky130_fd_sc_hd__mux4_1_1/a_27_413# VDD 0.12fF
C1532 ota_v2_0/in ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# 0.05fF
C1533 ota_v2_0/ip ota_v2_0/on 1.37fF
C1534 transmission_gate_21/in ota_v2_0/p2 0.06fF
C1535 transmission_gate_25/in ota_v2_0/p1_b 0.47fF
C1536 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/c1_n930_n880# 0.07fF
C1537 ota_v2_0/cm ota_v2_0/ota_v2_without_cmfb_0/bias_b 0.00fF
C1538 a_mux4_en_1/switch_5t_mux4_0/en_b a_mod_grp_ctrl_0 0.26fF
C1539 transmission_gate_30/out onebit_dac_0/out -0.18fF
C1540 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in -0.00fF
C1541 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# -0.00fF
C1542 VDD m2_74560_34230# 0.06fF
C1543 clock_v2_0/A clock_v2_0/p1d 0.80fF
C1544 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# VDD 1.87fF
C1545 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.01fF
C1546 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.04fF
C1547 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# -0.06fF
C1548 a_mux4_en_0/switch_5t_mux4_0/en_b a_mux4_en_0/switch_5t_mux4_1/in 0.00fF
C1549 a_mux4_en_0/switch_5t_mux4_3/a_300_216# a_mod_grp_ctrl_1 0.04fF
C1550 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.03fF
C1551 a_mux2_en_1/switch_5t_mux2_1/en a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in -0.01fF
C1552 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# 0.07fF
C1553 debug a_mux4_en_0/switch_5t_mux4_2/en_b 0.43fF
C1554 d_clk_grp_1_ctrl_0 ota_v2_0/p1_b 0.08fF
C1555 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VDD 0.06fF
C1556 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# -0.00fF
C1557 a_mux4_en_1/switch_5t_mux4_1/in a_mux4_en_1/transmission_gate_3/en_b 0.00fF
C1558 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C1559 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0.14fF
C1560 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C1561 a_mux2_en_0/switch_5t_mux2_1/in a_mux2_en_0/switch_5t_mux2_1/en -0.02fF
C1562 a_mux4_en_1/switch_5t_mux4_0/a_300_216# a_mod_grp_ctrl_1 0.04fF
C1563 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clk 0.00fF
C1564 a_mod_grp_ctrl_0 a_probe_2 3.71fF
C1565 transmission_gate_7/en clock_v2_0/Bd 0.28fF
C1566 sky130_fd_sc_hd__mux4_1_3/a_27_413# VDD 0.07fF
C1567 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.21fF
C1568 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/p1_b 0.00fF
C1569 transmission_gate_7/en clock_v2_0/B 4.11fF
C1570 a_mux4_en_0/in2 ota_v2_0/p2 0.00fF
C1571 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.12fF
C1572 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# a_mux2_en_0/in0 0.07fF
C1573 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# -0.00fF
C1574 sky130_fd_sc_hd__mux4_1_1/a_834_97# ota_v2_0/p2_b 0.00fF
C1575 a_mux4_en_0/switch_5t_mux4_0/in a_mod_grp_ctrl_0 0.00fF
C1576 sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210# 0.03fF
C1577 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# -0.01fF
C1578 sky130_fd_sc_hd__mux4_1_2/a_27_413# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C1579 transmission_gate_2/in transmission_gate_3/in 1.29fF
C1580 ota_v2_0/in clock_v2_0/p2d_b 0.21fF
C1581 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/X 0.02fF
C1582 sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C1583 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# ota_v2_0/on 0.65fF
C1584 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C1585 ota_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.00fF
C1586 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD 0.07fF
C1587 ota_v2_0/p2_b transmission_gate_25/in 0.43fF
C1588 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# -0.21fF
C1589 a_mux2_en_1/switch_5t_mux2_1/in ota_v2_0/op 0.05fF
C1590 debug a_mux4_en_1/switch_5t_mux4_2/in 0.18fF
C1591 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.00fF
C1592 a_mux4_en_1/in1 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# 0.23fF
C1593 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_v2_0/op 0.00fF
C1594 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y -0.00fF
C1595 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/c1_n930_n880# 0.07fF
C1596 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210# 0.03fF
C1597 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.02fF
C1598 transmission_gate_29/out ota_v2_0/in 0.21fF
C1599 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A -0.00fF
C1600 onebit_dac_1/v_b comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X 0.00fF
C1601 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# 0.03fF
C1602 debug a_mux4_en_1/in3 -0.00fF
C1603 ota_v2_0/sc_cmfb_0/transmission_gate_3/out VDD 2.63fF
C1604 a_mux4_en_0/switch_5t_mux4_0/in a_mux4_en_0/in1 0.00fF
C1605 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X -0.00fF
C1606 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.06fF
C1607 d_clk_grp_1_ctrl_0 ota_v2_0/p2_b 0.18fF
C1608 sky130_fd_sc_hd__mux4_1_2/X clock_v2_0/Bd_b 0.00fF
C1609 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.13fF
C1610 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# ota_v2_0/ota_v2_without_cmfb_0/bias_b -0.00fF
C1611 a_mux4_en_1/switch_5t_mux4_3/en a_mod_grp_ctrl_0 0.12fF
C1612 rst_n clock_v2_0/p1d 0.59fF
C1613 a_mux2_en_0/in1 clock_v2_0/Ad_b 1.47fF
C1614 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# transmission_gate_3/in 0.13fF
C1615 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in -0.01fF
C1616 debug a_mux4_en_0/switch_5t_mux4_3/a_300_216# 0.38fF
C1617 a_mux4_en_1/switch_5t_mux4_0/en a_mod_grp_ctrl_0 0.29fF
C1618 a_mux4_en_0/switch_5t_mux4_3/en a_mux4_en_0/switch_5t_mux4_2/en 0.00fF
C1619 sky130_fd_sc_hd__mux4_1_3/a_750_97# ota_v2_0/p1_b 0.13fF
C1620 a_mux2_en_0/in1 transmission_gate_21/in 0.00fF
C1621 clock_v2_0/B transmission_gate_3/in 2.15fF
C1622 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out ota_v2_0/p1_b 0.01fF
C1623 a_mux4_en_1/switch_5t_mux4_3/in a_mod_grp_ctrl_0 -0.00fF
C1624 sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C1625 ota_w_test_v2_0/on ota_v2_0/p2 0.00fF
C1626 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out -0.00fF
C1627 debug a_mux4_en_1/switch_5t_mux4_0/a_300_216# 0.13fF
C1628 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# -0.00fF
C1629 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/m3_n1030_n980# 0.09fF
C1630 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_218_47# 0.00fF
C1631 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/c1_n930_n880# VDD 3.45fF
C1632 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/c1_n930_n880# -0.01fF
C1633 a_mux4_en_1/switch_5t_mux4_0/in a_mux4_en_1/transmission_gate_3/en_b 0.00fF
C1634 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# 0.17fF
C1635 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# 0.07fF
C1636 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.00fF
C1637 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/X 0.00fF
C1638 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD 0.06fF
C1639 sky130_fd_sc_hd__mux4_1_0/a_923_363# ota_v2_0/p2_b 0.02fF
C1640 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C1641 ota_w_test_v2_0/in transmission_gate_2/in 0.09fF
C1642 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C1643 ota_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/p2 0.01fF
C1644 ota_w_test_v2_0/on ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.00fF
C1645 a_mux4_en_1/in2 a_mux4_en_0/in2 0.28fF
C1646 a_mod_grp_ctrl_0 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C1647 sky130_fd_sc_hd__mux4_1_2/X VDD 1.01fF
C1648 ota_v2_0/in transmission_gate_21/out 1.71fF
C1649 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# a_mux4_en_0/in1 0.00fF
C1650 a_mux4_en_0/switch_5t_mux4_0/en_b a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C1651 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/p1d 0.01fF
C1652 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# ota_v2_0/in 0.11fF
C1653 ota_v2_0/cm ota_v2_0/sc_cmfb_0/bias_a 0.00fF
C1654 a_probe_3 VDD 4.12fF
C1655 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/Ad_b 0.00fF
C1656 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# transmission_gate_2/in 0.09fF
C1657 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y VDD 0.47fF
C1658 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.01fF
C1659 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# 0.07fF
C1660 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VDD -0.00fF
C1661 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.03fF
C1662 a_mux4_en_1/in2 a_mux4_en_0/in1 0.23fF
C1663 ota_v2_0/cm ota_v2_0/ip 0.82fF
C1664 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/c1_n260_n210# 0.03fF
C1665 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C1666 transmission_gate_7/en ota_v2_0/op 0.10fF
C1667 transmission_gate_21/in ota_v2_0/on 0.07fF
C1668 transmission_gate_31/out clock_v2_0/p2d_b 0.50fF
C1669 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_3/en_b 1.20fF
C1670 sky130_fd_sc_hd__mux4_1_2/a_27_413# VDD 0.11fF
C1671 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# 0.03fF
C1672 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_1/en_b 0.41fF
C1673 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C1674 sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/c1_n930_n880# 0.07fF
C1675 clock_v2_0/p2d_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/c1_n260_n210# 0.02fF
C1676 clock_v2_0/p2d_b sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.07fF
C1677 clock_v2_0/p1d_b transmission_gate_7/en 0.61fF
C1678 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/B_b 0.00fF
C1679 clock_v2_0/p2d transmission_gate_7/en 0.57fF
C1680 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.13fF
C1681 a_mod_grp_ctrl_0 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_2/a_113_47# -0.00fF
C1682 in i_bias_1 0.16fF
C1683 ota_v2_0/p2_b sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.00fF
C1684 a_mux4_en_0/in0 transmission_gate_9/in 0.03fF
C1685 ota_w_test_v2_0/in clock_v2_0/B 0.12fF
C1686 ota_v2_0/p2_b ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out 0.01fF
C1687 a_mux2_en_1/switch_5t_mux2_1/en a_mux2_en_1/switch_5t_mux2_1/in -0.02fF
C1688 a_mux4_en_1/switch_5t_mux4_1/en a_mux4_en_1/switch_5t_mux4_2/en -0.00fF
C1689 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.02fF
C1690 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.02fF
C1691 rst_n clock_v2_0/A 0.30fF
C1692 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# -0.00fF
C1693 transmission_gate_29/out ip 0.02fF
C1694 a_mux4_en_1/switch_5t_mux4_3/en_b VDD 1.03fF
C1695 transmission_gate_7/en clock_v2_0/Ad 0.28fF
C1696 a_mux2_en_0/in0 ota_v2_0/p2 0.06fF
C1697 transmission_gate_23/in ota_v2_0/ip 1.08fF
C1698 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# -0.12fF
C1699 ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# ota_v2_0/ota_v2_without_cmfb_0/bias_b 0.00fF
C1700 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# -0.00fF
C1701 a_mux4_en_1/switch_5t_mux4_2/in a_mux4_en_1/in3 -0.00fF
C1702 a_mux4_en_1/switch_5t_mux4_2/en_b VDD 0.99fF
C1703 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C1704 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# 0.04fF
C1705 sky130_fd_sc_hd__mux4_1_3/a_193_413# ota_v2_0/p1_b 0.04fF
C1706 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C1707 transmission_gate_2/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/m3_n1030_n980# 0.09fF
C1708 a_mux4_en_1/in0 ota_v2_0/p2 0.02fF
C1709 transmission_gate_32/out in 0.11fF
C1710 in a_mux4_en_0/in0 0.28fF
C1711 sky130_fd_sc_hd__mux4_1_0/a_247_21# clock_v2_0/B_b 0.11fF
C1712 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C1713 sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C1714 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# clock_v2_0/p2d_b 0.02fF
C1715 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C1716 ota_v2_0/sc_cmfb_0/cmc ota_v2_0/ip 0.25fF
C1717 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C1718 a_mux2_en_0/in1 ota_w_test_v2_0/on 0.37fF
C1719 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# -0.00fF
C1720 d_probe_2 VDD 6.87fF
C1721 sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# -0.06fF
C1722 a_mux2_en_1/switch_5t_mux2_0/in a_mod_grp_ctrl_0 0.02fF
C1723 clock_v2_0/A_b clock_v2_0/Bd_b 0.48fF
C1724 clock_v2_0/B_b clock_v2_0/Bd_b 8.13fF
C1725 sky130_fd_sc_hd__mux4_1_0/a_247_21# ota_v2_0/p2 0.01fF
C1726 sky130_fd_sc_hd__clkinv_4_0/Y VDD 1.01fF
C1727 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in 0.00fF
C1728 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A -0.00fF
C1729 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.03fF
C1730 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/c1_n260_n210# 0.03fF
C1731 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X -0.00fF
C1732 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C1733 a_mux4_en_1/switch_5t_mux4_1/a_300_216# a_mod_grp_ctrl_0 0.24fF
C1734 sky130_fd_sc_hd__mux4_1_2/a_1290_413# VDD 0.07fF
C1735 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# -0.00fF
C1736 sky130_fd_sc_hd__mux4_1_2/a_757_363# clock_v2_0/Ad_b 0.00fF
C1737 ota_v2_0/ota_v2_without_cmfb_0/bias_d ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# 0.01fF
C1738 transmission_gate_7/en ota_v2_0/p1_b 0.83fF
C1739 sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980# 0.09fF
C1740 a_mux2_en_1/transmission_gate_1/en_b ota_v2_0/op 0.00fF
C1741 VDD a_mux4_en_0/switch_5t_mux4_2/a_300_216# 0.22fF
C1742 a_mux2_en_0/switch_5t_mux2_0/in a_mod_grp_ctrl_0 0.02fF
C1743 ota_v2_0/p2 clock_v2_0/Bd_b 0.96fF
C1744 sky130_fd_sc_hd__mux4_1_3/a_27_413# clock_v2_0/A -0.00fF
C1745 a_mux4_en_1/switch_5t_mux4_3/en_b a_mod_grp_ctrl_1 0.08fF
C1746 clock_v2_0/B_b VDD 2.64fF
C1747 clock_v2_0/A_b VDD 2.79fF
C1748 m5_41088_30705# transmission_gate_3/in 0.27fF
C1749 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# -0.00fF
C1750 a_mux4_en_1/switch_5t_mux4_0/en_b VDD 0.96fF
C1751 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_3/a_193_47# 0.01fF
C1752 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C1753 sky130_fd_sc_hd__mux4_1_2/X d_clk_grp_2_ctrl_1 0.00fF
C1754 a_mux4_en_1/switch_5t_mux4_2/en_b a_mod_grp_ctrl_1 0.08fF
C1755 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_v2_0/sc_cmfb_0/transmission_gate_4/out -0.00fF
C1756 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.02fF
C1757 sky130_fd_sc_hd__mux4_1_0/a_750_97# clock_v2_0/B 0.00fF
C1758 sky130_fd_sc_hd__mux4_1_2/a_923_363# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.01fF
C1759 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B -0.00fF
C1760 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.01fF
C1761 ota_v2_0/p2 VDD 9.46fF
C1762 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.00fF
C1763 transmission_gate_31/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980# 0.81fF
C1764 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD 0.01fF
C1765 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/p1d 0.00fF
C1766 ota_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p1 -0.00fF
C1767 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clk 0.00fF
C1768 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y -0.00fF
C1769 comparator_v2_0/li_940_3458# ota_v2_0/on 0.00fF
C1770 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/in3 0.00fF
C1771 a_mux4_en_1/in2 a_mux4_en_1/in0 1.41fF
C1772 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.00fF
C1773 a_mux2_en_0/in1 a_mux2_en_0/in0 3.69fF
C1774 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_0/en_b 0.45fF
C1775 ota_w_test_v2_0/op clock_v2_0/Ad_b 0.45fF
C1776 a_probe_2 VDD 4.15fF
C1777 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# ota_v2_0/in 0.25fF
C1778 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# -0.09fF
C1779 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_193_413# -0.00fF
C1780 ota_v2_0/in ota_v2_0/op 1.29fF
C1781 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.21fF
C1782 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_0/a_300_216# 0.61fF
C1783 ota_v2_0/p2_b transmission_gate_7/en 0.70fF
C1784 ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p1_b 0.00fF
C1785 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.04fF
C1786 a_mux4_en_0/switch_5t_mux4_0/in VDD 0.64fF
C1787 a_mux4_en_0/switch_5t_mux4_2/a_300_216# a_mod_grp_ctrl_1 0.04fF
C1788 comparator_v2_0/li_940_818# ota_v2_0/on 0.00fF
C1789 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C1790 a_mux4_en_0/switch_5t_mux4_0/en a_mux4_en_0/switch_5t_mux4_1/en -0.00fF
C1791 clock_v2_0/p2d ota_v2_0/in 0.14fF
C1792 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD 0.00fF
C1793 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.02fF
C1794 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C1795 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C1796 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C1797 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.02fF
C1798 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X -0.01fF
C1799 sky130_fd_sc_hd__mux4_1_0/a_27_413# VDD 0.11fF
C1800 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# VDD 0.28fF
C1801 a_mux4_en_1/switch_5t_mux4_0/en_b a_mod_grp_ctrl_1 0.14fF
C1802 debug a_mux4_en_1/switch_5t_mux4_3/en_b 1.02fF
C1803 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in VDD 0.94fF
C1804 onebit_dac_1/out i_bias_2 0.24fF
C1805 transmission_gate_23/in transmission_gate_21/in 0.25fF
C1806 ota_v2_0/ip ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# 0.09fF
C1807 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# transmission_gate_2/in 0.12fF
C1808 a_mux4_en_0/in2 ota_w_test_v2_0/op 0.56fF
C1809 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# -0.03fF
C1810 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# 0.04fF
C1811 debug a_mux4_en_1/switch_5t_mux4_2/en_b 0.30fF
C1812 sky130_fd_sc_hd__mux4_1_3/a_27_47# clock_v2_0/B 0.00fF
C1813 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# ota_v2_0/on 0.13fF
C1814 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C1815 a_mux2_en_0/in1 clock_v2_0/Bd_b 0.17fF
C1816 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VDD 0.74fF
C1817 d_probe_2 d_clk_grp_2_ctrl_1 0.03fF
C1818 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# 0.04fF
C1819 a_mux4_en_1/switch_5t_mux4_3/en VDD 0.13fF
C1820 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# VDD 1.92fF
C1821 a_mux4_en_0/in2 in 0.28fF
C1822 a_mux4_en_1/switch_5t_mux4_0/en VDD -0.04fF
C1823 sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/c1_n930_n880# -0.06fF
C1824 a_mux4_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# 0.10fF
C1825 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# -0.05fF
C1826 a_mux4_en_1/switch_5t_mux4_3/in VDD 0.61fF
C1827 a_mux4_en_1/in2 VDD 6.93fF
C1828 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_439_47# 0.00fF
C1829 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# ota_v2_0/in 0.04fF
C1830 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/c1_n260_n210# 0.03fF
C1831 a_mux4_en_1/switch_5t_mux4_3/en_b a_mux4_en_1/switch_5t_mux4_3/a_300_216# -0.00fF
C1832 sky130_fd_sc_hd__mux4_1_2/a_1290_413# d_clk_grp_2_ctrl_1 0.11fF
C1833 ota_v2_0/p2_b transmission_gate_3/in 0.19fF
C1834 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VDD -0.01fF
C1835 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C1836 in a_mux4_en_0/in1 0.29fF
C1837 ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p2_b 0.05fF
C1838 a_mux4_en_0/switch_5t_mux4_0/in a_mod_grp_ctrl_1 0.00fF
C1839 ota_v2_0/op m1_86360_35183# 0.02fF
C1840 transmission_gate_29/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.03fF
C1841 a_mux2_en_0/in1 VDD 13.11fF
C1842 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A VDD 0.15fF
C1843 sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C1844 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/Bd_b 0.14fF
C1845 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y VDD 0.14fF
C1846 clock_v2_0/A_b clock_v2_0/p1d 0.72fF
C1847 clock_v2_0/B_b clock_v2_0/p1d 0.95fF
C1848 debug a_mux4_en_0/switch_5t_mux4_2/a_300_216# 0.19fF
C1849 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# -0.01fF
C1850 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# 0.07fF
C1851 a_mux4_en_0/switch_5t_mux4_1/en a_mux4_en_0/switch_5t_mux4_2/en -0.00fF
C1852 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C1853 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1854 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_2/X 0.02fF
C1855 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/p1 0.01fF
C1856 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C1857 ota_v2_0/ip clock_v2_0/p2d_b 0.88fF
C1858 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/c1_n260_n210# 0.03fF
C1859 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C1860 sky130_fd_sc_hd__mux4_1_0/a_834_97# clock_v2_0/B_b 0.01fF
C1861 sky130_fd_sc_hd__mux4_1_0/a_277_47# d_clk_grp_1_ctrl_1 0.15fF
C1862 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C1863 sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C1864 transmission_gate_31/out clock_v2_0/p1d_b 0.33fF
C1865 onebit_dac_1/out a_mux4_en_1/in1 0.14fF
C1866 sky130_fd_sc_hd__mux4_1_3/X VDD 0.82fF
C1867 a_mux4_en_0/switch_5t_mux4_0/in a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C1868 a_mux4_en_1/switch_5t_mux4_0/en_b debug 0.16fF
C1869 ota_w_test_v2_0/on ota_w_test_v2_0/op 0.91fF
C1870 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/c1_n930_n880# 0.07fF
C1871 a_mux4_en_0/switch_5t_mux4_3/en_b VDD 2.67fF
C1872 ota_v2_0/p2 clock_v2_0/p1d 2.41fF
C1873 transmission_gate_31/out clock_v2_0/p2d 0.13fF
C1874 VDD a_mux4_en_0/switch_5t_mux4_1/en_b 0.96fF
C1875 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# -0.00fF
C1876 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# -0.04fF
C1877 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210# 0.03fF
C1878 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# 0.09fF
C1879 transmission_gate_2/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/m3_n1030_n980# 0.09fF
C1880 clock_v2_0/p1d_b ip 0.95fF
C1881 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/switch_5t_mux4_2/en -0.01fF
C1882 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VDD -0.01fF
C1883 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C1884 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.00fF
C1885 sky130_fd_sc_hd__mux4_1_2/a_750_97# VDD 0.16fF
C1886 transmission_gate_29/out ota_v2_0/ip 1.29fF
C1887 a_mux4_en_1/switch_5t_mux4_3/en a_mod_grp_ctrl_1 0.07fF
C1888 a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in a_mux2_en_0/switch_5t_mux2_1/en -0.01fF
C1889 a_mux2_en_1/switch_5t_mux2_1/en a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in -0.02fF
C1890 clock_v2_0/p2d ip 0.18fF
C1891 a_mux4_en_1/switch_5t_mux4_0/en a_mod_grp_ctrl_1 0.20fF
C1892 ota_v2_0/on VDD 13.59fF
C1893 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/p2d_b 0.00fF
C1894 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.12fF
C1895 a_mod_grp_ctrl_0 a_mux4_en_1/transmission_gate_3/en_b 0.00fF
C1896 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VDD 0.00fF
C1897 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# -0.01fF
C1898 transmission_gate_32/out clock_v2_0/p2d_b 3.27fF
C1899 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C1900 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A VDD 0.25fF
C1901 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.03fF
C1902 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/cm 0.01fF
C1903 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# -0.00fF
C1904 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# 0.07fF
C1905 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/on 1.42fF
C1906 a_mux4_en_1/switch_5t_mux4_3/en_b a_mux4_en_1/switch_5t_mux4_2/in -0.00fF
C1907 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C1908 onebit_dac_1/out transmission_gate_31/out 0.01fF
C1909 ota_v2_0/p1 a_mux4_en_0/in0 0.28fF
C1910 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.02fF
C1911 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y a_mod_grp_ctrl_1 0.00fF
C1912 debug a_mux4_en_0/switch_5t_mux4_0/in 0.65fF
C1913 a_mux4_en_1/switch_5t_mux4_2/in a_mux4_en_1/switch_5t_mux4_2/en_b -0.00fF
C1914 sky130_fd_sc_hd__mux4_1_0/a_27_413# clock_v2_0/p1d 0.00fF
C1915 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C1916 a_mux4_en_0/switch_5t_mux4_2/en_b a_mux4_en_0/switch_5t_mux4_2/a_300_216# -0.00fF
C1917 onebit_dac_1/out ip 0.17fF
C1918 transmission_gate_8/in ota_v2_0/p2 0.49fF
C1919 ota_v2_0/in ota_v2_0/p2_b 0.09fF
C1920 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# -0.13fF
C1921 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# -0.13fF
C1922 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C1923 d_probe_0 d_probe_1 1.24fF
C1924 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in VDD 1.43fF
C1925 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# -0.00fF
C1926 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C1927 ota_v2_0/in transmission_gate_25/in 1.07fF
C1928 ota_v2_0/ip transmission_gate_21/out 0.10fF
C1929 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in VDD 3.49fF
C1930 a_mux2_en_0/in0 transmission_gate_9/in 0.18fF
C1931 sky130_fd_sc_hd__mux4_1_3/a_757_363# VDD 0.03fF
C1932 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.00fF
C1933 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# ota_v2_0/ip 0.35fF
C1934 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# 0.03fF
C1935 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_2/en 0.13fF
C1936 clock_v2_0/B_b clock_v2_0/A 1.08fF
C1937 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VDD 0.09fF
C1938 sky130_fd_sc_hd__mux4_1_0/a_750_97# ota_v2_0/p1_b 0.00fF
C1939 ota_w_test_v2_0/ip transmission_gate_3/in 0.08fF
C1940 clock_v2_0/A_b clock_v2_0/A 19.60fF
C1941 a_mux4_en_0/switch_5t_mux4_3/en_b a_mod_grp_ctrl_1 0.07fF
C1942 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/p2 0.01fF
C1943 a_mux2_en_1/switch_5t_mux2_0/in VDD 0.41fF
C1944 a_mux4_en_0/switch_5t_mux4_1/en_b a_mod_grp_ctrl_1 0.08fF
C1945 sky130_fd_sc_hd__clkinv_4_1/Y d_probe_2 1.71fF
C1946 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# -0.14fF
C1947 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.03fF
C1948 sky130_fd_sc_hd__mux4_1_2/a_27_413# sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.01fF
C1949 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# 0.09fF
C1950 a_mux2_en_0/in0 ota_w_test_v2_0/op 0.25fF
C1951 ota_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/sc_cmfb_0/cmc -0.01fF
C1952 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# -0.21fF
C1953 sky130_fd_sc_hd__mux4_1_2/a_757_363# clock_v2_0/Bd_b 0.01fF
C1954 a_mux4_en_1/switch_5t_mux4_1/a_300_216# VDD 0.41fF
C1955 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_4_0/Y 0.09fF
C1956 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.00fF
C1957 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# transmission_gate_3/in 0.12fF
C1958 a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in 0.00fF
C1959 a_mux4_en_0/switch_5t_mux4_1/a_300_216# a_mod_grp_ctrl_0 0.60fF
C1960 ota_v2_0/p2 clock_v2_0/A 6.35fF
C1961 sky130_fd_sc_hd__mux4_1_0/a_193_413# ota_v2_0/p1 0.00fF
C1962 debug a_mux4_en_1/switch_5t_mux4_3/en 0.11fF
C1963 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.00fF
C1964 in a_mux2_en_0/in0 0.18fF
C1965 sky130_fd_sc_hd__mux4_1_3/a_834_97# VDD 0.01fF
C1966 a_mux2_en_0/switch_5t_mux2_0/in VDD 0.40fF
C1967 a_mux4_en_1/switch_5t_mux4_0/en debug 0.13fF
C1968 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.03fF
C1969 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_3/in -0.00fF
C1970 debug a_mux4_en_1/switch_5t_mux4_3/in 1.84fF
C1971 a_mux4_en_1/in2 debug 0.00fF
C1972 ota_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/op 0.01fF
C1973 a_mux2_en_0/in1 clock_v2_0/p1d 0.81fF
C1974 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A -0.00fF
C1975 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C1976 sky130_fd_sc_hd__clkinv_4_0/Y sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C1977 in a_mux4_en_1/in0 0.22fF
C1978 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/X 0.00fF
C1979 sky130_fd_sc_hd__mux4_1_2/a_757_363# VDD 0.06fF
C1980 a_mux4_en_0/in2 a_mux4_en_0/switch_5t_mux4_3/in -0.00fF
C1981 a_mux4_en_0/in0 transmission_gate_2/in 0.58fF
C1982 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# 0.03fF
C1983 transmission_gate_32/out transmission_gate_2/in 1.60fF
C1984 sky130_fd_sc_hd__mux4_1_3/a_923_363# ota_v2_0/p1_b 0.01fF
C1985 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1986 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# 0.03fF
C1987 a_mux4_en_1/switch_5t_mux4_3/en a_mux4_en_1/switch_5t_mux4_3/a_300_216# -0.00fF
C1988 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD 0.00fF
C1989 sky130_fd_sc_hd__mux4_1_1/a_1290_413# VDD 0.07fF
C1990 ota_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/sc_cmfb_0/cmc 0.00fF
C1991 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# -0.06fF
C1992 sky130_fd_sc_hd__mux4_1_0/a_750_97# ota_v2_0/p2_b 0.15fF
C1993 clock_v2_0/p2d_b clock_v2_0/Ad_b 1.15fF
C1994 sky130_fd_sc_hd__mux4_1_0/a_27_413# clock_v2_0/A 0.00fF
C1995 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C1996 ota_w_test_v2_0/op clock_v2_0/Bd_b 0.45fF
C1997 ota_w_test_v2_0/in ota_w_test_v2_0/ip 0.60fF
C1998 comparator_v2_0/li_n2324_818# ota_v2_0/on 0.02fF
C1999 transmission_gate_32/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980# 1.63fF
C2000 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C2001 transmission_gate_21/in clock_v2_0/p2d_b 0.45fF
C2002 a_mux4_en_0/switch_5t_mux4_0/en_b VDD 1.00fF
C2003 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# 0.07fF
C2004 debug a_mux4_en_0/switch_5t_mux4_3/en_b 1.22fF
C2005 clock_v2_0/A_b rst_n 0.28fF
C2006 rst_n clock_v2_0/B_b 0.29fF
C2007 sky130_fd_sc_hd__mux4_1_2/a_750_97# d_clk_grp_2_ctrl_1 0.09fF
C2008 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980# transmission_gate_2/in 0.12fF
C2009 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X VDD 0.05fF
C2010 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# 0.07fF
C2011 debug a_mux4_en_0/switch_5t_mux4_1/en_b 0.43fF
C2012 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VDD 0.00fF
C2013 sky130_fd_sc_hd__mux4_1_3/a_247_21# VDD 0.03fF
C2014 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C2015 a_mux4_en_1/switch_5t_mux4_1/a_300_216# a_mod_grp_ctrl_1 0.04fF
C2016 ota_v2_0/p1 clock_v2_0/Ad_b 1.08fF
C2017 d_clk_grp_1_ctrl_1 ota_v2_0/p1 0.01fF
C2018 VDD transmission_gate_9/in 0.30fF
C2019 a_mux4_en_0/switch_5t_mux4_0/a_300_216# VDD 0.22fF
C2020 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/switch_5t_mux4_0/a_300_216# -0.00fF
C2021 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C2022 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/c1_n930_n880# 0.07fF
C2023 transmission_gate_21/in ota_v2_0/p1 0.07fF
C2024 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VDD -0.00fF
C2025 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# 0.14fF
C2026 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# a_mux4_en_0/in1 -0.00fF
C2027 transmission_gate_29/out transmission_gate_21/in 1.05fF
C2028 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y -0.00fF
C2029 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.02fF
C2030 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# -0.10fF
C2031 rst_n ota_v2_0/p2 0.71fF
C2032 ota_w_test_v2_0/op VDD 9.68fF
C2033 ota_v2_0/cm VDD 6.74fF
C2034 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.20fF
C2035 sky130_fd_sc_hd__mux4_1_0/a_757_363# clock_v2_0/Ad_b 0.00fF
C2036 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VDD 0.09fF
C2037 sky130_fd_sc_hd__mux4_1_2/a_923_363# clock_v2_0/p2d_b 0.02fF
C2038 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__clkinv_4_0/Y 0.00fF
C2039 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C2040 sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# -0.12fF
C2041 ota_v2_0/cm ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# 0.00fF
C2042 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/c1_n930_n880# 0.07fF
C2043 in VDD 5.01fF
C2044 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/Bd 0.00fF
C2045 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.02fF
C2046 sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/c1_n930_n880# 0.07fF
C2047 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.02fF
C2048 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/B 0.00fF
C2049 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in a_mux2_en_0/switch_5t_mux2_1/en -0.02fF
C2050 ota_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p1_b -0.01fF
C2051 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/X 0.00fF
C2052 ota_v2_0/sc_cmfb_0/transmission_gate_7/in ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.00fF
C2053 a_mux4_en_0/in2 ota_v2_0/p1 -0.02fF
C2054 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_1478_413# -0.00fF
C2055 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# 0.03fF
C2056 sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C2057 ota_v2_0/p1 sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.00fF
C2058 transmission_gate_23/in VDD 0.82fF
C2059 a_mux4_en_1/in0 a_mux4_en_1/transmission_gate_3/en_b 0.03fF
C2060 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_1/X 0.05fF
C2061 transmission_gate_7/en transmission_gate_3/in 0.19fF
C2062 a_mux4_en_1/switch_5t_mux4_3/in a_mux4_en_1/switch_5t_mux4_2/in 0.00fF
C2063 a_mux4_en_0/switch_5t_mux4_0/en_b a_mod_grp_ctrl_1 0.14fF
C2064 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_3/a_757_363# 0.01fF
C2065 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.01fF
C2066 transmission_gate_21/in transmission_gate_21/out 0.33fF
C2067 a_mux4_en_1/in2 a_mux4_en_1/switch_5t_mux4_2/in 0.05fF
C2068 debug a_mux2_en_1/switch_5t_mux2_0/in -0.00fF
C2069 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# transmission_gate_21/in 0.03fF
C2070 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/op -2.00fF
C2071 a_mux4_en_0/switch_5t_mux4_3/en_b a_mux4_en_0/switch_5t_mux4_2/en_b 0.00fF
C2072 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.01fF
C2073 ota_v2_0/ota_v2_without_cmfb_0/bias_c ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# 0.00fF
C2074 a_mux4_en_0/switch_5t_mux4_2/en_b a_mux4_en_0/switch_5t_mux4_1/en_b 0.00fF
C2075 a_mux4_en_0/switch_5t_mux4_0/a_300_216# a_mod_grp_ctrl_1 0.04fF
C2076 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD 0.20fF
C2077 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.03fF
C2078 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# 0.07fF
C2079 transmission_gate_21/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210# 0.13fF
C2080 a_mux4_en_1/in2 a_mux4_en_1/in3 0.00fF
C2081 a_mux4_en_1/switch_5t_mux4_1/a_300_216# debug 0.13fF
C2082 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210# -0.06fF
C2083 sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# 0.07fF
C2084 transmission_gate_30/out in 0.03fF
C2085 ota_v2_0/sc_cmfb_0/cmc VDD 3.53fF
C2086 sky130_fd_sc_hd__mux4_1_0/a_1290_413# ota_v2_0/p2 0.00fF
C2087 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C2088 a_mux4_en_1/in2 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# 0.36fF
C2089 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.07fF
C2090 ota_v2_0/ip ota_v2_0/op 0.68fF
C2091 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# 0.12fF
C2092 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y VDD 0.33fF
C2093 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_3/a_27_47# -0.00fF
C2094 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C2095 a_mux2_en_0/switch_5t_mux2_0/in debug -0.00fF
C2096 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VDD 0.00fF
C2097 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.03fF
C2098 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.01fF
C2099 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.01fF
C2100 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_mux4_3/en 0.12fF
C2101 sky130_fd_sc_hd__mux4_1_3/a_27_413# ota_v2_0/p2 0.00fF
C2102 onebit_dac_1/out onebit_dac_1/v_b 0.52fF
C2103 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/sc_cmfb_0/cmc 0.27fF
C2104 a_mux4_en_1/switch_5t_mux4_0/en a_mux4_en_1/switch_5t_mux4_0/a_300_216# -0.00fF
C2105 a_mux4_en_1/in2 onebit_dac_0/out 0.10fF
C2106 clock_v2_0/p2d ota_v2_0/ip 0.14fF
C2107 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C2108 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.00fF
C2109 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_1290_413# -0.00fF
C2110 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C2111 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# -0.00fF
C2112 sky130_fd_sc_hd__mux4_1_1/a_923_363# VDD 0.01fF
C2113 sky130_fd_sc_hd__mux4_1_1/a_1290_413# clock_v2_0/p1d 0.00fF
C2114 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0.12fF
C2115 ota_v2_0/sc_cmfb_0/transmission_gate_6/in ota_v2_0/p2_b 0.04fF
C2116 a_mux4_en_0/switch_5t_mux4_1/en a_mux4_en_0/switch_5t_mux4_1/in -0.00fF
C2117 sky130_fd_sc_hd__mux4_1_2/a_834_97# clock_v2_0/Ad_b 0.00fF
C2118 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.00fF
C2119 ota_v2_0/ota_v2_without_cmfb_0/bias_d ota_v2_0/ota_v2_without_cmfb_0/bias_b -0.00fF
C2120 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VDD 0.08fF
C2121 sky130_fd_sc_hd__mux4_1_1/a_1290_413# d_clk_grp_2_ctrl_1 0.09fF
C2122 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# -0.26fF
C2123 clock_v2_0/Bd clock_v2_0/Ad_b 1.23fF
C2124 a_mux2_en_0/in1 onebit_dac_0/out 0.16fF
C2125 ota_w_test_v2_0/on ota_v2_0/p1 -0.03fF
C2126 clock_v2_0/B clock_v2_0/Ad_b 0.61fF
C2127 d_clk_grp_1_ctrl_1 clock_v2_0/B 0.01fF
C2128 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.09fF
C2129 a_mux2_en_0/in1 rst_n 0.45fF
C2130 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.13fF
C2131 sky130_fd_sc_hd__mux4_1_0/a_277_47# VDD 0.13fF
C2132 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# ota_v2_0/op 0.06fF
C2133 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/p1d_b 0.15fF
C2134 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A -0.00fF
C2135 transmission_gate_32/out clock_v2_0/p1d_b 0.31fF
C2136 ota_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/p1 0.01fF
C2137 VDD a_mux4_en_1/transmission_gate_3/en_b 0.73fF
C2138 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.02fF
C2139 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# 0.03fF
C2140 a_mux4_en_0/switch_5t_mux4_2/in a_mux4_en_0/switch_5t_mux4_1/in -0.00fF
C2141 debug a_mux4_en_0/switch_5t_mux4_0/en_b 0.43fF
C2142 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.01fF
C2143 transmission_gate_32/out clock_v2_0/p2d 0.13fF
C2144 a_mux4_en_0/switch_5t_mux4_3/en_b a_mux4_en_0/switch_5t_mux4_3/a_300_216# -0.00fF
C2145 onebit_dac_1/out i_bias_1 0.15fF
C2146 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.03fF
C2147 ota_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/p2 -0.00fF
C2148 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y VDD 0.33fF
C2149 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C2150 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.01fF
C2151 debug a_mux4_en_0/switch_5t_mux4_0/a_300_216# 0.19fF
C2152 d_clk_grp_2_ctrl_0 clock_v2_0/Ad_b 0.07fF
C2153 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.03fF
C2154 ota_v2_0/in transmission_gate_7/en 0.10fF
C2155 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# 0.12fF
C2156 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_mux4_2/a_300_216# 0.24fF
C2157 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/Ad 0.00fF
C2158 sky130_fd_sc_hd__mux4_1_1/a_193_413# d_clk_grp_2_ctrl_0 0.00fF
C2159 sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/c1_n260_n210# -0.14fF
C2160 ota_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# -0.00fF
C2161 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/p1_b -0.00fF
C2162 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# a_mux2_en_0/in1 0.01fF
C2163 a_mux4_en_1/switch_5t_mux4_3/en_b a_mux4_en_1/switch_5t_mux4_2/en_b 0.00fF
C2164 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/c1_n260_n210# -0.09fF
C2165 onebit_dac_0/out ota_v2_0/on 0.16fF
C2166 clock_v2_0/p2d sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C2167 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.11fF
C2168 rst_n ota_v2_0/on 0.42fF
C2169 in clock_v2_0/p1d 1.45fF
C2170 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C2171 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/p2d_b 0.00fF
C2172 a_mux4_en_1/switch_5t_mux4_2/en VDD 0.15fF
C2173 onebit_dac_1/out transmission_gate_32/out 0.02fF
C2174 onebit_dac_1/out a_mux4_en_0/in0 0.22fF
C2175 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X -0.00fF
C2176 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C2177 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0.01fF
C2178 ota_v2_0/sc_cmfb_0/transmission_gate_9/in ota_v2_0/p1 0.01fF
C2179 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C2180 transmission_gate_8/in transmission_gate_9/in 0.61fF
C2181 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C2182 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/Ad 0.01fF
C2183 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_1/X 0.00fF
C2184 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.11fF
C2185 d_probe_0 VDD 6.56fF
C2186 a_mux2_en_0/in0 ota_v2_0/p1 0.07fF
C2187 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/c1_n260_n210# ota_v2_0/on 0.09fF
C2188 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# ota_v2_0/op 0.03fF
C2189 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# 0.13fF
C2190 a_mux4_en_0/switch_5t_mux4_1/a_300_216# VDD 0.41fF
C2191 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.00fF
C2192 a_mux4_en_1/transmission_gate_3/en_b a_mod_grp_ctrl_1 0.00fF
C2193 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C2194 ota_v2_0/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.04fF
C2195 a_mux4_en_0/switch_5t_mux4_3/in VDD 0.55fF
C2196 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# -0.00fF
C2197 ota_v2_0/p2 sky130_fd_sc_hd__mux4_1_0/a_193_47# 0.01fF
C2198 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.08fF
C2199 ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# VDD 0.28fF
C2200 ota_v2_0/p1 a_mux4_en_1/in0 0.00fF
C2201 a_mux4_en_1/switch_5t_mux4_1/in a_mux4_en_1/switch_5t_mux4_1/en_b -0.00fF
C2202 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A -0.00fF
C2203 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# 0.09fF
C2204 a_mux4_en_0/in0 ota_v2_0/p1_b -0.01fF
C2205 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.11fF
C2206 sky130_fd_sc_hd__mux4_1_3/a_247_21# clock_v2_0/A 0.01fF
C2207 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.00fF
C2208 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A -0.01fF
C2209 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# 0.03fF
C2210 ota_v2_0/sc_cmfb_0/bias_a ota_v2_0/p2_b -0.00fF
C2211 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y VDD -0.00fF
C2212 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VDD 0.06fF
C2213 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.01fF
C2214 ota_w_test_v2_0/on clock_v2_0/Bd 0.64fF
C2215 clock_v2_0/p2d_b clock_v2_0/Bd_b 2.96fF
C2216 clock_v2_0/p2d sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/c1_n930_n880# 0.09fF
C2217 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# -0.13fF
C2218 sky130_fd_sc_hd__mux4_1_1/a_247_21# clock_v2_0/Ad 0.01fF
C2219 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_923_363# 0.01fF
C2220 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# ota_v2_0/ip 0.04fF
C2221 clock_v2_0/p1d_b clock_v2_0/Ad_b 2.74fF
C2222 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# ota_v2_0/in 0.03fF
C2223 a_mux4_en_1/switch_5t_mux4_2/en a_mod_grp_ctrl_1 0.08fF
C2224 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y -0.00fF
C2225 sky130_fd_sc_hd__mux4_1_1/a_193_413# clock_v2_0/p1d_b 0.07fF
C2226 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_1/a_1290_413# 0.00fF
C2227 ota_v2_0/ip ota_v2_0/p2_b 0.16fF
C2228 clock_v2_0/p2d clock_v2_0/Ad_b 1.46fF
C2229 clock_v2_0/p1d_b transmission_gate_21/in 0.24fF
C2230 a_mux2_en_0/in0 transmission_gate_21/out 0.16fF
C2231 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# 0.03fF
C2232 ota_v2_0/p1 clock_v2_0/Bd_b 1.77fF
C2233 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C2234 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VDD -0.00fF
C2235 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C2236 d_probe_1 sky130_fd_sc_hd__clkinv_4_3/Y 0.08fF
C2237 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C2238 sky130_fd_sc_hd__mux4_1_1/a_193_413# clock_v2_0/p2d 0.00fF
C2239 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/c1_n930_n880# 0.07fF
C2240 sky130_fd_sc_hd__mux4_1_3/a_668_97# VDD 0.00fF
C2241 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.03fF
C2242 clock_v2_0/p2d transmission_gate_21/in 0.49fF
C2243 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210# ota_v2_0/op 0.03fF
C2244 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# ota_v2_0/ota_v2_without_cmfb_0/bias_b 0.00fF
C2245 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/Ad_b 0.00fF
C2246 sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C2247 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/c1_n260_n210# 0.02fF
C2248 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980# transmission_gate_2/in 0.09fF
C2249 a_mux4_en_0/switch_5t_mux4_1/a_300_216# a_mod_grp_ctrl_1 0.04fF
C2250 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.00fF
C2251 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_v2_0/ota_v2_without_cmfb_0/bias_b -0.00fF
C2252 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C2253 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C2254 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C2255 clock_v2_0/Ad clock_v2_0/Ad_b 19.78fF
C2256 a_mux2_en_0/in0 transmission_gate_2/in -13.49fF
C2257 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# 0.04fF
C2258 clock_v2_0/p2d_b VDD 11.34fF
C2259 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.07fF
C2260 clock_v2_0/p2d sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# 0.09fF
C2261 sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# 0.13fF
C2262 clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y VDD 0.13fF
C2263 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# 0.25fF
C2264 debug a_mux4_en_1/transmission_gate_3/en_b -0.01fF
C2265 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.03fF
C2266 a_mux4_en_0/in0 ota_v2_0/p2_b 0.07fF
C2267 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C2268 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A -0.00fF
C2269 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# -0.01fF
C2270 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# 0.07fF
C2271 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_0/a_113_47# a_mux4_en_0/switch_5t_mux4_3/en_b -0.00fF
C2272 ota_v2_0/p1 VDD 13.84fF
C2273 sky130_fd_sc_hd__mux4_1_1/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C2274 clock_v2_0/A_b clock_v2_0/B_b 0.92fF
C2275 ota_v2_0/sc_cmfb_0/transmission_gate_3/out ota_v2_0/on -0.01fF
C2276 transmission_gate_29/out VDD 0.66fF
C2277 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# 0.07fF
C2278 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# 0.07fF
C2279 sky130_fd_sc_hd__mux4_1_0/a_757_363# VDD 0.09fF
C2280 transmission_gate_31/out transmission_gate_3/in 1.55fF
C2281 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.00fF
C2282 in a_mux4_en_1/in3 0.03fF
C2283 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VDD -0.00fF
C2284 a_mux2_en_0/in0 clock_v2_0/Bd 0.19fF
C2285 clock_v2_0/A_b ota_v2_0/p2 1.76fF
C2286 ota_v2_0/p2 clock_v2_0/B_b 1.43fF
C2287 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/a_1478_413# -0.00fF
C2288 transmission_gate_30/out clock_v2_0/p2d_b 0.32fF
C2289 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# ota_v2_0/ota_v2_without_cmfb_0/bias_b 0.02fF
C2290 a_mux4_en_1/switch_5t_mux4_3/en a_mux4_en_1/switch_5t_mux4_3/en_b 0.00fF
C2291 a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# 0.07fF
C2292 a_mux4_en_1/switch_5t_mux4_1/en a_mux4_en_1/switch_5t_mux4_1/en_b -0.00fF
C2293 debug a_mux4_en_1/switch_5t_mux4_2/en 0.12fF
C2294 ota_v2_0/p1_b clock_v2_0/Ad_b 1.14fF
C2295 sky130_fd_sc_hd__mux4_1_0/a_27_47# VDD 0.01fF
C2296 ota_v2_0/cm rst_n 0.94fF
C2297 d_clk_grp_1_ctrl_1 ota_v2_0/p1_b 0.13fF
C2298 sky130_fd_sc_hd__mux4_1_0/a_193_413# ota_v2_0/p2_b 0.07fF
C2299 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C2300 a_mux4_en_1/switch_5t_mux4_3/in a_mux4_en_1/switch_5t_mux4_3/en_b 0.00fF
C2301 transmission_gate_21/in ota_v2_0/p1_b 0.05fF
C2302 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# 0.03fF
C2303 onebit_dac_1/out a_mux4_en_0/in2 0.23fF
C2304 in onebit_dac_0/out 0.17fF
C2305 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.00fF
C2306 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# -0.00fF
C2307 sky130_fd_sc_hd__mux4_1_3/a_1478_413# VDD 0.08fF
C2308 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.00fF
C2309 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C2310 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_w_test_v2_0/ip 0.09fF
C2311 transmission_gate_30/out transmission_gate_29/out 0.41fF
C2312 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C2313 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.00fF
C2314 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.04fF
C2315 transmission_gate_21/out VDD 0.80fF
C2316 debug a_mux4_en_0/switch_5t_mux4_1/a_300_216# 0.19fF
C2317 a_mod_grp_ctrl_0 a_mux2_en_0/switch_5t_mux2_1/en 0.13fF
C2318 onebit_dac_1/out a_mux4_en_0/in1 0.25fF
C2319 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.06fF
C2320 sky130_fd_sc_hd__mux4_1_0/a_247_21# clock_v2_0/B 0.01fF
C2321 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# 0.07fF
C2322 a_mux4_en_0/switch_5t_mux4_3/en VDD 0.13fF
C2323 debug a_mux4_en_0/switch_5t_mux4_3/in 2.22fF
C2324 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00fF
C2325 a_mux2_en_1/switch_5t_mux2_1/en a_mod_grp_ctrl_0 0.13fF
C2326 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C2327 a_mux4_en_1/switch_5t_mux4_2/en_b a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C2328 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C2329 transmission_gate_2/in VDD 3.39fF
C2330 sky130_fd_sc_hd__mux4_1_2/a_834_97# clock_v2_0/Bd_b 0.01fF
C2331 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.03fF
C2332 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.02fF
C2333 a_mux4_en_0/in2 ota_v2_0/p1_b -0.02fF
C2334 clock_v2_0/B clock_v2_0/Bd_b 4.77fF
C2335 clock_v2_0/Bd clock_v2_0/Bd_b 19.82fF
C2336 ota_w_test_v2_0/op m2_74560_34230# 0.29fF
C2337 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# ota_v2_0/in 0.32fF
C2338 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y -0.00fF
C2339 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C2340 sky130_fd_sc_hd__mux4_1_3/a_1290_413# ota_v2_0/p1_b -0.00fF
C2341 ota_v2_0/op comparator_v2_0/li_940_3458# 0.00fF
C2342 a_mux4_en_0/in2 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.07fF
C2343 ota_v2_0/in m1_86360_35183# 0.00fF
C2344 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A -0.00fF
C2345 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C2346 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/Ad_b 0.01fF
C2347 sky130_fd_sc_hd__mux4_1_0/a_27_413# ota_v2_0/p2 0.01fF
C2348 ota_w_test_v2_0/on clock_v2_0/Ad 0.57fF
C2349 a_mux4_en_0/switch_5t_mux4_1/en a_mod_grp_ctrl_0 0.13fF
C2350 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C2351 transmission_gate_30/out transmission_gate_21/out 1.16fF
C2352 ota_v2_0/p2_b clock_v2_0/Ad_b 1.06fF
C2353 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# VDD 1.86fF
C2354 d_clk_grp_1_ctrl_1 ota_v2_0/p2_b 0.13fF
C2355 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C2356 ota_v2_0/p2 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in 0.01fF
C2357 a_mux4_en_1/switch_5t_mux4_2/in a_mux4_en_1/transmission_gate_3/en_b 0.00fF
C2358 transmission_gate_21/in ota_v2_0/p2_b 0.05fF
C2359 ota_v2_0/sc_cmfb_0/transmission_gate_4/out VDD 0.53fF
C2360 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/switch_5t_mux4_0/en -0.02fF
C2361 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C2362 sky130_fd_sc_hd__mux4_1_2/a_834_97# VDD 0.01fF
C2363 sky130_fd_sc_hd__mux4_1_1/a_757_363# clock_v2_0/p2d_b 0.00fF
C2364 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# 0.13fF
C2365 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C2366 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# 0.03fF
C2367 clock_v2_0/p2d_b clock_v2_0/p1d 0.81fF
C2368 transmission_gate_21/in transmission_gate_25/in 0.50fF
C2369 d_clk_grp_2_ctrl_0 clock_v2_0/Bd_b 0.14fF
C2370 clock_v2_0/Bd VDD 2.23fF
C2371 comparator_v2_0/li_940_818# ota_v2_0/op 0.00fF
C2372 sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/c1_n930_n880# 0.07fF
C2373 clock_v2_0/B VDD 2.70fF
C2374 a_mux4_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# 0.19fF
C2375 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# -0.04fF
C2376 a_mux4_en_1/in3 a_mux4_en_1/transmission_gate_3/en_b -0.00fF
C2377 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__clkinv_4_0/Y 0.02fF
C2378 clock_v2_0/p2d_b d_clk_grp_2_ctrl_1 0.13fF
C2379 a_mux4_en_0/switch_5t_mux4_2/in a_mod_grp_ctrl_0 0.00fF
C2380 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# ota_v2_0/ip 0.09fF
C2381 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# 0.09fF
C2382 a_mux4_en_1/switch_5t_mux4_2/a_300_216# VDD 0.22fF
C2383 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X -0.00fF
C2384 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C2385 ota_v2_0/p1 clock_v2_0/p1d 8.74fF
C2386 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# -0.06fF
C2387 a_mux4_en_0/switch_5t_mux4_3/en a_mod_grp_ctrl_1 0.07fF
C2388 d_clk_grp_1_ctrl_0 d_probe_1 0.15fF
C2389 d_clk_grp_1_ctrl_0 clock_v2_0/Ad_b 0.03fF
C2390 d_probe_3 VDD 7.02fF
C2391 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD 0.07fF
C2392 d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 3.05fF
C2393 transmission_gate_29/out clock_v2_0/p1d 0.15fF
C2394 a_mux4_en_1/switch_5t_mux4_0/en_b a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C2395 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# ota_v2_0/on 0.03fF
C2396 a_mux4_en_1/switch_5t_mux4_3/en_b a_mux4_en_1/sky130_fd_sc_hd__nand2_1_0/a_113_47# -0.00fF
C2397 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VDD 0.07fF
C2398 sky130_fd_sc_hd__mux4_1_2/a_27_47# VDD 0.01fF
C2399 clock_v2_0/p1d_b sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.05fF
C2400 sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.03fF
C2401 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.00fF
C2402 a_mux4_en_1/switch_5t_mux4_2/in a_mux4_en_1/switch_5t_mux4_2/en 0.00fF
C2403 a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in a_mod_grp_ctrl_0 0.01fF
C2404 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.00fF
C2405 d_clk_grp_2_ctrl_0 VDD 6.77fF
C2406 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# 0.01fF
C2407 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# 0.03fF
C2408 clock_v2_0/p1d_b a_mux2_en_0/in0 0.73fF
C2409 a_mux2_en_0/in1 ota_v2_0/p2 0.06fF
C2410 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C2411 clock_v2_0/A_b sky130_fd_sc_hd__mux4_1_3/X 0.00fF
C2412 ota_w_test_v2_0/on ota_v2_0/p1_b -0.01fF
C2413 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B VDD 0.00fF
C2414 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.11fF
C2415 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VDD 0.00fF
C2416 sky130_fd_sc_hd__mux4_1_3/a_277_47# VDD 0.08fF
C2417 sky130_fd_sc_hd__mux4_1_2/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.05fF
C2418 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/c1_n260_n210# 0.13fF
C2419 ota_v2_0/sc_cmfb_0/transmission_gate_8/in ota_v2_0/p1_b 0.00fF
C2420 a_mux4_en_1/in2 a_mux4_en_0/switch_5t_mux4_0/in 0.08fF
C2421 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/Ad -0.00fF
C2422 a_mux2_en_0/switch_5t_mux2_1/in a_mod_grp_ctrl_0 -0.00fF
C2423 a_mux4_en_1/in1 ip 0.18fF
C2424 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# 0.07fF
C2425 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# -0.21fF
C2426 a_mux2_en_0/in0 clock_v2_0/Ad 0.23fF
C2427 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# -0.10fF
C2428 sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.00fF
C2429 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X -0.00fF
C2430 transmission_gate_8/in ota_v2_0/p1 0.52fF
C2431 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# 0.03fF
C2432 transmission_gate_21/out clock_v2_0/p1d 0.18fF
C2433 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.02fF
C2434 onebit_dac_1/out a_mux2_en_0/in0 0.41fF
C2435 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C2436 a_mux4_en_1/switch_5t_mux4_2/a_300_216# a_mod_grp_ctrl_1 0.04fF
C2437 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0.00fF
C2438 a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/c1_n930_n880# 0.07fF
C2439 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# 0.03fF
C2440 ota_v2_0/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.03fF
C2441 ota_v2_0/p2 ota_v2_0/on 0.08fF
C2442 m5_41088_30705# VSS 2.80fF $ **FLOATING
C2443 m2_74560_34230# VSS 0.14fF $ **FLOATING
C2444 m2_72825_34855# VSS 0.11fF $ **FLOATING
C2445 m1_86360_35183# VSS 0.13fF $ **FLOATING
C2446 transmission_gate_30/out VSS -5.50fF
C2447 ip VSS 79.30fF
C2448 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# VSS 0.63fF
C2449 sky130_fd_pr__cap_mim_m3_1_CGPBWM_17/m3_n1030_n980# VSS 2.79fF
C2450 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# VSS 0.63fF
C2451 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# VSS 2.79fF
C2452 sky130_fd_pr__cap_mim_m3_1_CGPBWM_36/m3_n1030_n980# VSS 2.79fF
C2453 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# VSS 2.79fF
C2454 sky130_fd_pr__cap_mim_m3_1_CGPBWM_35/m3_n1030_n980# VSS 2.79fF
C2455 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# VSS 2.79fF
C2456 comparator_v2_0/li_940_3458# VSS -1566.64fF
C2457 comparator_v2_0/li_940_818# VSS -2215.58fF
C2458 ota_v2_0/on VSS -321.94fF
C2459 comparator_v2_0/li_n2324_818# VSS -3688.45fF
C2460 ota_v2_0/op VSS -402.32fF
C2461 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A VSS -3.23fF
C2462 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A VSS -131.69fF
C2463 ota_v2_0/p1_b VSS 490.77fF
C2464 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# VSS 0.15fF
C2465 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# VSS 0.15fF
C2466 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X VSS 43.25fF
C2467 comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.06fF
C2468 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X VSS 23.78fF
C2469 comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.06fF
C2470 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# VSS 2.79fF
C2471 sky130_fd_pr__cap_mim_m3_1_CGPBWM_23/m3_n1030_n980# VSS 2.79fF
C2472 sky130_fd_pr__cap_mim_m3_1_CGPBWM_12/m3_n1030_n980# VSS 2.79fF
C2473 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# VSS 4.59fF
C2474 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# VSS 3.91fF
C2475 sky130_fd_pr__cap_mim_m3_1_CGPBWM_22/m3_n1030_n980# VSS 2.79fF
C2476 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/c1_n930_n880# VSS 0.03fF
C2477 sky130_fd_pr__cap_mim_m3_1_CGPBWM_11/m3_n1030_n980# VSS 2.79fF
C2478 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# VSS 2.79fF
C2479 sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/c1_n930_n880# VSS 4.57fF
C2480 sky130_fd_pr__cap_mim_m3_1_CGPBWM_21/m3_n1030_n980# VSS 3.91fF
C2481 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# VSS 2.79fF
C2482 sky130_fd_pr__cap_mim_m3_1_CGPBWM_20/m3_n1030_n980# VSS 2.79fF
C2483 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# VSS 2.79fF
C2484 sky130_fd_pr__cap_mim_m3_1_CGPBWM_30/m3_n1030_n980# VSS 2.79fF
C2485 a_mux4_en_1/switch_5t_mux4_2/a_300_216# VSS 3.07fF
C2486 a_mux4_en_1/switch_5t_mux4_1/en VSS 9.03fF
C2487 a_mux4_en_1/switch_5t_mux4_1/a_300_216# VSS 2.89fF
C2488 a_mux4_en_1/switch_5t_mux4_0/a_300_216# VSS 2.86fF
C2489 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y VSS 41.77fF
C2490 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y VSS 14.40fF
C2491 a_mux4_en_1/switch_5t_mux4_0/en_b VSS 16.44fF
C2492 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS -0.00fF
C2493 a_mux4_en_1/switch_5t_mux4_1/en_b VSS 15.98fF
C2494 a_mux4_en_1/switch_5t_mux4_3/in VSS 8.05fF
C2495 a_mux4_en_1/in3 VSS 1.44fF
C2496 a_mux4_en_1/switch_5t_mux4_2/in VSS 3.70fF
C2497 a_mux4_en_1/transmission_gate_3/en_b VSS -3.70fF
C2498 a_mux4_en_1/switch_5t_mux4_1/in VSS 2.81fF
C2499 a_mux4_en_1/switch_5t_mux4_0/in VSS 3.59fF
C2500 a_mux4_en_1/switch_5t_mux4_3/en VSS 5.03fF
C2501 a_mux4_en_1/switch_5t_mux4_3/en_b VSS 7.15fF
C2502 a_mux4_en_1/switch_5t_mux4_2/en VSS 10.22fF
C2503 a_mux4_en_1/switch_5t_mux4_2/en_b VSS 12.59fF
C2504 a_mux4_en_1/switch_5t_mux4_0/en VSS 4.74fF
C2505 a_probe_3 VSS 45.76fF
C2506 a_mux4_en_1/switch_5t_mux4_3/a_300_216# VSS 8.49fF
C2507 a_mux4_en_0/switch_5t_mux4_2/a_300_216# VSS 4.53fF
C2508 a_mux4_en_0/switch_5t_mux4_1/en VSS 9.03fF
C2509 a_mux4_en_0/switch_5t_mux4_1/a_300_216# VSS 4.53fF
C2510 a_mux4_en_0/switch_5t_mux4_0/a_300_216# VSS 3.14fF
C2511 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y VSS 41.77fF
C2512 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y VSS 14.40fF
C2513 a_mux4_en_0/switch_5t_mux4_0/en_b VSS 16.51fF
C2514 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS -0.00fF
C2515 a_mux4_en_0/switch_5t_mux4_1/en_b VSS 16.41fF
C2516 a_mod_grp_ctrl_1 VSS 113.84fF
C2517 debug VSS 129.31fF
C2518 a_mux4_en_0/switch_5t_mux4_3/in VSS 9.27fF
C2519 a_mux4_en_0/in3 VSS 1.44fF
C2520 a_mux4_en_0/switch_5t_mux4_2/in VSS 5.32fF
C2521 a_mux4_en_0/transmission_gate_3/en_b VSS -3.70fF
C2522 a_mux4_en_0/switch_5t_mux4_1/in VSS 4.41fF
C2523 a_mux4_en_0/switch_5t_mux4_0/in VSS 3.78fF
C2524 a_mux4_en_0/switch_5t_mux4_3/en VSS 5.11fF
C2525 a_mux4_en_0/switch_5t_mux4_3/en_b VSS 7.48fF
C2526 a_mux4_en_0/switch_5t_mux4_2/en VSS 10.10fF
C2527 a_mux4_en_0/switch_5t_mux4_2/en_b VSS 12.59fF
C2528 a_mux4_en_0/switch_5t_mux4_0/en VSS 4.73fF
C2529 a_probe_2 VSS 46.50fF
C2530 a_mux4_en_0/switch_5t_mux4_3/a_300_216# VSS 9.79fF
C2531 transmission_gate_8/in VSS 7.29fF
C2532 transmission_gate_2/in VSS 46.07fF
C2533 transmission_gate_3/in VSS 23.08fF
C2534 transmission_gate_9/in VSS -0.93fF
C2535 ota_w_test_v2_0/ip VSS -54.00fF
C2536 sky130_fd_pr__cap_mim_m3_1_CGPBWM_6/m3_n1030_n980# VSS 2.79fF
C2537 clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y VSS 29.20fF
C2538 clk VSS 26.54fF
C2539 clock_v2_0/p1d VSS 83.49fF
C2540 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_10/a_110_47# VSS 1.28fF
C2541 clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B VSS 19.01fF
C2542 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y VSS 21.31fF
C2543 clock_v2_0/Bd_b VSS 77.44fF
C2544 clock_v2_0/Ad_b VSS 74.46fF
C2545 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S VSS -2.96fF
C2546 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/X VSS 22.21fF
C2547 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_439_47# VSS 0.00fF
C2548 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_218_47# VSS 0.00fF
C2549 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21# VSS 0.16fF
C2550 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# VSS 0.11fF
C2551 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B VSS 38.37fF
C2552 clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y VSS 20.80fF
C2553 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A VSS 32.40fF
C2554 clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A VSS 28.71fF
C2555 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS 8.67fF
C2556 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# VSS 0.10fF
C2557 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# VSS 0.18fF
C2558 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# VSS 0.18fF
C2559 clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y VSS 27.29fF
C2560 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A VSS 21.60fF
C2561 clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A VSS 19.30fF
C2562 clock_v2_0/sky130_fd_sc_hd__nand2_1_2/B VSS 10.42fF
C2563 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS 8.05fF
C2564 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# VSS 0.10fF
C2565 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# VSS 0.18fF
C2566 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# VSS 0.18fF
C2567 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS 25.52fF
C2568 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# VSS 0.10fF
C2569 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# VSS 0.18fF
C2570 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# VSS 0.18fF
C2571 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS 21.56fF
C2572 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# VSS 0.10fF
C2573 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# VSS 0.18fF
C2574 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# VSS 0.18fF
C2575 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y VSS 19.50fF
C2576 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_9/a_110_47# VSS 1.28fF
C2577 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A VSS 32.94fF
C2578 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/B VSS 12.62fF
C2579 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS 20.02fF
C2580 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# VSS 0.10fF
C2581 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# VSS 0.18fF
C2582 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# VSS 0.18fF
C2583 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS 23.77fF
C2584 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# VSS 0.10fF
C2585 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# VSS 0.18fF
C2586 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# VSS 0.18fF
C2587 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS 9.64fF
C2588 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# VSS 0.10fF
C2589 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# VSS 0.18fF
C2590 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# VSS 0.18fF
C2591 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS 19.34fF
C2592 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS 26.12fF
C2593 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# VSS 0.10fF
C2594 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# VSS 0.18fF
C2595 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# VSS 0.18fF
C2596 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS 14.09fF
C2597 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# VSS 0.10fF
C2598 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# VSS 0.18fF
C2599 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# VSS 0.18fF
C2600 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_8/a_110_47# VSS 1.28fF
C2601 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A VSS 27.90fF
C2602 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS 20.17fF
C2603 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# VSS 0.10fF
C2604 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# VSS 0.18fF
C2605 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# VSS 0.18fF
C2606 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS 23.06fF
C2607 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# VSS 0.10fF
C2608 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# VSS 0.18fF
C2609 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# VSS 0.18fF
C2610 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS 20.10fF
C2611 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# VSS 0.10fF
C2612 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# VSS 0.18fF
C2613 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# VSS 0.18fF
C2614 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# VSS 0.10fF
C2615 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# VSS 0.18fF
C2616 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# VSS 0.18fF
C2617 clock_v2_0/A VSS 128.64fF
C2618 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# VSS 1.28fF
C2619 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS 9.14fF
C2620 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# VSS 0.10fF
C2621 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# VSS 0.18fF
C2622 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# VSS 0.18fF
C2623 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS 25.49fF
C2624 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# VSS 0.10fF
C2625 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# VSS 0.18fF
C2626 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# VSS 0.18fF
C2627 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS 20.06fF
C2628 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# VSS 0.10fF
C2629 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# VSS 0.18fF
C2630 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# VSS 0.18fF
C2631 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS 13.27fF
C2632 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# VSS 0.10fF
C2633 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# VSS 0.18fF
C2634 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# VSS 0.18fF
C2635 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS 15.71fF
C2636 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# VSS 0.10fF
C2637 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# VSS 0.18fF
C2638 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# VSS 0.18fF
C2639 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS 14.89fF
C2640 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# VSS 0.10fF
C2641 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# VSS 0.18fF
C2642 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# VSS 0.18fF
C2643 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS 19.88fF
C2644 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# VSS 0.10fF
C2645 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# VSS 0.18fF
C2646 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# VSS 0.18fF
C2647 clock_v2_0/A_b VSS 24.28fF
C2648 clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y VSS 19.50fF
C2649 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_6/a_110_47# VSS 1.28fF
C2650 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS 31.10fF
C2651 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS 23.44fF
C2652 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# VSS 0.10fF
C2653 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# VSS 0.18fF
C2654 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# VSS 0.18fF
C2655 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS 10.79fF
C2656 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS 4.15fF
C2657 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# VSS 0.10fF
C2658 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# VSS 0.18fF
C2659 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# VSS 0.18fF
C2660 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS 14.02fF
C2661 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS 15.02fF
C2662 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# VSS 0.10fF
C2663 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# VSS 0.18fF
C2664 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# VSS 0.18fF
C2665 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS 41.04fF
C2666 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# VSS 0.10fF
C2667 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# VSS 0.18fF
C2668 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# VSS 0.18fF
C2669 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# VSS 0.10fF
C2670 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# VSS 0.18fF
C2671 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# VSS 0.18fF
C2672 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS 15.97fF
C2673 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS 14.02fF
C2674 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# VSS 0.10fF
C2675 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# VSS 0.18fF
C2676 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# VSS 0.18fF
C2677 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS 20.25fF
C2678 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# VSS 0.10fF
C2679 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# VSS 0.18fF
C2680 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# VSS 0.18fF
C2681 clock_v2_0/Ad VSS 62.74fF
C2682 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_5/a_110_47# VSS 1.28fF
C2683 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# VSS 0.10fF
C2684 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# VSS 0.18fF
C2685 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# VSS 0.18fF
C2686 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS 39.79fF
C2687 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# VSS 0.10fF
C2688 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# VSS 0.18fF
C2689 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# VSS 0.18fF
C2690 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS 20.08fF
C2691 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# VSS 0.10fF
C2692 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# VSS 0.18fF
C2693 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# VSS 0.18fF
C2694 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS 9.17fF
C2695 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# VSS 0.10fF
C2696 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# VSS 0.18fF
C2697 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# VSS 0.18fF
C2698 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B VSS 37.80fF
C2699 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# VSS 0.17fF
C2700 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# VSS 0.31fF
C2701 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# VSS 0.18fF
C2702 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# VSS 0.10fF
C2703 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# VSS 0.18fF
C2704 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# VSS 0.18fF
C2705 clock_v2_0/sky130_fd_sc_hd__nand2_1_0/A VSS 17.43fF
C2706 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS 14.10fF
C2707 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# VSS 0.10fF
C2708 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# VSS 0.18fF
C2709 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# VSS 0.18fF
C2710 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS 19.92fF
C2711 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# VSS 0.10fF
C2712 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# VSS 0.18fF
C2713 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# VSS 0.18fF
C2714 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# VSS 0.10fF
C2715 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# VSS 0.18fF
C2716 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# VSS 0.18fF
C2717 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_4/a_110_47# VSS 1.28fF
C2718 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS 14.88fF
C2719 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# VSS 0.10fF
C2720 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# VSS 0.18fF
C2721 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# VSS 0.18fF
C2722 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS 23.36fF
C2723 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# VSS 0.10fF
C2724 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# VSS 0.18fF
C2725 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# VSS 0.18fF
C2726 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS 15.70fF
C2727 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# VSS 0.10fF
C2728 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# VSS 0.18fF
C2729 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# VSS 0.18fF
C2730 VDD VSS -37429.17fF
C2731 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS 10.93fF
C2732 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# VSS 0.10fF
C2733 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# VSS 0.18fF
C2734 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# VSS 0.18fF
C2735 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS 19.62fF
C2736 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# VSS 0.10fF
C2737 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# VSS 0.18fF
C2738 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# VSS 0.18fF
C2739 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# VSS 0.10fF
C2740 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# VSS 0.18fF
C2741 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# VSS 0.49fF
C2742 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS 15.70fF
C2743 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# VSS 0.10fF
C2744 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# VSS 0.18fF
C2745 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# VSS 0.18fF
C2746 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS 14.06fF
C2747 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# VSS 0.10fF
C2748 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# VSS 0.18fF
C2749 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# VSS 0.18fF
C2750 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS 18.40fF
C2751 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# VSS 0.10fF
C2752 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# VSS 0.18fF
C2753 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# VSS 0.18fF
C2754 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS 20.91fF
C2755 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# VSS 0.10fF
C2756 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# VSS 0.18fF
C2757 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# VSS 0.18fF
C2758 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VSS 1.28fF
C2759 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS 20.23fF
C2760 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# VSS 0.10fF
C2761 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# VSS 0.18fF
C2762 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# VSS 0.18fF
C2763 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS 14.02fF
C2764 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS 15.02fF
C2765 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# VSS 0.10fF
C2766 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# VSS 0.18fF
C2767 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# VSS 0.18fF
C2768 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS 11.17fF
C2769 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS 6.68fF
C2770 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# VSS 0.10fF
C2771 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# VSS 0.18fF
C2772 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# VSS 0.18fF
C2773 clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y VSS 1.34fF
C2774 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# VSS 0.10fF
C2775 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# VSS 0.18fF
C2776 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# VSS 0.18fF
C2777 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# VSS 0.10fF
C2778 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# VSS 0.18fF
C2779 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# VSS 0.18fF
C2780 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS 15.73fF
C2781 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS 19.85fF
C2782 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# VSS 0.10fF
C2783 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# VSS 0.18fF
C2784 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# VSS 0.18fF
C2785 clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y VSS 34.58fF
C2786 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# VSS 0.10fF
C2787 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# VSS 0.18fF
C2788 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# VSS 0.18fF
C2789 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# VSS 0.10fF
C2790 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# VSS 0.18fF
C2791 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# VSS 0.18fF
C2792 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS 9.06fF
C2793 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# VSS 0.10fF
C2794 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# VSS 0.18fF
C2795 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# VSS 0.18fF
C2796 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS 25.87fF
C2797 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS 20.02fF
C2798 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# VSS 0.10fF
C2799 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# VSS 0.18fF
C2800 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# VSS 0.18fF
C2801 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS 38.55fF
C2802 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# VSS 0.10fF
C2803 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# VSS 0.18fF
C2804 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# VSS 0.18fF
C2805 clock_v2_0/B_b VSS 56.90fF
C2806 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y VSS 37.82fF
C2807 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_2/a_110_47# VSS 1.28fF
C2808 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS 14.10fF
C2809 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# VSS 0.10fF
C2810 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# VSS 0.18fF
C2811 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# VSS 0.18fF
C2812 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# VSS 0.10fF
C2813 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# VSS 0.18fF
C2814 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# VSS 0.24fF
C2815 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS 14.09fF
C2816 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# VSS 0.10fF
C2817 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# VSS 0.18fF
C2818 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# VSS 0.18fF
C2819 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B VSS 50.37fF
C2820 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VSS 0.16fF
C2821 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VSS 0.57fF
C2822 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# VSS 0.18fF
C2823 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS 19.55fF
C2824 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS 15.56fF
C2825 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# VSS 0.10fF
C2826 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# VSS 0.18fF
C2827 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# VSS 0.18fF
C2828 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS 25.49fF
C2829 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# VSS 0.10fF
C2830 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# VSS 0.18fF
C2831 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# VSS 0.18fF
C2832 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS 47.14fF
C2833 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# VSS 0.10fF
C2834 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# VSS 0.18fF
C2835 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# VSS 0.18fF
C2836 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS 9.16fF
C2837 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# VSS 0.10fF
C2838 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# VSS 0.18fF
C2839 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# VSS 0.18fF
C2840 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS 23.33fF
C2841 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# VSS 0.10fF
C2842 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# VSS 0.18fF
C2843 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# VSS 0.18fF
C2844 clock_v2_0/Bd VSS 50.99fF
C2845 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_1/a_110_47# VSS 1.28fF
C2846 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS 35.19fF
C2847 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# VSS 0.10fF
C2848 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# VSS 0.18fF
C2849 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# VSS 0.18fF
C2850 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS 15.70fF
C2851 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# VSS 0.10fF
C2852 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# VSS 0.18fF
C2853 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# VSS 0.18fF
C2854 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS 14.13fF
C2855 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# VSS 0.10fF
C2856 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# VSS 0.18fF
C2857 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# VSS 0.18fF
C2858 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS 12.08fF
C2859 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# VSS 0.10fF
C2860 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# VSS 0.18fF
C2861 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# VSS 0.18fF
C2862 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS 14.52fF
C2863 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VSS 0.10fF
C2864 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VSS 0.18fF
C2865 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VSS 0.18fF
C2866 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B VSS 50.31fF
C2867 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# VSS 0.17fF
C2868 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# VSS 0.53fF
C2869 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# VSS 0.18fF
C2870 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS 14.10fF
C2871 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# VSS 0.10fF
C2872 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# VSS 0.18fF
C2873 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# VSS 0.18fF
C2874 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS 20.02fF
C2875 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# VSS 0.10fF
C2876 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# VSS 0.18fF
C2877 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# VSS 0.18fF
C2878 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# VSS 0.10fF
C2879 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# VSS 0.18fF
C2880 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# VSS 0.18fF
C2881 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS 34.82fF
C2882 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# VSS 0.10fF
C2883 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# VSS 0.18fF
C2884 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# VSS 0.18fF
C2885 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS 8.19fF
C2886 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# VSS 0.10fF
C2887 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# VSS 0.18fF
C2888 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# VSS 0.18fF
C2889 clock_v2_0/B VSS 88.14fF
C2890 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_0/a_110_47# VSS 1.28fF
C2891 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS 22.31fF
C2892 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# VSS 0.10fF
C2893 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# VSS 0.18fF
C2894 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# VSS 0.18fF
C2895 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# VSS 0.10fF
C2896 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# VSS 0.18fF
C2897 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# VSS 0.18fF
C2898 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS 51.40fF
C2899 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# VSS 0.10fF
C2900 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# VSS 0.18fF
C2901 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# VSS 0.18fF
C2902 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# VSS 0.10fF
C2903 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# VSS 0.18fF
C2904 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# VSS 0.18fF
C2905 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS 14.77fF
C2906 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# VSS 0.10fF
C2907 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# VSS 0.18fF
C2908 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# VSS 0.18fF
C2909 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS 41.03fF
C2910 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# VSS 0.10fF
C2911 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# VSS 0.18fF
C2912 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# VSS 0.18fF
C2913 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS 20.08fF
C2914 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# VSS 0.10fF
C2915 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# VSS 0.18fF
C2916 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# VSS 0.18fF
C2917 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS 23.37fF
C2918 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# VSS 0.10fF
C2919 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# VSS 0.18fF
C2920 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# VSS 0.18fF
C2921 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS 41.72fF
C2922 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# VSS 0.10fF
C2923 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# VSS 0.18fF
C2924 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# VSS 0.18fF
C2925 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS 21.03fF
C2926 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# VSS 0.10fF
C2927 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# VSS 0.18fF
C2928 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# VSS 0.18fF
C2929 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS 19.88fF
C2930 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# VSS 0.10fF
C2931 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# VSS 0.18fF
C2932 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# VSS 0.18fF
C2933 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS 10.62fF
C2934 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y VSS 27.38fF
C2935 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# VSS 0.10fF
C2936 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# VSS 0.18fF
C2937 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VSS 0.48fF
C2938 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS 14.04fF
C2939 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS 14.52fF
C2940 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# VSS 0.10fF
C2941 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# VSS 0.18fF
C2942 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# VSS 0.18fF
C2943 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS 14.44fF
C2944 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# VSS 0.10fF
C2945 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# VSS 0.18fF
C2946 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# VSS 0.18fF
C2947 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS 23.77fF
C2948 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# VSS 0.10fF
C2949 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# VSS 0.18fF
C2950 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# VSS 0.18fF
C2951 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS 20.06fF
C2952 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# VSS 0.10fF
C2953 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# VSS 0.18fF
C2954 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# VSS 0.18fF
C2955 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS 41.37fF
C2956 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# VSS 0.10fF
C2957 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# VSS 0.18fF
C2958 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# VSS 0.18fF
C2959 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS 20.10fF
C2960 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# VSS 0.10fF
C2961 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# VSS 0.18fF
C2962 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# VSS 0.18fF
C2963 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS 19.92fF
C2964 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# VSS 0.10fF
C2965 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# VSS 0.18fF
C2966 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# VSS 0.18fF
C2967 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS 23.77fF
C2968 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# VSS 0.10fF
C2969 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# VSS 0.18fF
C2970 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# VSS 0.18fF
C2971 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# VSS 0.10fF
C2972 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# VSS 0.18fF
C2973 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# VSS 0.18fF
C2974 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A VSS 48.85fF
C2975 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D VSS 7.04fF
C2976 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_381_47# VSS 0.03fF
C2977 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# VSS 0.09fF
C2978 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413# VSS 0.12fF
C2979 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# VSS 0.24fF
C2980 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# VSS 0.11fF
C2981 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# VSS 0.12fF
C2982 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VSS 0.21fF
C2983 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VSS 0.31fF
C2984 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS 20.23fF
C2985 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# VSS 0.10fF
C2986 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# VSS 0.18fF
C2987 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# VSS 0.18fF
C2988 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS 13.88fF
C2989 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# VSS 0.10fF
C2990 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# VSS 0.18fF
C2991 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# VSS 0.18fF
C2992 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS 13.23fF
C2993 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# VSS 0.10fF
C2994 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# VSS 0.18fF
C2995 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# VSS 0.18fF
C2996 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS 9.06fF
C2997 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# VSS 0.10fF
C2998 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# VSS 0.18fF
C2999 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# VSS 0.18fF
C3000 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS 0.05fF
C3001 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VSS 0.03fF
C3002 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VSS 0.09fF
C3003 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VSS 0.12fF
C3004 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VSS 0.24fF
C3005 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VSS 0.11fF
C3006 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VSS 0.12fF
C3007 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VSS 0.21fF
C3008 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VSS 0.31fF
C3009 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS 14.69fF
C3010 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS 10.20fF
C3011 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# VSS 0.10fF
C3012 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# VSS 0.18fF
C3013 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# VSS 0.18fF
C3014 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS 20.18fF
C3015 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# VSS 0.10fF
C3016 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# VSS 0.18fF
C3017 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# VSS 0.18fF
C3018 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS 9.17fF
C3019 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# VSS 0.10fF
C3020 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# VSS 0.18fF
C3021 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# VSS 0.18fF
C3022 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS 20.16fF
C3023 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# VSS 0.10fF
C3024 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# VSS 0.18fF
C3025 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# VSS 0.18fF
C3026 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS 34.93fF
C3027 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# VSS 0.10fF
C3028 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# VSS 0.18fF
C3029 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# VSS 0.18fF
C3030 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y VSS 55.55fF
C3031 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y VSS 92.52fF
C3032 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS 40.80fF
C3033 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# VSS 0.10fF
C3034 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# VSS 0.18fF
C3035 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# VSS 0.18fF
C3036 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS 13.27fF
C3037 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VSS 0.10fF
C3038 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VSS 0.18fF
C3039 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VSS 0.18fF
C3040 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS 13.28fF
C3041 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VSS 0.10fF
C3042 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VSS 0.18fF
C3043 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VSS 0.18fF
C3044 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS 34.61fF
C3045 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VSS 0.10fF
C3046 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VSS 0.18fF
C3047 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VSS 0.18fF
C3048 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS 47.27fF
C3049 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VSS 0.10fF
C3050 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VSS 0.18fF
C3051 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VSS 0.18fF
C3052 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS 39.64fF
C3053 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VSS 0.10fF
C3054 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VSS 0.18fF
C3055 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VSS 0.18fF
C3056 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A VSS 54.21fF
C3057 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y VSS 73.28fF
C3058 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS 19.98fF
C3059 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VSS 0.10fF
C3060 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VSS 0.18fF
C3061 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VSS 0.18fF
C3062 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y VSS 46.35fF
C3063 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS 20.75fF
C3064 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VSS 0.10fF
C3065 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VSS 0.18fF
C3066 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VSS 0.18fF
C3067 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47# VSS 0.06fF
C3068 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A VSS 91.96fF
C3069 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VSS 0.10fF
C3070 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VSS 0.18fF
C3071 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VSS 0.18fF
C3072 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y VSS 45.02fF
C3073 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47# VSS 0.06fF
C3074 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y VSS 45.11fF
C3075 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.06fF
C3076 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B VSS 50.40fF
C3077 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VSS 0.17fF
C3078 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VSS 0.31fF
C3079 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VSS 0.18fF
C3080 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.06fF
C3081 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS 14.51fF
C3082 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VSS 0.10fF
C3083 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VSS 0.18fF
C3084 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VSS 0.18fF
C3085 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VSS 1.28fF
C3086 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS 14.76fF
C3087 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS 10.62fF
C3088 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VSS 0.10fF
C3089 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VSS 0.18fF
C3090 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VSS 0.18fF
C3091 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A VSS 66.86fF
C3092 clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y VSS 19.57fF
C3093 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VSS 1.28fF
C3094 clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y VSS 27.32fF
C3095 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VSS 0.10fF
C3096 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VSS 0.18fF
C3097 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VSS 0.25fF
C3098 clock_v2_0/p2d VSS 65.36fF
C3099 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VSS 1.28fF
C3100 clock_v2_0/p2d_b VSS 52.59fF
C3101 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VSS 1.28fF
C3102 clock_v2_0/p1d_b VSS 78.65fF
C3103 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VSS 1.28fF
C3104 ota_w_test_v2_0/in VSS -33.01fF
C3105 sky130_fd_sc_hd__mux4_1_3/X VSS 19.72fF
C3106 d_clk_grp_1_ctrl_1 VSS 96.55fF
C3107 d_clk_grp_1_ctrl_0 VSS 47.94fF
C3108 sky130_fd_sc_hd__mux4_1_3/a_834_97# VSS 0.04fF
C3109 sky130_fd_sc_hd__mux4_1_3/a_668_97# VSS 0.04fF
C3110 sky130_fd_sc_hd__mux4_1_3/a_193_47# VSS 0.00fF
C3111 sky130_fd_sc_hd__mux4_1_3/a_27_47# VSS 0.11fF
C3112 sky130_fd_sc_hd__mux4_1_3/a_1478_413# VSS 0.20fF
C3113 sky130_fd_sc_hd__mux4_1_3/a_1290_413# VSS 0.21fF
C3114 sky130_fd_sc_hd__mux4_1_3/a_750_97# VSS 0.10fF
C3115 sky130_fd_sc_hd__mux4_1_3/a_757_363# VSS 0.01fF
C3116 sky130_fd_sc_hd__mux4_1_3/a_277_47# VSS 0.15fF
C3117 sky130_fd_sc_hd__mux4_1_3/a_247_21# VSS 0.31fF
C3118 sky130_fd_sc_hd__mux4_1_3/a_193_413# VSS 0.01fF
C3119 sky130_fd_sc_hd__mux4_1_3/a_27_413# VSS 0.01fF
C3120 sky130_fd_pr__cap_mim_m3_1_CGPBWM_5/m3_n1030_n980# VSS 2.79fF
C3121 sky130_fd_sc_hd__mux4_1_2/X VSS 19.94fF
C3122 sky130_fd_sc_hd__mux4_1_2/a_834_97# VSS 0.04fF
C3123 sky130_fd_sc_hd__mux4_1_2/a_668_97# VSS 0.04fF
C3124 sky130_fd_sc_hd__mux4_1_2/a_193_47# VSS 0.00fF
C3125 sky130_fd_sc_hd__mux4_1_2/a_27_47# VSS 0.12fF
C3126 sky130_fd_sc_hd__mux4_1_2/a_1478_413# VSS 0.19fF
C3127 sky130_fd_sc_hd__mux4_1_2/a_1290_413# VSS 0.19fF
C3128 sky130_fd_sc_hd__mux4_1_2/a_750_97# VSS 0.06fF
C3129 sky130_fd_sc_hd__mux4_1_2/a_757_363# VSS 0.00fF
C3130 sky130_fd_sc_hd__mux4_1_2/a_277_47# VSS 0.15fF
C3131 sky130_fd_sc_hd__mux4_1_2/a_247_21# VSS 0.30fF
C3132 sky130_fd_sc_hd__mux4_1_2/a_27_413# VSS 0.00fF
C3133 sky130_fd_pr__cap_mim_m3_1_CEWQ64_16/m3_n360_n310# VSS 0.63fF
C3134 sky130_fd_sc_hd__mux4_1_1/X VSS 18.13fF
C3135 d_clk_grp_2_ctrl_1 VSS 97.71fF
C3136 d_clk_grp_2_ctrl_0 VSS 46.39fF
C3137 sky130_fd_sc_hd__mux4_1_1/a_834_97# VSS 0.04fF
C3138 sky130_fd_sc_hd__mux4_1_1/a_668_97# VSS 0.04fF
C3139 sky130_fd_sc_hd__mux4_1_1/a_193_47# VSS 0.00fF
C3140 sky130_fd_sc_hd__mux4_1_1/a_27_47# VSS 0.12fF
C3141 sky130_fd_sc_hd__mux4_1_1/a_1478_413# VSS 0.21fF
C3142 sky130_fd_sc_hd__mux4_1_1/a_1290_413# VSS 0.20fF
C3143 sky130_fd_sc_hd__mux4_1_1/a_750_97# VSS 0.10fF
C3144 sky130_fd_sc_hd__mux4_1_1/a_757_363# VSS 0.01fF
C3145 sky130_fd_sc_hd__mux4_1_1/a_277_47# VSS 0.16fF
C3146 sky130_fd_sc_hd__mux4_1_1/a_247_21# VSS 0.30fF
C3147 sky130_fd_sc_hd__mux4_1_1/a_193_413# VSS 0.01fF
C3148 sky130_fd_sc_hd__mux4_1_1/a_27_413# VSS 0.01fF
C3149 sky130_fd_pr__cap_mim_m3_1_CEWQ64_59/m3_n360_n310# VSS 0.63fF
C3150 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/c1_n260_n210# VSS 0.60fF
C3151 sky130_fd_pr__cap_mim_m3_1_CEWQ64_48/m3_n360_n310# VSS 0.91fF
C3152 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# VSS 0.63fF
C3153 sky130_fd_sc_hd__mux4_1_0/X VSS 18.32fF
C3154 sky130_fd_sc_hd__mux4_1_0/a_834_97# VSS 0.04fF
C3155 sky130_fd_sc_hd__mux4_1_0/a_668_97# VSS 0.05fF
C3156 sky130_fd_sc_hd__mux4_1_0/a_193_47# VSS 0.00fF
C3157 sky130_fd_sc_hd__mux4_1_0/a_27_47# VSS 0.13fF
C3158 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VSS 0.21fF
C3159 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VSS 0.21fF
C3160 sky130_fd_sc_hd__mux4_1_0/a_750_97# VSS 0.11fF
C3161 sky130_fd_sc_hd__mux4_1_0/a_757_363# VSS 0.01fF
C3162 sky130_fd_sc_hd__mux4_1_0/a_277_47# VSS 0.19fF
C3163 sky130_fd_sc_hd__mux4_1_0/a_247_21# VSS 0.32fF
C3164 sky130_fd_sc_hd__mux4_1_0/a_193_413# VSS 0.01fF
C3165 sky130_fd_sc_hd__mux4_1_0/a_27_413# VSS 0.02fF
C3166 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# VSS 0.63fF
C3167 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# VSS 0.63fF
C3168 a_mux2_en_1/switch_5t_mux2_0/in VSS 1.10fF
C3169 a_mux2_en_1/transmission_gate_1/en_b VSS -1.21fF
C3170 a_mux2_en_1/switch_5t_mux2_1/in VSS -1.20fF
C3171 a_mux2_en_1/switch_5t_mux2_1/en VSS 12.01fF
C3172 a_mux2_en_1/switch_5t_mux2_1/transmission_gate_1/in VSS 2.73fF
C3173 a_probe_1 VSS 38.37fF
C3174 a_mux2_en_1/switch_5t_mux2_0/transmission_gate_1/in VSS 2.04fF
C3175 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# VSS 2.14fF
C3176 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 2.19fF
C3177 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# VSS 2.14fF
C3178 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 2.19fF
C3179 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# VSS 0.96fF
C3180 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.99fF
C3181 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# VSS 1.96fF
C3182 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 2.27fF
C3183 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C3184 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# VSS 2.14fF
C3185 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 2.19fF
C3186 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C3187 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C3188 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C3189 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# VSS 2.02fF
C3190 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.95fF
C3191 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_9/in VSS 3.89fF
C3192 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# VSS 2.16fF
C3193 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 2.17fF
C3194 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.32fF
C3195 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.32fF
C3196 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# VSS 0.89fF
C3197 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.96fF
C3198 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# VSS 0.96fF
C3199 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.98fF
C3200 ota_v2_0/p2 VSS 461.71fF
C3201 ota_v2_0/p2_b VSS 155.55fF
C3202 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.32fF
C3203 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# VSS 0.91fF
C3204 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 2.10fF
C3205 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.32fF
C3206 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# VSS 0.94fF
C3207 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.92fF
C3208 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# VSS 0.86fF
C3209 ota_w_test_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.89fF
C3210 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_3/out VSS 1.77fF
C3211 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_8/in VSS 1.57fF
C3212 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_6/in VSS -13.54fF
C3213 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_7/in VSS 8.59fF
C3214 a_mux4_en_0/in0 VSS 9.86fF
C3215 ota_v2_0/p1 VSS 275.51fF
C3216 ota_w_test_v2_0/op VSS 10.13fF
C3217 ota_w_test_v2_0/sc_cmfb_0/transmission_gate_4/out VSS -4.30fF
C3218 ota_w_test_v2_0/on VSS -47.99fF
C3219 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C3220 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF
C3221 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_18877_3928# VSS 0.07fF
C3222 ota_w_test_v2_0/ota_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C3223 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11121_570# VSS 9.29fF
C3224 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_11122_5650# VSS -32.46fF
C3225 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8434_570# VSS 9.95fF
C3226 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_8436_5651# VSS 7.31fF
C3227 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -341.49fF
C3228 a_mux4_en_0/in1 VSS -360.62fF
C3229 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C3230 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.86fF
C3231 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C3232 i_bias_1 VSS -26.00fF
C3233 a_mux4_en_1/in1 VSS -146.28fF
C3234 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C3235 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C3236 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C3237 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C3238 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C3239 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C3240 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C3241 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C3242 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.13fF
C3243 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C3244 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C3245 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C3246 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.14fF
C3247 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C3248 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C3249 a_mux4_en_1/in2 VSS -231.76fF
C3250 ota_w_test_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 5.34fF
C3251 a_mux4_en_1/in0 VSS -310.57fF
C3252 ota_w_test_v2_0/ota_v2_without_cmfb_0/li_14138_570# VSS 37.42fF
C3253 a_mux4_en_0/in2 VSS -128.31fF
C3254 sky130_fd_pr__cap_mim_m3_1_CEWQ64_68/m3_n360_n310# VSS 0.63fF
C3255 sky130_fd_pr__cap_mim_m3_1_CEWQ64_57/m3_n360_n310# VSS 0.63fF
C3256 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# VSS 0.63fF
C3257 sky130_fd_pr__cap_mim_m3_1_CEWQ64_13/m3_n360_n310# VSS 0.63fF
C3258 onebit_dac_1/out VSS 52.54fF
C3259 a_mux2_en_0/switch_5t_mux2_0/in VSS 1.10fF
C3260 a_mux2_en_0/transmission_gate_1/en_b VSS -1.22fF
C3261 a_mux2_en_0/switch_5t_mux2_1/in VSS -1.20fF
C3262 a_mux2_en_0/switch_5t_mux2_1/en VSS 19.50fF
C3263 a_mod_grp_ctrl_0 VSS 129.38fF
C3264 a_mux2_en_0/switch_5t_mux2_1/transmission_gate_1/in VSS 2.08fF
C3265 a_probe_0 VSS 41.79fF
C3266 a_mux2_en_0/switch_5t_mux2_0/transmission_gate_1/in VSS 2.48fF
C3267 transmission_gate_29/out VSS -24.80fF
C3268 in VSS 84.02fF
C3269 sky130_fd_sc_hd__clkinv_4_3/Y VSS 55.49fF
C3270 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# VSS 2.79fF
C3271 sky130_fd_pr__cap_mim_m3_1_CEWQ64_67/m3_n360_n310# VSS 0.63fF
C3272 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# VSS 0.63fF
C3273 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# VSS 0.63fF
C3274 onebit_dac_1/v_b VSS 22.76fF
C3275 op VSS 50.58fF
C3276 onebit_dac_0/out VSS 44.26fF
C3277 sky130_fd_sc_hd__clkinv_4_2/Y VSS 55.96fF
C3278 sky130_fd_pr__cap_mim_m3_1_CEWQ64_66/m3_n360_n310# VSS 0.63fF
C3279 sky130_fd_pr__cap_mim_m3_1_CEWQ64_44/m3_n360_n310# VSS 0.63fF
C3280 sky130_fd_pr__cap_mim_m3_1_CEWQ64_11/m3_n360_n310# VSS 0.63fF
C3281 d_probe_0 VSS -76.06fF
C3282 transmission_gate_7/en VSS -32.71fF
C3283 rst_n VSS -5.73fF
C3284 sky130_fd_sc_hd__clkinv_4_1/Y VSS 56.91fF
C3285 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# VSS 0.63fF
C3286 d_probe_3 VSS -77.54fF
C3287 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# VSS 0.63fF
C3288 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# VSS 0.63fF
C3289 sky130_fd_pr__cap_mim_m3_1_CEWQ64_21/m3_n360_n310# VSS 0.63fF
C3290 ota_v2_0/in VSS 4.75fF
C3291 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# VSS 0.63fF
C3292 sky130_fd_sc_hd__clkinv_4_0/Y VSS 55.43fF
C3293 sky130_fd_pr__cap_mim_m3_1_CEWQ64_64/m3_n360_n310# VSS 0.63fF
C3294 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/c1_n260_n210# VSS 0.58fF
C3295 sky130_fd_pr__cap_mim_m3_1_CEWQ64_20/m3_n360_n310# VSS 0.89fF
C3296 d_probe_2 VSS -76.73fF
C3297 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# VSS 0.63fF
C3298 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# VSS 1.97fF
C3299 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 2.18fF
C3300 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# VSS 2.15fF
C3301 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 2.20fF
C3302 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# VSS 0.94fF
C3303 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.97fF
C3304 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# VSS 2.15fF
C3305 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 2.14fF
C3306 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C3307 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# VSS 1.97fF
C3308 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 2.33fF
C3309 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C3310 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C3311 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C3312 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# VSS 2.02fF
C3313 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.77fF
C3314 ota_v2_0/sc_cmfb_0/transmission_gate_9/in VSS 3.28fF
C3315 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# VSS 2.16fF
C3316 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 2.16fF
C3317 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C3318 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C3319 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# VSS 0.82fF
C3320 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.94fF
C3321 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# VSS 0.94fF
C3322 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.98fF
C3323 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C3324 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# VSS 0.96fF
C3325 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.96fF
C3326 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C3327 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# VSS 0.87fF
C3328 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 2.05fF
C3329 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# VSS 0.85fF
C3330 ota_v2_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.93fF
C3331 ota_v2_0/sc_cmfb_0/transmission_gate_3/out VSS 1.83fF
C3332 ota_v2_0/sc_cmfb_0/transmission_gate_8/in VSS 1.62fF
C3333 ota_v2_0/sc_cmfb_0/transmission_gate_6/in VSS -14.07fF
C3334 ota_v2_0/sc_cmfb_0/transmission_gate_7/in VSS 8.55fF
C3335 ota_v2_0/cm VSS 46.31fF
C3336 ota_v2_0/sc_cmfb_0/transmission_gate_4/out VSS -4.30fF
C3337 ota_v2_0/ota_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C3338 ota_v2_0/ota_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF
C3339 ota_v2_0/ota_v2_without_cmfb_0/m1_18877_3928# VSS 0.05fF
C3340 ota_v2_0/ota_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C3341 ota_v2_0/ota_v2_without_cmfb_0/li_11121_570# VSS 9.30fF
C3342 ota_v2_0/ota_v2_without_cmfb_0/li_11122_5650# VSS -32.42fF
C3343 ota_v2_0/ota_v2_without_cmfb_0/li_8434_570# VSS 9.95fF
C3344 ota_v2_0/ota_v2_without_cmfb_0/li_8436_5651# VSS 6.76fF
C3345 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -341.42fF
C3346 ota_v2_0/ota_v2_without_cmfb_0/bias_b VSS -358.51fF
C3347 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C3348 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.85fF
C3349 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C3350 i_bias_2 VSS -19.47fF
C3351 ota_v2_0/ota_v2_without_cmfb_0/bias_c VSS -126.27fF
C3352 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C3353 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C3354 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C3355 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C3356 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C3357 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C3358 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C3359 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C3360 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.13fF
C3361 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C3362 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C3363 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C3364 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.14fF
C3365 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C3366 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C3367 ota_v2_0/ota_v2_without_cmfb_0/bias_d VSS -235.44fF
C3368 ota_v2_0/ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 4.88fF
C3369 ota_v2_0/sc_cmfb_0/bias_a VSS -319.96fF
C3370 ota_v2_0/ota_v2_without_cmfb_0/li_14138_570# VSS 38.28fF
C3371 ota_v2_0/sc_cmfb_0/cmc VSS -132.28fF
C3372 d_probe_1 VSS -75.79fF
C3373 sky130_fd_pr__cap_mim_m3_1_CEWQ64_63/m3_n360_n310# VSS 0.63fF
C3374 a_mux2_en_0/in1 VSS 54.37fF
C3375 transmission_gate_25/in VSS 4.03fF
C3376 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# VSS 0.63fF
C3377 sky130_fd_pr__cap_mim_m3_1_CEWQ64_62/m3_n360_n310# VSS 0.63fF
C3378 sky130_fd_pr__cap_mim_m3_1_CEWQ64_40/m3_n360_n310# VSS 0.63fF
C3379 a_mux2_en_0/in0 VSS 31.93fF
C3380 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# VSS 0.63fF
C3381 sky130_fd_pr__cap_mim_m3_1_CEWQ64_61/m3_n360_n310# VSS 0.63fF
C3382 transmission_gate_31/out VSS 7.53fF
C3383 ota_v2_0/ip VSS -3.60fF
C3384 transmission_gate_23/in VSS -30.33fF
C3385 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# VSS 0.63fF
C3386 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# VSS 0.63fF
C3387 sky130_fd_pr__cap_mim_m3_1_CEWQ64_60/m3_n360_n310# VSS 0.63fF
C3388 transmission_gate_32/out VSS 7.78fF
C3389 transmission_gate_21/out VSS -13.82fF
C3390 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# VSS 0.63fF
C3391 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# VSS 2.79fF
C3392 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# VSS 0.63fF
C3393 transmission_gate_21/in VSS -3.17fF
C3394 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# VSS 2.79fF
C3395 sky130_fd_pr__cap_mim_m3_1_CGPBWM_18/m3_n1030_n980# VSS 2.79fF
C3396 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# VSS 0.63fF
.ends

