magic
tech sky130A
magscale 1 2
timestamp 1653694315
<< nwell >>
rect -2098 7664 -804 8314
rect 6902 7664 8196 8314
rect -2098 5864 -804 6514
rect 6902 5864 8196 6514
rect -2098 4064 -804 4714
rect 6902 4064 8196 4714
rect -2098 2264 -804 2914
rect 6902 2264 8196 2914
rect -2098 464 -804 1114
rect 6902 464 8196 1114
rect -2098 -1336 -804 -686
rect 6902 -1336 8196 -686
<< pwell >>
rect -2098 7200 -804 7662
rect 6902 7200 8196 7662
rect -2098 5400 -804 5862
rect 6902 5400 8196 5862
rect -2098 3600 -804 4062
rect 6902 3600 8196 4062
rect -2098 1800 -804 2262
rect 6902 1800 8196 2262
rect -2098 0 -804 462
rect 6902 0 8196 462
rect -2098 -1800 -804 -1338
rect 6902 -1800 8196 -1338
<< nmos >>
rect -1898 7410 -1868 7514
rect -1802 7410 -1772 7514
rect -1706 7410 -1676 7514
rect -1610 7410 -1580 7514
rect -1514 7410 -1484 7514
rect -1418 7410 -1388 7514
rect -1322 7410 -1292 7514
rect -1226 7410 -1196 7514
rect -1130 7410 -1100 7514
rect -1034 7410 -1004 7514
rect 7102 7410 7132 7514
rect 7198 7410 7228 7514
rect 7294 7410 7324 7514
rect 7390 7410 7420 7514
rect 7486 7410 7516 7514
rect 7582 7410 7612 7514
rect 7678 7410 7708 7514
rect 7774 7410 7804 7514
rect 7870 7410 7900 7514
rect 7966 7410 7996 7514
rect -1898 5610 -1868 5714
rect -1802 5610 -1772 5714
rect -1706 5610 -1676 5714
rect -1610 5610 -1580 5714
rect -1514 5610 -1484 5714
rect -1418 5610 -1388 5714
rect -1322 5610 -1292 5714
rect -1226 5610 -1196 5714
rect -1130 5610 -1100 5714
rect -1034 5610 -1004 5714
rect 7102 5610 7132 5714
rect 7198 5610 7228 5714
rect 7294 5610 7324 5714
rect 7390 5610 7420 5714
rect 7486 5610 7516 5714
rect 7582 5610 7612 5714
rect 7678 5610 7708 5714
rect 7774 5610 7804 5714
rect 7870 5610 7900 5714
rect 7966 5610 7996 5714
rect -1898 3810 -1868 3914
rect -1802 3810 -1772 3914
rect -1706 3810 -1676 3914
rect -1610 3810 -1580 3914
rect -1514 3810 -1484 3914
rect -1418 3810 -1388 3914
rect -1322 3810 -1292 3914
rect -1226 3810 -1196 3914
rect -1130 3810 -1100 3914
rect -1034 3810 -1004 3914
rect 7102 3810 7132 3914
rect 7198 3810 7228 3914
rect 7294 3810 7324 3914
rect 7390 3810 7420 3914
rect 7486 3810 7516 3914
rect 7582 3810 7612 3914
rect 7678 3810 7708 3914
rect 7774 3810 7804 3914
rect 7870 3810 7900 3914
rect 7966 3810 7996 3914
rect -1898 2010 -1868 2114
rect -1802 2010 -1772 2114
rect -1706 2010 -1676 2114
rect -1610 2010 -1580 2114
rect -1514 2010 -1484 2114
rect -1418 2010 -1388 2114
rect -1322 2010 -1292 2114
rect -1226 2010 -1196 2114
rect -1130 2010 -1100 2114
rect -1034 2010 -1004 2114
rect 7102 2010 7132 2114
rect 7198 2010 7228 2114
rect 7294 2010 7324 2114
rect 7390 2010 7420 2114
rect 7486 2010 7516 2114
rect 7582 2010 7612 2114
rect 7678 2010 7708 2114
rect 7774 2010 7804 2114
rect 7870 2010 7900 2114
rect 7966 2010 7996 2114
rect -1898 210 -1868 314
rect -1802 210 -1772 314
rect -1706 210 -1676 314
rect -1610 210 -1580 314
rect -1514 210 -1484 314
rect -1418 210 -1388 314
rect -1322 210 -1292 314
rect -1226 210 -1196 314
rect -1130 210 -1100 314
rect -1034 210 -1004 314
rect 7102 210 7132 314
rect 7198 210 7228 314
rect 7294 210 7324 314
rect 7390 210 7420 314
rect 7486 210 7516 314
rect 7582 210 7612 314
rect 7678 210 7708 314
rect 7774 210 7804 314
rect 7870 210 7900 314
rect 7966 210 7996 314
rect -1898 -1590 -1868 -1486
rect -1802 -1590 -1772 -1486
rect -1706 -1590 -1676 -1486
rect -1610 -1590 -1580 -1486
rect -1514 -1590 -1484 -1486
rect -1418 -1590 -1388 -1486
rect -1322 -1590 -1292 -1486
rect -1226 -1590 -1196 -1486
rect -1130 -1590 -1100 -1486
rect -1034 -1590 -1004 -1486
rect 7102 -1590 7132 -1486
rect 7198 -1590 7228 -1486
rect 7294 -1590 7324 -1486
rect 7390 -1590 7420 -1486
rect 7486 -1590 7516 -1486
rect 7582 -1590 7612 -1486
rect 7678 -1590 7708 -1486
rect 7774 -1590 7804 -1486
rect 7870 -1590 7900 -1486
rect 7966 -1590 7996 -1486
<< pmos >>
rect -1898 7822 -1868 8094
rect -1802 7822 -1772 8094
rect -1706 7822 -1676 8094
rect -1610 7822 -1580 8094
rect -1514 7822 -1484 8094
rect -1418 7822 -1388 8094
rect -1322 7822 -1292 8094
rect -1226 7822 -1196 8094
rect -1130 7822 -1100 8094
rect -1034 7822 -1004 8094
rect 7102 7822 7132 8094
rect 7198 7822 7228 8094
rect 7294 7822 7324 8094
rect 7390 7822 7420 8094
rect 7486 7822 7516 8094
rect 7582 7822 7612 8094
rect 7678 7822 7708 8094
rect 7774 7822 7804 8094
rect 7870 7822 7900 8094
rect 7966 7822 7996 8094
rect -1898 6022 -1868 6294
rect -1802 6022 -1772 6294
rect -1706 6022 -1676 6294
rect -1610 6022 -1580 6294
rect -1514 6022 -1484 6294
rect -1418 6022 -1388 6294
rect -1322 6022 -1292 6294
rect -1226 6022 -1196 6294
rect -1130 6022 -1100 6294
rect -1034 6022 -1004 6294
rect 7102 6022 7132 6294
rect 7198 6022 7228 6294
rect 7294 6022 7324 6294
rect 7390 6022 7420 6294
rect 7486 6022 7516 6294
rect 7582 6022 7612 6294
rect 7678 6022 7708 6294
rect 7774 6022 7804 6294
rect 7870 6022 7900 6294
rect 7966 6022 7996 6294
rect -1898 4222 -1868 4494
rect -1802 4222 -1772 4494
rect -1706 4222 -1676 4494
rect -1610 4222 -1580 4494
rect -1514 4222 -1484 4494
rect -1418 4222 -1388 4494
rect -1322 4222 -1292 4494
rect -1226 4222 -1196 4494
rect -1130 4222 -1100 4494
rect -1034 4222 -1004 4494
rect 7102 4222 7132 4494
rect 7198 4222 7228 4494
rect 7294 4222 7324 4494
rect 7390 4222 7420 4494
rect 7486 4222 7516 4494
rect 7582 4222 7612 4494
rect 7678 4222 7708 4494
rect 7774 4222 7804 4494
rect 7870 4222 7900 4494
rect 7966 4222 7996 4494
rect -1898 2422 -1868 2694
rect -1802 2422 -1772 2694
rect -1706 2422 -1676 2694
rect -1610 2422 -1580 2694
rect -1514 2422 -1484 2694
rect -1418 2422 -1388 2694
rect -1322 2422 -1292 2694
rect -1226 2422 -1196 2694
rect -1130 2422 -1100 2694
rect -1034 2422 -1004 2694
rect 7102 2422 7132 2694
rect 7198 2422 7228 2694
rect 7294 2422 7324 2694
rect 7390 2422 7420 2694
rect 7486 2422 7516 2694
rect 7582 2422 7612 2694
rect 7678 2422 7708 2694
rect 7774 2422 7804 2694
rect 7870 2422 7900 2694
rect 7966 2422 7996 2694
rect -1898 622 -1868 894
rect -1802 622 -1772 894
rect -1706 622 -1676 894
rect -1610 622 -1580 894
rect -1514 622 -1484 894
rect -1418 622 -1388 894
rect -1322 622 -1292 894
rect -1226 622 -1196 894
rect -1130 622 -1100 894
rect -1034 622 -1004 894
rect 7102 622 7132 894
rect 7198 622 7228 894
rect 7294 622 7324 894
rect 7390 622 7420 894
rect 7486 622 7516 894
rect 7582 622 7612 894
rect 7678 622 7708 894
rect 7774 622 7804 894
rect 7870 622 7900 894
rect 7966 622 7996 894
rect -1898 -1178 -1868 -906
rect -1802 -1178 -1772 -906
rect -1706 -1178 -1676 -906
rect -1610 -1178 -1580 -906
rect -1514 -1178 -1484 -906
rect -1418 -1178 -1388 -906
rect -1322 -1178 -1292 -906
rect -1226 -1178 -1196 -906
rect -1130 -1178 -1100 -906
rect -1034 -1178 -1004 -906
rect 7102 -1178 7132 -906
rect 7198 -1178 7228 -906
rect 7294 -1178 7324 -906
rect 7390 -1178 7420 -906
rect 7486 -1178 7516 -906
rect 7582 -1178 7612 -906
rect 7678 -1178 7708 -906
rect 7774 -1178 7804 -906
rect 7870 -1178 7900 -906
rect 7966 -1178 7996 -906
<< ndiff >>
rect -1960 7502 -1898 7514
rect -1960 7422 -1948 7502
rect -1914 7422 -1898 7502
rect -1960 7410 -1898 7422
rect -1868 7502 -1802 7514
rect -1868 7422 -1852 7502
rect -1818 7422 -1802 7502
rect -1868 7410 -1802 7422
rect -1772 7502 -1706 7514
rect -1772 7422 -1756 7502
rect -1722 7422 -1706 7502
rect -1772 7410 -1706 7422
rect -1676 7502 -1610 7514
rect -1676 7422 -1660 7502
rect -1626 7422 -1610 7502
rect -1676 7410 -1610 7422
rect -1580 7502 -1514 7514
rect -1580 7422 -1564 7502
rect -1530 7422 -1514 7502
rect -1580 7410 -1514 7422
rect -1484 7502 -1418 7514
rect -1484 7422 -1468 7502
rect -1434 7422 -1418 7502
rect -1484 7410 -1418 7422
rect -1388 7502 -1322 7514
rect -1388 7422 -1372 7502
rect -1338 7422 -1322 7502
rect -1388 7410 -1322 7422
rect -1292 7502 -1226 7514
rect -1292 7422 -1276 7502
rect -1242 7422 -1226 7502
rect -1292 7410 -1226 7422
rect -1196 7502 -1130 7514
rect -1196 7422 -1180 7502
rect -1146 7422 -1130 7502
rect -1196 7410 -1130 7422
rect -1100 7502 -1034 7514
rect -1100 7422 -1084 7502
rect -1050 7422 -1034 7502
rect -1100 7410 -1034 7422
rect -1004 7502 -942 7514
rect -1004 7422 -988 7502
rect -954 7422 -942 7502
rect -1004 7410 -942 7422
rect 7040 7502 7102 7514
rect 7040 7422 7052 7502
rect 7086 7422 7102 7502
rect 7040 7410 7102 7422
rect 7132 7502 7198 7514
rect 7132 7422 7148 7502
rect 7182 7422 7198 7502
rect 7132 7410 7198 7422
rect 7228 7502 7294 7514
rect 7228 7422 7244 7502
rect 7278 7422 7294 7502
rect 7228 7410 7294 7422
rect 7324 7502 7390 7514
rect 7324 7422 7340 7502
rect 7374 7422 7390 7502
rect 7324 7410 7390 7422
rect 7420 7502 7486 7514
rect 7420 7422 7436 7502
rect 7470 7422 7486 7502
rect 7420 7410 7486 7422
rect 7516 7502 7582 7514
rect 7516 7422 7532 7502
rect 7566 7422 7582 7502
rect 7516 7410 7582 7422
rect 7612 7502 7678 7514
rect 7612 7422 7628 7502
rect 7662 7422 7678 7502
rect 7612 7410 7678 7422
rect 7708 7502 7774 7514
rect 7708 7422 7724 7502
rect 7758 7422 7774 7502
rect 7708 7410 7774 7422
rect 7804 7502 7870 7514
rect 7804 7422 7820 7502
rect 7854 7422 7870 7502
rect 7804 7410 7870 7422
rect 7900 7502 7966 7514
rect 7900 7422 7916 7502
rect 7950 7422 7966 7502
rect 7900 7410 7966 7422
rect 7996 7502 8058 7514
rect 7996 7422 8012 7502
rect 8046 7422 8058 7502
rect 7996 7410 8058 7422
rect -1960 5702 -1898 5714
rect -1960 5622 -1948 5702
rect -1914 5622 -1898 5702
rect -1960 5610 -1898 5622
rect -1868 5702 -1802 5714
rect -1868 5622 -1852 5702
rect -1818 5622 -1802 5702
rect -1868 5610 -1802 5622
rect -1772 5702 -1706 5714
rect -1772 5622 -1756 5702
rect -1722 5622 -1706 5702
rect -1772 5610 -1706 5622
rect -1676 5702 -1610 5714
rect -1676 5622 -1660 5702
rect -1626 5622 -1610 5702
rect -1676 5610 -1610 5622
rect -1580 5702 -1514 5714
rect -1580 5622 -1564 5702
rect -1530 5622 -1514 5702
rect -1580 5610 -1514 5622
rect -1484 5702 -1418 5714
rect -1484 5622 -1468 5702
rect -1434 5622 -1418 5702
rect -1484 5610 -1418 5622
rect -1388 5702 -1322 5714
rect -1388 5622 -1372 5702
rect -1338 5622 -1322 5702
rect -1388 5610 -1322 5622
rect -1292 5702 -1226 5714
rect -1292 5622 -1276 5702
rect -1242 5622 -1226 5702
rect -1292 5610 -1226 5622
rect -1196 5702 -1130 5714
rect -1196 5622 -1180 5702
rect -1146 5622 -1130 5702
rect -1196 5610 -1130 5622
rect -1100 5702 -1034 5714
rect -1100 5622 -1084 5702
rect -1050 5622 -1034 5702
rect -1100 5610 -1034 5622
rect -1004 5702 -942 5714
rect -1004 5622 -988 5702
rect -954 5622 -942 5702
rect -1004 5610 -942 5622
rect 7040 5702 7102 5714
rect 7040 5622 7052 5702
rect 7086 5622 7102 5702
rect 7040 5610 7102 5622
rect 7132 5702 7198 5714
rect 7132 5622 7148 5702
rect 7182 5622 7198 5702
rect 7132 5610 7198 5622
rect 7228 5702 7294 5714
rect 7228 5622 7244 5702
rect 7278 5622 7294 5702
rect 7228 5610 7294 5622
rect 7324 5702 7390 5714
rect 7324 5622 7340 5702
rect 7374 5622 7390 5702
rect 7324 5610 7390 5622
rect 7420 5702 7486 5714
rect 7420 5622 7436 5702
rect 7470 5622 7486 5702
rect 7420 5610 7486 5622
rect 7516 5702 7582 5714
rect 7516 5622 7532 5702
rect 7566 5622 7582 5702
rect 7516 5610 7582 5622
rect 7612 5702 7678 5714
rect 7612 5622 7628 5702
rect 7662 5622 7678 5702
rect 7612 5610 7678 5622
rect 7708 5702 7774 5714
rect 7708 5622 7724 5702
rect 7758 5622 7774 5702
rect 7708 5610 7774 5622
rect 7804 5702 7870 5714
rect 7804 5622 7820 5702
rect 7854 5622 7870 5702
rect 7804 5610 7870 5622
rect 7900 5702 7966 5714
rect 7900 5622 7916 5702
rect 7950 5622 7966 5702
rect 7900 5610 7966 5622
rect 7996 5702 8058 5714
rect 7996 5622 8012 5702
rect 8046 5622 8058 5702
rect 7996 5610 8058 5622
rect -1960 3902 -1898 3914
rect -1960 3822 -1948 3902
rect -1914 3822 -1898 3902
rect -1960 3810 -1898 3822
rect -1868 3902 -1802 3914
rect -1868 3822 -1852 3902
rect -1818 3822 -1802 3902
rect -1868 3810 -1802 3822
rect -1772 3902 -1706 3914
rect -1772 3822 -1756 3902
rect -1722 3822 -1706 3902
rect -1772 3810 -1706 3822
rect -1676 3902 -1610 3914
rect -1676 3822 -1660 3902
rect -1626 3822 -1610 3902
rect -1676 3810 -1610 3822
rect -1580 3902 -1514 3914
rect -1580 3822 -1564 3902
rect -1530 3822 -1514 3902
rect -1580 3810 -1514 3822
rect -1484 3902 -1418 3914
rect -1484 3822 -1468 3902
rect -1434 3822 -1418 3902
rect -1484 3810 -1418 3822
rect -1388 3902 -1322 3914
rect -1388 3822 -1372 3902
rect -1338 3822 -1322 3902
rect -1388 3810 -1322 3822
rect -1292 3902 -1226 3914
rect -1292 3822 -1276 3902
rect -1242 3822 -1226 3902
rect -1292 3810 -1226 3822
rect -1196 3902 -1130 3914
rect -1196 3822 -1180 3902
rect -1146 3822 -1130 3902
rect -1196 3810 -1130 3822
rect -1100 3902 -1034 3914
rect -1100 3822 -1084 3902
rect -1050 3822 -1034 3902
rect -1100 3810 -1034 3822
rect -1004 3902 -942 3914
rect -1004 3822 -988 3902
rect -954 3822 -942 3902
rect -1004 3810 -942 3822
rect 7040 3902 7102 3914
rect 7040 3822 7052 3902
rect 7086 3822 7102 3902
rect 7040 3810 7102 3822
rect 7132 3902 7198 3914
rect 7132 3822 7148 3902
rect 7182 3822 7198 3902
rect 7132 3810 7198 3822
rect 7228 3902 7294 3914
rect 7228 3822 7244 3902
rect 7278 3822 7294 3902
rect 7228 3810 7294 3822
rect 7324 3902 7390 3914
rect 7324 3822 7340 3902
rect 7374 3822 7390 3902
rect 7324 3810 7390 3822
rect 7420 3902 7486 3914
rect 7420 3822 7436 3902
rect 7470 3822 7486 3902
rect 7420 3810 7486 3822
rect 7516 3902 7582 3914
rect 7516 3822 7532 3902
rect 7566 3822 7582 3902
rect 7516 3810 7582 3822
rect 7612 3902 7678 3914
rect 7612 3822 7628 3902
rect 7662 3822 7678 3902
rect 7612 3810 7678 3822
rect 7708 3902 7774 3914
rect 7708 3822 7724 3902
rect 7758 3822 7774 3902
rect 7708 3810 7774 3822
rect 7804 3902 7870 3914
rect 7804 3822 7820 3902
rect 7854 3822 7870 3902
rect 7804 3810 7870 3822
rect 7900 3902 7966 3914
rect 7900 3822 7916 3902
rect 7950 3822 7966 3902
rect 7900 3810 7966 3822
rect 7996 3902 8058 3914
rect 7996 3822 8012 3902
rect 8046 3822 8058 3902
rect 7996 3810 8058 3822
rect -1960 2102 -1898 2114
rect -1960 2022 -1948 2102
rect -1914 2022 -1898 2102
rect -1960 2010 -1898 2022
rect -1868 2102 -1802 2114
rect -1868 2022 -1852 2102
rect -1818 2022 -1802 2102
rect -1868 2010 -1802 2022
rect -1772 2102 -1706 2114
rect -1772 2022 -1756 2102
rect -1722 2022 -1706 2102
rect -1772 2010 -1706 2022
rect -1676 2102 -1610 2114
rect -1676 2022 -1660 2102
rect -1626 2022 -1610 2102
rect -1676 2010 -1610 2022
rect -1580 2102 -1514 2114
rect -1580 2022 -1564 2102
rect -1530 2022 -1514 2102
rect -1580 2010 -1514 2022
rect -1484 2102 -1418 2114
rect -1484 2022 -1468 2102
rect -1434 2022 -1418 2102
rect -1484 2010 -1418 2022
rect -1388 2102 -1322 2114
rect -1388 2022 -1372 2102
rect -1338 2022 -1322 2102
rect -1388 2010 -1322 2022
rect -1292 2102 -1226 2114
rect -1292 2022 -1276 2102
rect -1242 2022 -1226 2102
rect -1292 2010 -1226 2022
rect -1196 2102 -1130 2114
rect -1196 2022 -1180 2102
rect -1146 2022 -1130 2102
rect -1196 2010 -1130 2022
rect -1100 2102 -1034 2114
rect -1100 2022 -1084 2102
rect -1050 2022 -1034 2102
rect -1100 2010 -1034 2022
rect -1004 2102 -942 2114
rect -1004 2022 -988 2102
rect -954 2022 -942 2102
rect -1004 2010 -942 2022
rect 7040 2102 7102 2114
rect 7040 2022 7052 2102
rect 7086 2022 7102 2102
rect 7040 2010 7102 2022
rect 7132 2102 7198 2114
rect 7132 2022 7148 2102
rect 7182 2022 7198 2102
rect 7132 2010 7198 2022
rect 7228 2102 7294 2114
rect 7228 2022 7244 2102
rect 7278 2022 7294 2102
rect 7228 2010 7294 2022
rect 7324 2102 7390 2114
rect 7324 2022 7340 2102
rect 7374 2022 7390 2102
rect 7324 2010 7390 2022
rect 7420 2102 7486 2114
rect 7420 2022 7436 2102
rect 7470 2022 7486 2102
rect 7420 2010 7486 2022
rect 7516 2102 7582 2114
rect 7516 2022 7532 2102
rect 7566 2022 7582 2102
rect 7516 2010 7582 2022
rect 7612 2102 7678 2114
rect 7612 2022 7628 2102
rect 7662 2022 7678 2102
rect 7612 2010 7678 2022
rect 7708 2102 7774 2114
rect 7708 2022 7724 2102
rect 7758 2022 7774 2102
rect 7708 2010 7774 2022
rect 7804 2102 7870 2114
rect 7804 2022 7820 2102
rect 7854 2022 7870 2102
rect 7804 2010 7870 2022
rect 7900 2102 7966 2114
rect 7900 2022 7916 2102
rect 7950 2022 7966 2102
rect 7900 2010 7966 2022
rect 7996 2102 8058 2114
rect 7996 2022 8012 2102
rect 8046 2022 8058 2102
rect 7996 2010 8058 2022
rect -1960 302 -1898 314
rect -1960 222 -1948 302
rect -1914 222 -1898 302
rect -1960 210 -1898 222
rect -1868 302 -1802 314
rect -1868 222 -1852 302
rect -1818 222 -1802 302
rect -1868 210 -1802 222
rect -1772 302 -1706 314
rect -1772 222 -1756 302
rect -1722 222 -1706 302
rect -1772 210 -1706 222
rect -1676 302 -1610 314
rect -1676 222 -1660 302
rect -1626 222 -1610 302
rect -1676 210 -1610 222
rect -1580 302 -1514 314
rect -1580 222 -1564 302
rect -1530 222 -1514 302
rect -1580 210 -1514 222
rect -1484 302 -1418 314
rect -1484 222 -1468 302
rect -1434 222 -1418 302
rect -1484 210 -1418 222
rect -1388 302 -1322 314
rect -1388 222 -1372 302
rect -1338 222 -1322 302
rect -1388 210 -1322 222
rect -1292 302 -1226 314
rect -1292 222 -1276 302
rect -1242 222 -1226 302
rect -1292 210 -1226 222
rect -1196 302 -1130 314
rect -1196 222 -1180 302
rect -1146 222 -1130 302
rect -1196 210 -1130 222
rect -1100 302 -1034 314
rect -1100 222 -1084 302
rect -1050 222 -1034 302
rect -1100 210 -1034 222
rect -1004 302 -942 314
rect -1004 222 -988 302
rect -954 222 -942 302
rect -1004 210 -942 222
rect 7040 302 7102 314
rect 7040 222 7052 302
rect 7086 222 7102 302
rect 7040 210 7102 222
rect 7132 302 7198 314
rect 7132 222 7148 302
rect 7182 222 7198 302
rect 7132 210 7198 222
rect 7228 302 7294 314
rect 7228 222 7244 302
rect 7278 222 7294 302
rect 7228 210 7294 222
rect 7324 302 7390 314
rect 7324 222 7340 302
rect 7374 222 7390 302
rect 7324 210 7390 222
rect 7420 302 7486 314
rect 7420 222 7436 302
rect 7470 222 7486 302
rect 7420 210 7486 222
rect 7516 302 7582 314
rect 7516 222 7532 302
rect 7566 222 7582 302
rect 7516 210 7582 222
rect 7612 302 7678 314
rect 7612 222 7628 302
rect 7662 222 7678 302
rect 7612 210 7678 222
rect 7708 302 7774 314
rect 7708 222 7724 302
rect 7758 222 7774 302
rect 7708 210 7774 222
rect 7804 302 7870 314
rect 7804 222 7820 302
rect 7854 222 7870 302
rect 7804 210 7870 222
rect 7900 302 7966 314
rect 7900 222 7916 302
rect 7950 222 7966 302
rect 7900 210 7966 222
rect 7996 302 8058 314
rect 7996 222 8012 302
rect 8046 222 8058 302
rect 7996 210 8058 222
rect -1960 -1498 -1898 -1486
rect -1960 -1578 -1948 -1498
rect -1914 -1578 -1898 -1498
rect -1960 -1590 -1898 -1578
rect -1868 -1498 -1802 -1486
rect -1868 -1578 -1852 -1498
rect -1818 -1578 -1802 -1498
rect -1868 -1590 -1802 -1578
rect -1772 -1498 -1706 -1486
rect -1772 -1578 -1756 -1498
rect -1722 -1578 -1706 -1498
rect -1772 -1590 -1706 -1578
rect -1676 -1498 -1610 -1486
rect -1676 -1578 -1660 -1498
rect -1626 -1578 -1610 -1498
rect -1676 -1590 -1610 -1578
rect -1580 -1498 -1514 -1486
rect -1580 -1578 -1564 -1498
rect -1530 -1578 -1514 -1498
rect -1580 -1590 -1514 -1578
rect -1484 -1498 -1418 -1486
rect -1484 -1578 -1468 -1498
rect -1434 -1578 -1418 -1498
rect -1484 -1590 -1418 -1578
rect -1388 -1498 -1322 -1486
rect -1388 -1578 -1372 -1498
rect -1338 -1578 -1322 -1498
rect -1388 -1590 -1322 -1578
rect -1292 -1498 -1226 -1486
rect -1292 -1578 -1276 -1498
rect -1242 -1578 -1226 -1498
rect -1292 -1590 -1226 -1578
rect -1196 -1498 -1130 -1486
rect -1196 -1578 -1180 -1498
rect -1146 -1578 -1130 -1498
rect -1196 -1590 -1130 -1578
rect -1100 -1498 -1034 -1486
rect -1100 -1578 -1084 -1498
rect -1050 -1578 -1034 -1498
rect -1100 -1590 -1034 -1578
rect -1004 -1498 -942 -1486
rect -1004 -1578 -988 -1498
rect -954 -1578 -942 -1498
rect -1004 -1590 -942 -1578
rect 7040 -1498 7102 -1486
rect 7040 -1578 7052 -1498
rect 7086 -1578 7102 -1498
rect 7040 -1590 7102 -1578
rect 7132 -1498 7198 -1486
rect 7132 -1578 7148 -1498
rect 7182 -1578 7198 -1498
rect 7132 -1590 7198 -1578
rect 7228 -1498 7294 -1486
rect 7228 -1578 7244 -1498
rect 7278 -1578 7294 -1498
rect 7228 -1590 7294 -1578
rect 7324 -1498 7390 -1486
rect 7324 -1578 7340 -1498
rect 7374 -1578 7390 -1498
rect 7324 -1590 7390 -1578
rect 7420 -1498 7486 -1486
rect 7420 -1578 7436 -1498
rect 7470 -1578 7486 -1498
rect 7420 -1590 7486 -1578
rect 7516 -1498 7582 -1486
rect 7516 -1578 7532 -1498
rect 7566 -1578 7582 -1498
rect 7516 -1590 7582 -1578
rect 7612 -1498 7678 -1486
rect 7612 -1578 7628 -1498
rect 7662 -1578 7678 -1498
rect 7612 -1590 7678 -1578
rect 7708 -1498 7774 -1486
rect 7708 -1578 7724 -1498
rect 7758 -1578 7774 -1498
rect 7708 -1590 7774 -1578
rect 7804 -1498 7870 -1486
rect 7804 -1578 7820 -1498
rect 7854 -1578 7870 -1498
rect 7804 -1590 7870 -1578
rect 7900 -1498 7966 -1486
rect 7900 -1578 7916 -1498
rect 7950 -1578 7966 -1498
rect 7900 -1590 7966 -1578
rect 7996 -1498 8058 -1486
rect 7996 -1578 8012 -1498
rect 8046 -1578 8058 -1498
rect 7996 -1590 8058 -1578
<< pdiff >>
rect -1960 8082 -1898 8094
rect -1960 7834 -1948 8082
rect -1914 7834 -1898 8082
rect -1960 7822 -1898 7834
rect -1868 8082 -1802 8094
rect -1868 7834 -1852 8082
rect -1818 7834 -1802 8082
rect -1868 7822 -1802 7834
rect -1772 8082 -1706 8094
rect -1772 7834 -1756 8082
rect -1722 7834 -1706 8082
rect -1772 7822 -1706 7834
rect -1676 8082 -1610 8094
rect -1676 7834 -1660 8082
rect -1626 7834 -1610 8082
rect -1676 7822 -1610 7834
rect -1580 8082 -1514 8094
rect -1580 7834 -1564 8082
rect -1530 7834 -1514 8082
rect -1580 7822 -1514 7834
rect -1484 8082 -1418 8094
rect -1484 7834 -1468 8082
rect -1434 7834 -1418 8082
rect -1484 7822 -1418 7834
rect -1388 8082 -1322 8094
rect -1388 7834 -1372 8082
rect -1338 7834 -1322 8082
rect -1388 7822 -1322 7834
rect -1292 8082 -1226 8094
rect -1292 7834 -1276 8082
rect -1242 7834 -1226 8082
rect -1292 7822 -1226 7834
rect -1196 8082 -1130 8094
rect -1196 7834 -1180 8082
rect -1146 7834 -1130 8082
rect -1196 7822 -1130 7834
rect -1100 8082 -1034 8094
rect -1100 7834 -1084 8082
rect -1050 7834 -1034 8082
rect -1100 7822 -1034 7834
rect -1004 8082 -942 8094
rect -1004 7834 -988 8082
rect -954 7834 -942 8082
rect -1004 7822 -942 7834
rect 7040 8082 7102 8094
rect 7040 7834 7052 8082
rect 7086 7834 7102 8082
rect 7040 7822 7102 7834
rect 7132 8082 7198 8094
rect 7132 7834 7148 8082
rect 7182 7834 7198 8082
rect 7132 7822 7198 7834
rect 7228 8082 7294 8094
rect 7228 7834 7244 8082
rect 7278 7834 7294 8082
rect 7228 7822 7294 7834
rect 7324 8082 7390 8094
rect 7324 7834 7340 8082
rect 7374 7834 7390 8082
rect 7324 7822 7390 7834
rect 7420 8082 7486 8094
rect 7420 7834 7436 8082
rect 7470 7834 7486 8082
rect 7420 7822 7486 7834
rect 7516 8082 7582 8094
rect 7516 7834 7532 8082
rect 7566 7834 7582 8082
rect 7516 7822 7582 7834
rect 7612 8082 7678 8094
rect 7612 7834 7628 8082
rect 7662 7834 7678 8082
rect 7612 7822 7678 7834
rect 7708 8082 7774 8094
rect 7708 7834 7724 8082
rect 7758 7834 7774 8082
rect 7708 7822 7774 7834
rect 7804 8082 7870 8094
rect 7804 7834 7820 8082
rect 7854 7834 7870 8082
rect 7804 7822 7870 7834
rect 7900 8082 7966 8094
rect 7900 7834 7916 8082
rect 7950 7834 7966 8082
rect 7900 7822 7966 7834
rect 7996 8082 8058 8094
rect 7996 7834 8012 8082
rect 8046 7834 8058 8082
rect 7996 7822 8058 7834
rect -1960 6282 -1898 6294
rect -1960 6034 -1948 6282
rect -1914 6034 -1898 6282
rect -1960 6022 -1898 6034
rect -1868 6282 -1802 6294
rect -1868 6034 -1852 6282
rect -1818 6034 -1802 6282
rect -1868 6022 -1802 6034
rect -1772 6282 -1706 6294
rect -1772 6034 -1756 6282
rect -1722 6034 -1706 6282
rect -1772 6022 -1706 6034
rect -1676 6282 -1610 6294
rect -1676 6034 -1660 6282
rect -1626 6034 -1610 6282
rect -1676 6022 -1610 6034
rect -1580 6282 -1514 6294
rect -1580 6034 -1564 6282
rect -1530 6034 -1514 6282
rect -1580 6022 -1514 6034
rect -1484 6282 -1418 6294
rect -1484 6034 -1468 6282
rect -1434 6034 -1418 6282
rect -1484 6022 -1418 6034
rect -1388 6282 -1322 6294
rect -1388 6034 -1372 6282
rect -1338 6034 -1322 6282
rect -1388 6022 -1322 6034
rect -1292 6282 -1226 6294
rect -1292 6034 -1276 6282
rect -1242 6034 -1226 6282
rect -1292 6022 -1226 6034
rect -1196 6282 -1130 6294
rect -1196 6034 -1180 6282
rect -1146 6034 -1130 6282
rect -1196 6022 -1130 6034
rect -1100 6282 -1034 6294
rect -1100 6034 -1084 6282
rect -1050 6034 -1034 6282
rect -1100 6022 -1034 6034
rect -1004 6282 -942 6294
rect -1004 6034 -988 6282
rect -954 6034 -942 6282
rect -1004 6022 -942 6034
rect 7040 6282 7102 6294
rect 7040 6034 7052 6282
rect 7086 6034 7102 6282
rect 7040 6022 7102 6034
rect 7132 6282 7198 6294
rect 7132 6034 7148 6282
rect 7182 6034 7198 6282
rect 7132 6022 7198 6034
rect 7228 6282 7294 6294
rect 7228 6034 7244 6282
rect 7278 6034 7294 6282
rect 7228 6022 7294 6034
rect 7324 6282 7390 6294
rect 7324 6034 7340 6282
rect 7374 6034 7390 6282
rect 7324 6022 7390 6034
rect 7420 6282 7486 6294
rect 7420 6034 7436 6282
rect 7470 6034 7486 6282
rect 7420 6022 7486 6034
rect 7516 6282 7582 6294
rect 7516 6034 7532 6282
rect 7566 6034 7582 6282
rect 7516 6022 7582 6034
rect 7612 6282 7678 6294
rect 7612 6034 7628 6282
rect 7662 6034 7678 6282
rect 7612 6022 7678 6034
rect 7708 6282 7774 6294
rect 7708 6034 7724 6282
rect 7758 6034 7774 6282
rect 7708 6022 7774 6034
rect 7804 6282 7870 6294
rect 7804 6034 7820 6282
rect 7854 6034 7870 6282
rect 7804 6022 7870 6034
rect 7900 6282 7966 6294
rect 7900 6034 7916 6282
rect 7950 6034 7966 6282
rect 7900 6022 7966 6034
rect 7996 6282 8058 6294
rect 7996 6034 8012 6282
rect 8046 6034 8058 6282
rect 7996 6022 8058 6034
rect -1960 4482 -1898 4494
rect -1960 4234 -1948 4482
rect -1914 4234 -1898 4482
rect -1960 4222 -1898 4234
rect -1868 4482 -1802 4494
rect -1868 4234 -1852 4482
rect -1818 4234 -1802 4482
rect -1868 4222 -1802 4234
rect -1772 4482 -1706 4494
rect -1772 4234 -1756 4482
rect -1722 4234 -1706 4482
rect -1772 4222 -1706 4234
rect -1676 4482 -1610 4494
rect -1676 4234 -1660 4482
rect -1626 4234 -1610 4482
rect -1676 4222 -1610 4234
rect -1580 4482 -1514 4494
rect -1580 4234 -1564 4482
rect -1530 4234 -1514 4482
rect -1580 4222 -1514 4234
rect -1484 4482 -1418 4494
rect -1484 4234 -1468 4482
rect -1434 4234 -1418 4482
rect -1484 4222 -1418 4234
rect -1388 4482 -1322 4494
rect -1388 4234 -1372 4482
rect -1338 4234 -1322 4482
rect -1388 4222 -1322 4234
rect -1292 4482 -1226 4494
rect -1292 4234 -1276 4482
rect -1242 4234 -1226 4482
rect -1292 4222 -1226 4234
rect -1196 4482 -1130 4494
rect -1196 4234 -1180 4482
rect -1146 4234 -1130 4482
rect -1196 4222 -1130 4234
rect -1100 4482 -1034 4494
rect -1100 4234 -1084 4482
rect -1050 4234 -1034 4482
rect -1100 4222 -1034 4234
rect -1004 4482 -942 4494
rect -1004 4234 -988 4482
rect -954 4234 -942 4482
rect -1004 4222 -942 4234
rect 7040 4482 7102 4494
rect 7040 4234 7052 4482
rect 7086 4234 7102 4482
rect 7040 4222 7102 4234
rect 7132 4482 7198 4494
rect 7132 4234 7148 4482
rect 7182 4234 7198 4482
rect 7132 4222 7198 4234
rect 7228 4482 7294 4494
rect 7228 4234 7244 4482
rect 7278 4234 7294 4482
rect 7228 4222 7294 4234
rect 7324 4482 7390 4494
rect 7324 4234 7340 4482
rect 7374 4234 7390 4482
rect 7324 4222 7390 4234
rect 7420 4482 7486 4494
rect 7420 4234 7436 4482
rect 7470 4234 7486 4482
rect 7420 4222 7486 4234
rect 7516 4482 7582 4494
rect 7516 4234 7532 4482
rect 7566 4234 7582 4482
rect 7516 4222 7582 4234
rect 7612 4482 7678 4494
rect 7612 4234 7628 4482
rect 7662 4234 7678 4482
rect 7612 4222 7678 4234
rect 7708 4482 7774 4494
rect 7708 4234 7724 4482
rect 7758 4234 7774 4482
rect 7708 4222 7774 4234
rect 7804 4482 7870 4494
rect 7804 4234 7820 4482
rect 7854 4234 7870 4482
rect 7804 4222 7870 4234
rect 7900 4482 7966 4494
rect 7900 4234 7916 4482
rect 7950 4234 7966 4482
rect 7900 4222 7966 4234
rect 7996 4482 8058 4494
rect 7996 4234 8012 4482
rect 8046 4234 8058 4482
rect 7996 4222 8058 4234
rect -1960 2682 -1898 2694
rect -1960 2434 -1948 2682
rect -1914 2434 -1898 2682
rect -1960 2422 -1898 2434
rect -1868 2682 -1802 2694
rect -1868 2434 -1852 2682
rect -1818 2434 -1802 2682
rect -1868 2422 -1802 2434
rect -1772 2682 -1706 2694
rect -1772 2434 -1756 2682
rect -1722 2434 -1706 2682
rect -1772 2422 -1706 2434
rect -1676 2682 -1610 2694
rect -1676 2434 -1660 2682
rect -1626 2434 -1610 2682
rect -1676 2422 -1610 2434
rect -1580 2682 -1514 2694
rect -1580 2434 -1564 2682
rect -1530 2434 -1514 2682
rect -1580 2422 -1514 2434
rect -1484 2682 -1418 2694
rect -1484 2434 -1468 2682
rect -1434 2434 -1418 2682
rect -1484 2422 -1418 2434
rect -1388 2682 -1322 2694
rect -1388 2434 -1372 2682
rect -1338 2434 -1322 2682
rect -1388 2422 -1322 2434
rect -1292 2682 -1226 2694
rect -1292 2434 -1276 2682
rect -1242 2434 -1226 2682
rect -1292 2422 -1226 2434
rect -1196 2682 -1130 2694
rect -1196 2434 -1180 2682
rect -1146 2434 -1130 2682
rect -1196 2422 -1130 2434
rect -1100 2682 -1034 2694
rect -1100 2434 -1084 2682
rect -1050 2434 -1034 2682
rect -1100 2422 -1034 2434
rect -1004 2682 -942 2694
rect -1004 2434 -988 2682
rect -954 2434 -942 2682
rect -1004 2422 -942 2434
rect 7040 2682 7102 2694
rect 7040 2434 7052 2682
rect 7086 2434 7102 2682
rect 7040 2422 7102 2434
rect 7132 2682 7198 2694
rect 7132 2434 7148 2682
rect 7182 2434 7198 2682
rect 7132 2422 7198 2434
rect 7228 2682 7294 2694
rect 7228 2434 7244 2682
rect 7278 2434 7294 2682
rect 7228 2422 7294 2434
rect 7324 2682 7390 2694
rect 7324 2434 7340 2682
rect 7374 2434 7390 2682
rect 7324 2422 7390 2434
rect 7420 2682 7486 2694
rect 7420 2434 7436 2682
rect 7470 2434 7486 2682
rect 7420 2422 7486 2434
rect 7516 2682 7582 2694
rect 7516 2434 7532 2682
rect 7566 2434 7582 2682
rect 7516 2422 7582 2434
rect 7612 2682 7678 2694
rect 7612 2434 7628 2682
rect 7662 2434 7678 2682
rect 7612 2422 7678 2434
rect 7708 2682 7774 2694
rect 7708 2434 7724 2682
rect 7758 2434 7774 2682
rect 7708 2422 7774 2434
rect 7804 2682 7870 2694
rect 7804 2434 7820 2682
rect 7854 2434 7870 2682
rect 7804 2422 7870 2434
rect 7900 2682 7966 2694
rect 7900 2434 7916 2682
rect 7950 2434 7966 2682
rect 7900 2422 7966 2434
rect 7996 2682 8058 2694
rect 7996 2434 8012 2682
rect 8046 2434 8058 2682
rect 7996 2422 8058 2434
rect -1960 882 -1898 894
rect -1960 634 -1948 882
rect -1914 634 -1898 882
rect -1960 622 -1898 634
rect -1868 882 -1802 894
rect -1868 634 -1852 882
rect -1818 634 -1802 882
rect -1868 622 -1802 634
rect -1772 882 -1706 894
rect -1772 634 -1756 882
rect -1722 634 -1706 882
rect -1772 622 -1706 634
rect -1676 882 -1610 894
rect -1676 634 -1660 882
rect -1626 634 -1610 882
rect -1676 622 -1610 634
rect -1580 882 -1514 894
rect -1580 634 -1564 882
rect -1530 634 -1514 882
rect -1580 622 -1514 634
rect -1484 882 -1418 894
rect -1484 634 -1468 882
rect -1434 634 -1418 882
rect -1484 622 -1418 634
rect -1388 882 -1322 894
rect -1388 634 -1372 882
rect -1338 634 -1322 882
rect -1388 622 -1322 634
rect -1292 882 -1226 894
rect -1292 634 -1276 882
rect -1242 634 -1226 882
rect -1292 622 -1226 634
rect -1196 882 -1130 894
rect -1196 634 -1180 882
rect -1146 634 -1130 882
rect -1196 622 -1130 634
rect -1100 882 -1034 894
rect -1100 634 -1084 882
rect -1050 634 -1034 882
rect -1100 622 -1034 634
rect -1004 882 -942 894
rect -1004 634 -988 882
rect -954 634 -942 882
rect -1004 622 -942 634
rect 7040 882 7102 894
rect 7040 634 7052 882
rect 7086 634 7102 882
rect 7040 622 7102 634
rect 7132 882 7198 894
rect 7132 634 7148 882
rect 7182 634 7198 882
rect 7132 622 7198 634
rect 7228 882 7294 894
rect 7228 634 7244 882
rect 7278 634 7294 882
rect 7228 622 7294 634
rect 7324 882 7390 894
rect 7324 634 7340 882
rect 7374 634 7390 882
rect 7324 622 7390 634
rect 7420 882 7486 894
rect 7420 634 7436 882
rect 7470 634 7486 882
rect 7420 622 7486 634
rect 7516 882 7582 894
rect 7516 634 7532 882
rect 7566 634 7582 882
rect 7516 622 7582 634
rect 7612 882 7678 894
rect 7612 634 7628 882
rect 7662 634 7678 882
rect 7612 622 7678 634
rect 7708 882 7774 894
rect 7708 634 7724 882
rect 7758 634 7774 882
rect 7708 622 7774 634
rect 7804 882 7870 894
rect 7804 634 7820 882
rect 7854 634 7870 882
rect 7804 622 7870 634
rect 7900 882 7966 894
rect 7900 634 7916 882
rect 7950 634 7966 882
rect 7900 622 7966 634
rect 7996 882 8058 894
rect 7996 634 8012 882
rect 8046 634 8058 882
rect 7996 622 8058 634
rect -1960 -918 -1898 -906
rect -1960 -1166 -1948 -918
rect -1914 -1166 -1898 -918
rect -1960 -1178 -1898 -1166
rect -1868 -918 -1802 -906
rect -1868 -1166 -1852 -918
rect -1818 -1166 -1802 -918
rect -1868 -1178 -1802 -1166
rect -1772 -918 -1706 -906
rect -1772 -1166 -1756 -918
rect -1722 -1166 -1706 -918
rect -1772 -1178 -1706 -1166
rect -1676 -918 -1610 -906
rect -1676 -1166 -1660 -918
rect -1626 -1166 -1610 -918
rect -1676 -1178 -1610 -1166
rect -1580 -918 -1514 -906
rect -1580 -1166 -1564 -918
rect -1530 -1166 -1514 -918
rect -1580 -1178 -1514 -1166
rect -1484 -918 -1418 -906
rect -1484 -1166 -1468 -918
rect -1434 -1166 -1418 -918
rect -1484 -1178 -1418 -1166
rect -1388 -918 -1322 -906
rect -1388 -1166 -1372 -918
rect -1338 -1166 -1322 -918
rect -1388 -1178 -1322 -1166
rect -1292 -918 -1226 -906
rect -1292 -1166 -1276 -918
rect -1242 -1166 -1226 -918
rect -1292 -1178 -1226 -1166
rect -1196 -918 -1130 -906
rect -1196 -1166 -1180 -918
rect -1146 -1166 -1130 -918
rect -1196 -1178 -1130 -1166
rect -1100 -918 -1034 -906
rect -1100 -1166 -1084 -918
rect -1050 -1166 -1034 -918
rect -1100 -1178 -1034 -1166
rect -1004 -918 -942 -906
rect -1004 -1166 -988 -918
rect -954 -1166 -942 -918
rect -1004 -1178 -942 -1166
rect 7040 -918 7102 -906
rect 7040 -1166 7052 -918
rect 7086 -1166 7102 -918
rect 7040 -1178 7102 -1166
rect 7132 -918 7198 -906
rect 7132 -1166 7148 -918
rect 7182 -1166 7198 -918
rect 7132 -1178 7198 -1166
rect 7228 -918 7294 -906
rect 7228 -1166 7244 -918
rect 7278 -1166 7294 -918
rect 7228 -1178 7294 -1166
rect 7324 -918 7390 -906
rect 7324 -1166 7340 -918
rect 7374 -1166 7390 -918
rect 7324 -1178 7390 -1166
rect 7420 -918 7486 -906
rect 7420 -1166 7436 -918
rect 7470 -1166 7486 -918
rect 7420 -1178 7486 -1166
rect 7516 -918 7582 -906
rect 7516 -1166 7532 -918
rect 7566 -1166 7582 -918
rect 7516 -1178 7582 -1166
rect 7612 -918 7678 -906
rect 7612 -1166 7628 -918
rect 7662 -1166 7678 -918
rect 7612 -1178 7678 -1166
rect 7708 -918 7774 -906
rect 7708 -1166 7724 -918
rect 7758 -1166 7774 -918
rect 7708 -1178 7774 -1166
rect 7804 -918 7870 -906
rect 7804 -1166 7820 -918
rect 7854 -1166 7870 -918
rect 7804 -1178 7870 -1166
rect 7900 -918 7966 -906
rect 7900 -1166 7916 -918
rect 7950 -1166 7966 -918
rect 7900 -1178 7966 -1166
rect 7996 -918 8058 -906
rect 7996 -1166 8012 -918
rect 8046 -1166 8058 -918
rect 7996 -1178 8058 -1166
<< ndiffc >>
rect -1948 7422 -1914 7502
rect -1852 7422 -1818 7502
rect -1756 7422 -1722 7502
rect -1660 7422 -1626 7502
rect -1564 7422 -1530 7502
rect -1468 7422 -1434 7502
rect -1372 7422 -1338 7502
rect -1276 7422 -1242 7502
rect -1180 7422 -1146 7502
rect -1084 7422 -1050 7502
rect -988 7422 -954 7502
rect 7052 7422 7086 7502
rect 7148 7422 7182 7502
rect 7244 7422 7278 7502
rect 7340 7422 7374 7502
rect 7436 7422 7470 7502
rect 7532 7422 7566 7502
rect 7628 7422 7662 7502
rect 7724 7422 7758 7502
rect 7820 7422 7854 7502
rect 7916 7422 7950 7502
rect 8012 7422 8046 7502
rect -1948 5622 -1914 5702
rect -1852 5622 -1818 5702
rect -1756 5622 -1722 5702
rect -1660 5622 -1626 5702
rect -1564 5622 -1530 5702
rect -1468 5622 -1434 5702
rect -1372 5622 -1338 5702
rect -1276 5622 -1242 5702
rect -1180 5622 -1146 5702
rect -1084 5622 -1050 5702
rect -988 5622 -954 5702
rect 7052 5622 7086 5702
rect 7148 5622 7182 5702
rect 7244 5622 7278 5702
rect 7340 5622 7374 5702
rect 7436 5622 7470 5702
rect 7532 5622 7566 5702
rect 7628 5622 7662 5702
rect 7724 5622 7758 5702
rect 7820 5622 7854 5702
rect 7916 5622 7950 5702
rect 8012 5622 8046 5702
rect -1948 3822 -1914 3902
rect -1852 3822 -1818 3902
rect -1756 3822 -1722 3902
rect -1660 3822 -1626 3902
rect -1564 3822 -1530 3902
rect -1468 3822 -1434 3902
rect -1372 3822 -1338 3902
rect -1276 3822 -1242 3902
rect -1180 3822 -1146 3902
rect -1084 3822 -1050 3902
rect -988 3822 -954 3902
rect 7052 3822 7086 3902
rect 7148 3822 7182 3902
rect 7244 3822 7278 3902
rect 7340 3822 7374 3902
rect 7436 3822 7470 3902
rect 7532 3822 7566 3902
rect 7628 3822 7662 3902
rect 7724 3822 7758 3902
rect 7820 3822 7854 3902
rect 7916 3822 7950 3902
rect 8012 3822 8046 3902
rect -1948 2022 -1914 2102
rect -1852 2022 -1818 2102
rect -1756 2022 -1722 2102
rect -1660 2022 -1626 2102
rect -1564 2022 -1530 2102
rect -1468 2022 -1434 2102
rect -1372 2022 -1338 2102
rect -1276 2022 -1242 2102
rect -1180 2022 -1146 2102
rect -1084 2022 -1050 2102
rect -988 2022 -954 2102
rect 7052 2022 7086 2102
rect 7148 2022 7182 2102
rect 7244 2022 7278 2102
rect 7340 2022 7374 2102
rect 7436 2022 7470 2102
rect 7532 2022 7566 2102
rect 7628 2022 7662 2102
rect 7724 2022 7758 2102
rect 7820 2022 7854 2102
rect 7916 2022 7950 2102
rect 8012 2022 8046 2102
rect -1948 222 -1914 302
rect -1852 222 -1818 302
rect -1756 222 -1722 302
rect -1660 222 -1626 302
rect -1564 222 -1530 302
rect -1468 222 -1434 302
rect -1372 222 -1338 302
rect -1276 222 -1242 302
rect -1180 222 -1146 302
rect -1084 222 -1050 302
rect -988 222 -954 302
rect 7052 222 7086 302
rect 7148 222 7182 302
rect 7244 222 7278 302
rect 7340 222 7374 302
rect 7436 222 7470 302
rect 7532 222 7566 302
rect 7628 222 7662 302
rect 7724 222 7758 302
rect 7820 222 7854 302
rect 7916 222 7950 302
rect 8012 222 8046 302
rect -1948 -1578 -1914 -1498
rect -1852 -1578 -1818 -1498
rect -1756 -1578 -1722 -1498
rect -1660 -1578 -1626 -1498
rect -1564 -1578 -1530 -1498
rect -1468 -1578 -1434 -1498
rect -1372 -1578 -1338 -1498
rect -1276 -1578 -1242 -1498
rect -1180 -1578 -1146 -1498
rect -1084 -1578 -1050 -1498
rect -988 -1578 -954 -1498
rect 7052 -1578 7086 -1498
rect 7148 -1578 7182 -1498
rect 7244 -1578 7278 -1498
rect 7340 -1578 7374 -1498
rect 7436 -1578 7470 -1498
rect 7532 -1578 7566 -1498
rect 7628 -1578 7662 -1498
rect 7724 -1578 7758 -1498
rect 7820 -1578 7854 -1498
rect 7916 -1578 7950 -1498
rect 8012 -1578 8046 -1498
<< pdiffc >>
rect -1948 7834 -1914 8082
rect -1852 7834 -1818 8082
rect -1756 7834 -1722 8082
rect -1660 7834 -1626 8082
rect -1564 7834 -1530 8082
rect -1468 7834 -1434 8082
rect -1372 7834 -1338 8082
rect -1276 7834 -1242 8082
rect -1180 7834 -1146 8082
rect -1084 7834 -1050 8082
rect -988 7834 -954 8082
rect 7052 7834 7086 8082
rect 7148 7834 7182 8082
rect 7244 7834 7278 8082
rect 7340 7834 7374 8082
rect 7436 7834 7470 8082
rect 7532 7834 7566 8082
rect 7628 7834 7662 8082
rect 7724 7834 7758 8082
rect 7820 7834 7854 8082
rect 7916 7834 7950 8082
rect 8012 7834 8046 8082
rect -1948 6034 -1914 6282
rect -1852 6034 -1818 6282
rect -1756 6034 -1722 6282
rect -1660 6034 -1626 6282
rect -1564 6034 -1530 6282
rect -1468 6034 -1434 6282
rect -1372 6034 -1338 6282
rect -1276 6034 -1242 6282
rect -1180 6034 -1146 6282
rect -1084 6034 -1050 6282
rect -988 6034 -954 6282
rect 7052 6034 7086 6282
rect 7148 6034 7182 6282
rect 7244 6034 7278 6282
rect 7340 6034 7374 6282
rect 7436 6034 7470 6282
rect 7532 6034 7566 6282
rect 7628 6034 7662 6282
rect 7724 6034 7758 6282
rect 7820 6034 7854 6282
rect 7916 6034 7950 6282
rect 8012 6034 8046 6282
rect -1948 4234 -1914 4482
rect -1852 4234 -1818 4482
rect -1756 4234 -1722 4482
rect -1660 4234 -1626 4482
rect -1564 4234 -1530 4482
rect -1468 4234 -1434 4482
rect -1372 4234 -1338 4482
rect -1276 4234 -1242 4482
rect -1180 4234 -1146 4482
rect -1084 4234 -1050 4482
rect -988 4234 -954 4482
rect 7052 4234 7086 4482
rect 7148 4234 7182 4482
rect 7244 4234 7278 4482
rect 7340 4234 7374 4482
rect 7436 4234 7470 4482
rect 7532 4234 7566 4482
rect 7628 4234 7662 4482
rect 7724 4234 7758 4482
rect 7820 4234 7854 4482
rect 7916 4234 7950 4482
rect 8012 4234 8046 4482
rect -1948 2434 -1914 2682
rect -1852 2434 -1818 2682
rect -1756 2434 -1722 2682
rect -1660 2434 -1626 2682
rect -1564 2434 -1530 2682
rect -1468 2434 -1434 2682
rect -1372 2434 -1338 2682
rect -1276 2434 -1242 2682
rect -1180 2434 -1146 2682
rect -1084 2434 -1050 2682
rect -988 2434 -954 2682
rect 7052 2434 7086 2682
rect 7148 2434 7182 2682
rect 7244 2434 7278 2682
rect 7340 2434 7374 2682
rect 7436 2434 7470 2682
rect 7532 2434 7566 2682
rect 7628 2434 7662 2682
rect 7724 2434 7758 2682
rect 7820 2434 7854 2682
rect 7916 2434 7950 2682
rect 8012 2434 8046 2682
rect -1948 634 -1914 882
rect -1852 634 -1818 882
rect -1756 634 -1722 882
rect -1660 634 -1626 882
rect -1564 634 -1530 882
rect -1468 634 -1434 882
rect -1372 634 -1338 882
rect -1276 634 -1242 882
rect -1180 634 -1146 882
rect -1084 634 -1050 882
rect -988 634 -954 882
rect 7052 634 7086 882
rect 7148 634 7182 882
rect 7244 634 7278 882
rect 7340 634 7374 882
rect 7436 634 7470 882
rect 7532 634 7566 882
rect 7628 634 7662 882
rect 7724 634 7758 882
rect 7820 634 7854 882
rect 7916 634 7950 882
rect 8012 634 8046 882
rect -1948 -1166 -1914 -918
rect -1852 -1166 -1818 -918
rect -1756 -1166 -1722 -918
rect -1660 -1166 -1626 -918
rect -1564 -1166 -1530 -918
rect -1468 -1166 -1434 -918
rect -1372 -1166 -1338 -918
rect -1276 -1166 -1242 -918
rect -1180 -1166 -1146 -918
rect -1084 -1166 -1050 -918
rect -988 -1166 -954 -918
rect 7052 -1166 7086 -918
rect 7148 -1166 7182 -918
rect 7244 -1166 7278 -918
rect 7340 -1166 7374 -918
rect 7436 -1166 7470 -918
rect 7532 -1166 7566 -918
rect 7628 -1166 7662 -918
rect 7724 -1166 7758 -918
rect 7820 -1166 7854 -918
rect 7916 -1166 7950 -918
rect 8012 -1166 8046 -918
<< psubdiff >>
rect -2062 7592 -1966 7626
rect -936 7592 -840 7626
rect -2062 7530 -2028 7592
rect -874 7530 -840 7592
rect -2062 7270 -2028 7332
rect -874 7270 -840 7332
rect -2062 7236 -1966 7270
rect -936 7236 -840 7270
rect 6938 7592 7034 7626
rect 8064 7592 8160 7626
rect 6938 7530 6972 7592
rect 8126 7530 8160 7592
rect 6938 7270 6972 7332
rect 8126 7270 8160 7332
rect 6938 7236 7034 7270
rect 8064 7236 8160 7270
rect -2062 5792 -1966 5826
rect -936 5792 -840 5826
rect -2062 5730 -2028 5792
rect -874 5730 -840 5792
rect -2062 5470 -2028 5532
rect -874 5470 -840 5532
rect -2062 5436 -1966 5470
rect -936 5436 -840 5470
rect 6938 5792 7034 5826
rect 8064 5792 8160 5826
rect 6938 5730 6972 5792
rect 8126 5730 8160 5792
rect 6938 5470 6972 5532
rect 8126 5470 8160 5532
rect 6938 5436 7034 5470
rect 8064 5436 8160 5470
rect -2062 3992 -1966 4026
rect -936 3992 -840 4026
rect -2062 3930 -2028 3992
rect -874 3930 -840 3992
rect -2062 3670 -2028 3732
rect -874 3670 -840 3732
rect -2062 3636 -1966 3670
rect -936 3636 -840 3670
rect 6938 3992 7034 4026
rect 8064 3992 8160 4026
rect 6938 3930 6972 3992
rect 8126 3930 8160 3992
rect 6938 3670 6972 3732
rect 8126 3670 8160 3732
rect 6938 3636 7034 3670
rect 8064 3636 8160 3670
rect -2062 2192 -1966 2226
rect -936 2192 -840 2226
rect -2062 2130 -2028 2192
rect -874 2130 -840 2192
rect -2062 1870 -2028 1932
rect -874 1870 -840 1932
rect -2062 1836 -1966 1870
rect -936 1836 -840 1870
rect 6938 2192 7034 2226
rect 8064 2192 8160 2226
rect 6938 2130 6972 2192
rect 8126 2130 8160 2192
rect 6938 1870 6972 1932
rect 8126 1870 8160 1932
rect 6938 1836 7034 1870
rect 8064 1836 8160 1870
rect -2062 392 -1966 426
rect -936 392 -840 426
rect -2062 330 -2028 392
rect -874 330 -840 392
rect -2062 70 -2028 132
rect -874 70 -840 132
rect -2062 36 -1966 70
rect -936 36 -840 70
rect 6938 392 7034 426
rect 8064 392 8160 426
rect 6938 330 6972 392
rect 8126 330 8160 392
rect 6938 70 6972 132
rect 8126 70 8160 132
rect 6938 36 7034 70
rect 8064 36 8160 70
rect -2062 -1408 -1966 -1374
rect -936 -1408 -840 -1374
rect -2062 -1470 -2028 -1408
rect -874 -1470 -840 -1408
rect -2062 -1730 -2028 -1668
rect -874 -1730 -840 -1668
rect -2062 -1764 -1966 -1730
rect -936 -1764 -840 -1730
rect 6938 -1408 7034 -1374
rect 8064 -1408 8160 -1374
rect 6938 -1470 6972 -1408
rect 8126 -1470 8160 -1408
rect 6938 -1730 6972 -1668
rect 8126 -1730 8160 -1668
rect 6938 -1764 7034 -1730
rect 8064 -1764 8160 -1730
<< nsubdiff >>
rect -2062 8244 -1966 8278
rect -936 8244 -840 8278
rect -2062 8182 -2028 8244
rect -874 8182 -840 8244
rect -2062 7734 -2028 7796
rect -874 7734 -840 7796
rect -2062 7700 -1966 7734
rect -936 7700 -840 7734
rect 6938 8244 7034 8278
rect 8064 8244 8160 8278
rect 6938 8182 6972 8244
rect 8126 8182 8160 8244
rect 6938 7734 6972 7796
rect 8126 7734 8160 7796
rect 6938 7700 7034 7734
rect 8064 7700 8160 7734
rect -2062 6444 -1966 6478
rect -936 6444 -840 6478
rect -2062 6382 -2028 6444
rect -874 6382 -840 6444
rect -2062 5934 -2028 5996
rect -874 5934 -840 5996
rect -2062 5900 -1966 5934
rect -936 5900 -840 5934
rect 6938 6444 7034 6478
rect 8064 6444 8160 6478
rect 6938 6382 6972 6444
rect 8126 6382 8160 6444
rect 6938 5934 6972 5996
rect 8126 5934 8160 5996
rect 6938 5900 7034 5934
rect 8064 5900 8160 5934
rect -2062 4644 -1966 4678
rect -936 4644 -840 4678
rect -2062 4582 -2028 4644
rect -874 4582 -840 4644
rect -2062 4134 -2028 4196
rect -874 4134 -840 4196
rect -2062 4100 -1966 4134
rect -936 4100 -840 4134
rect 6938 4644 7034 4678
rect 8064 4644 8160 4678
rect 6938 4582 6972 4644
rect 8126 4582 8160 4644
rect 6938 4134 6972 4196
rect 8126 4134 8160 4196
rect 6938 4100 7034 4134
rect 8064 4100 8160 4134
rect -2062 2844 -1966 2878
rect -936 2844 -840 2878
rect -2062 2782 -2028 2844
rect -874 2782 -840 2844
rect -2062 2334 -2028 2396
rect -874 2334 -840 2396
rect -2062 2300 -1966 2334
rect -936 2300 -840 2334
rect 6938 2844 7034 2878
rect 8064 2844 8160 2878
rect 6938 2782 6972 2844
rect 8126 2782 8160 2844
rect 6938 2334 6972 2396
rect 8126 2334 8160 2396
rect 6938 2300 7034 2334
rect 8064 2300 8160 2334
rect -2062 1044 -1966 1078
rect -936 1044 -840 1078
rect -2062 982 -2028 1044
rect -874 982 -840 1044
rect -2062 534 -2028 596
rect -874 534 -840 596
rect -2062 500 -1966 534
rect -936 500 -840 534
rect 6938 1044 7034 1078
rect 8064 1044 8160 1078
rect 6938 982 6972 1044
rect 8126 982 8160 1044
rect 6938 534 6972 596
rect 8126 534 8160 596
rect 6938 500 7034 534
rect 8064 500 8160 534
rect -2062 -756 -1966 -722
rect -936 -756 -840 -722
rect -2062 -818 -2028 -756
rect -874 -818 -840 -756
rect -2062 -1266 -2028 -1204
rect -874 -1266 -840 -1204
rect -2062 -1300 -1966 -1266
rect -936 -1300 -840 -1266
rect 6938 -756 7034 -722
rect 8064 -756 8160 -722
rect 6938 -818 6972 -756
rect 8126 -818 8160 -756
rect 6938 -1266 6972 -1204
rect 8126 -1266 8160 -1204
rect 6938 -1300 7034 -1266
rect 8064 -1300 8160 -1266
<< psubdiffcont >>
rect -1966 7592 -936 7626
rect -2062 7332 -2028 7530
rect -874 7332 -840 7530
rect -1966 7236 -936 7270
rect 7034 7592 8064 7626
rect 6938 7332 6972 7530
rect 8126 7332 8160 7530
rect 7034 7236 8064 7270
rect -1966 5792 -936 5826
rect -2062 5532 -2028 5730
rect -874 5532 -840 5730
rect -1966 5436 -936 5470
rect 7034 5792 8064 5826
rect 6938 5532 6972 5730
rect 8126 5532 8160 5730
rect 7034 5436 8064 5470
rect -1966 3992 -936 4026
rect -2062 3732 -2028 3930
rect -874 3732 -840 3930
rect -1966 3636 -936 3670
rect 7034 3992 8064 4026
rect 6938 3732 6972 3930
rect 8126 3732 8160 3930
rect 7034 3636 8064 3670
rect -1966 2192 -936 2226
rect -2062 1932 -2028 2130
rect -874 1932 -840 2130
rect -1966 1836 -936 1870
rect 7034 2192 8064 2226
rect 6938 1932 6972 2130
rect 8126 1932 8160 2130
rect 7034 1836 8064 1870
rect -1966 392 -936 426
rect -2062 132 -2028 330
rect -874 132 -840 330
rect -1966 36 -936 70
rect 7034 392 8064 426
rect 6938 132 6972 330
rect 8126 132 8160 330
rect 7034 36 8064 70
rect -1966 -1408 -936 -1374
rect -2062 -1668 -2028 -1470
rect -874 -1668 -840 -1470
rect -1966 -1764 -936 -1730
rect 7034 -1408 8064 -1374
rect 6938 -1668 6972 -1470
rect 8126 -1668 8160 -1470
rect 7034 -1764 8064 -1730
<< nsubdiffcont >>
rect -1966 8244 -936 8278
rect -2062 7796 -2028 8182
rect -874 7796 -840 8182
rect -1966 7700 -936 7734
rect 7034 8244 8064 8278
rect 6938 7796 6972 8182
rect 8126 7796 8160 8182
rect 7034 7700 8064 7734
rect -1966 6444 -936 6478
rect -2062 5996 -2028 6382
rect -874 5996 -840 6382
rect -1966 5900 -936 5934
rect 7034 6444 8064 6478
rect 6938 5996 6972 6382
rect 8126 5996 8160 6382
rect 7034 5900 8064 5934
rect -1966 4644 -936 4678
rect -2062 4196 -2028 4582
rect -874 4196 -840 4582
rect -1966 4100 -936 4134
rect 7034 4644 8064 4678
rect 6938 4196 6972 4582
rect 8126 4196 8160 4582
rect 7034 4100 8064 4134
rect -1966 2844 -936 2878
rect -2062 2396 -2028 2782
rect -874 2396 -840 2782
rect -1966 2300 -936 2334
rect 7034 2844 8064 2878
rect 6938 2396 6972 2782
rect 8126 2396 8160 2782
rect 7034 2300 8064 2334
rect -1966 1044 -936 1078
rect -2062 596 -2028 982
rect -874 596 -840 982
rect -1966 500 -936 534
rect 7034 1044 8064 1078
rect 6938 596 6972 982
rect 8126 596 8160 982
rect 7034 500 8064 534
rect -1966 -756 -936 -722
rect -2062 -1204 -2028 -818
rect -874 -1204 -840 -818
rect -1966 -1300 -936 -1266
rect 7034 -756 8064 -722
rect 6938 -1204 6972 -818
rect 8126 -1204 8160 -818
rect 7034 -1300 8064 -1266
<< poly >>
rect -1964 8176 -938 8192
rect -1964 8142 -1948 8176
rect -1914 8142 -1756 8176
rect -1722 8142 -1564 8176
rect -1530 8142 -1372 8176
rect -1338 8142 -1180 8176
rect -1146 8142 -988 8176
rect -954 8142 -938 8176
rect -1964 8126 -938 8142
rect -1898 8094 -1868 8126
rect -1802 8094 -1772 8126
rect -1706 8094 -1676 8126
rect -1610 8094 -1580 8126
rect -1514 8094 -1484 8126
rect -1418 8094 -1388 8126
rect -1322 8094 -1292 8126
rect -1226 8094 -1196 8126
rect -1130 8094 -1100 8126
rect -1034 8094 -1004 8126
rect -1898 7796 -1868 7822
rect -1802 7796 -1772 7822
rect -1706 7796 -1676 7822
rect -1610 7796 -1580 7822
rect -1514 7796 -1484 7822
rect -1418 7796 -1388 7822
rect -1322 7796 -1292 7822
rect -1226 7796 -1196 7822
rect -1130 7796 -1100 7822
rect -1034 7796 -1004 7822
rect 7036 8176 8062 8192
rect 7036 8142 7052 8176
rect 7086 8142 7244 8176
rect 7278 8142 7436 8176
rect 7470 8142 7628 8176
rect 7662 8142 7820 8176
rect 7854 8142 8012 8176
rect 8046 8142 8062 8176
rect 7036 8126 8062 8142
rect 7102 8094 7132 8126
rect 7198 8094 7228 8126
rect 7294 8094 7324 8126
rect 7390 8094 7420 8126
rect 7486 8094 7516 8126
rect 7582 8094 7612 8126
rect 7678 8094 7708 8126
rect 7774 8094 7804 8126
rect 7870 8094 7900 8126
rect 7966 8094 7996 8126
rect 7102 7796 7132 7822
rect 7198 7796 7228 7822
rect 7294 7796 7324 7822
rect 7390 7796 7420 7822
rect 7486 7796 7516 7822
rect 7582 7796 7612 7822
rect 7678 7796 7708 7822
rect 7774 7796 7804 7822
rect 7870 7796 7900 7822
rect 7966 7796 7996 7822
rect -1898 7514 -1868 7540
rect -1802 7514 -1772 7540
rect -1706 7514 -1676 7540
rect -1610 7514 -1580 7540
rect -1514 7514 -1484 7540
rect -1418 7514 -1388 7540
rect -1322 7514 -1292 7540
rect -1226 7514 -1196 7540
rect -1130 7514 -1100 7540
rect -1034 7514 -1004 7540
rect -1898 7388 -1868 7410
rect -1802 7388 -1772 7410
rect -1706 7388 -1676 7410
rect -1610 7388 -1580 7410
rect -1514 7388 -1484 7410
rect -1418 7388 -1388 7410
rect -1322 7388 -1292 7410
rect -1226 7388 -1196 7410
rect -1130 7388 -1100 7410
rect -1034 7388 -1004 7410
rect -1964 7368 -938 7388
rect -1964 7334 -1948 7368
rect -1914 7334 -1756 7368
rect -1722 7334 -1564 7368
rect -1530 7334 -1372 7368
rect -1338 7334 -1180 7368
rect -1146 7334 -988 7368
rect -954 7334 -938 7368
rect -1964 7322 -938 7334
rect 7102 7514 7132 7540
rect 7198 7514 7228 7540
rect 7294 7514 7324 7540
rect 7390 7514 7420 7540
rect 7486 7514 7516 7540
rect 7582 7514 7612 7540
rect 7678 7514 7708 7540
rect 7774 7514 7804 7540
rect 7870 7514 7900 7540
rect 7966 7514 7996 7540
rect 7102 7388 7132 7410
rect 7198 7388 7228 7410
rect 7294 7388 7324 7410
rect 7390 7388 7420 7410
rect 7486 7388 7516 7410
rect 7582 7388 7612 7410
rect 7678 7388 7708 7410
rect 7774 7388 7804 7410
rect 7870 7388 7900 7410
rect 7966 7388 7996 7410
rect 7036 7368 8062 7388
rect 7036 7334 7052 7368
rect 7086 7334 7244 7368
rect 7278 7334 7436 7368
rect 7470 7334 7628 7368
rect 7662 7334 7820 7368
rect 7854 7334 8012 7368
rect 8046 7334 8062 7368
rect 7036 7322 8062 7334
rect -1964 6376 -938 6392
rect -1964 6342 -1948 6376
rect -1914 6342 -1756 6376
rect -1722 6342 -1564 6376
rect -1530 6342 -1372 6376
rect -1338 6342 -1180 6376
rect -1146 6342 -988 6376
rect -954 6342 -938 6376
rect -1964 6326 -938 6342
rect -1898 6294 -1868 6326
rect -1802 6294 -1772 6326
rect -1706 6294 -1676 6326
rect -1610 6294 -1580 6326
rect -1514 6294 -1484 6326
rect -1418 6294 -1388 6326
rect -1322 6294 -1292 6326
rect -1226 6294 -1196 6326
rect -1130 6294 -1100 6326
rect -1034 6294 -1004 6326
rect -1898 5996 -1868 6022
rect -1802 5996 -1772 6022
rect -1706 5996 -1676 6022
rect -1610 5996 -1580 6022
rect -1514 5996 -1484 6022
rect -1418 5996 -1388 6022
rect -1322 5996 -1292 6022
rect -1226 5996 -1196 6022
rect -1130 5996 -1100 6022
rect -1034 5996 -1004 6022
rect 7036 6376 8062 6392
rect 7036 6342 7052 6376
rect 7086 6342 7244 6376
rect 7278 6342 7436 6376
rect 7470 6342 7628 6376
rect 7662 6342 7820 6376
rect 7854 6342 8012 6376
rect 8046 6342 8062 6376
rect 7036 6326 8062 6342
rect 7102 6294 7132 6326
rect 7198 6294 7228 6326
rect 7294 6294 7324 6326
rect 7390 6294 7420 6326
rect 7486 6294 7516 6326
rect 7582 6294 7612 6326
rect 7678 6294 7708 6326
rect 7774 6294 7804 6326
rect 7870 6294 7900 6326
rect 7966 6294 7996 6326
rect 7102 5996 7132 6022
rect 7198 5996 7228 6022
rect 7294 5996 7324 6022
rect 7390 5996 7420 6022
rect 7486 5996 7516 6022
rect 7582 5996 7612 6022
rect 7678 5996 7708 6022
rect 7774 5996 7804 6022
rect 7870 5996 7900 6022
rect 7966 5996 7996 6022
rect -1898 5714 -1868 5740
rect -1802 5714 -1772 5740
rect -1706 5714 -1676 5740
rect -1610 5714 -1580 5740
rect -1514 5714 -1484 5740
rect -1418 5714 -1388 5740
rect -1322 5714 -1292 5740
rect -1226 5714 -1196 5740
rect -1130 5714 -1100 5740
rect -1034 5714 -1004 5740
rect -1898 5588 -1868 5610
rect -1802 5588 -1772 5610
rect -1706 5588 -1676 5610
rect -1610 5588 -1580 5610
rect -1514 5588 -1484 5610
rect -1418 5588 -1388 5610
rect -1322 5588 -1292 5610
rect -1226 5588 -1196 5610
rect -1130 5588 -1100 5610
rect -1034 5588 -1004 5610
rect -1964 5568 -938 5588
rect -1964 5534 -1948 5568
rect -1914 5534 -1756 5568
rect -1722 5534 -1564 5568
rect -1530 5534 -1372 5568
rect -1338 5534 -1180 5568
rect -1146 5534 -988 5568
rect -954 5534 -938 5568
rect -1964 5522 -938 5534
rect 7102 5714 7132 5740
rect 7198 5714 7228 5740
rect 7294 5714 7324 5740
rect 7390 5714 7420 5740
rect 7486 5714 7516 5740
rect 7582 5714 7612 5740
rect 7678 5714 7708 5740
rect 7774 5714 7804 5740
rect 7870 5714 7900 5740
rect 7966 5714 7996 5740
rect 7102 5588 7132 5610
rect 7198 5588 7228 5610
rect 7294 5588 7324 5610
rect 7390 5588 7420 5610
rect 7486 5588 7516 5610
rect 7582 5588 7612 5610
rect 7678 5588 7708 5610
rect 7774 5588 7804 5610
rect 7870 5588 7900 5610
rect 7966 5588 7996 5610
rect 7036 5568 8062 5588
rect 7036 5534 7052 5568
rect 7086 5534 7244 5568
rect 7278 5534 7436 5568
rect 7470 5534 7628 5568
rect 7662 5534 7820 5568
rect 7854 5534 8012 5568
rect 8046 5534 8062 5568
rect 7036 5522 8062 5534
rect -1964 4576 -938 4592
rect -1964 4542 -1948 4576
rect -1914 4542 -1756 4576
rect -1722 4542 -1564 4576
rect -1530 4542 -1372 4576
rect -1338 4542 -1180 4576
rect -1146 4542 -988 4576
rect -954 4542 -938 4576
rect -1964 4526 -938 4542
rect -1898 4494 -1868 4526
rect -1802 4494 -1772 4526
rect -1706 4494 -1676 4526
rect -1610 4494 -1580 4526
rect -1514 4494 -1484 4526
rect -1418 4494 -1388 4526
rect -1322 4494 -1292 4526
rect -1226 4494 -1196 4526
rect -1130 4494 -1100 4526
rect -1034 4494 -1004 4526
rect -1898 4196 -1868 4222
rect -1802 4196 -1772 4222
rect -1706 4196 -1676 4222
rect -1610 4196 -1580 4222
rect -1514 4196 -1484 4222
rect -1418 4196 -1388 4222
rect -1322 4196 -1292 4222
rect -1226 4196 -1196 4222
rect -1130 4196 -1100 4222
rect -1034 4196 -1004 4222
rect 7036 4576 8062 4592
rect 7036 4542 7052 4576
rect 7086 4542 7244 4576
rect 7278 4542 7436 4576
rect 7470 4542 7628 4576
rect 7662 4542 7820 4576
rect 7854 4542 8012 4576
rect 8046 4542 8062 4576
rect 7036 4526 8062 4542
rect 7102 4494 7132 4526
rect 7198 4494 7228 4526
rect 7294 4494 7324 4526
rect 7390 4494 7420 4526
rect 7486 4494 7516 4526
rect 7582 4494 7612 4526
rect 7678 4494 7708 4526
rect 7774 4494 7804 4526
rect 7870 4494 7900 4526
rect 7966 4494 7996 4526
rect 7102 4196 7132 4222
rect 7198 4196 7228 4222
rect 7294 4196 7324 4222
rect 7390 4196 7420 4222
rect 7486 4196 7516 4222
rect 7582 4196 7612 4222
rect 7678 4196 7708 4222
rect 7774 4196 7804 4222
rect 7870 4196 7900 4222
rect 7966 4196 7996 4222
rect -1898 3914 -1868 3940
rect -1802 3914 -1772 3940
rect -1706 3914 -1676 3940
rect -1610 3914 -1580 3940
rect -1514 3914 -1484 3940
rect -1418 3914 -1388 3940
rect -1322 3914 -1292 3940
rect -1226 3914 -1196 3940
rect -1130 3914 -1100 3940
rect -1034 3914 -1004 3940
rect -1898 3788 -1868 3810
rect -1802 3788 -1772 3810
rect -1706 3788 -1676 3810
rect -1610 3788 -1580 3810
rect -1514 3788 -1484 3810
rect -1418 3788 -1388 3810
rect -1322 3788 -1292 3810
rect -1226 3788 -1196 3810
rect -1130 3788 -1100 3810
rect -1034 3788 -1004 3810
rect -1964 3768 -938 3788
rect -1964 3734 -1948 3768
rect -1914 3734 -1756 3768
rect -1722 3734 -1564 3768
rect -1530 3734 -1372 3768
rect -1338 3734 -1180 3768
rect -1146 3734 -988 3768
rect -954 3734 -938 3768
rect -1964 3722 -938 3734
rect 7102 3914 7132 3940
rect 7198 3914 7228 3940
rect 7294 3914 7324 3940
rect 7390 3914 7420 3940
rect 7486 3914 7516 3940
rect 7582 3914 7612 3940
rect 7678 3914 7708 3940
rect 7774 3914 7804 3940
rect 7870 3914 7900 3940
rect 7966 3914 7996 3940
rect 7102 3788 7132 3810
rect 7198 3788 7228 3810
rect 7294 3788 7324 3810
rect 7390 3788 7420 3810
rect 7486 3788 7516 3810
rect 7582 3788 7612 3810
rect 7678 3788 7708 3810
rect 7774 3788 7804 3810
rect 7870 3788 7900 3810
rect 7966 3788 7996 3810
rect 7036 3768 8062 3788
rect 7036 3734 7052 3768
rect 7086 3734 7244 3768
rect 7278 3734 7436 3768
rect 7470 3734 7628 3768
rect 7662 3734 7820 3768
rect 7854 3734 8012 3768
rect 8046 3734 8062 3768
rect 7036 3722 8062 3734
rect -1964 2776 -938 2792
rect -1964 2742 -1948 2776
rect -1914 2742 -1756 2776
rect -1722 2742 -1564 2776
rect -1530 2742 -1372 2776
rect -1338 2742 -1180 2776
rect -1146 2742 -988 2776
rect -954 2742 -938 2776
rect -1964 2726 -938 2742
rect -1898 2694 -1868 2726
rect -1802 2694 -1772 2726
rect -1706 2694 -1676 2726
rect -1610 2694 -1580 2726
rect -1514 2694 -1484 2726
rect -1418 2694 -1388 2726
rect -1322 2694 -1292 2726
rect -1226 2694 -1196 2726
rect -1130 2694 -1100 2726
rect -1034 2694 -1004 2726
rect -1898 2396 -1868 2422
rect -1802 2396 -1772 2422
rect -1706 2396 -1676 2422
rect -1610 2396 -1580 2422
rect -1514 2396 -1484 2422
rect -1418 2396 -1388 2422
rect -1322 2396 -1292 2422
rect -1226 2396 -1196 2422
rect -1130 2396 -1100 2422
rect -1034 2396 -1004 2422
rect 7036 2776 8062 2792
rect 7036 2742 7052 2776
rect 7086 2742 7244 2776
rect 7278 2742 7436 2776
rect 7470 2742 7628 2776
rect 7662 2742 7820 2776
rect 7854 2742 8012 2776
rect 8046 2742 8062 2776
rect 7036 2726 8062 2742
rect 7102 2694 7132 2726
rect 7198 2694 7228 2726
rect 7294 2694 7324 2726
rect 7390 2694 7420 2726
rect 7486 2694 7516 2726
rect 7582 2694 7612 2726
rect 7678 2694 7708 2726
rect 7774 2694 7804 2726
rect 7870 2694 7900 2726
rect 7966 2694 7996 2726
rect 7102 2396 7132 2422
rect 7198 2396 7228 2422
rect 7294 2396 7324 2422
rect 7390 2396 7420 2422
rect 7486 2396 7516 2422
rect 7582 2396 7612 2422
rect 7678 2396 7708 2422
rect 7774 2396 7804 2422
rect 7870 2396 7900 2422
rect 7966 2396 7996 2422
rect -1898 2114 -1868 2140
rect -1802 2114 -1772 2140
rect -1706 2114 -1676 2140
rect -1610 2114 -1580 2140
rect -1514 2114 -1484 2140
rect -1418 2114 -1388 2140
rect -1322 2114 -1292 2140
rect -1226 2114 -1196 2140
rect -1130 2114 -1100 2140
rect -1034 2114 -1004 2140
rect -1898 1988 -1868 2010
rect -1802 1988 -1772 2010
rect -1706 1988 -1676 2010
rect -1610 1988 -1580 2010
rect -1514 1988 -1484 2010
rect -1418 1988 -1388 2010
rect -1322 1988 -1292 2010
rect -1226 1988 -1196 2010
rect -1130 1988 -1100 2010
rect -1034 1988 -1004 2010
rect -1964 1968 -938 1988
rect -1964 1934 -1948 1968
rect -1914 1934 -1756 1968
rect -1722 1934 -1564 1968
rect -1530 1934 -1372 1968
rect -1338 1934 -1180 1968
rect -1146 1934 -988 1968
rect -954 1934 -938 1968
rect -1964 1922 -938 1934
rect 7102 2114 7132 2140
rect 7198 2114 7228 2140
rect 7294 2114 7324 2140
rect 7390 2114 7420 2140
rect 7486 2114 7516 2140
rect 7582 2114 7612 2140
rect 7678 2114 7708 2140
rect 7774 2114 7804 2140
rect 7870 2114 7900 2140
rect 7966 2114 7996 2140
rect 7102 1988 7132 2010
rect 7198 1988 7228 2010
rect 7294 1988 7324 2010
rect 7390 1988 7420 2010
rect 7486 1988 7516 2010
rect 7582 1988 7612 2010
rect 7678 1988 7708 2010
rect 7774 1988 7804 2010
rect 7870 1988 7900 2010
rect 7966 1988 7996 2010
rect 7036 1968 8062 1988
rect 7036 1934 7052 1968
rect 7086 1934 7244 1968
rect 7278 1934 7436 1968
rect 7470 1934 7628 1968
rect 7662 1934 7820 1968
rect 7854 1934 8012 1968
rect 8046 1934 8062 1968
rect 7036 1922 8062 1934
rect -1964 976 -938 992
rect -1964 942 -1948 976
rect -1914 942 -1756 976
rect -1722 942 -1564 976
rect -1530 942 -1372 976
rect -1338 942 -1180 976
rect -1146 942 -988 976
rect -954 942 -938 976
rect -1964 926 -938 942
rect -1898 894 -1868 926
rect -1802 894 -1772 926
rect -1706 894 -1676 926
rect -1610 894 -1580 926
rect -1514 894 -1484 926
rect -1418 894 -1388 926
rect -1322 894 -1292 926
rect -1226 894 -1196 926
rect -1130 894 -1100 926
rect -1034 894 -1004 926
rect -1898 596 -1868 622
rect -1802 596 -1772 622
rect -1706 596 -1676 622
rect -1610 596 -1580 622
rect -1514 596 -1484 622
rect -1418 596 -1388 622
rect -1322 596 -1292 622
rect -1226 596 -1196 622
rect -1130 596 -1100 622
rect -1034 596 -1004 622
rect 7036 976 8062 992
rect 7036 942 7052 976
rect 7086 942 7244 976
rect 7278 942 7436 976
rect 7470 942 7628 976
rect 7662 942 7820 976
rect 7854 942 8012 976
rect 8046 942 8062 976
rect 7036 926 8062 942
rect 7102 894 7132 926
rect 7198 894 7228 926
rect 7294 894 7324 926
rect 7390 894 7420 926
rect 7486 894 7516 926
rect 7582 894 7612 926
rect 7678 894 7708 926
rect 7774 894 7804 926
rect 7870 894 7900 926
rect 7966 894 7996 926
rect 7102 596 7132 622
rect 7198 596 7228 622
rect 7294 596 7324 622
rect 7390 596 7420 622
rect 7486 596 7516 622
rect 7582 596 7612 622
rect 7678 596 7708 622
rect 7774 596 7804 622
rect 7870 596 7900 622
rect 7966 596 7996 622
rect -1898 314 -1868 340
rect -1802 314 -1772 340
rect -1706 314 -1676 340
rect -1610 314 -1580 340
rect -1514 314 -1484 340
rect -1418 314 -1388 340
rect -1322 314 -1292 340
rect -1226 314 -1196 340
rect -1130 314 -1100 340
rect -1034 314 -1004 340
rect -1898 188 -1868 210
rect -1802 188 -1772 210
rect -1706 188 -1676 210
rect -1610 188 -1580 210
rect -1514 188 -1484 210
rect -1418 188 -1388 210
rect -1322 188 -1292 210
rect -1226 188 -1196 210
rect -1130 188 -1100 210
rect -1034 188 -1004 210
rect -1964 168 -938 188
rect -1964 134 -1948 168
rect -1914 134 -1756 168
rect -1722 134 -1564 168
rect -1530 134 -1372 168
rect -1338 134 -1180 168
rect -1146 134 -988 168
rect -954 134 -938 168
rect -1964 122 -938 134
rect 7102 314 7132 340
rect 7198 314 7228 340
rect 7294 314 7324 340
rect 7390 314 7420 340
rect 7486 314 7516 340
rect 7582 314 7612 340
rect 7678 314 7708 340
rect 7774 314 7804 340
rect 7870 314 7900 340
rect 7966 314 7996 340
rect 7102 188 7132 210
rect 7198 188 7228 210
rect 7294 188 7324 210
rect 7390 188 7420 210
rect 7486 188 7516 210
rect 7582 188 7612 210
rect 7678 188 7708 210
rect 7774 188 7804 210
rect 7870 188 7900 210
rect 7966 188 7996 210
rect 7036 168 8062 188
rect 7036 134 7052 168
rect 7086 134 7244 168
rect 7278 134 7436 168
rect 7470 134 7628 168
rect 7662 134 7820 168
rect 7854 134 8012 168
rect 8046 134 8062 168
rect 7036 122 8062 134
rect -1964 -824 -938 -808
rect -1964 -858 -1948 -824
rect -1914 -858 -1756 -824
rect -1722 -858 -1564 -824
rect -1530 -858 -1372 -824
rect -1338 -858 -1180 -824
rect -1146 -858 -988 -824
rect -954 -858 -938 -824
rect -1964 -874 -938 -858
rect -1898 -906 -1868 -874
rect -1802 -906 -1772 -874
rect -1706 -906 -1676 -874
rect -1610 -906 -1580 -874
rect -1514 -906 -1484 -874
rect -1418 -906 -1388 -874
rect -1322 -906 -1292 -874
rect -1226 -906 -1196 -874
rect -1130 -906 -1100 -874
rect -1034 -906 -1004 -874
rect -1898 -1204 -1868 -1178
rect -1802 -1204 -1772 -1178
rect -1706 -1204 -1676 -1178
rect -1610 -1204 -1580 -1178
rect -1514 -1204 -1484 -1178
rect -1418 -1204 -1388 -1178
rect -1322 -1204 -1292 -1178
rect -1226 -1204 -1196 -1178
rect -1130 -1204 -1100 -1178
rect -1034 -1204 -1004 -1178
rect 7036 -824 8062 -808
rect 7036 -858 7052 -824
rect 7086 -858 7244 -824
rect 7278 -858 7436 -824
rect 7470 -858 7628 -824
rect 7662 -858 7820 -824
rect 7854 -858 8012 -824
rect 8046 -858 8062 -824
rect 7036 -874 8062 -858
rect 7102 -906 7132 -874
rect 7198 -906 7228 -874
rect 7294 -906 7324 -874
rect 7390 -906 7420 -874
rect 7486 -906 7516 -874
rect 7582 -906 7612 -874
rect 7678 -906 7708 -874
rect 7774 -906 7804 -874
rect 7870 -906 7900 -874
rect 7966 -906 7996 -874
rect 7102 -1204 7132 -1178
rect 7198 -1204 7228 -1178
rect 7294 -1204 7324 -1178
rect 7390 -1204 7420 -1178
rect 7486 -1204 7516 -1178
rect 7582 -1204 7612 -1178
rect 7678 -1204 7708 -1178
rect 7774 -1204 7804 -1178
rect 7870 -1204 7900 -1178
rect 7966 -1204 7996 -1178
rect -1898 -1486 -1868 -1460
rect -1802 -1486 -1772 -1460
rect -1706 -1486 -1676 -1460
rect -1610 -1486 -1580 -1460
rect -1514 -1486 -1484 -1460
rect -1418 -1486 -1388 -1460
rect -1322 -1486 -1292 -1460
rect -1226 -1486 -1196 -1460
rect -1130 -1486 -1100 -1460
rect -1034 -1486 -1004 -1460
rect -1898 -1612 -1868 -1590
rect -1802 -1612 -1772 -1590
rect -1706 -1612 -1676 -1590
rect -1610 -1612 -1580 -1590
rect -1514 -1612 -1484 -1590
rect -1418 -1612 -1388 -1590
rect -1322 -1612 -1292 -1590
rect -1226 -1612 -1196 -1590
rect -1130 -1612 -1100 -1590
rect -1034 -1612 -1004 -1590
rect -1964 -1632 -938 -1612
rect -1964 -1666 -1948 -1632
rect -1914 -1666 -1756 -1632
rect -1722 -1666 -1564 -1632
rect -1530 -1666 -1372 -1632
rect -1338 -1666 -1180 -1632
rect -1146 -1666 -988 -1632
rect -954 -1666 -938 -1632
rect -1964 -1678 -938 -1666
rect 7102 -1486 7132 -1460
rect 7198 -1486 7228 -1460
rect 7294 -1486 7324 -1460
rect 7390 -1486 7420 -1460
rect 7486 -1486 7516 -1460
rect 7582 -1486 7612 -1460
rect 7678 -1486 7708 -1460
rect 7774 -1486 7804 -1460
rect 7870 -1486 7900 -1460
rect 7966 -1486 7996 -1460
rect 7102 -1612 7132 -1590
rect 7198 -1612 7228 -1590
rect 7294 -1612 7324 -1590
rect 7390 -1612 7420 -1590
rect 7486 -1612 7516 -1590
rect 7582 -1612 7612 -1590
rect 7678 -1612 7708 -1590
rect 7774 -1612 7804 -1590
rect 7870 -1612 7900 -1590
rect 7966 -1612 7996 -1590
rect 7036 -1632 8062 -1612
rect 7036 -1666 7052 -1632
rect 7086 -1666 7244 -1632
rect 7278 -1666 7436 -1632
rect 7470 -1666 7628 -1632
rect 7662 -1666 7820 -1632
rect 7854 -1666 8012 -1632
rect 8046 -1666 8062 -1632
rect 7036 -1678 8062 -1666
<< polycont >>
rect -1948 8142 -1914 8176
rect -1756 8142 -1722 8176
rect -1564 8142 -1530 8176
rect -1372 8142 -1338 8176
rect -1180 8142 -1146 8176
rect -988 8142 -954 8176
rect 7052 8142 7086 8176
rect 7244 8142 7278 8176
rect 7436 8142 7470 8176
rect 7628 8142 7662 8176
rect 7820 8142 7854 8176
rect 8012 8142 8046 8176
rect -1948 7334 -1914 7368
rect -1756 7334 -1722 7368
rect -1564 7334 -1530 7368
rect -1372 7334 -1338 7368
rect -1180 7334 -1146 7368
rect -988 7334 -954 7368
rect 7052 7334 7086 7368
rect 7244 7334 7278 7368
rect 7436 7334 7470 7368
rect 7628 7334 7662 7368
rect 7820 7334 7854 7368
rect 8012 7334 8046 7368
rect -1948 6342 -1914 6376
rect -1756 6342 -1722 6376
rect -1564 6342 -1530 6376
rect -1372 6342 -1338 6376
rect -1180 6342 -1146 6376
rect -988 6342 -954 6376
rect 7052 6342 7086 6376
rect 7244 6342 7278 6376
rect 7436 6342 7470 6376
rect 7628 6342 7662 6376
rect 7820 6342 7854 6376
rect 8012 6342 8046 6376
rect -1948 5534 -1914 5568
rect -1756 5534 -1722 5568
rect -1564 5534 -1530 5568
rect -1372 5534 -1338 5568
rect -1180 5534 -1146 5568
rect -988 5534 -954 5568
rect 7052 5534 7086 5568
rect 7244 5534 7278 5568
rect 7436 5534 7470 5568
rect 7628 5534 7662 5568
rect 7820 5534 7854 5568
rect 8012 5534 8046 5568
rect -1948 4542 -1914 4576
rect -1756 4542 -1722 4576
rect -1564 4542 -1530 4576
rect -1372 4542 -1338 4576
rect -1180 4542 -1146 4576
rect -988 4542 -954 4576
rect 7052 4542 7086 4576
rect 7244 4542 7278 4576
rect 7436 4542 7470 4576
rect 7628 4542 7662 4576
rect 7820 4542 7854 4576
rect 8012 4542 8046 4576
rect -1948 3734 -1914 3768
rect -1756 3734 -1722 3768
rect -1564 3734 -1530 3768
rect -1372 3734 -1338 3768
rect -1180 3734 -1146 3768
rect -988 3734 -954 3768
rect 7052 3734 7086 3768
rect 7244 3734 7278 3768
rect 7436 3734 7470 3768
rect 7628 3734 7662 3768
rect 7820 3734 7854 3768
rect 8012 3734 8046 3768
rect -1948 2742 -1914 2776
rect -1756 2742 -1722 2776
rect -1564 2742 -1530 2776
rect -1372 2742 -1338 2776
rect -1180 2742 -1146 2776
rect -988 2742 -954 2776
rect 7052 2742 7086 2776
rect 7244 2742 7278 2776
rect 7436 2742 7470 2776
rect 7628 2742 7662 2776
rect 7820 2742 7854 2776
rect 8012 2742 8046 2776
rect -1948 1934 -1914 1968
rect -1756 1934 -1722 1968
rect -1564 1934 -1530 1968
rect -1372 1934 -1338 1968
rect -1180 1934 -1146 1968
rect -988 1934 -954 1968
rect 7052 1934 7086 1968
rect 7244 1934 7278 1968
rect 7436 1934 7470 1968
rect 7628 1934 7662 1968
rect 7820 1934 7854 1968
rect 8012 1934 8046 1968
rect -1948 942 -1914 976
rect -1756 942 -1722 976
rect -1564 942 -1530 976
rect -1372 942 -1338 976
rect -1180 942 -1146 976
rect -988 942 -954 976
rect 7052 942 7086 976
rect 7244 942 7278 976
rect 7436 942 7470 976
rect 7628 942 7662 976
rect 7820 942 7854 976
rect 8012 942 8046 976
rect -1948 134 -1914 168
rect -1756 134 -1722 168
rect -1564 134 -1530 168
rect -1372 134 -1338 168
rect -1180 134 -1146 168
rect -988 134 -954 168
rect 7052 134 7086 168
rect 7244 134 7278 168
rect 7436 134 7470 168
rect 7628 134 7662 168
rect 7820 134 7854 168
rect 8012 134 8046 168
rect -1948 -858 -1914 -824
rect -1756 -858 -1722 -824
rect -1564 -858 -1530 -824
rect -1372 -858 -1338 -824
rect -1180 -858 -1146 -824
rect -988 -858 -954 -824
rect 7052 -858 7086 -824
rect 7244 -858 7278 -824
rect 7436 -858 7470 -824
rect 7628 -858 7662 -824
rect 7820 -858 7854 -824
rect 8012 -858 8046 -824
rect -1948 -1666 -1914 -1632
rect -1756 -1666 -1722 -1632
rect -1564 -1666 -1530 -1632
rect -1372 -1666 -1338 -1632
rect -1180 -1666 -1146 -1632
rect -988 -1666 -954 -1632
rect 7052 -1666 7086 -1632
rect 7244 -1666 7278 -1632
rect 7436 -1666 7470 -1632
rect 7628 -1666 7662 -1632
rect 7820 -1666 7854 -1632
rect 8012 -1666 8046 -1632
<< locali >>
rect -2062 8244 -1966 8278
rect -936 8244 -840 8278
rect -2062 8182 -2028 8244
rect -874 8182 -840 8244
rect -1964 8142 -1948 8176
rect -1914 8142 -1898 8176
rect -1772 8142 -1756 8176
rect -1722 8142 -1706 8176
rect -1580 8142 -1564 8176
rect -1530 8142 -1514 8176
rect -1388 8142 -1372 8176
rect -1338 8142 -1322 8176
rect -1196 8142 -1180 8176
rect -1146 8142 -1130 8176
rect -1004 8142 -988 8176
rect -954 8142 -938 8176
rect -1948 8082 -1914 8098
rect -1948 7818 -1914 7834
rect -1852 8082 -1818 8098
rect -1852 7818 -1818 7834
rect -1756 8082 -1722 8098
rect -1756 7818 -1722 7834
rect -1660 8082 -1626 8098
rect -1660 7818 -1626 7834
rect -1564 8082 -1530 8098
rect -1564 7818 -1530 7834
rect -1468 8082 -1434 8098
rect -1468 7818 -1434 7834
rect -1372 8082 -1338 8098
rect -1372 7818 -1338 7834
rect -1276 8082 -1242 8098
rect -1276 7818 -1242 7834
rect -1180 8082 -1146 8098
rect -1180 7818 -1146 7834
rect -1084 8082 -1050 8098
rect -1084 7818 -1050 7834
rect -988 8082 -954 8098
rect -988 7818 -954 7834
rect -2062 7734 -2028 7796
rect -874 7734 -840 7796
rect -2062 7700 -1966 7734
rect -936 7700 -840 7734
rect 6938 8244 7034 8278
rect 8064 8244 8160 8278
rect 6938 8182 6972 8244
rect 8126 8182 8160 8244
rect 7036 8142 7052 8176
rect 7086 8142 7102 8176
rect 7228 8142 7244 8176
rect 7278 8142 7294 8176
rect 7420 8142 7436 8176
rect 7470 8142 7486 8176
rect 7612 8142 7628 8176
rect 7662 8142 7678 8176
rect 7804 8142 7820 8176
rect 7854 8142 7870 8176
rect 7996 8142 8012 8176
rect 8046 8142 8062 8176
rect 7052 8082 7086 8098
rect 7052 7818 7086 7834
rect 7148 8082 7182 8098
rect 7148 7818 7182 7834
rect 7244 8082 7278 8098
rect 7244 7818 7278 7834
rect 7340 8082 7374 8098
rect 7340 7818 7374 7834
rect 7436 8082 7470 8098
rect 7436 7818 7470 7834
rect 7532 8082 7566 8098
rect 7532 7818 7566 7834
rect 7628 8082 7662 8098
rect 7628 7818 7662 7834
rect 7724 8082 7758 8098
rect 7724 7818 7758 7834
rect 7820 8082 7854 8098
rect 7820 7818 7854 7834
rect 7916 8082 7950 8098
rect 7916 7818 7950 7834
rect 8012 8082 8046 8098
rect 8012 7818 8046 7834
rect 6938 7734 6972 7796
rect 8126 7734 8160 7796
rect 6938 7700 7034 7734
rect 8064 7700 8160 7734
rect -2062 7592 -1966 7626
rect -936 7592 -840 7626
rect -2062 7532 -2028 7592
rect -874 7530 -840 7592
rect -1948 7502 -1914 7518
rect -1948 7406 -1914 7422
rect -1852 7502 -1818 7518
rect -1852 7406 -1818 7422
rect -1756 7502 -1722 7518
rect -1756 7406 -1722 7422
rect -1660 7502 -1626 7518
rect -1660 7406 -1626 7422
rect -1564 7502 -1530 7518
rect -1564 7406 -1530 7422
rect -1468 7502 -1434 7518
rect -1468 7406 -1434 7422
rect -1372 7502 -1338 7518
rect -1372 7406 -1338 7422
rect -1276 7502 -1242 7518
rect -1276 7406 -1242 7422
rect -1180 7502 -1146 7518
rect -1180 7406 -1146 7422
rect -1084 7502 -1050 7518
rect -1084 7406 -1050 7422
rect -988 7502 -954 7518
rect -988 7406 -954 7422
rect -1964 7334 -1948 7368
rect -1914 7334 -1898 7368
rect -1772 7334 -1756 7368
rect -1722 7334 -1706 7368
rect -1580 7334 -1564 7368
rect -1530 7334 -1514 7368
rect -1388 7334 -1372 7368
rect -1338 7334 -1322 7368
rect -1196 7334 -1180 7368
rect -1146 7334 -1130 7368
rect -1004 7334 -988 7368
rect -954 7334 -938 7368
rect -2062 7270 -2028 7332
rect -874 7270 -840 7332
rect -2062 7236 -1966 7270
rect -936 7236 -840 7270
rect 6938 7592 7034 7626
rect 8064 7592 8160 7626
rect 6938 7532 6972 7592
rect 8126 7530 8160 7592
rect 7052 7502 7086 7518
rect 7052 7406 7086 7422
rect 7148 7502 7182 7518
rect 7148 7406 7182 7422
rect 7244 7502 7278 7518
rect 7244 7406 7278 7422
rect 7340 7502 7374 7518
rect 7340 7406 7374 7422
rect 7436 7502 7470 7518
rect 7436 7406 7470 7422
rect 7532 7502 7566 7518
rect 7532 7406 7566 7422
rect 7628 7502 7662 7518
rect 7628 7406 7662 7422
rect 7724 7502 7758 7518
rect 7724 7406 7758 7422
rect 7820 7502 7854 7518
rect 7820 7406 7854 7422
rect 7916 7502 7950 7518
rect 7916 7406 7950 7422
rect 8012 7502 8046 7518
rect 8012 7406 8046 7422
rect 7036 7334 7052 7368
rect 7086 7334 7102 7368
rect 7228 7334 7244 7368
rect 7278 7334 7294 7368
rect 7420 7334 7436 7368
rect 7470 7334 7486 7368
rect 7612 7334 7628 7368
rect 7662 7334 7678 7368
rect 7804 7334 7820 7368
rect 7854 7334 7870 7368
rect 7996 7334 8012 7368
rect 8046 7334 8062 7368
rect 6938 7270 6972 7332
rect 8126 7270 8160 7332
rect 6938 7236 7034 7270
rect 8064 7236 8160 7270
rect -2062 6444 -1966 6478
rect -936 6444 -840 6478
rect -2062 6382 -2028 6444
rect -874 6382 -840 6444
rect -1964 6342 -1948 6376
rect -1914 6342 -1898 6376
rect -1772 6342 -1756 6376
rect -1722 6342 -1706 6376
rect -1580 6342 -1564 6376
rect -1530 6342 -1514 6376
rect -1388 6342 -1372 6376
rect -1338 6342 -1322 6376
rect -1196 6342 -1180 6376
rect -1146 6342 -1130 6376
rect -1004 6342 -988 6376
rect -954 6342 -938 6376
rect -1948 6282 -1914 6298
rect -1948 6018 -1914 6034
rect -1852 6282 -1818 6298
rect -1852 6018 -1818 6034
rect -1756 6282 -1722 6298
rect -1756 6018 -1722 6034
rect -1660 6282 -1626 6298
rect -1660 6018 -1626 6034
rect -1564 6282 -1530 6298
rect -1564 6018 -1530 6034
rect -1468 6282 -1434 6298
rect -1468 6018 -1434 6034
rect -1372 6282 -1338 6298
rect -1372 6018 -1338 6034
rect -1276 6282 -1242 6298
rect -1276 6018 -1242 6034
rect -1180 6282 -1146 6298
rect -1180 6018 -1146 6034
rect -1084 6282 -1050 6298
rect -1084 6018 -1050 6034
rect -988 6282 -954 6298
rect -988 6018 -954 6034
rect -2062 5934 -2028 5996
rect -874 5934 -840 5996
rect -2062 5900 -1966 5934
rect -936 5900 -840 5934
rect 6938 6444 7034 6478
rect 8064 6444 8160 6478
rect 6938 6382 6972 6444
rect 8126 6382 8160 6444
rect 7036 6342 7052 6376
rect 7086 6342 7102 6376
rect 7228 6342 7244 6376
rect 7278 6342 7294 6376
rect 7420 6342 7436 6376
rect 7470 6342 7486 6376
rect 7612 6342 7628 6376
rect 7662 6342 7678 6376
rect 7804 6342 7820 6376
rect 7854 6342 7870 6376
rect 7996 6342 8012 6376
rect 8046 6342 8062 6376
rect 7052 6282 7086 6298
rect 7052 6018 7086 6034
rect 7148 6282 7182 6298
rect 7148 6018 7182 6034
rect 7244 6282 7278 6298
rect 7244 6018 7278 6034
rect 7340 6282 7374 6298
rect 7340 6018 7374 6034
rect 7436 6282 7470 6298
rect 7436 6018 7470 6034
rect 7532 6282 7566 6298
rect 7532 6018 7566 6034
rect 7628 6282 7662 6298
rect 7628 6018 7662 6034
rect 7724 6282 7758 6298
rect 7724 6018 7758 6034
rect 7820 6282 7854 6298
rect 7820 6018 7854 6034
rect 7916 6282 7950 6298
rect 7916 6018 7950 6034
rect 8012 6282 8046 6298
rect 8012 6018 8046 6034
rect 6938 5934 6972 5996
rect 8126 5934 8160 5996
rect 6938 5900 7034 5934
rect 8064 5900 8160 5934
rect -2062 5792 -1966 5826
rect -936 5792 -840 5826
rect -2062 5732 -2028 5792
rect -874 5730 -840 5792
rect -1948 5702 -1914 5718
rect -1948 5606 -1914 5622
rect -1852 5702 -1818 5718
rect -1852 5606 -1818 5622
rect -1756 5702 -1722 5718
rect -1756 5606 -1722 5622
rect -1660 5702 -1626 5718
rect -1660 5606 -1626 5622
rect -1564 5702 -1530 5718
rect -1564 5606 -1530 5622
rect -1468 5702 -1434 5718
rect -1468 5606 -1434 5622
rect -1372 5702 -1338 5718
rect -1372 5606 -1338 5622
rect -1276 5702 -1242 5718
rect -1276 5606 -1242 5622
rect -1180 5702 -1146 5718
rect -1180 5606 -1146 5622
rect -1084 5702 -1050 5718
rect -1084 5606 -1050 5622
rect -988 5702 -954 5718
rect -988 5606 -954 5622
rect -1964 5534 -1948 5568
rect -1914 5534 -1898 5568
rect -1772 5534 -1756 5568
rect -1722 5534 -1706 5568
rect -1580 5534 -1564 5568
rect -1530 5534 -1514 5568
rect -1388 5534 -1372 5568
rect -1338 5534 -1322 5568
rect -1196 5534 -1180 5568
rect -1146 5534 -1130 5568
rect -1004 5534 -988 5568
rect -954 5534 -938 5568
rect -2062 5470 -2028 5532
rect -874 5470 -840 5532
rect -2062 5436 -1966 5470
rect -936 5436 -840 5470
rect 6938 5792 7034 5826
rect 8064 5792 8160 5826
rect 6938 5732 6972 5792
rect 8126 5730 8160 5792
rect 7052 5702 7086 5718
rect 7052 5606 7086 5622
rect 7148 5702 7182 5718
rect 7148 5606 7182 5622
rect 7244 5702 7278 5718
rect 7244 5606 7278 5622
rect 7340 5702 7374 5718
rect 7340 5606 7374 5622
rect 7436 5702 7470 5718
rect 7436 5606 7470 5622
rect 7532 5702 7566 5718
rect 7532 5606 7566 5622
rect 7628 5702 7662 5718
rect 7628 5606 7662 5622
rect 7724 5702 7758 5718
rect 7724 5606 7758 5622
rect 7820 5702 7854 5718
rect 7820 5606 7854 5622
rect 7916 5702 7950 5718
rect 7916 5606 7950 5622
rect 8012 5702 8046 5718
rect 8012 5606 8046 5622
rect 7036 5534 7052 5568
rect 7086 5534 7102 5568
rect 7228 5534 7244 5568
rect 7278 5534 7294 5568
rect 7420 5534 7436 5568
rect 7470 5534 7486 5568
rect 7612 5534 7628 5568
rect 7662 5534 7678 5568
rect 7804 5534 7820 5568
rect 7854 5534 7870 5568
rect 7996 5534 8012 5568
rect 8046 5534 8062 5568
rect 6938 5470 6972 5532
rect 8126 5470 8160 5532
rect 6938 5436 7034 5470
rect 8064 5436 8160 5470
rect -2062 4644 -1966 4678
rect -936 4644 -840 4678
rect -2062 4582 -2028 4644
rect -874 4582 -840 4644
rect -1964 4542 -1948 4576
rect -1914 4542 -1898 4576
rect -1772 4542 -1756 4576
rect -1722 4542 -1706 4576
rect -1580 4542 -1564 4576
rect -1530 4542 -1514 4576
rect -1388 4542 -1372 4576
rect -1338 4542 -1322 4576
rect -1196 4542 -1180 4576
rect -1146 4542 -1130 4576
rect -1004 4542 -988 4576
rect -954 4542 -938 4576
rect -1948 4482 -1914 4498
rect -1948 4218 -1914 4234
rect -1852 4482 -1818 4498
rect -1852 4218 -1818 4234
rect -1756 4482 -1722 4498
rect -1756 4218 -1722 4234
rect -1660 4482 -1626 4498
rect -1660 4218 -1626 4234
rect -1564 4482 -1530 4498
rect -1564 4218 -1530 4234
rect -1468 4482 -1434 4498
rect -1468 4218 -1434 4234
rect -1372 4482 -1338 4498
rect -1372 4218 -1338 4234
rect -1276 4482 -1242 4498
rect -1276 4218 -1242 4234
rect -1180 4482 -1146 4498
rect -1180 4218 -1146 4234
rect -1084 4482 -1050 4498
rect -1084 4218 -1050 4234
rect -988 4482 -954 4498
rect -988 4218 -954 4234
rect -2062 4134 -2028 4196
rect -874 4134 -840 4196
rect -2062 4100 -1966 4134
rect -936 4100 -840 4134
rect 6938 4644 7034 4678
rect 8064 4644 8160 4678
rect 6938 4582 6972 4644
rect 8126 4582 8160 4644
rect 7036 4542 7052 4576
rect 7086 4542 7102 4576
rect 7228 4542 7244 4576
rect 7278 4542 7294 4576
rect 7420 4542 7436 4576
rect 7470 4542 7486 4576
rect 7612 4542 7628 4576
rect 7662 4542 7678 4576
rect 7804 4542 7820 4576
rect 7854 4542 7870 4576
rect 7996 4542 8012 4576
rect 8046 4542 8062 4576
rect 7052 4482 7086 4498
rect 7052 4218 7086 4234
rect 7148 4482 7182 4498
rect 7148 4218 7182 4234
rect 7244 4482 7278 4498
rect 7244 4218 7278 4234
rect 7340 4482 7374 4498
rect 7340 4218 7374 4234
rect 7436 4482 7470 4498
rect 7436 4218 7470 4234
rect 7532 4482 7566 4498
rect 7532 4218 7566 4234
rect 7628 4482 7662 4498
rect 7628 4218 7662 4234
rect 7724 4482 7758 4498
rect 7724 4218 7758 4234
rect 7820 4482 7854 4498
rect 7820 4218 7854 4234
rect 7916 4482 7950 4498
rect 7916 4218 7950 4234
rect 8012 4482 8046 4498
rect 8012 4218 8046 4234
rect 6938 4134 6972 4196
rect 8126 4134 8160 4196
rect 6938 4100 7034 4134
rect 8064 4100 8160 4134
rect -2062 3992 -1966 4026
rect -936 3992 -840 4026
rect -2062 3932 -2028 3992
rect -874 3930 -840 3992
rect -1948 3902 -1914 3918
rect -1948 3806 -1914 3822
rect -1852 3902 -1818 3918
rect -1852 3806 -1818 3822
rect -1756 3902 -1722 3918
rect -1756 3806 -1722 3822
rect -1660 3902 -1626 3918
rect -1660 3806 -1626 3822
rect -1564 3902 -1530 3918
rect -1564 3806 -1530 3822
rect -1468 3902 -1434 3918
rect -1468 3806 -1434 3822
rect -1372 3902 -1338 3918
rect -1372 3806 -1338 3822
rect -1276 3902 -1242 3918
rect -1276 3806 -1242 3822
rect -1180 3902 -1146 3918
rect -1180 3806 -1146 3822
rect -1084 3902 -1050 3918
rect -1084 3806 -1050 3822
rect -988 3902 -954 3918
rect -988 3806 -954 3822
rect -1964 3734 -1948 3768
rect -1914 3734 -1898 3768
rect -1772 3734 -1756 3768
rect -1722 3734 -1706 3768
rect -1580 3734 -1564 3768
rect -1530 3734 -1514 3768
rect -1388 3734 -1372 3768
rect -1338 3734 -1322 3768
rect -1196 3734 -1180 3768
rect -1146 3734 -1130 3768
rect -1004 3734 -988 3768
rect -954 3734 -938 3768
rect -2062 3670 -2028 3732
rect -874 3670 -840 3732
rect -2062 3636 -1966 3670
rect -936 3636 -840 3670
rect 6938 3992 7034 4026
rect 8064 3992 8160 4026
rect 6938 3932 6972 3992
rect 8126 3930 8160 3992
rect 7052 3902 7086 3918
rect 7052 3806 7086 3822
rect 7148 3902 7182 3918
rect 7148 3806 7182 3822
rect 7244 3902 7278 3918
rect 7244 3806 7278 3822
rect 7340 3902 7374 3918
rect 7340 3806 7374 3822
rect 7436 3902 7470 3918
rect 7436 3806 7470 3822
rect 7532 3902 7566 3918
rect 7532 3806 7566 3822
rect 7628 3902 7662 3918
rect 7628 3806 7662 3822
rect 7724 3902 7758 3918
rect 7724 3806 7758 3822
rect 7820 3902 7854 3918
rect 7820 3806 7854 3822
rect 7916 3902 7950 3918
rect 7916 3806 7950 3822
rect 8012 3902 8046 3918
rect 8012 3806 8046 3822
rect 7036 3734 7052 3768
rect 7086 3734 7102 3768
rect 7228 3734 7244 3768
rect 7278 3734 7294 3768
rect 7420 3734 7436 3768
rect 7470 3734 7486 3768
rect 7612 3734 7628 3768
rect 7662 3734 7678 3768
rect 7804 3734 7820 3768
rect 7854 3734 7870 3768
rect 7996 3734 8012 3768
rect 8046 3734 8062 3768
rect 6938 3670 6972 3732
rect 8126 3670 8160 3732
rect 6938 3636 7034 3670
rect 8064 3636 8160 3670
rect -2062 2844 -1966 2878
rect -936 2844 -840 2878
rect -2062 2782 -2028 2844
rect -874 2782 -840 2844
rect -1964 2742 -1948 2776
rect -1914 2742 -1898 2776
rect -1772 2742 -1756 2776
rect -1722 2742 -1706 2776
rect -1580 2742 -1564 2776
rect -1530 2742 -1514 2776
rect -1388 2742 -1372 2776
rect -1338 2742 -1322 2776
rect -1196 2742 -1180 2776
rect -1146 2742 -1130 2776
rect -1004 2742 -988 2776
rect -954 2742 -938 2776
rect -1948 2682 -1914 2698
rect -1948 2418 -1914 2434
rect -1852 2682 -1818 2698
rect -1852 2418 -1818 2434
rect -1756 2682 -1722 2698
rect -1756 2418 -1722 2434
rect -1660 2682 -1626 2698
rect -1660 2418 -1626 2434
rect -1564 2682 -1530 2698
rect -1564 2418 -1530 2434
rect -1468 2682 -1434 2698
rect -1468 2418 -1434 2434
rect -1372 2682 -1338 2698
rect -1372 2418 -1338 2434
rect -1276 2682 -1242 2698
rect -1276 2418 -1242 2434
rect -1180 2682 -1146 2698
rect -1180 2418 -1146 2434
rect -1084 2682 -1050 2698
rect -1084 2418 -1050 2434
rect -988 2682 -954 2698
rect -988 2418 -954 2434
rect -2062 2334 -2028 2396
rect -874 2334 -840 2396
rect -2062 2300 -1966 2334
rect -936 2300 -840 2334
rect 6938 2844 7034 2878
rect 8064 2844 8160 2878
rect 6938 2782 6972 2844
rect 8126 2782 8160 2844
rect 7036 2742 7052 2776
rect 7086 2742 7102 2776
rect 7228 2742 7244 2776
rect 7278 2742 7294 2776
rect 7420 2742 7436 2776
rect 7470 2742 7486 2776
rect 7612 2742 7628 2776
rect 7662 2742 7678 2776
rect 7804 2742 7820 2776
rect 7854 2742 7870 2776
rect 7996 2742 8012 2776
rect 8046 2742 8062 2776
rect 7052 2682 7086 2698
rect 7052 2418 7086 2434
rect 7148 2682 7182 2698
rect 7148 2418 7182 2434
rect 7244 2682 7278 2698
rect 7244 2418 7278 2434
rect 7340 2682 7374 2698
rect 7340 2418 7374 2434
rect 7436 2682 7470 2698
rect 7436 2418 7470 2434
rect 7532 2682 7566 2698
rect 7532 2418 7566 2434
rect 7628 2682 7662 2698
rect 7628 2418 7662 2434
rect 7724 2682 7758 2698
rect 7724 2418 7758 2434
rect 7820 2682 7854 2698
rect 7820 2418 7854 2434
rect 7916 2682 7950 2698
rect 7916 2418 7950 2434
rect 8012 2682 8046 2698
rect 8012 2418 8046 2434
rect 6938 2334 6972 2396
rect 8126 2334 8160 2396
rect 6938 2300 7034 2334
rect 8064 2300 8160 2334
rect -2062 2192 -1966 2226
rect -936 2192 -840 2226
rect -2062 2132 -2028 2192
rect -874 2130 -840 2192
rect -1948 2102 -1914 2118
rect -1948 2006 -1914 2022
rect -1852 2102 -1818 2118
rect -1852 2006 -1818 2022
rect -1756 2102 -1722 2118
rect -1756 2006 -1722 2022
rect -1660 2102 -1626 2118
rect -1660 2006 -1626 2022
rect -1564 2102 -1530 2118
rect -1564 2006 -1530 2022
rect -1468 2102 -1434 2118
rect -1468 2006 -1434 2022
rect -1372 2102 -1338 2118
rect -1372 2006 -1338 2022
rect -1276 2102 -1242 2118
rect -1276 2006 -1242 2022
rect -1180 2102 -1146 2118
rect -1180 2006 -1146 2022
rect -1084 2102 -1050 2118
rect -1084 2006 -1050 2022
rect -988 2102 -954 2118
rect -988 2006 -954 2022
rect -1964 1934 -1948 1968
rect -1914 1934 -1898 1968
rect -1772 1934 -1756 1968
rect -1722 1934 -1706 1968
rect -1580 1934 -1564 1968
rect -1530 1934 -1514 1968
rect -1388 1934 -1372 1968
rect -1338 1934 -1322 1968
rect -1196 1934 -1180 1968
rect -1146 1934 -1130 1968
rect -1004 1934 -988 1968
rect -954 1934 -938 1968
rect -2062 1870 -2028 1932
rect -874 1870 -840 1932
rect -2062 1836 -1966 1870
rect -936 1836 -840 1870
rect 6938 2192 7034 2226
rect 8064 2192 8160 2226
rect 6938 2132 6972 2192
rect 8126 2130 8160 2192
rect 7052 2102 7086 2118
rect 7052 2006 7086 2022
rect 7148 2102 7182 2118
rect 7148 2006 7182 2022
rect 7244 2102 7278 2118
rect 7244 2006 7278 2022
rect 7340 2102 7374 2118
rect 7340 2006 7374 2022
rect 7436 2102 7470 2118
rect 7436 2006 7470 2022
rect 7532 2102 7566 2118
rect 7532 2006 7566 2022
rect 7628 2102 7662 2118
rect 7628 2006 7662 2022
rect 7724 2102 7758 2118
rect 7724 2006 7758 2022
rect 7820 2102 7854 2118
rect 7820 2006 7854 2022
rect 7916 2102 7950 2118
rect 7916 2006 7950 2022
rect 8012 2102 8046 2118
rect 8012 2006 8046 2022
rect 7036 1934 7052 1968
rect 7086 1934 7102 1968
rect 7228 1934 7244 1968
rect 7278 1934 7294 1968
rect 7420 1934 7436 1968
rect 7470 1934 7486 1968
rect 7612 1934 7628 1968
rect 7662 1934 7678 1968
rect 7804 1934 7820 1968
rect 7854 1934 7870 1968
rect 7996 1934 8012 1968
rect 8046 1934 8062 1968
rect 6938 1870 6972 1932
rect 8126 1870 8160 1932
rect 6938 1836 7034 1870
rect 8064 1836 8160 1870
rect -2062 1044 -1966 1078
rect -936 1044 -840 1078
rect -2062 982 -2028 1044
rect -874 982 -840 1044
rect -1964 942 -1948 976
rect -1914 942 -1898 976
rect -1772 942 -1756 976
rect -1722 942 -1706 976
rect -1580 942 -1564 976
rect -1530 942 -1514 976
rect -1388 942 -1372 976
rect -1338 942 -1322 976
rect -1196 942 -1180 976
rect -1146 942 -1130 976
rect -1004 942 -988 976
rect -954 942 -938 976
rect -1948 882 -1914 898
rect -1948 618 -1914 634
rect -1852 882 -1818 898
rect -1852 618 -1818 634
rect -1756 882 -1722 898
rect -1756 618 -1722 634
rect -1660 882 -1626 898
rect -1660 618 -1626 634
rect -1564 882 -1530 898
rect -1564 618 -1530 634
rect -1468 882 -1434 898
rect -1468 618 -1434 634
rect -1372 882 -1338 898
rect -1372 618 -1338 634
rect -1276 882 -1242 898
rect -1276 618 -1242 634
rect -1180 882 -1146 898
rect -1180 618 -1146 634
rect -1084 882 -1050 898
rect -1084 618 -1050 634
rect -988 882 -954 898
rect -988 618 -954 634
rect -2062 534 -2028 596
rect -874 534 -840 596
rect -2062 500 -1966 534
rect -936 500 -840 534
rect 6938 1044 7034 1078
rect 8064 1044 8160 1078
rect 6938 982 6972 1044
rect 8126 982 8160 1044
rect 7036 942 7052 976
rect 7086 942 7102 976
rect 7228 942 7244 976
rect 7278 942 7294 976
rect 7420 942 7436 976
rect 7470 942 7486 976
rect 7612 942 7628 976
rect 7662 942 7678 976
rect 7804 942 7820 976
rect 7854 942 7870 976
rect 7996 942 8012 976
rect 8046 942 8062 976
rect 7052 882 7086 898
rect 7052 618 7086 634
rect 7148 882 7182 898
rect 7148 618 7182 634
rect 7244 882 7278 898
rect 7244 618 7278 634
rect 7340 882 7374 898
rect 7340 618 7374 634
rect 7436 882 7470 898
rect 7436 618 7470 634
rect 7532 882 7566 898
rect 7532 618 7566 634
rect 7628 882 7662 898
rect 7628 618 7662 634
rect 7724 882 7758 898
rect 7724 618 7758 634
rect 7820 882 7854 898
rect 7820 618 7854 634
rect 7916 882 7950 898
rect 7916 618 7950 634
rect 8012 882 8046 898
rect 8012 618 8046 634
rect 6938 534 6972 596
rect 8126 534 8160 596
rect 6938 500 7034 534
rect 8064 500 8160 534
rect -2062 392 -1966 426
rect -936 392 -840 426
rect -2062 332 -2028 392
rect -874 330 -840 392
rect -1948 302 -1914 318
rect -1948 206 -1914 222
rect -1852 302 -1818 318
rect -1852 206 -1818 222
rect -1756 302 -1722 318
rect -1756 206 -1722 222
rect -1660 302 -1626 318
rect -1660 206 -1626 222
rect -1564 302 -1530 318
rect -1564 206 -1530 222
rect -1468 302 -1434 318
rect -1468 206 -1434 222
rect -1372 302 -1338 318
rect -1372 206 -1338 222
rect -1276 302 -1242 318
rect -1276 206 -1242 222
rect -1180 302 -1146 318
rect -1180 206 -1146 222
rect -1084 302 -1050 318
rect -1084 206 -1050 222
rect -988 302 -954 318
rect -988 206 -954 222
rect -1964 134 -1948 168
rect -1914 134 -1898 168
rect -1772 134 -1756 168
rect -1722 134 -1706 168
rect -1580 134 -1564 168
rect -1530 134 -1514 168
rect -1388 134 -1372 168
rect -1338 134 -1322 168
rect -1196 134 -1180 168
rect -1146 134 -1130 168
rect -1004 134 -988 168
rect -954 134 -938 168
rect -2062 70 -2028 132
rect -874 70 -840 132
rect -2062 36 -1966 70
rect -936 36 -840 70
rect 6938 392 7034 426
rect 8064 392 8160 426
rect 6938 332 6972 392
rect 8126 330 8160 392
rect 7052 302 7086 318
rect 7052 206 7086 222
rect 7148 302 7182 318
rect 7148 206 7182 222
rect 7244 302 7278 318
rect 7244 206 7278 222
rect 7340 302 7374 318
rect 7340 206 7374 222
rect 7436 302 7470 318
rect 7436 206 7470 222
rect 7532 302 7566 318
rect 7532 206 7566 222
rect 7628 302 7662 318
rect 7628 206 7662 222
rect 7724 302 7758 318
rect 7724 206 7758 222
rect 7820 302 7854 318
rect 7820 206 7854 222
rect 7916 302 7950 318
rect 7916 206 7950 222
rect 8012 302 8046 318
rect 8012 206 8046 222
rect 7036 134 7052 168
rect 7086 134 7102 168
rect 7228 134 7244 168
rect 7278 134 7294 168
rect 7420 134 7436 168
rect 7470 134 7486 168
rect 7612 134 7628 168
rect 7662 134 7678 168
rect 7804 134 7820 168
rect 7854 134 7870 168
rect 7996 134 8012 168
rect 8046 134 8062 168
rect 6938 70 6972 132
rect 8126 70 8160 132
rect 6938 36 7034 70
rect 8064 36 8160 70
rect -2062 -756 -1966 -722
rect -936 -756 -840 -722
rect -2062 -818 -2028 -756
rect -874 -818 -840 -756
rect -1964 -858 -1948 -824
rect -1914 -858 -1898 -824
rect -1772 -858 -1756 -824
rect -1722 -858 -1706 -824
rect -1580 -858 -1564 -824
rect -1530 -858 -1514 -824
rect -1388 -858 -1372 -824
rect -1338 -858 -1322 -824
rect -1196 -858 -1180 -824
rect -1146 -858 -1130 -824
rect -1004 -858 -988 -824
rect -954 -858 -938 -824
rect -1948 -918 -1914 -902
rect -1948 -1182 -1914 -1166
rect -1852 -918 -1818 -902
rect -1852 -1182 -1818 -1166
rect -1756 -918 -1722 -902
rect -1756 -1182 -1722 -1166
rect -1660 -918 -1626 -902
rect -1660 -1182 -1626 -1166
rect -1564 -918 -1530 -902
rect -1564 -1182 -1530 -1166
rect -1468 -918 -1434 -902
rect -1468 -1182 -1434 -1166
rect -1372 -918 -1338 -902
rect -1372 -1182 -1338 -1166
rect -1276 -918 -1242 -902
rect -1276 -1182 -1242 -1166
rect -1180 -918 -1146 -902
rect -1180 -1182 -1146 -1166
rect -1084 -918 -1050 -902
rect -1084 -1182 -1050 -1166
rect -988 -918 -954 -902
rect -988 -1182 -954 -1166
rect -2062 -1266 -2028 -1204
rect -874 -1266 -840 -1204
rect -2062 -1300 -1966 -1266
rect -936 -1300 -840 -1266
rect 6938 -756 7034 -722
rect 8064 -756 8160 -722
rect 6938 -818 6972 -756
rect 8126 -818 8160 -756
rect 7036 -858 7052 -824
rect 7086 -858 7102 -824
rect 7228 -858 7244 -824
rect 7278 -858 7294 -824
rect 7420 -858 7436 -824
rect 7470 -858 7486 -824
rect 7612 -858 7628 -824
rect 7662 -858 7678 -824
rect 7804 -858 7820 -824
rect 7854 -858 7870 -824
rect 7996 -858 8012 -824
rect 8046 -858 8062 -824
rect 7052 -918 7086 -902
rect 7052 -1182 7086 -1166
rect 7148 -918 7182 -902
rect 7148 -1182 7182 -1166
rect 7244 -918 7278 -902
rect 7244 -1182 7278 -1166
rect 7340 -918 7374 -902
rect 7340 -1182 7374 -1166
rect 7436 -918 7470 -902
rect 7436 -1182 7470 -1166
rect 7532 -918 7566 -902
rect 7532 -1182 7566 -1166
rect 7628 -918 7662 -902
rect 7628 -1182 7662 -1166
rect 7724 -918 7758 -902
rect 7724 -1182 7758 -1166
rect 7820 -918 7854 -902
rect 7820 -1182 7854 -1166
rect 7916 -918 7950 -902
rect 7916 -1182 7950 -1166
rect 8012 -918 8046 -902
rect 8012 -1182 8046 -1166
rect 6938 -1266 6972 -1204
rect 8126 -1266 8160 -1204
rect 6938 -1300 7034 -1266
rect 8064 -1300 8160 -1266
rect -2062 -1408 -1966 -1374
rect -936 -1408 -840 -1374
rect -2062 -1468 -2028 -1408
rect -874 -1470 -840 -1408
rect -1948 -1498 -1914 -1482
rect -1948 -1594 -1914 -1578
rect -1852 -1498 -1818 -1482
rect -1852 -1594 -1818 -1578
rect -1756 -1498 -1722 -1482
rect -1756 -1594 -1722 -1578
rect -1660 -1498 -1626 -1482
rect -1660 -1594 -1626 -1578
rect -1564 -1498 -1530 -1482
rect -1564 -1594 -1530 -1578
rect -1468 -1498 -1434 -1482
rect -1468 -1594 -1434 -1578
rect -1372 -1498 -1338 -1482
rect -1372 -1594 -1338 -1578
rect -1276 -1498 -1242 -1482
rect -1276 -1594 -1242 -1578
rect -1180 -1498 -1146 -1482
rect -1180 -1594 -1146 -1578
rect -1084 -1498 -1050 -1482
rect -1084 -1594 -1050 -1578
rect -988 -1498 -954 -1482
rect -988 -1594 -954 -1578
rect -1964 -1666 -1948 -1632
rect -1914 -1666 -1898 -1632
rect -1772 -1666 -1756 -1632
rect -1722 -1666 -1706 -1632
rect -1580 -1666 -1564 -1632
rect -1530 -1666 -1514 -1632
rect -1388 -1666 -1372 -1632
rect -1338 -1666 -1322 -1632
rect -1196 -1666 -1180 -1632
rect -1146 -1666 -1130 -1632
rect -1004 -1666 -988 -1632
rect -954 -1666 -938 -1632
rect -2062 -1730 -2028 -1668
rect -874 -1730 -840 -1668
rect -2062 -1764 -1966 -1730
rect -936 -1764 -840 -1730
rect 6938 -1408 7034 -1374
rect 8064 -1408 8160 -1374
rect 6938 -1468 6972 -1408
rect 8126 -1470 8160 -1408
rect 7052 -1498 7086 -1482
rect 7052 -1594 7086 -1578
rect 7148 -1498 7182 -1482
rect 7148 -1594 7182 -1578
rect 7244 -1498 7278 -1482
rect 7244 -1594 7278 -1578
rect 7340 -1498 7374 -1482
rect 7340 -1594 7374 -1578
rect 7436 -1498 7470 -1482
rect 7436 -1594 7470 -1578
rect 7532 -1498 7566 -1482
rect 7532 -1594 7566 -1578
rect 7628 -1498 7662 -1482
rect 7628 -1594 7662 -1578
rect 7724 -1498 7758 -1482
rect 7724 -1594 7758 -1578
rect 7820 -1498 7854 -1482
rect 7820 -1594 7854 -1578
rect 7916 -1498 7950 -1482
rect 7916 -1594 7950 -1578
rect 8012 -1498 8046 -1482
rect 8012 -1594 8046 -1578
rect 7036 -1666 7052 -1632
rect 7086 -1666 7102 -1632
rect 7228 -1666 7244 -1632
rect 7278 -1666 7294 -1632
rect 7420 -1666 7436 -1632
rect 7470 -1666 7486 -1632
rect 7612 -1666 7628 -1632
rect 7662 -1666 7678 -1632
rect 7804 -1666 7820 -1632
rect 7854 -1666 7870 -1632
rect 7996 -1666 8012 -1632
rect 8046 -1666 8062 -1632
rect 6938 -1730 6972 -1668
rect 8126 -1730 8160 -1668
rect 6938 -1764 7034 -1730
rect 8064 -1764 8160 -1730
<< viali >>
rect -2062 7796 -2028 8182
rect -1948 8142 -1914 8176
rect -1756 8142 -1722 8176
rect -1564 8142 -1530 8176
rect -1372 8142 -1338 8176
rect -1180 8142 -1146 8176
rect -988 8142 -954 8176
rect -1948 7834 -1914 8082
rect -1852 7834 -1818 8082
rect -1756 7834 -1722 8082
rect -1660 7834 -1626 8082
rect -1564 7834 -1530 8082
rect -1468 7834 -1434 8082
rect -1372 7834 -1338 8082
rect -1276 7834 -1242 8082
rect -1180 7834 -1146 8082
rect -1084 7834 -1050 8082
rect -988 7834 -954 8082
rect 6938 7796 6972 8182
rect 7052 8142 7086 8176
rect 7244 8142 7278 8176
rect 7436 8142 7470 8176
rect 7628 8142 7662 8176
rect 7820 8142 7854 8176
rect 8012 8142 8046 8176
rect 7052 7834 7086 8082
rect 7148 7834 7182 8082
rect 7244 7834 7278 8082
rect 7340 7834 7374 8082
rect 7436 7834 7470 8082
rect 7532 7834 7566 8082
rect 7628 7834 7662 8082
rect 7724 7834 7758 8082
rect 7820 7834 7854 8082
rect 7916 7834 7950 8082
rect 8012 7834 8046 8082
rect -2062 7530 -2028 7532
rect -2062 7332 -2028 7530
rect -1948 7422 -1914 7502
rect -1852 7422 -1818 7502
rect -1756 7422 -1722 7502
rect -1660 7422 -1626 7502
rect -1564 7422 -1530 7502
rect -1468 7422 -1434 7502
rect -1372 7422 -1338 7502
rect -1276 7422 -1242 7502
rect -1180 7422 -1146 7502
rect -1084 7422 -1050 7502
rect -988 7422 -954 7502
rect -1948 7334 -1914 7368
rect -1756 7334 -1722 7368
rect -1564 7334 -1530 7368
rect -1372 7334 -1338 7368
rect -1180 7334 -1146 7368
rect -988 7334 -954 7368
rect 6938 7530 6972 7532
rect 6938 7332 6972 7530
rect 7052 7422 7086 7502
rect 7148 7422 7182 7502
rect 7244 7422 7278 7502
rect 7340 7422 7374 7502
rect 7436 7422 7470 7502
rect 7532 7422 7566 7502
rect 7628 7422 7662 7502
rect 7724 7422 7758 7502
rect 7820 7422 7854 7502
rect 7916 7422 7950 7502
rect 8012 7422 8046 7502
rect 7052 7334 7086 7368
rect 7244 7334 7278 7368
rect 7436 7334 7470 7368
rect 7628 7334 7662 7368
rect 7820 7334 7854 7368
rect 8012 7334 8046 7368
rect -2062 5996 -2028 6382
rect -1948 6342 -1914 6376
rect -1756 6342 -1722 6376
rect -1564 6342 -1530 6376
rect -1372 6342 -1338 6376
rect -1180 6342 -1146 6376
rect -988 6342 -954 6376
rect -1948 6034 -1914 6282
rect -1852 6034 -1818 6282
rect -1756 6034 -1722 6282
rect -1660 6034 -1626 6282
rect -1564 6034 -1530 6282
rect -1468 6034 -1434 6282
rect -1372 6034 -1338 6282
rect -1276 6034 -1242 6282
rect -1180 6034 -1146 6282
rect -1084 6034 -1050 6282
rect -988 6034 -954 6282
rect 6938 5996 6972 6382
rect 7052 6342 7086 6376
rect 7244 6342 7278 6376
rect 7436 6342 7470 6376
rect 7628 6342 7662 6376
rect 7820 6342 7854 6376
rect 8012 6342 8046 6376
rect 7052 6034 7086 6282
rect 7148 6034 7182 6282
rect 7244 6034 7278 6282
rect 7340 6034 7374 6282
rect 7436 6034 7470 6282
rect 7532 6034 7566 6282
rect 7628 6034 7662 6282
rect 7724 6034 7758 6282
rect 7820 6034 7854 6282
rect 7916 6034 7950 6282
rect 8012 6034 8046 6282
rect -2062 5730 -2028 5732
rect -2062 5532 -2028 5730
rect -1948 5622 -1914 5702
rect -1852 5622 -1818 5702
rect -1756 5622 -1722 5702
rect -1660 5622 -1626 5702
rect -1564 5622 -1530 5702
rect -1468 5622 -1434 5702
rect -1372 5622 -1338 5702
rect -1276 5622 -1242 5702
rect -1180 5622 -1146 5702
rect -1084 5622 -1050 5702
rect -988 5622 -954 5702
rect -1948 5534 -1914 5568
rect -1756 5534 -1722 5568
rect -1564 5534 -1530 5568
rect -1372 5534 -1338 5568
rect -1180 5534 -1146 5568
rect -988 5534 -954 5568
rect 6938 5730 6972 5732
rect 6938 5532 6972 5730
rect 7052 5622 7086 5702
rect 7148 5622 7182 5702
rect 7244 5622 7278 5702
rect 7340 5622 7374 5702
rect 7436 5622 7470 5702
rect 7532 5622 7566 5702
rect 7628 5622 7662 5702
rect 7724 5622 7758 5702
rect 7820 5622 7854 5702
rect 7916 5622 7950 5702
rect 8012 5622 8046 5702
rect 7052 5534 7086 5568
rect 7244 5534 7278 5568
rect 7436 5534 7470 5568
rect 7628 5534 7662 5568
rect 7820 5534 7854 5568
rect 8012 5534 8046 5568
rect -2062 4196 -2028 4582
rect -1948 4542 -1914 4576
rect -1756 4542 -1722 4576
rect -1564 4542 -1530 4576
rect -1372 4542 -1338 4576
rect -1180 4542 -1146 4576
rect -988 4542 -954 4576
rect -1948 4234 -1914 4482
rect -1852 4234 -1818 4482
rect -1756 4234 -1722 4482
rect -1660 4234 -1626 4482
rect -1564 4234 -1530 4482
rect -1468 4234 -1434 4482
rect -1372 4234 -1338 4482
rect -1276 4234 -1242 4482
rect -1180 4234 -1146 4482
rect -1084 4234 -1050 4482
rect -988 4234 -954 4482
rect 6938 4196 6972 4582
rect 7052 4542 7086 4576
rect 7244 4542 7278 4576
rect 7436 4542 7470 4576
rect 7628 4542 7662 4576
rect 7820 4542 7854 4576
rect 8012 4542 8046 4576
rect 7052 4234 7086 4482
rect 7148 4234 7182 4482
rect 7244 4234 7278 4482
rect 7340 4234 7374 4482
rect 7436 4234 7470 4482
rect 7532 4234 7566 4482
rect 7628 4234 7662 4482
rect 7724 4234 7758 4482
rect 7820 4234 7854 4482
rect 7916 4234 7950 4482
rect 8012 4234 8046 4482
rect -2062 3930 -2028 3932
rect -2062 3732 -2028 3930
rect -1948 3822 -1914 3902
rect -1852 3822 -1818 3902
rect -1756 3822 -1722 3902
rect -1660 3822 -1626 3902
rect -1564 3822 -1530 3902
rect -1468 3822 -1434 3902
rect -1372 3822 -1338 3902
rect -1276 3822 -1242 3902
rect -1180 3822 -1146 3902
rect -1084 3822 -1050 3902
rect -988 3822 -954 3902
rect -1948 3734 -1914 3768
rect -1756 3734 -1722 3768
rect -1564 3734 -1530 3768
rect -1372 3734 -1338 3768
rect -1180 3734 -1146 3768
rect -988 3734 -954 3768
rect 6938 3930 6972 3932
rect 6938 3732 6972 3930
rect 7052 3822 7086 3902
rect 7148 3822 7182 3902
rect 7244 3822 7278 3902
rect 7340 3822 7374 3902
rect 7436 3822 7470 3902
rect 7532 3822 7566 3902
rect 7628 3822 7662 3902
rect 7724 3822 7758 3902
rect 7820 3822 7854 3902
rect 7916 3822 7950 3902
rect 8012 3822 8046 3902
rect 7052 3734 7086 3768
rect 7244 3734 7278 3768
rect 7436 3734 7470 3768
rect 7628 3734 7662 3768
rect 7820 3734 7854 3768
rect 8012 3734 8046 3768
rect -2062 2396 -2028 2782
rect -1948 2742 -1914 2776
rect -1756 2742 -1722 2776
rect -1564 2742 -1530 2776
rect -1372 2742 -1338 2776
rect -1180 2742 -1146 2776
rect -988 2742 -954 2776
rect -1948 2434 -1914 2682
rect -1852 2434 -1818 2682
rect -1756 2434 -1722 2682
rect -1660 2434 -1626 2682
rect -1564 2434 -1530 2682
rect -1468 2434 -1434 2682
rect -1372 2434 -1338 2682
rect -1276 2434 -1242 2682
rect -1180 2434 -1146 2682
rect -1084 2434 -1050 2682
rect -988 2434 -954 2682
rect 6938 2396 6972 2782
rect 7052 2742 7086 2776
rect 7244 2742 7278 2776
rect 7436 2742 7470 2776
rect 7628 2742 7662 2776
rect 7820 2742 7854 2776
rect 8012 2742 8046 2776
rect 7052 2434 7086 2682
rect 7148 2434 7182 2682
rect 7244 2434 7278 2682
rect 7340 2434 7374 2682
rect 7436 2434 7470 2682
rect 7532 2434 7566 2682
rect 7628 2434 7662 2682
rect 7724 2434 7758 2682
rect 7820 2434 7854 2682
rect 7916 2434 7950 2682
rect 8012 2434 8046 2682
rect -2062 2130 -2028 2132
rect -2062 1932 -2028 2130
rect -1948 2022 -1914 2102
rect -1852 2022 -1818 2102
rect -1756 2022 -1722 2102
rect -1660 2022 -1626 2102
rect -1564 2022 -1530 2102
rect -1468 2022 -1434 2102
rect -1372 2022 -1338 2102
rect -1276 2022 -1242 2102
rect -1180 2022 -1146 2102
rect -1084 2022 -1050 2102
rect -988 2022 -954 2102
rect -1948 1934 -1914 1968
rect -1756 1934 -1722 1968
rect -1564 1934 -1530 1968
rect -1372 1934 -1338 1968
rect -1180 1934 -1146 1968
rect -988 1934 -954 1968
rect 6938 2130 6972 2132
rect 6938 1932 6972 2130
rect 7052 2022 7086 2102
rect 7148 2022 7182 2102
rect 7244 2022 7278 2102
rect 7340 2022 7374 2102
rect 7436 2022 7470 2102
rect 7532 2022 7566 2102
rect 7628 2022 7662 2102
rect 7724 2022 7758 2102
rect 7820 2022 7854 2102
rect 7916 2022 7950 2102
rect 8012 2022 8046 2102
rect 7052 1934 7086 1968
rect 7244 1934 7278 1968
rect 7436 1934 7470 1968
rect 7628 1934 7662 1968
rect 7820 1934 7854 1968
rect 8012 1934 8046 1968
rect -2062 596 -2028 982
rect -1948 942 -1914 976
rect -1756 942 -1722 976
rect -1564 942 -1530 976
rect -1372 942 -1338 976
rect -1180 942 -1146 976
rect -988 942 -954 976
rect -1948 634 -1914 882
rect -1852 634 -1818 882
rect -1756 634 -1722 882
rect -1660 634 -1626 882
rect -1564 634 -1530 882
rect -1468 634 -1434 882
rect -1372 634 -1338 882
rect -1276 634 -1242 882
rect -1180 634 -1146 882
rect -1084 634 -1050 882
rect -988 634 -954 882
rect 6938 596 6972 982
rect 7052 942 7086 976
rect 7244 942 7278 976
rect 7436 942 7470 976
rect 7628 942 7662 976
rect 7820 942 7854 976
rect 8012 942 8046 976
rect 7052 634 7086 882
rect 7148 634 7182 882
rect 7244 634 7278 882
rect 7340 634 7374 882
rect 7436 634 7470 882
rect 7532 634 7566 882
rect 7628 634 7662 882
rect 7724 634 7758 882
rect 7820 634 7854 882
rect 7916 634 7950 882
rect 8012 634 8046 882
rect -2062 330 -2028 332
rect -2062 132 -2028 330
rect -1948 222 -1914 302
rect -1852 222 -1818 302
rect -1756 222 -1722 302
rect -1660 222 -1626 302
rect -1564 222 -1530 302
rect -1468 222 -1434 302
rect -1372 222 -1338 302
rect -1276 222 -1242 302
rect -1180 222 -1146 302
rect -1084 222 -1050 302
rect -988 222 -954 302
rect -1948 134 -1914 168
rect -1756 134 -1722 168
rect -1564 134 -1530 168
rect -1372 134 -1338 168
rect -1180 134 -1146 168
rect -988 134 -954 168
rect 6938 330 6972 332
rect 6938 132 6972 330
rect 7052 222 7086 302
rect 7148 222 7182 302
rect 7244 222 7278 302
rect 7340 222 7374 302
rect 7436 222 7470 302
rect 7532 222 7566 302
rect 7628 222 7662 302
rect 7724 222 7758 302
rect 7820 222 7854 302
rect 7916 222 7950 302
rect 8012 222 8046 302
rect 7052 134 7086 168
rect 7244 134 7278 168
rect 7436 134 7470 168
rect 7628 134 7662 168
rect 7820 134 7854 168
rect 8012 134 8046 168
rect -2062 -1204 -2028 -818
rect -1948 -858 -1914 -824
rect -1756 -858 -1722 -824
rect -1564 -858 -1530 -824
rect -1372 -858 -1338 -824
rect -1180 -858 -1146 -824
rect -988 -858 -954 -824
rect -1948 -1166 -1914 -918
rect -1852 -1166 -1818 -918
rect -1756 -1166 -1722 -918
rect -1660 -1166 -1626 -918
rect -1564 -1166 -1530 -918
rect -1468 -1166 -1434 -918
rect -1372 -1166 -1338 -918
rect -1276 -1166 -1242 -918
rect -1180 -1166 -1146 -918
rect -1084 -1166 -1050 -918
rect -988 -1166 -954 -918
rect 6938 -1204 6972 -818
rect 7052 -858 7086 -824
rect 7244 -858 7278 -824
rect 7436 -858 7470 -824
rect 7628 -858 7662 -824
rect 7820 -858 7854 -824
rect 8012 -858 8046 -824
rect 7052 -1166 7086 -918
rect 7148 -1166 7182 -918
rect 7244 -1166 7278 -918
rect 7340 -1166 7374 -918
rect 7436 -1166 7470 -918
rect 7532 -1166 7566 -918
rect 7628 -1166 7662 -918
rect 7724 -1166 7758 -918
rect 7820 -1166 7854 -918
rect 7916 -1166 7950 -918
rect 8012 -1166 8046 -918
rect -2062 -1470 -2028 -1468
rect -2062 -1668 -2028 -1470
rect -1948 -1578 -1914 -1498
rect -1852 -1578 -1818 -1498
rect -1756 -1578 -1722 -1498
rect -1660 -1578 -1626 -1498
rect -1564 -1578 -1530 -1498
rect -1468 -1578 -1434 -1498
rect -1372 -1578 -1338 -1498
rect -1276 -1578 -1242 -1498
rect -1180 -1578 -1146 -1498
rect -1084 -1578 -1050 -1498
rect -988 -1578 -954 -1498
rect -1948 -1666 -1914 -1632
rect -1756 -1666 -1722 -1632
rect -1564 -1666 -1530 -1632
rect -1372 -1666 -1338 -1632
rect -1180 -1666 -1146 -1632
rect -988 -1666 -954 -1632
rect 6938 -1470 6972 -1468
rect 6938 -1668 6972 -1470
rect 7052 -1578 7086 -1498
rect 7148 -1578 7182 -1498
rect 7244 -1578 7278 -1498
rect 7340 -1578 7374 -1498
rect 7436 -1578 7470 -1498
rect 7532 -1578 7566 -1498
rect 7628 -1578 7662 -1498
rect 7724 -1578 7758 -1498
rect 7820 -1578 7854 -1498
rect 7916 -1578 7950 -1498
rect 8012 -1578 8046 -1498
rect 7052 -1666 7086 -1632
rect 7244 -1666 7278 -1632
rect 7436 -1666 7470 -1632
rect 7628 -1666 7662 -1632
rect 7820 -1666 7854 -1632
rect 8012 -1666 8046 -1632
<< metal1 >>
rect -2068 8182 -2022 8360
rect -1852 8244 -770 8278
rect -2068 7796 -2062 8182
rect -2028 7796 -2022 8182
rect -1967 8134 -1957 8186
rect -1905 8134 -1895 8186
rect -1852 8094 -1818 8244
rect -1775 8134 -1765 8186
rect -1713 8134 -1703 8186
rect -1660 8094 -1626 8244
rect -1583 8134 -1573 8186
rect -1521 8134 -1511 8186
rect -1468 8094 -1434 8244
rect -1391 8134 -1381 8186
rect -1329 8134 -1319 8186
rect -1276 8094 -1242 8244
rect -1200 8134 -1190 8186
rect -1138 8134 -1128 8186
rect -1084 8094 -1050 8244
rect -1007 8134 -997 8186
rect -945 8134 -935 8186
rect -1954 8082 -1908 8094
rect -1954 7834 -1948 8082
rect -1914 7834 -1908 8082
rect -1954 7822 -1908 7834
rect -1858 8082 -1812 8094
rect -1858 7834 -1852 8082
rect -1818 7834 -1812 8082
rect -1858 7822 -1812 7834
rect -1762 8082 -1716 8094
rect -1762 7834 -1756 8082
rect -1722 7834 -1716 8082
rect -1762 7822 -1716 7834
rect -1666 8082 -1620 8094
rect -1666 7834 -1660 8082
rect -1626 7834 -1620 8082
rect -1666 7822 -1620 7834
rect -1570 8082 -1524 8094
rect -1570 7834 -1564 8082
rect -1530 7834 -1524 8082
rect -1570 7822 -1524 7834
rect -1474 8082 -1428 8094
rect -1474 7834 -1468 8082
rect -1434 7834 -1428 8082
rect -1474 7822 -1428 7834
rect -1378 8082 -1332 8094
rect -1378 7834 -1372 8082
rect -1338 7834 -1332 8082
rect -1378 7822 -1332 7834
rect -1282 8082 -1236 8094
rect -1282 7834 -1276 8082
rect -1242 7834 -1236 8082
rect -1282 7822 -1236 7834
rect -1186 8082 -1140 8094
rect -1186 7834 -1180 8082
rect -1146 7834 -1140 8082
rect -1186 7822 -1140 7834
rect -1090 8082 -1044 8094
rect -1090 7834 -1084 8082
rect -1050 7834 -1044 8082
rect -1090 7822 -1044 7834
rect -994 8082 -948 8094
rect -994 7834 -988 8082
rect -954 7834 -948 8082
rect -994 7822 -948 7834
rect -2068 7784 -2022 7796
rect -1948 7681 -1914 7822
rect -1756 7681 -1722 7822
rect -1564 7681 -1530 7822
rect -1372 7681 -1338 7822
rect -1180 7681 -1146 7822
rect -988 7695 -954 7822
rect -1032 7681 -1022 7695
rect -3494 7647 -1022 7681
rect -3494 -1319 -3419 7647
rect -2068 7532 -2022 7544
rect -2068 7332 -2062 7532
rect -2028 7332 -2022 7532
rect -1948 7514 -1914 7647
rect -1756 7514 -1722 7647
rect -1564 7514 -1530 7647
rect -1372 7514 -1338 7647
rect -1180 7514 -1146 7647
rect -1032 7631 -1022 7647
rect -958 7631 -948 7695
rect -804 7681 -770 8244
rect -730 8134 -720 8186
rect -668 8134 -641 8186
rect 6932 8182 6978 8360
rect 7148 8244 8230 8278
rect 6932 7796 6938 8182
rect 6972 7796 6978 8182
rect 7033 8134 7043 8186
rect 7095 8134 7105 8186
rect 7148 8094 7182 8244
rect 7225 8134 7235 8186
rect 7287 8134 7297 8186
rect 7340 8094 7374 8244
rect 7417 8134 7427 8186
rect 7479 8134 7489 8186
rect 7532 8094 7566 8244
rect 7609 8134 7619 8186
rect 7671 8134 7681 8186
rect 7724 8094 7758 8244
rect 7800 8134 7810 8186
rect 7862 8134 7872 8186
rect 7916 8094 7950 8244
rect 7993 8134 8003 8186
rect 8055 8134 8065 8186
rect 7046 8082 7092 8094
rect 7046 7834 7052 8082
rect 7086 7834 7092 8082
rect 7046 7822 7092 7834
rect 7142 8082 7188 8094
rect 7142 7834 7148 8082
rect 7182 7834 7188 8082
rect 7142 7822 7188 7834
rect 7238 8082 7284 8094
rect 7238 7834 7244 8082
rect 7278 7834 7284 8082
rect 7238 7822 7284 7834
rect 7334 8082 7380 8094
rect 7334 7834 7340 8082
rect 7374 7834 7380 8082
rect 7334 7822 7380 7834
rect 7430 8082 7476 8094
rect 7430 7834 7436 8082
rect 7470 7834 7476 8082
rect 7430 7822 7476 7834
rect 7526 8082 7572 8094
rect 7526 7834 7532 8082
rect 7566 7834 7572 8082
rect 7526 7822 7572 7834
rect 7622 8082 7668 8094
rect 7622 7834 7628 8082
rect 7662 7834 7668 8082
rect 7622 7822 7668 7834
rect 7718 8082 7764 8094
rect 7718 7834 7724 8082
rect 7758 7834 7764 8082
rect 7718 7822 7764 7834
rect 7814 8082 7860 8094
rect 7814 7834 7820 8082
rect 7854 7834 7860 8082
rect 7814 7822 7860 7834
rect 7910 8082 7956 8094
rect 7910 7834 7916 8082
rect 7950 7834 7956 8082
rect 7910 7822 7956 7834
rect 8006 8082 8052 8094
rect 8006 7834 8012 8082
rect 8046 7834 8052 8082
rect 8006 7822 8052 7834
rect 6932 7784 6978 7796
rect -485 7681 2411 7697
rect -804 7647 2411 7681
rect -988 7514 -954 7631
rect -1954 7502 -1908 7514
rect -1954 7422 -1948 7502
rect -1914 7422 -1908 7502
rect -1954 7410 -1908 7422
rect -1858 7502 -1812 7514
rect -1858 7422 -1852 7502
rect -1818 7422 -1812 7502
rect -1858 7410 -1812 7422
rect -1762 7502 -1716 7514
rect -1762 7422 -1756 7502
rect -1722 7422 -1716 7502
rect -1762 7410 -1716 7422
rect -1666 7502 -1620 7514
rect -1666 7422 -1660 7502
rect -1626 7422 -1620 7502
rect -1666 7410 -1620 7422
rect -1570 7502 -1524 7514
rect -1570 7422 -1564 7502
rect -1530 7422 -1524 7502
rect -1570 7410 -1524 7422
rect -1474 7502 -1428 7514
rect -1474 7422 -1468 7502
rect -1434 7422 -1428 7502
rect -1474 7410 -1428 7422
rect -1378 7502 -1332 7514
rect -1378 7422 -1372 7502
rect -1338 7422 -1332 7502
rect -1378 7410 -1332 7422
rect -1282 7502 -1236 7514
rect -1282 7422 -1276 7502
rect -1242 7422 -1236 7502
rect -1282 7410 -1236 7422
rect -1186 7502 -1140 7514
rect -1186 7422 -1180 7502
rect -1146 7422 -1140 7502
rect -1186 7410 -1140 7422
rect -1090 7502 -1044 7514
rect -1090 7422 -1084 7502
rect -1050 7422 -1044 7502
rect -1090 7410 -1044 7422
rect -994 7502 -948 7514
rect -994 7422 -988 7502
rect -954 7422 -948 7502
rect -994 7410 -948 7422
rect -1964 7378 -1898 7382
rect -2068 7160 -2022 7332
rect -1967 7326 -1957 7378
rect -1905 7326 -1895 7378
rect -1964 7322 -1898 7326
rect -1852 7270 -1818 7410
rect -1772 7378 -1706 7382
rect -1775 7326 -1765 7378
rect -1713 7326 -1703 7378
rect -1772 7322 -1706 7326
rect -1660 7270 -1626 7410
rect -1580 7379 -1514 7382
rect -1582 7327 -1572 7379
rect -1520 7327 -1510 7379
rect -1580 7322 -1514 7327
rect -1468 7270 -1434 7410
rect -1388 7379 -1322 7382
rect -1390 7327 -1380 7379
rect -1328 7327 -1318 7379
rect -1388 7322 -1322 7327
rect -1276 7270 -1242 7410
rect -1196 7379 -1130 7382
rect -1198 7327 -1188 7379
rect -1136 7327 -1126 7379
rect -1196 7322 -1130 7327
rect -1084 7270 -1050 7410
rect -1004 7379 -938 7382
rect -1007 7327 -997 7379
rect -945 7327 -935 7379
rect -1004 7322 -938 7327
rect -804 7270 -770 7647
rect -485 7633 2411 7647
rect 6681 7633 6691 7697
rect 6755 7681 6765 7697
rect 7052 7681 7086 7822
rect 7244 7681 7278 7822
rect 7436 7681 7470 7822
rect 7628 7681 7662 7822
rect 7820 7681 7854 7822
rect 8012 7681 8046 7822
rect 6755 7647 8046 7681
rect 6755 7633 6765 7647
rect -730 7327 -720 7379
rect -668 7327 -641 7379
rect -1852 7236 -770 7270
rect -2068 6382 -2022 6560
rect -1852 6444 -770 6478
rect -2068 5996 -2062 6382
rect -2028 5996 -2022 6382
rect -1967 6334 -1957 6386
rect -1905 6334 -1895 6386
rect -1852 6294 -1818 6444
rect -1775 6334 -1765 6386
rect -1713 6334 -1703 6386
rect -1660 6294 -1626 6444
rect -1583 6334 -1573 6386
rect -1521 6334 -1511 6386
rect -1468 6294 -1434 6444
rect -1391 6334 -1381 6386
rect -1329 6334 -1319 6386
rect -1276 6294 -1242 6444
rect -1200 6334 -1190 6386
rect -1138 6334 -1128 6386
rect -1084 6294 -1050 6444
rect -1007 6334 -997 6386
rect -945 6334 -935 6386
rect -1954 6282 -1908 6294
rect -1954 6034 -1948 6282
rect -1914 6034 -1908 6282
rect -1954 6022 -1908 6034
rect -1858 6282 -1812 6294
rect -1858 6034 -1852 6282
rect -1818 6034 -1812 6282
rect -1858 6022 -1812 6034
rect -1762 6282 -1716 6294
rect -1762 6034 -1756 6282
rect -1722 6034 -1716 6282
rect -1762 6022 -1716 6034
rect -1666 6282 -1620 6294
rect -1666 6034 -1660 6282
rect -1626 6034 -1620 6282
rect -1666 6022 -1620 6034
rect -1570 6282 -1524 6294
rect -1570 6034 -1564 6282
rect -1530 6034 -1524 6282
rect -1570 6022 -1524 6034
rect -1474 6282 -1428 6294
rect -1474 6034 -1468 6282
rect -1434 6034 -1428 6282
rect -1474 6022 -1428 6034
rect -1378 6282 -1332 6294
rect -1378 6034 -1372 6282
rect -1338 6034 -1332 6282
rect -1378 6022 -1332 6034
rect -1282 6282 -1236 6294
rect -1282 6034 -1276 6282
rect -1242 6034 -1236 6282
rect -1282 6022 -1236 6034
rect -1186 6282 -1140 6294
rect -1186 6034 -1180 6282
rect -1146 6034 -1140 6282
rect -1186 6022 -1140 6034
rect -1090 6282 -1044 6294
rect -1090 6034 -1084 6282
rect -1050 6034 -1044 6282
rect -1090 6022 -1044 6034
rect -994 6282 -948 6294
rect -994 6034 -988 6282
rect -954 6034 -948 6282
rect -994 6022 -948 6034
rect -2068 5984 -2022 5996
rect -1948 5881 -1914 6022
rect -1756 5881 -1722 6022
rect -1564 5881 -1530 6022
rect -1372 5881 -1338 6022
rect -1180 5881 -1146 6022
rect -988 5895 -954 6022
rect -1038 5881 -1028 5895
rect -2886 5847 -1028 5881
rect -2886 481 -2811 5847
rect -2068 5732 -2022 5744
rect -2068 5532 -2062 5732
rect -2028 5532 -2022 5732
rect -1948 5714 -1914 5847
rect -1756 5714 -1722 5847
rect -1564 5714 -1530 5847
rect -1372 5714 -1338 5847
rect -1180 5714 -1146 5847
rect -1038 5831 -1028 5847
rect -964 5831 -954 5895
rect -988 5714 -954 5831
rect -804 5881 -770 6444
rect 1618 6412 1628 6476
rect 1692 6412 1702 6476
rect -730 6334 -720 6386
rect -668 6334 -641 6386
rect -487 5881 -477 5893
rect -804 5847 -477 5881
rect -1954 5702 -1908 5714
rect -1954 5622 -1948 5702
rect -1914 5622 -1908 5702
rect -1954 5610 -1908 5622
rect -1858 5702 -1812 5714
rect -1858 5622 -1852 5702
rect -1818 5622 -1812 5702
rect -1858 5610 -1812 5622
rect -1762 5702 -1716 5714
rect -1762 5622 -1756 5702
rect -1722 5622 -1716 5702
rect -1762 5610 -1716 5622
rect -1666 5702 -1620 5714
rect -1666 5622 -1660 5702
rect -1626 5622 -1620 5702
rect -1666 5610 -1620 5622
rect -1570 5702 -1524 5714
rect -1570 5622 -1564 5702
rect -1530 5622 -1524 5702
rect -1570 5610 -1524 5622
rect -1474 5702 -1428 5714
rect -1474 5622 -1468 5702
rect -1434 5622 -1428 5702
rect -1474 5610 -1428 5622
rect -1378 5702 -1332 5714
rect -1378 5622 -1372 5702
rect -1338 5622 -1332 5702
rect -1378 5610 -1332 5622
rect -1282 5702 -1236 5714
rect -1282 5622 -1276 5702
rect -1242 5622 -1236 5702
rect -1282 5610 -1236 5622
rect -1186 5702 -1140 5714
rect -1186 5622 -1180 5702
rect -1146 5622 -1140 5702
rect -1186 5610 -1140 5622
rect -1090 5702 -1044 5714
rect -1090 5622 -1084 5702
rect -1050 5622 -1044 5702
rect -1090 5610 -1044 5622
rect -994 5702 -948 5714
rect -994 5622 -988 5702
rect -954 5622 -948 5702
rect -994 5610 -948 5622
rect -1964 5578 -1898 5582
rect -2068 5360 -2022 5532
rect -1967 5526 -1957 5578
rect -1905 5526 -1895 5578
rect -1964 5522 -1898 5526
rect -1852 5470 -1818 5610
rect -1772 5578 -1706 5582
rect -1775 5526 -1765 5578
rect -1713 5526 -1703 5578
rect -1772 5522 -1706 5526
rect -1660 5470 -1626 5610
rect -1580 5579 -1514 5582
rect -1582 5527 -1572 5579
rect -1520 5527 -1510 5579
rect -1580 5522 -1514 5527
rect -1468 5470 -1434 5610
rect -1388 5579 -1322 5582
rect -1390 5527 -1380 5579
rect -1328 5527 -1318 5579
rect -1388 5522 -1322 5527
rect -1276 5470 -1242 5610
rect -1196 5579 -1130 5582
rect -1198 5527 -1188 5579
rect -1136 5527 -1126 5579
rect -1196 5522 -1130 5527
rect -1084 5470 -1050 5610
rect -1004 5579 -938 5582
rect -1007 5527 -997 5579
rect -945 5527 -935 5579
rect -1004 5522 -938 5527
rect -804 5470 -770 5847
rect -487 5829 -477 5847
rect -413 5829 -403 5893
rect -730 5527 -720 5579
rect -668 5527 -641 5579
rect -1852 5436 -770 5470
rect -2068 4582 -2022 4760
rect -1852 4644 -770 4678
rect -2068 4196 -2062 4582
rect -2028 4196 -2022 4582
rect -1967 4534 -1957 4586
rect -1905 4534 -1895 4586
rect -1852 4494 -1818 4644
rect -1775 4534 -1765 4586
rect -1713 4534 -1703 4586
rect -1660 4494 -1626 4644
rect -1583 4534 -1573 4586
rect -1521 4534 -1511 4586
rect -1468 4494 -1434 4644
rect -1391 4534 -1381 4586
rect -1329 4534 -1319 4586
rect -1276 4494 -1242 4644
rect -1200 4534 -1190 4586
rect -1138 4534 -1128 4586
rect -1084 4494 -1050 4644
rect -1007 4534 -997 4586
rect -945 4534 -935 4586
rect -1954 4482 -1908 4494
rect -1954 4234 -1948 4482
rect -1914 4234 -1908 4482
rect -1954 4222 -1908 4234
rect -1858 4482 -1812 4494
rect -1858 4234 -1852 4482
rect -1818 4234 -1812 4482
rect -1858 4222 -1812 4234
rect -1762 4482 -1716 4494
rect -1762 4234 -1756 4482
rect -1722 4234 -1716 4482
rect -1762 4222 -1716 4234
rect -1666 4482 -1620 4494
rect -1666 4234 -1660 4482
rect -1626 4234 -1620 4482
rect -1666 4222 -1620 4234
rect -1570 4482 -1524 4494
rect -1570 4234 -1564 4482
rect -1530 4234 -1524 4482
rect -1570 4222 -1524 4234
rect -1474 4482 -1428 4494
rect -1474 4234 -1468 4482
rect -1434 4234 -1428 4482
rect -1474 4222 -1428 4234
rect -1378 4482 -1332 4494
rect -1378 4234 -1372 4482
rect -1338 4234 -1332 4482
rect -1378 4222 -1332 4234
rect -1282 4482 -1236 4494
rect -1282 4234 -1276 4482
rect -1242 4234 -1236 4482
rect -1282 4222 -1236 4234
rect -1186 4482 -1140 4494
rect -1186 4234 -1180 4482
rect -1146 4234 -1140 4482
rect -1186 4222 -1140 4234
rect -1090 4482 -1044 4494
rect -1090 4234 -1084 4482
rect -1050 4234 -1044 4482
rect -1090 4222 -1044 4234
rect -994 4482 -948 4494
rect -994 4234 -988 4482
rect -954 4234 -948 4482
rect -994 4222 -948 4234
rect -2068 4184 -2022 4196
rect -1948 4081 -1914 4222
rect -1756 4081 -1722 4222
rect -1564 4081 -1530 4222
rect -1372 4081 -1338 4222
rect -1180 4081 -1146 4222
rect -988 4095 -954 4222
rect -1034 4081 -1024 4095
rect -2428 4047 -1024 4081
rect -2428 2281 -2353 4047
rect -2068 3932 -2022 3944
rect -2068 3732 -2062 3932
rect -2028 3732 -2022 3932
rect -1948 3914 -1914 4047
rect -1756 3914 -1722 4047
rect -1564 3914 -1530 4047
rect -1372 3914 -1338 4047
rect -1180 3914 -1146 4047
rect -1034 4031 -1024 4047
rect -960 4031 -950 4095
rect -804 4081 -770 4644
rect -730 4534 -720 4586
rect -668 4534 -641 4586
rect -444 4081 -434 4094
rect -804 4047 -434 4081
rect -988 3914 -954 4031
rect -1954 3902 -1908 3914
rect -1954 3822 -1948 3902
rect -1914 3822 -1908 3902
rect -1954 3810 -1908 3822
rect -1858 3902 -1812 3914
rect -1858 3822 -1852 3902
rect -1818 3822 -1812 3902
rect -1858 3810 -1812 3822
rect -1762 3902 -1716 3914
rect -1762 3822 -1756 3902
rect -1722 3822 -1716 3902
rect -1762 3810 -1716 3822
rect -1666 3902 -1620 3914
rect -1666 3822 -1660 3902
rect -1626 3822 -1620 3902
rect -1666 3810 -1620 3822
rect -1570 3902 -1524 3914
rect -1570 3822 -1564 3902
rect -1530 3822 -1524 3902
rect -1570 3810 -1524 3822
rect -1474 3902 -1428 3914
rect -1474 3822 -1468 3902
rect -1434 3822 -1428 3902
rect -1474 3810 -1428 3822
rect -1378 3902 -1332 3914
rect -1378 3822 -1372 3902
rect -1338 3822 -1332 3902
rect -1378 3810 -1332 3822
rect -1282 3902 -1236 3914
rect -1282 3822 -1276 3902
rect -1242 3822 -1236 3902
rect -1282 3810 -1236 3822
rect -1186 3902 -1140 3914
rect -1186 3822 -1180 3902
rect -1146 3822 -1140 3902
rect -1186 3810 -1140 3822
rect -1090 3902 -1044 3914
rect -1090 3822 -1084 3902
rect -1050 3822 -1044 3902
rect -1090 3810 -1044 3822
rect -994 3902 -948 3914
rect -994 3822 -988 3902
rect -954 3822 -948 3902
rect -994 3810 -948 3822
rect -1964 3778 -1898 3782
rect -2068 3560 -2022 3732
rect -1967 3726 -1957 3778
rect -1905 3726 -1895 3778
rect -1964 3722 -1898 3726
rect -1852 3670 -1818 3810
rect -1772 3778 -1706 3782
rect -1775 3726 -1765 3778
rect -1713 3726 -1703 3778
rect -1772 3722 -1706 3726
rect -1660 3670 -1626 3810
rect -1580 3779 -1514 3782
rect -1582 3727 -1572 3779
rect -1520 3727 -1510 3779
rect -1580 3722 -1514 3727
rect -1468 3670 -1434 3810
rect -1388 3779 -1322 3782
rect -1390 3727 -1380 3779
rect -1328 3727 -1318 3779
rect -1388 3722 -1322 3727
rect -1276 3670 -1242 3810
rect -1196 3779 -1130 3782
rect -1198 3727 -1188 3779
rect -1136 3727 -1126 3779
rect -1196 3722 -1130 3727
rect -1084 3670 -1050 3810
rect -1004 3779 -938 3782
rect -1007 3727 -997 3779
rect -945 3727 -935 3779
rect -1004 3722 -938 3727
rect -804 3670 -770 4047
rect -444 4030 -434 4047
rect -370 4030 -360 4094
rect 1628 3846 1692 6412
rect 2347 4563 2411 7633
rect 6932 7532 6978 7544
rect 6932 7332 6938 7532
rect 6972 7332 6978 7532
rect 7052 7514 7086 7647
rect 7244 7514 7278 7647
rect 7436 7514 7470 7647
rect 7628 7514 7662 7647
rect 7820 7514 7854 7647
rect 8012 7514 8046 7647
rect 8196 7681 8230 8244
rect 8270 8134 8280 8186
rect 8332 8134 8359 8186
rect 8196 7647 9310 7681
rect 7046 7502 7092 7514
rect 7046 7422 7052 7502
rect 7086 7422 7092 7502
rect 7046 7410 7092 7422
rect 7142 7502 7188 7514
rect 7142 7422 7148 7502
rect 7182 7422 7188 7502
rect 7142 7410 7188 7422
rect 7238 7502 7284 7514
rect 7238 7422 7244 7502
rect 7278 7422 7284 7502
rect 7238 7410 7284 7422
rect 7334 7502 7380 7514
rect 7334 7422 7340 7502
rect 7374 7422 7380 7502
rect 7334 7410 7380 7422
rect 7430 7502 7476 7514
rect 7430 7422 7436 7502
rect 7470 7422 7476 7502
rect 7430 7410 7476 7422
rect 7526 7502 7572 7514
rect 7526 7422 7532 7502
rect 7566 7422 7572 7502
rect 7526 7410 7572 7422
rect 7622 7502 7668 7514
rect 7622 7422 7628 7502
rect 7662 7422 7668 7502
rect 7622 7410 7668 7422
rect 7718 7502 7764 7514
rect 7718 7422 7724 7502
rect 7758 7422 7764 7502
rect 7718 7410 7764 7422
rect 7814 7502 7860 7514
rect 7814 7422 7820 7502
rect 7854 7422 7860 7502
rect 7814 7410 7860 7422
rect 7910 7502 7956 7514
rect 7910 7422 7916 7502
rect 7950 7422 7956 7502
rect 7910 7410 7956 7422
rect 8006 7502 8052 7514
rect 8006 7422 8012 7502
rect 8046 7422 8052 7502
rect 8006 7410 8052 7422
rect 7036 7378 7102 7382
rect 6932 7160 6978 7332
rect 7033 7326 7043 7378
rect 7095 7326 7105 7378
rect 7036 7322 7102 7326
rect 7148 7270 7182 7410
rect 7228 7378 7294 7382
rect 7225 7326 7235 7378
rect 7287 7326 7297 7378
rect 7228 7322 7294 7326
rect 7340 7270 7374 7410
rect 7420 7379 7486 7382
rect 7418 7327 7428 7379
rect 7480 7327 7490 7379
rect 7420 7322 7486 7327
rect 7532 7270 7566 7410
rect 7612 7379 7678 7382
rect 7610 7327 7620 7379
rect 7672 7327 7682 7379
rect 7612 7322 7678 7327
rect 7724 7270 7758 7410
rect 7804 7379 7870 7382
rect 7802 7327 7812 7379
rect 7864 7327 7874 7379
rect 7804 7322 7870 7327
rect 7916 7270 7950 7410
rect 7996 7379 8062 7382
rect 7993 7327 8003 7379
rect 8055 7327 8065 7379
rect 7996 7322 8062 7327
rect 8196 7270 8230 7647
rect 8270 7327 8280 7379
rect 8332 7327 8359 7379
rect 7148 7236 8230 7270
rect 6932 6382 6978 6560
rect 7148 6444 8230 6478
rect 6932 5996 6938 6382
rect 6972 5996 6978 6382
rect 7033 6334 7043 6386
rect 7095 6334 7105 6386
rect 7148 6294 7182 6444
rect 7225 6334 7235 6386
rect 7287 6334 7297 6386
rect 7340 6294 7374 6444
rect 7417 6334 7427 6386
rect 7479 6334 7489 6386
rect 7532 6294 7566 6444
rect 7609 6334 7619 6386
rect 7671 6334 7681 6386
rect 7724 6294 7758 6444
rect 7800 6334 7810 6386
rect 7862 6334 7872 6386
rect 7916 6294 7950 6444
rect 7993 6334 8003 6386
rect 8055 6334 8065 6386
rect 7046 6282 7092 6294
rect 7046 6034 7052 6282
rect 7086 6034 7092 6282
rect 7046 6022 7092 6034
rect 7142 6282 7188 6294
rect 7142 6034 7148 6282
rect 7182 6034 7188 6282
rect 7142 6022 7188 6034
rect 7238 6282 7284 6294
rect 7238 6034 7244 6282
rect 7278 6034 7284 6282
rect 7238 6022 7284 6034
rect 7334 6282 7380 6294
rect 7334 6034 7340 6282
rect 7374 6034 7380 6282
rect 7334 6022 7380 6034
rect 7430 6282 7476 6294
rect 7430 6034 7436 6282
rect 7470 6034 7476 6282
rect 7430 6022 7476 6034
rect 7526 6282 7572 6294
rect 7526 6034 7532 6282
rect 7566 6034 7572 6282
rect 7526 6022 7572 6034
rect 7622 6282 7668 6294
rect 7622 6034 7628 6282
rect 7662 6034 7668 6282
rect 7622 6022 7668 6034
rect 7718 6282 7764 6294
rect 7718 6034 7724 6282
rect 7758 6034 7764 6282
rect 7718 6022 7764 6034
rect 7814 6282 7860 6294
rect 7814 6034 7820 6282
rect 7854 6034 7860 6282
rect 7814 6022 7860 6034
rect 7910 6282 7956 6294
rect 7910 6034 7916 6282
rect 7950 6034 7956 6282
rect 7910 6022 7956 6034
rect 8006 6282 8052 6294
rect 8006 6034 8012 6282
rect 8046 6034 8052 6282
rect 8006 6022 8052 6034
rect 6932 5984 6978 5996
rect 6694 5831 6704 5895
rect 6768 5881 6778 5895
rect 7052 5881 7086 6022
rect 7244 5881 7278 6022
rect 7436 5881 7470 6022
rect 7628 5881 7662 6022
rect 7820 5881 7854 6022
rect 8012 5881 8046 6022
rect 6768 5847 8046 5881
rect 6768 5831 6778 5847
rect 6932 5732 6978 5744
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 6932 5532 6938 5732
rect 6972 5532 6978 5732
rect 7052 5714 7086 5847
rect 7244 5714 7278 5847
rect 7436 5714 7470 5847
rect 7628 5714 7662 5847
rect 7820 5714 7854 5847
rect 8012 5714 8046 5847
rect 8196 5881 8230 6444
rect 8270 6334 8280 6386
rect 8332 6334 8359 6386
rect 8196 5847 8799 5881
rect 7046 5702 7092 5714
rect 7046 5622 7052 5702
rect 7086 5622 7092 5702
rect 7046 5610 7092 5622
rect 7142 5702 7188 5714
rect 7142 5622 7148 5702
rect 7182 5622 7188 5702
rect 7142 5610 7188 5622
rect 7238 5702 7284 5714
rect 7238 5622 7244 5702
rect 7278 5622 7284 5702
rect 7238 5610 7284 5622
rect 7334 5702 7380 5714
rect 7334 5622 7340 5702
rect 7374 5622 7380 5702
rect 7334 5610 7380 5622
rect 7430 5702 7476 5714
rect 7430 5622 7436 5702
rect 7470 5622 7476 5702
rect 7430 5610 7476 5622
rect 7526 5702 7572 5714
rect 7526 5622 7532 5702
rect 7566 5622 7572 5702
rect 7526 5610 7572 5622
rect 7622 5702 7668 5714
rect 7622 5622 7628 5702
rect 7662 5622 7668 5702
rect 7622 5610 7668 5622
rect 7718 5702 7764 5714
rect 7718 5622 7724 5702
rect 7758 5622 7764 5702
rect 7718 5610 7764 5622
rect 7814 5702 7860 5714
rect 7814 5622 7820 5702
rect 7854 5622 7860 5702
rect 7814 5610 7860 5622
rect 7910 5702 7956 5714
rect 7910 5622 7916 5702
rect 7950 5622 7956 5702
rect 7910 5610 7956 5622
rect 8006 5702 8052 5714
rect 8006 5622 8012 5702
rect 8046 5622 8052 5702
rect 8006 5610 8052 5622
rect 7036 5578 7102 5582
rect 3157 5084 3221 5494
rect 6932 5360 6978 5532
rect 7033 5526 7043 5578
rect 7095 5526 7105 5578
rect 7036 5522 7102 5526
rect 7148 5470 7182 5610
rect 7228 5578 7294 5582
rect 7225 5526 7235 5578
rect 7287 5526 7297 5578
rect 7228 5522 7294 5526
rect 7340 5470 7374 5610
rect 7420 5579 7486 5582
rect 7418 5527 7428 5579
rect 7480 5527 7490 5579
rect 7420 5522 7486 5527
rect 7532 5470 7566 5610
rect 7612 5579 7678 5582
rect 7610 5527 7620 5579
rect 7672 5527 7682 5579
rect 7612 5522 7678 5527
rect 7724 5470 7758 5610
rect 7804 5579 7870 5582
rect 7802 5527 7812 5579
rect 7864 5527 7874 5579
rect 7804 5522 7870 5527
rect 7916 5470 7950 5610
rect 7996 5579 8062 5582
rect 7993 5527 8003 5579
rect 8055 5527 8065 5579
rect 7996 5522 8062 5527
rect 8196 5470 8230 5847
rect 8270 5527 8280 5579
rect 8332 5527 8359 5579
rect 7148 5436 8230 5470
rect 3147 5020 3157 5084
rect 3221 5020 3231 5084
rect 3831 4928 6166 4932
rect 3758 4864 3768 4928
rect 3832 4868 6166 4928
rect 6230 4868 6240 4932
rect 3832 4864 3842 4868
rect 6932 4582 6978 4760
rect 7148 4644 8230 4678
rect 2347 4499 3106 4563
rect 3170 4499 3180 4563
rect 4874 4326 5207 4390
rect 5271 4326 5281 4390
rect 3298 4148 3308 4212
rect 3372 4148 3382 4212
rect 3308 4085 3372 4148
rect 1628 3782 1866 3846
rect -730 3727 -720 3779
rect -668 3727 -641 3779
rect -1852 3636 -770 3670
rect 323 3419 333 3483
rect 397 3419 1631 3483
rect 1695 3419 1705 3483
rect 1802 3154 1866 3782
rect 323 3090 333 3154
rect 397 3090 1866 3154
rect -2068 2782 -2022 2960
rect -1852 2844 -770 2878
rect -2068 2396 -2062 2782
rect -2028 2396 -2022 2782
rect -1967 2734 -1957 2786
rect -1905 2734 -1895 2786
rect -1852 2694 -1818 2844
rect -1775 2734 -1765 2786
rect -1713 2734 -1703 2786
rect -1660 2694 -1626 2844
rect -1583 2734 -1573 2786
rect -1521 2734 -1511 2786
rect -1468 2694 -1434 2844
rect -1391 2734 -1381 2786
rect -1329 2734 -1319 2786
rect -1276 2694 -1242 2844
rect -1200 2734 -1190 2786
rect -1138 2734 -1128 2786
rect -1084 2694 -1050 2844
rect -1007 2734 -997 2786
rect -945 2734 -935 2786
rect -1954 2682 -1908 2694
rect -1954 2434 -1948 2682
rect -1914 2434 -1908 2682
rect -1954 2422 -1908 2434
rect -1858 2682 -1812 2694
rect -1858 2434 -1852 2682
rect -1818 2434 -1812 2682
rect -1858 2422 -1812 2434
rect -1762 2682 -1716 2694
rect -1762 2434 -1756 2682
rect -1722 2434 -1716 2682
rect -1762 2422 -1716 2434
rect -1666 2682 -1620 2694
rect -1666 2434 -1660 2682
rect -1626 2434 -1620 2682
rect -1666 2422 -1620 2434
rect -1570 2682 -1524 2694
rect -1570 2434 -1564 2682
rect -1530 2434 -1524 2682
rect -1570 2422 -1524 2434
rect -1474 2682 -1428 2694
rect -1474 2434 -1468 2682
rect -1434 2434 -1428 2682
rect -1474 2422 -1428 2434
rect -1378 2682 -1332 2694
rect -1378 2434 -1372 2682
rect -1338 2434 -1332 2682
rect -1378 2422 -1332 2434
rect -1282 2682 -1236 2694
rect -1282 2434 -1276 2682
rect -1242 2434 -1236 2682
rect -1282 2422 -1236 2434
rect -1186 2682 -1140 2694
rect -1186 2434 -1180 2682
rect -1146 2434 -1140 2682
rect -1186 2422 -1140 2434
rect -1090 2682 -1044 2694
rect -1090 2434 -1084 2682
rect -1050 2434 -1044 2682
rect -1090 2422 -1044 2434
rect -994 2682 -948 2694
rect -994 2434 -988 2682
rect -954 2434 -948 2682
rect -994 2422 -948 2434
rect -2068 2384 -2022 2396
rect -1948 2281 -1914 2422
rect -1756 2281 -1722 2422
rect -1564 2281 -1530 2422
rect -1372 2281 -1338 2422
rect -1180 2281 -1146 2422
rect -988 2295 -954 2422
rect -1037 2281 -1027 2295
rect -2428 2247 -1027 2281
rect -2068 2132 -2022 2144
rect -2068 1932 -2062 2132
rect -2028 1932 -2022 2132
rect -1948 2114 -1914 2247
rect -1756 2114 -1722 2247
rect -1564 2114 -1530 2247
rect -1372 2114 -1338 2247
rect -1180 2114 -1146 2247
rect -1037 2231 -1027 2247
rect -963 2231 -953 2295
rect -804 2281 -770 2844
rect -730 2734 -720 2786
rect -668 2734 -641 2786
rect -444 2281 -434 2291
rect -804 2247 -434 2281
rect -988 2114 -954 2231
rect -1954 2102 -1908 2114
rect -1954 2022 -1948 2102
rect -1914 2022 -1908 2102
rect -1954 2010 -1908 2022
rect -1858 2102 -1812 2114
rect -1858 2022 -1852 2102
rect -1818 2022 -1812 2102
rect -1858 2010 -1812 2022
rect -1762 2102 -1716 2114
rect -1762 2022 -1756 2102
rect -1722 2022 -1716 2102
rect -1762 2010 -1716 2022
rect -1666 2102 -1620 2114
rect -1666 2022 -1660 2102
rect -1626 2022 -1620 2102
rect -1666 2010 -1620 2022
rect -1570 2102 -1524 2114
rect -1570 2022 -1564 2102
rect -1530 2022 -1524 2102
rect -1570 2010 -1524 2022
rect -1474 2102 -1428 2114
rect -1474 2022 -1468 2102
rect -1434 2022 -1428 2102
rect -1474 2010 -1428 2022
rect -1378 2102 -1332 2114
rect -1378 2022 -1372 2102
rect -1338 2022 -1332 2102
rect -1378 2010 -1332 2022
rect -1282 2102 -1236 2114
rect -1282 2022 -1276 2102
rect -1242 2022 -1236 2102
rect -1282 2010 -1236 2022
rect -1186 2102 -1140 2114
rect -1186 2022 -1180 2102
rect -1146 2022 -1140 2102
rect -1186 2010 -1140 2022
rect -1090 2102 -1044 2114
rect -1090 2022 -1084 2102
rect -1050 2022 -1044 2102
rect -1090 2010 -1044 2022
rect -994 2102 -948 2114
rect -994 2022 -988 2102
rect -954 2022 -948 2102
rect -994 2010 -948 2022
rect -1964 1978 -1898 1982
rect -2068 1760 -2022 1932
rect -1967 1926 -1957 1978
rect -1905 1926 -1895 1978
rect -1964 1922 -1898 1926
rect -1852 1870 -1818 2010
rect -1772 1978 -1706 1982
rect -1775 1926 -1765 1978
rect -1713 1926 -1703 1978
rect -1772 1922 -1706 1926
rect -1660 1870 -1626 2010
rect -1580 1979 -1514 1982
rect -1582 1927 -1572 1979
rect -1520 1927 -1510 1979
rect -1580 1922 -1514 1927
rect -1468 1870 -1434 2010
rect -1388 1979 -1322 1982
rect -1390 1927 -1380 1979
rect -1328 1927 -1318 1979
rect -1388 1922 -1322 1927
rect -1276 1870 -1242 2010
rect -1196 1979 -1130 1982
rect -1198 1927 -1188 1979
rect -1136 1927 -1126 1979
rect -1196 1922 -1130 1927
rect -1084 1870 -1050 2010
rect -1004 1979 -938 1982
rect -1007 1927 -997 1979
rect -945 1927 -935 1979
rect -1004 1922 -938 1927
rect -804 1870 -770 2247
rect -444 2227 -434 2247
rect -370 2227 -360 2291
rect 3308 2223 3371 4085
rect 4874 3642 4938 4326
rect 6932 4196 6938 4582
rect 6972 4196 6978 4582
rect 7033 4534 7043 4586
rect 7095 4534 7105 4586
rect 7148 4494 7182 4644
rect 7225 4534 7235 4586
rect 7287 4534 7297 4586
rect 7340 4494 7374 4644
rect 7417 4534 7427 4586
rect 7479 4534 7489 4586
rect 7532 4494 7566 4644
rect 7609 4534 7619 4586
rect 7671 4534 7681 4586
rect 7724 4494 7758 4644
rect 7800 4534 7810 4586
rect 7862 4534 7872 4586
rect 7916 4494 7950 4644
rect 7993 4534 8003 4586
rect 8055 4534 8065 4586
rect 7046 4482 7092 4494
rect 7046 4234 7052 4482
rect 7086 4234 7092 4482
rect 7046 4222 7092 4234
rect 7142 4482 7188 4494
rect 7142 4234 7148 4482
rect 7182 4234 7188 4482
rect 7142 4222 7188 4234
rect 7238 4482 7284 4494
rect 7238 4234 7244 4482
rect 7278 4234 7284 4482
rect 7238 4222 7284 4234
rect 7334 4482 7380 4494
rect 7334 4234 7340 4482
rect 7374 4234 7380 4482
rect 7334 4222 7380 4234
rect 7430 4482 7476 4494
rect 7430 4234 7436 4482
rect 7470 4234 7476 4482
rect 7430 4222 7476 4234
rect 7526 4482 7572 4494
rect 7526 4234 7532 4482
rect 7566 4234 7572 4482
rect 7526 4222 7572 4234
rect 7622 4482 7668 4494
rect 7622 4234 7628 4482
rect 7662 4234 7668 4482
rect 7622 4222 7668 4234
rect 7718 4482 7764 4494
rect 7718 4234 7724 4482
rect 7758 4234 7764 4482
rect 7718 4222 7764 4234
rect 7814 4482 7860 4494
rect 7814 4234 7820 4482
rect 7854 4234 7860 4482
rect 7814 4222 7860 4234
rect 7910 4482 7956 4494
rect 7910 4234 7916 4482
rect 7950 4234 7956 4482
rect 7910 4222 7956 4234
rect 8006 4482 8052 4494
rect 8006 4234 8012 4482
rect 8046 4234 8052 4482
rect 8006 4222 8052 4234
rect 6932 4184 6978 4196
rect 6749 4031 6759 4095
rect 6823 4081 6833 4095
rect 7052 4081 7086 4222
rect 7244 4081 7278 4222
rect 7436 4081 7470 4222
rect 7628 4081 7662 4222
rect 7820 4081 7854 4222
rect 8012 4081 8046 4222
rect 6823 4047 8046 4081
rect 6823 4031 6833 4047
rect 6932 3932 6978 3944
rect 6932 3732 6938 3932
rect 6972 3732 6978 3932
rect 7052 3914 7086 4047
rect 7244 3914 7278 4047
rect 7436 3914 7470 4047
rect 7628 3914 7662 4047
rect 7820 3914 7854 4047
rect 8012 3914 8046 4047
rect 8196 4081 8230 4644
rect 8270 4534 8280 4586
rect 8332 4534 8359 4586
rect 8724 4081 8799 5847
rect 8196 4047 8799 4081
rect 7046 3902 7092 3914
rect 7046 3822 7052 3902
rect 7086 3822 7092 3902
rect 7046 3810 7092 3822
rect 7142 3902 7188 3914
rect 7142 3822 7148 3902
rect 7182 3822 7188 3902
rect 7142 3810 7188 3822
rect 7238 3902 7284 3914
rect 7238 3822 7244 3902
rect 7278 3822 7284 3902
rect 7238 3810 7284 3822
rect 7334 3902 7380 3914
rect 7334 3822 7340 3902
rect 7374 3822 7380 3902
rect 7334 3810 7380 3822
rect 7430 3902 7476 3914
rect 7430 3822 7436 3902
rect 7470 3822 7476 3902
rect 7430 3810 7476 3822
rect 7526 3902 7572 3914
rect 7526 3822 7532 3902
rect 7566 3822 7572 3902
rect 7526 3810 7572 3822
rect 7622 3902 7668 3914
rect 7622 3822 7628 3902
rect 7662 3822 7668 3902
rect 7622 3810 7668 3822
rect 7718 3902 7764 3914
rect 7718 3822 7724 3902
rect 7758 3822 7764 3902
rect 7718 3810 7764 3822
rect 7814 3902 7860 3914
rect 7814 3822 7820 3902
rect 7854 3822 7860 3902
rect 7814 3810 7860 3822
rect 7910 3902 7956 3914
rect 7910 3822 7916 3902
rect 7950 3822 7956 3902
rect 7910 3810 7956 3822
rect 8006 3902 8052 3914
rect 8006 3822 8012 3902
rect 8046 3822 8052 3902
rect 8006 3810 8052 3822
rect 7036 3778 7102 3782
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 6932 3560 6978 3732
rect 7033 3726 7043 3778
rect 7095 3726 7105 3778
rect 7036 3722 7102 3726
rect 7148 3670 7182 3810
rect 7228 3778 7294 3782
rect 7225 3726 7235 3778
rect 7287 3726 7297 3778
rect 7228 3722 7294 3726
rect 7340 3670 7374 3810
rect 7420 3779 7486 3782
rect 7418 3727 7428 3779
rect 7480 3727 7490 3779
rect 7420 3722 7486 3727
rect 7532 3670 7566 3810
rect 7612 3779 7678 3782
rect 7610 3727 7620 3779
rect 7672 3727 7682 3779
rect 7612 3722 7678 3727
rect 7724 3670 7758 3810
rect 7804 3779 7870 3782
rect 7802 3727 7812 3779
rect 7864 3727 7874 3779
rect 7804 3722 7870 3727
rect 7916 3670 7950 3810
rect 7996 3779 8062 3782
rect 7993 3727 8003 3779
rect 8055 3727 8065 3779
rect 7996 3722 8062 3727
rect 8196 3670 8230 4047
rect 8270 3727 8280 3779
rect 8332 3727 8359 3779
rect 7148 3636 8230 3670
rect 6932 2782 6978 2960
rect 7148 2844 8230 2878
rect 6932 2396 6938 2782
rect 6972 2396 6978 2782
rect 7033 2734 7043 2786
rect 7095 2734 7105 2786
rect 7148 2694 7182 2844
rect 7225 2734 7235 2786
rect 7287 2734 7297 2786
rect 7340 2694 7374 2844
rect 7417 2734 7427 2786
rect 7479 2734 7489 2786
rect 7532 2694 7566 2844
rect 7609 2734 7619 2786
rect 7671 2734 7681 2786
rect 7724 2694 7758 2844
rect 7800 2734 7810 2786
rect 7862 2734 7872 2786
rect 7916 2694 7950 2844
rect 7993 2734 8003 2786
rect 8055 2734 8065 2786
rect 7046 2682 7092 2694
rect 7046 2434 7052 2682
rect 7086 2434 7092 2682
rect 7046 2422 7092 2434
rect 7142 2682 7188 2694
rect 7142 2434 7148 2682
rect 7182 2434 7188 2682
rect 7142 2422 7188 2434
rect 7238 2682 7284 2694
rect 7238 2434 7244 2682
rect 7278 2434 7284 2682
rect 7238 2422 7284 2434
rect 7334 2682 7380 2694
rect 7334 2434 7340 2682
rect 7374 2434 7380 2682
rect 7334 2422 7380 2434
rect 7430 2682 7476 2694
rect 7430 2434 7436 2682
rect 7470 2434 7476 2682
rect 7430 2422 7476 2434
rect 7526 2682 7572 2694
rect 7526 2434 7532 2682
rect 7566 2434 7572 2682
rect 7526 2422 7572 2434
rect 7622 2682 7668 2694
rect 7622 2434 7628 2682
rect 7662 2434 7668 2682
rect 7622 2422 7668 2434
rect 7718 2682 7764 2694
rect 7718 2434 7724 2682
rect 7758 2434 7764 2682
rect 7718 2422 7764 2434
rect 7814 2682 7860 2694
rect 7814 2434 7820 2682
rect 7854 2434 7860 2682
rect 7814 2422 7860 2434
rect 7910 2682 7956 2694
rect 7910 2434 7916 2682
rect 7950 2434 7956 2682
rect 7910 2422 7956 2434
rect 8006 2682 8052 2694
rect 8006 2434 8012 2682
rect 8046 2434 8052 2682
rect 8006 2422 8052 2434
rect 6932 2384 6978 2396
rect 6754 2233 6764 2297
rect 6828 2281 6838 2297
rect 7052 2281 7086 2422
rect 7244 2281 7278 2422
rect 7436 2281 7470 2422
rect 7628 2281 7662 2422
rect 7820 2281 7854 2422
rect 8012 2281 8046 2422
rect 6828 2247 8046 2281
rect 6828 2233 6838 2247
rect 3298 2159 3308 2223
rect 3372 2159 3382 2223
rect 6932 2132 6978 2144
rect -730 1927 -720 1979
rect -668 1927 -641 1979
rect 6932 1932 6938 2132
rect 6972 1932 6978 2132
rect 7052 2114 7086 2247
rect 7244 2114 7278 2247
rect 7436 2114 7470 2247
rect 7628 2114 7662 2247
rect 7820 2114 7854 2247
rect 8012 2114 8046 2247
rect 8196 2281 8230 2844
rect 8270 2734 8280 2786
rect 8332 2734 8359 2786
rect 8724 2281 8799 4047
rect 8196 2247 8799 2281
rect 7046 2102 7092 2114
rect 7046 2022 7052 2102
rect 7086 2022 7092 2102
rect 7046 2010 7092 2022
rect 7142 2102 7188 2114
rect 7142 2022 7148 2102
rect 7182 2022 7188 2102
rect 7142 2010 7188 2022
rect 7238 2102 7284 2114
rect 7238 2022 7244 2102
rect 7278 2022 7284 2102
rect 7238 2010 7284 2022
rect 7334 2102 7380 2114
rect 7334 2022 7340 2102
rect 7374 2022 7380 2102
rect 7334 2010 7380 2022
rect 7430 2102 7476 2114
rect 7430 2022 7436 2102
rect 7470 2022 7476 2102
rect 7430 2010 7476 2022
rect 7526 2102 7572 2114
rect 7526 2022 7532 2102
rect 7566 2022 7572 2102
rect 7526 2010 7572 2022
rect 7622 2102 7668 2114
rect 7622 2022 7628 2102
rect 7662 2022 7668 2102
rect 7622 2010 7668 2022
rect 7718 2102 7764 2114
rect 7718 2022 7724 2102
rect 7758 2022 7764 2102
rect 7718 2010 7764 2022
rect 7814 2102 7860 2114
rect 7814 2022 7820 2102
rect 7854 2022 7860 2102
rect 7814 2010 7860 2022
rect 7910 2102 7956 2114
rect 7910 2022 7916 2102
rect 7950 2022 7956 2102
rect 7910 2010 7956 2022
rect 8006 2102 8052 2114
rect 8006 2022 8012 2102
rect 8046 2022 8052 2102
rect 8006 2010 8052 2022
rect 7036 1978 7102 1982
rect -1852 1836 -770 1870
rect 6932 1760 6978 1932
rect 7033 1926 7043 1978
rect 7095 1926 7105 1978
rect 7036 1922 7102 1926
rect 7148 1870 7182 2010
rect 7228 1978 7294 1982
rect 7225 1926 7235 1978
rect 7287 1926 7297 1978
rect 7228 1922 7294 1926
rect 7340 1870 7374 2010
rect 7420 1979 7486 1982
rect 7418 1927 7428 1979
rect 7480 1927 7490 1979
rect 7420 1922 7486 1927
rect 7532 1870 7566 2010
rect 7612 1979 7678 1982
rect 7610 1927 7620 1979
rect 7672 1927 7682 1979
rect 7612 1922 7678 1927
rect 7724 1870 7758 2010
rect 7804 1979 7870 1982
rect 7802 1927 7812 1979
rect 7864 1927 7874 1979
rect 7804 1922 7870 1927
rect 7916 1870 7950 2010
rect 7996 1979 8062 1982
rect 7993 1927 8003 1979
rect 8055 1927 8065 1979
rect 7996 1922 8062 1927
rect 8196 1870 8230 2247
rect 8270 1927 8280 1979
rect 8332 1927 8359 1979
rect 7148 1836 8230 1870
rect -364 1576 2330 1640
rect 2394 1576 2404 1640
rect -2068 982 -2022 1160
rect -1852 1044 -770 1078
rect -2068 596 -2062 982
rect -2028 596 -2022 982
rect -1967 934 -1957 986
rect -1905 934 -1895 986
rect -1852 894 -1818 1044
rect -1775 934 -1765 986
rect -1713 934 -1703 986
rect -1660 894 -1626 1044
rect -1583 934 -1573 986
rect -1521 934 -1511 986
rect -1468 894 -1434 1044
rect -1391 934 -1381 986
rect -1329 934 -1319 986
rect -1276 894 -1242 1044
rect -1200 934 -1190 986
rect -1138 934 -1128 986
rect -1084 894 -1050 1044
rect -1007 934 -997 986
rect -945 934 -935 986
rect -1954 882 -1908 894
rect -1954 634 -1948 882
rect -1914 634 -1908 882
rect -1954 622 -1908 634
rect -1858 882 -1812 894
rect -1858 634 -1852 882
rect -1818 634 -1812 882
rect -1858 622 -1812 634
rect -1762 882 -1716 894
rect -1762 634 -1756 882
rect -1722 634 -1716 882
rect -1762 622 -1716 634
rect -1666 882 -1620 894
rect -1666 634 -1660 882
rect -1626 634 -1620 882
rect -1666 622 -1620 634
rect -1570 882 -1524 894
rect -1570 634 -1564 882
rect -1530 634 -1524 882
rect -1570 622 -1524 634
rect -1474 882 -1428 894
rect -1474 634 -1468 882
rect -1434 634 -1428 882
rect -1474 622 -1428 634
rect -1378 882 -1332 894
rect -1378 634 -1372 882
rect -1338 634 -1332 882
rect -1378 622 -1332 634
rect -1282 882 -1236 894
rect -1282 634 -1276 882
rect -1242 634 -1236 882
rect -1282 622 -1236 634
rect -1186 882 -1140 894
rect -1186 634 -1180 882
rect -1146 634 -1140 882
rect -1186 622 -1140 634
rect -1090 882 -1044 894
rect -1090 634 -1084 882
rect -1050 634 -1044 882
rect -1090 622 -1044 634
rect -994 882 -948 894
rect -994 634 -988 882
rect -954 634 -948 882
rect -994 622 -948 634
rect -2068 584 -2022 596
rect -1948 481 -1914 622
rect -1756 481 -1722 622
rect -1564 481 -1530 622
rect -1372 481 -1338 622
rect -1180 481 -1146 622
rect -988 497 -954 622
rect -1030 481 -1020 497
rect -2886 447 -1020 481
rect -2068 332 -2022 344
rect -2068 132 -2062 332
rect -2028 132 -2022 332
rect -1948 314 -1914 447
rect -1756 314 -1722 447
rect -1564 314 -1530 447
rect -1372 314 -1338 447
rect -1180 314 -1146 447
rect -1030 433 -1020 447
rect -956 433 -946 497
rect -804 481 -770 1044
rect -730 934 -720 986
rect -668 934 -641 986
rect -364 481 -300 1576
rect 3592 1462 3602 1526
rect 3666 1462 6152 1526
rect 6216 1462 6226 1526
rect 160 1277 170 1341
rect 234 1277 4326 1341
rect 4390 1277 4400 1341
rect 6932 982 6978 1160
rect 7148 1044 8230 1078
rect 6932 596 6938 982
rect 6972 596 6978 982
rect 7033 934 7043 986
rect 7095 934 7105 986
rect 7148 894 7182 1044
rect 7225 934 7235 986
rect 7287 934 7297 986
rect 7340 894 7374 1044
rect 7417 934 7427 986
rect 7479 934 7489 986
rect 7532 894 7566 1044
rect 7609 934 7619 986
rect 7671 934 7681 986
rect 7724 894 7758 1044
rect 7800 934 7810 986
rect 7862 934 7872 986
rect 7916 894 7950 1044
rect 7993 934 8003 986
rect 8055 934 8065 986
rect 7046 882 7092 894
rect 7046 634 7052 882
rect 7086 634 7092 882
rect 7046 622 7092 634
rect 7142 882 7188 894
rect 7142 634 7148 882
rect 7182 634 7188 882
rect 7142 622 7188 634
rect 7238 882 7284 894
rect 7238 634 7244 882
rect 7278 634 7284 882
rect 7238 622 7284 634
rect 7334 882 7380 894
rect 7334 634 7340 882
rect 7374 634 7380 882
rect 7334 622 7380 634
rect 7430 882 7476 894
rect 7430 634 7436 882
rect 7470 634 7476 882
rect 7430 622 7476 634
rect 7526 882 7572 894
rect 7526 634 7532 882
rect 7566 634 7572 882
rect 7526 622 7572 634
rect 7622 882 7668 894
rect 7622 634 7628 882
rect 7662 634 7668 882
rect 7622 622 7668 634
rect 7718 882 7764 894
rect 7718 634 7724 882
rect 7758 634 7764 882
rect 7718 622 7764 634
rect 7814 882 7860 894
rect 7814 634 7820 882
rect 7854 634 7860 882
rect 7814 622 7860 634
rect 7910 882 7956 894
rect 7910 634 7916 882
rect 7950 634 7956 882
rect 7910 622 7956 634
rect 8006 882 8052 894
rect 8006 634 8012 882
rect 8046 634 8052 882
rect 8006 622 8052 634
rect 6932 584 6978 596
rect -804 447 -300 481
rect -988 314 -954 433
rect -1954 302 -1908 314
rect -1954 222 -1948 302
rect -1914 222 -1908 302
rect -1954 210 -1908 222
rect -1858 302 -1812 314
rect -1858 222 -1852 302
rect -1818 222 -1812 302
rect -1858 210 -1812 222
rect -1762 302 -1716 314
rect -1762 222 -1756 302
rect -1722 222 -1716 302
rect -1762 210 -1716 222
rect -1666 302 -1620 314
rect -1666 222 -1660 302
rect -1626 222 -1620 302
rect -1666 210 -1620 222
rect -1570 302 -1524 314
rect -1570 222 -1564 302
rect -1530 222 -1524 302
rect -1570 210 -1524 222
rect -1474 302 -1428 314
rect -1474 222 -1468 302
rect -1434 222 -1428 302
rect -1474 210 -1428 222
rect -1378 302 -1332 314
rect -1378 222 -1372 302
rect -1338 222 -1332 302
rect -1378 210 -1332 222
rect -1282 302 -1236 314
rect -1282 222 -1276 302
rect -1242 222 -1236 302
rect -1282 210 -1236 222
rect -1186 302 -1140 314
rect -1186 222 -1180 302
rect -1146 222 -1140 302
rect -1186 210 -1140 222
rect -1090 302 -1044 314
rect -1090 222 -1084 302
rect -1050 222 -1044 302
rect -1090 210 -1044 222
rect -994 302 -948 314
rect -994 222 -988 302
rect -954 222 -948 302
rect -994 210 -948 222
rect -1964 178 -1898 182
rect -2068 -40 -2022 132
rect -1967 126 -1957 178
rect -1905 126 -1895 178
rect -1964 122 -1898 126
rect -1852 70 -1818 210
rect -1772 178 -1706 182
rect -1775 126 -1765 178
rect -1713 126 -1703 178
rect -1772 122 -1706 126
rect -1660 70 -1626 210
rect -1580 179 -1514 182
rect -1582 127 -1572 179
rect -1520 127 -1510 179
rect -1580 122 -1514 127
rect -1468 70 -1434 210
rect -1388 179 -1322 182
rect -1390 127 -1380 179
rect -1328 127 -1318 179
rect -1388 122 -1322 127
rect -1276 70 -1242 210
rect -1196 179 -1130 182
rect -1198 127 -1188 179
rect -1136 127 -1126 179
rect -1196 122 -1130 127
rect -1084 70 -1050 210
rect -1004 179 -938 182
rect -1007 127 -997 179
rect -945 127 -935 179
rect -1004 122 -938 127
rect -804 70 -770 447
rect -364 446 -300 447
rect 6690 429 6700 493
rect 6764 481 6774 493
rect 7052 481 7086 622
rect 7244 481 7278 622
rect 7436 481 7470 622
rect 7628 481 7662 622
rect 7820 481 7854 622
rect 8012 481 8046 622
rect 6764 447 8046 481
rect 6764 429 6774 447
rect 6932 332 6978 344
rect -730 127 -720 179
rect -668 127 -641 179
rect 6932 132 6938 332
rect 6972 132 6978 332
rect 7052 314 7086 447
rect 7244 314 7278 447
rect 7436 314 7470 447
rect 7628 314 7662 447
rect 7820 314 7854 447
rect 8012 314 8046 447
rect 8196 481 8230 1044
rect 8270 934 8280 986
rect 8332 934 8359 986
rect 8724 481 8799 2247
rect 8196 447 8799 481
rect 7046 302 7092 314
rect 7046 222 7052 302
rect 7086 222 7092 302
rect 7046 210 7092 222
rect 7142 302 7188 314
rect 7142 222 7148 302
rect 7182 222 7188 302
rect 7142 210 7188 222
rect 7238 302 7284 314
rect 7238 222 7244 302
rect 7278 222 7284 302
rect 7238 210 7284 222
rect 7334 302 7380 314
rect 7334 222 7340 302
rect 7374 222 7380 302
rect 7334 210 7380 222
rect 7430 302 7476 314
rect 7430 222 7436 302
rect 7470 222 7476 302
rect 7430 210 7476 222
rect 7526 302 7572 314
rect 7526 222 7532 302
rect 7566 222 7572 302
rect 7526 210 7572 222
rect 7622 302 7668 314
rect 7622 222 7628 302
rect 7662 222 7668 302
rect 7622 210 7668 222
rect 7718 302 7764 314
rect 7718 222 7724 302
rect 7758 222 7764 302
rect 7718 210 7764 222
rect 7814 302 7860 314
rect 7814 222 7820 302
rect 7854 222 7860 302
rect 7814 210 7860 222
rect 7910 302 7956 314
rect 7910 222 7916 302
rect 7950 222 7956 302
rect 7910 210 7956 222
rect 8006 302 8052 314
rect 8006 222 8012 302
rect 8046 222 8052 302
rect 8006 210 8052 222
rect 7036 178 7102 182
rect -1852 36 -770 70
rect 6932 -40 6978 132
rect 7033 126 7043 178
rect 7095 126 7105 178
rect 7036 122 7102 126
rect 7148 70 7182 210
rect 7228 178 7294 182
rect 7225 126 7235 178
rect 7287 126 7297 178
rect 7228 122 7294 126
rect 7340 70 7374 210
rect 7420 179 7486 182
rect 7418 127 7428 179
rect 7480 127 7490 179
rect 7420 122 7486 127
rect 7532 70 7566 210
rect 7612 179 7678 182
rect 7610 127 7620 179
rect 7672 127 7682 179
rect 7612 122 7678 127
rect 7724 70 7758 210
rect 7804 179 7870 182
rect 7802 127 7812 179
rect 7864 127 7874 179
rect 7804 122 7870 127
rect 7916 70 7950 210
rect 7996 179 8062 182
rect 7993 127 8003 179
rect 8055 127 8065 179
rect 7996 122 8062 127
rect 8196 70 8230 447
rect 8270 127 8280 179
rect 8332 127 8359 179
rect 7148 36 8230 70
rect -2068 -818 -2022 -640
rect -1852 -756 -770 -722
rect -2068 -1204 -2062 -818
rect -2028 -1204 -2022 -818
rect -1967 -866 -1957 -814
rect -1905 -866 -1895 -814
rect -1852 -906 -1818 -756
rect -1775 -866 -1765 -814
rect -1713 -866 -1703 -814
rect -1660 -906 -1626 -756
rect -1583 -866 -1573 -814
rect -1521 -866 -1511 -814
rect -1468 -906 -1434 -756
rect -1391 -866 -1381 -814
rect -1329 -866 -1319 -814
rect -1276 -906 -1242 -756
rect -1200 -866 -1190 -814
rect -1138 -866 -1128 -814
rect -1084 -906 -1050 -756
rect -1007 -866 -997 -814
rect -945 -866 -935 -814
rect -1954 -918 -1908 -906
rect -1954 -1166 -1948 -918
rect -1914 -1166 -1908 -918
rect -1954 -1178 -1908 -1166
rect -1858 -918 -1812 -906
rect -1858 -1166 -1852 -918
rect -1818 -1166 -1812 -918
rect -1858 -1178 -1812 -1166
rect -1762 -918 -1716 -906
rect -1762 -1166 -1756 -918
rect -1722 -1166 -1716 -918
rect -1762 -1178 -1716 -1166
rect -1666 -918 -1620 -906
rect -1666 -1166 -1660 -918
rect -1626 -1166 -1620 -918
rect -1666 -1178 -1620 -1166
rect -1570 -918 -1524 -906
rect -1570 -1166 -1564 -918
rect -1530 -1166 -1524 -918
rect -1570 -1178 -1524 -1166
rect -1474 -918 -1428 -906
rect -1474 -1166 -1468 -918
rect -1434 -1166 -1428 -918
rect -1474 -1178 -1428 -1166
rect -1378 -918 -1332 -906
rect -1378 -1166 -1372 -918
rect -1338 -1166 -1332 -918
rect -1378 -1178 -1332 -1166
rect -1282 -918 -1236 -906
rect -1282 -1166 -1276 -918
rect -1242 -1166 -1236 -918
rect -1282 -1178 -1236 -1166
rect -1186 -918 -1140 -906
rect -1186 -1166 -1180 -918
rect -1146 -1166 -1140 -918
rect -1186 -1178 -1140 -1166
rect -1090 -918 -1044 -906
rect -1090 -1166 -1084 -918
rect -1050 -1166 -1044 -918
rect -1090 -1178 -1044 -1166
rect -994 -918 -948 -906
rect -994 -1166 -988 -918
rect -954 -1166 -948 -918
rect -994 -1178 -948 -1166
rect -2068 -1216 -2022 -1204
rect -1948 -1319 -1914 -1178
rect -1756 -1319 -1722 -1178
rect -1564 -1319 -1530 -1178
rect -1372 -1319 -1338 -1178
rect -1180 -1319 -1146 -1178
rect -988 -1304 -954 -1178
rect -1029 -1319 -1019 -1304
rect -3494 -1353 -1019 -1319
rect -2068 -1468 -2022 -1456
rect -2068 -1668 -2062 -1468
rect -2028 -1668 -2022 -1468
rect -1948 -1486 -1914 -1353
rect -1756 -1486 -1722 -1353
rect -1564 -1486 -1530 -1353
rect -1372 -1486 -1338 -1353
rect -1180 -1486 -1146 -1353
rect -1029 -1368 -1019 -1353
rect -955 -1368 -945 -1304
rect -804 -1319 -770 -756
rect -730 -866 -720 -814
rect -668 -866 -641 -814
rect 6932 -818 6978 -640
rect 7148 -756 8230 -722
rect 6932 -1204 6938 -818
rect 6972 -1204 6978 -818
rect 7033 -866 7043 -814
rect 7095 -866 7105 -814
rect 7148 -906 7182 -756
rect 7225 -866 7235 -814
rect 7287 -866 7297 -814
rect 7340 -906 7374 -756
rect 7417 -866 7427 -814
rect 7479 -866 7489 -814
rect 7532 -906 7566 -756
rect 7609 -866 7619 -814
rect 7671 -866 7681 -814
rect 7724 -906 7758 -756
rect 7800 -866 7810 -814
rect 7862 -866 7872 -814
rect 7916 -906 7950 -756
rect 7993 -866 8003 -814
rect 8055 -866 8065 -814
rect 7046 -918 7092 -906
rect 7046 -1166 7052 -918
rect 7086 -1166 7092 -918
rect 7046 -1178 7092 -1166
rect 7142 -918 7188 -906
rect 7142 -1166 7148 -918
rect 7182 -1166 7188 -918
rect 7142 -1178 7188 -1166
rect 7238 -918 7284 -906
rect 7238 -1166 7244 -918
rect 7278 -1166 7284 -918
rect 7238 -1178 7284 -1166
rect 7334 -918 7380 -906
rect 7334 -1166 7340 -918
rect 7374 -1166 7380 -918
rect 7334 -1178 7380 -1166
rect 7430 -918 7476 -906
rect 7430 -1166 7436 -918
rect 7470 -1166 7476 -918
rect 7430 -1178 7476 -1166
rect 7526 -918 7572 -906
rect 7526 -1166 7532 -918
rect 7566 -1166 7572 -918
rect 7526 -1178 7572 -1166
rect 7622 -918 7668 -906
rect 7622 -1166 7628 -918
rect 7662 -1166 7668 -918
rect 7622 -1178 7668 -1166
rect 7718 -918 7764 -906
rect 7718 -1166 7724 -918
rect 7758 -1166 7764 -918
rect 7718 -1178 7764 -1166
rect 7814 -918 7860 -906
rect 7814 -1166 7820 -918
rect 7854 -1166 7860 -918
rect 7814 -1178 7860 -1166
rect 7910 -918 7956 -906
rect 7910 -1166 7916 -918
rect 7950 -1166 7956 -918
rect 7910 -1178 7956 -1166
rect 8006 -918 8052 -906
rect 8006 -1166 8012 -918
rect 8046 -1166 8052 -918
rect 8006 -1178 8052 -1166
rect 6932 -1216 6978 -1204
rect -512 -1319 -502 -1301
rect -804 -1353 -502 -1319
rect -988 -1486 -954 -1368
rect -1954 -1498 -1908 -1486
rect -1954 -1578 -1948 -1498
rect -1914 -1578 -1908 -1498
rect -1954 -1590 -1908 -1578
rect -1858 -1498 -1812 -1486
rect -1858 -1578 -1852 -1498
rect -1818 -1578 -1812 -1498
rect -1858 -1590 -1812 -1578
rect -1762 -1498 -1716 -1486
rect -1762 -1578 -1756 -1498
rect -1722 -1578 -1716 -1498
rect -1762 -1590 -1716 -1578
rect -1666 -1498 -1620 -1486
rect -1666 -1578 -1660 -1498
rect -1626 -1578 -1620 -1498
rect -1666 -1590 -1620 -1578
rect -1570 -1498 -1524 -1486
rect -1570 -1578 -1564 -1498
rect -1530 -1578 -1524 -1498
rect -1570 -1590 -1524 -1578
rect -1474 -1498 -1428 -1486
rect -1474 -1578 -1468 -1498
rect -1434 -1578 -1428 -1498
rect -1474 -1590 -1428 -1578
rect -1378 -1498 -1332 -1486
rect -1378 -1578 -1372 -1498
rect -1338 -1578 -1332 -1498
rect -1378 -1590 -1332 -1578
rect -1282 -1498 -1236 -1486
rect -1282 -1578 -1276 -1498
rect -1242 -1578 -1236 -1498
rect -1282 -1590 -1236 -1578
rect -1186 -1498 -1140 -1486
rect -1186 -1578 -1180 -1498
rect -1146 -1578 -1140 -1498
rect -1186 -1590 -1140 -1578
rect -1090 -1498 -1044 -1486
rect -1090 -1578 -1084 -1498
rect -1050 -1578 -1044 -1498
rect -1090 -1590 -1044 -1578
rect -994 -1498 -948 -1486
rect -994 -1578 -988 -1498
rect -954 -1578 -948 -1498
rect -994 -1590 -948 -1578
rect -1964 -1622 -1898 -1618
rect -2068 -1840 -2022 -1668
rect -1967 -1674 -1957 -1622
rect -1905 -1674 -1895 -1622
rect -1964 -1678 -1898 -1674
rect -1852 -1730 -1818 -1590
rect -1772 -1622 -1706 -1618
rect -1775 -1674 -1765 -1622
rect -1713 -1674 -1703 -1622
rect -1772 -1678 -1706 -1674
rect -1660 -1730 -1626 -1590
rect -1580 -1621 -1514 -1618
rect -1582 -1673 -1572 -1621
rect -1520 -1673 -1510 -1621
rect -1580 -1678 -1514 -1673
rect -1468 -1730 -1434 -1590
rect -1388 -1621 -1322 -1618
rect -1390 -1673 -1380 -1621
rect -1328 -1673 -1318 -1621
rect -1388 -1678 -1322 -1673
rect -1276 -1730 -1242 -1590
rect -1196 -1621 -1130 -1618
rect -1198 -1673 -1188 -1621
rect -1136 -1673 -1126 -1621
rect -1196 -1678 -1130 -1673
rect -1084 -1730 -1050 -1590
rect -1004 -1621 -938 -1618
rect -1007 -1673 -997 -1621
rect -945 -1673 -935 -1621
rect -1004 -1678 -938 -1673
rect -804 -1730 -770 -1353
rect -512 -1365 -502 -1353
rect -438 -1365 -428 -1301
rect 6708 -1363 6718 -1299
rect 6782 -1319 6792 -1299
rect 7052 -1319 7086 -1178
rect 7244 -1319 7278 -1178
rect 7436 -1319 7470 -1178
rect 7628 -1319 7662 -1178
rect 7820 -1319 7854 -1178
rect 8012 -1319 8046 -1178
rect 6782 -1353 8046 -1319
rect 6782 -1363 6792 -1353
rect 6932 -1468 6978 -1456
rect -730 -1673 -720 -1621
rect -668 -1673 -641 -1621
rect 6932 -1668 6938 -1468
rect 6972 -1668 6978 -1468
rect 7052 -1486 7086 -1353
rect 7244 -1486 7278 -1353
rect 7436 -1486 7470 -1353
rect 7628 -1486 7662 -1353
rect 7820 -1486 7854 -1353
rect 8012 -1486 8046 -1353
rect 8196 -1319 8230 -756
rect 8270 -866 8280 -814
rect 8332 -866 8359 -814
rect 9235 -1319 9310 7647
rect 8196 -1353 9310 -1319
rect 7046 -1498 7092 -1486
rect 7046 -1578 7052 -1498
rect 7086 -1578 7092 -1498
rect 7046 -1590 7092 -1578
rect 7142 -1498 7188 -1486
rect 7142 -1578 7148 -1498
rect 7182 -1578 7188 -1498
rect 7142 -1590 7188 -1578
rect 7238 -1498 7284 -1486
rect 7238 -1578 7244 -1498
rect 7278 -1578 7284 -1498
rect 7238 -1590 7284 -1578
rect 7334 -1498 7380 -1486
rect 7334 -1578 7340 -1498
rect 7374 -1578 7380 -1498
rect 7334 -1590 7380 -1578
rect 7430 -1498 7476 -1486
rect 7430 -1578 7436 -1498
rect 7470 -1578 7476 -1498
rect 7430 -1590 7476 -1578
rect 7526 -1498 7572 -1486
rect 7526 -1578 7532 -1498
rect 7566 -1578 7572 -1498
rect 7526 -1590 7572 -1578
rect 7622 -1498 7668 -1486
rect 7622 -1578 7628 -1498
rect 7662 -1578 7668 -1498
rect 7622 -1590 7668 -1578
rect 7718 -1498 7764 -1486
rect 7718 -1578 7724 -1498
rect 7758 -1578 7764 -1498
rect 7718 -1590 7764 -1578
rect 7814 -1498 7860 -1486
rect 7814 -1578 7820 -1498
rect 7854 -1578 7860 -1498
rect 7814 -1590 7860 -1578
rect 7910 -1498 7956 -1486
rect 7910 -1578 7916 -1498
rect 7950 -1578 7956 -1498
rect 7910 -1590 7956 -1578
rect 8006 -1498 8052 -1486
rect 8006 -1578 8012 -1498
rect 8046 -1578 8052 -1498
rect 8006 -1590 8052 -1578
rect 7036 -1622 7102 -1618
rect -1852 -1764 -770 -1730
rect 6932 -1840 6978 -1668
rect 7033 -1674 7043 -1622
rect 7095 -1674 7105 -1622
rect 7036 -1678 7102 -1674
rect 7148 -1730 7182 -1590
rect 7228 -1622 7294 -1618
rect 7225 -1674 7235 -1622
rect 7287 -1674 7297 -1622
rect 7228 -1678 7294 -1674
rect 7340 -1730 7374 -1590
rect 7420 -1621 7486 -1618
rect 7418 -1673 7428 -1621
rect 7480 -1673 7490 -1621
rect 7420 -1678 7486 -1673
rect 7532 -1730 7566 -1590
rect 7612 -1621 7678 -1618
rect 7610 -1673 7620 -1621
rect 7672 -1673 7682 -1621
rect 7612 -1678 7678 -1673
rect 7724 -1730 7758 -1590
rect 7804 -1621 7870 -1618
rect 7802 -1673 7812 -1621
rect 7864 -1673 7874 -1621
rect 7804 -1678 7870 -1673
rect 7916 -1730 7950 -1590
rect 7996 -1621 8062 -1618
rect 7993 -1673 8003 -1621
rect 8055 -1673 8065 -1621
rect 7996 -1678 8062 -1673
rect 8196 -1730 8230 -1353
rect 8270 -1673 8280 -1621
rect 8332 -1673 8359 -1621
rect 7148 -1764 8230 -1730
<< via1 >>
rect -1957 8176 -1905 8186
rect -1957 8142 -1948 8176
rect -1948 8142 -1914 8176
rect -1914 8142 -1905 8176
rect -1957 8134 -1905 8142
rect -1765 8176 -1713 8186
rect -1765 8142 -1756 8176
rect -1756 8142 -1722 8176
rect -1722 8142 -1713 8176
rect -1765 8134 -1713 8142
rect -1573 8176 -1521 8186
rect -1573 8142 -1564 8176
rect -1564 8142 -1530 8176
rect -1530 8142 -1521 8176
rect -1573 8134 -1521 8142
rect -1381 8176 -1329 8186
rect -1381 8142 -1372 8176
rect -1372 8142 -1338 8176
rect -1338 8142 -1329 8176
rect -1381 8134 -1329 8142
rect -1190 8176 -1138 8186
rect -1190 8142 -1180 8176
rect -1180 8142 -1146 8176
rect -1146 8142 -1138 8176
rect -1190 8134 -1138 8142
rect -997 8176 -945 8186
rect -997 8142 -988 8176
rect -988 8142 -954 8176
rect -954 8142 -945 8176
rect -997 8134 -945 8142
rect -1022 7631 -958 7695
rect -720 8134 -668 8186
rect 7043 8176 7095 8186
rect 7043 8142 7052 8176
rect 7052 8142 7086 8176
rect 7086 8142 7095 8176
rect 7043 8134 7095 8142
rect 7235 8176 7287 8186
rect 7235 8142 7244 8176
rect 7244 8142 7278 8176
rect 7278 8142 7287 8176
rect 7235 8134 7287 8142
rect 7427 8176 7479 8186
rect 7427 8142 7436 8176
rect 7436 8142 7470 8176
rect 7470 8142 7479 8176
rect 7427 8134 7479 8142
rect 7619 8176 7671 8186
rect 7619 8142 7628 8176
rect 7628 8142 7662 8176
rect 7662 8142 7671 8176
rect 7619 8134 7671 8142
rect 7810 8176 7862 8186
rect 7810 8142 7820 8176
rect 7820 8142 7854 8176
rect 7854 8142 7862 8176
rect 7810 8134 7862 8142
rect 8003 8176 8055 8186
rect 8003 8142 8012 8176
rect 8012 8142 8046 8176
rect 8046 8142 8055 8176
rect 8003 8134 8055 8142
rect -1957 7368 -1905 7378
rect -1957 7334 -1948 7368
rect -1948 7334 -1914 7368
rect -1914 7334 -1905 7368
rect -1957 7326 -1905 7334
rect -1765 7368 -1713 7378
rect -1765 7334 -1756 7368
rect -1756 7334 -1722 7368
rect -1722 7334 -1713 7368
rect -1765 7326 -1713 7334
rect -1572 7368 -1520 7379
rect -1572 7334 -1564 7368
rect -1564 7334 -1530 7368
rect -1530 7334 -1520 7368
rect -1572 7327 -1520 7334
rect -1380 7368 -1328 7379
rect -1380 7334 -1372 7368
rect -1372 7334 -1338 7368
rect -1338 7334 -1328 7368
rect -1380 7327 -1328 7334
rect -1188 7368 -1136 7379
rect -1188 7334 -1180 7368
rect -1180 7334 -1146 7368
rect -1146 7334 -1136 7368
rect -1188 7327 -1136 7334
rect -997 7368 -945 7379
rect -997 7334 -988 7368
rect -988 7334 -954 7368
rect -954 7334 -945 7368
rect -997 7327 -945 7334
rect 6691 7633 6755 7697
rect -720 7327 -668 7379
rect -1957 6376 -1905 6386
rect -1957 6342 -1948 6376
rect -1948 6342 -1914 6376
rect -1914 6342 -1905 6376
rect -1957 6334 -1905 6342
rect -1765 6376 -1713 6386
rect -1765 6342 -1756 6376
rect -1756 6342 -1722 6376
rect -1722 6342 -1713 6376
rect -1765 6334 -1713 6342
rect -1573 6376 -1521 6386
rect -1573 6342 -1564 6376
rect -1564 6342 -1530 6376
rect -1530 6342 -1521 6376
rect -1573 6334 -1521 6342
rect -1381 6376 -1329 6386
rect -1381 6342 -1372 6376
rect -1372 6342 -1338 6376
rect -1338 6342 -1329 6376
rect -1381 6334 -1329 6342
rect -1190 6376 -1138 6386
rect -1190 6342 -1180 6376
rect -1180 6342 -1146 6376
rect -1146 6342 -1138 6376
rect -1190 6334 -1138 6342
rect -997 6376 -945 6386
rect -997 6342 -988 6376
rect -988 6342 -954 6376
rect -954 6342 -945 6376
rect -997 6334 -945 6342
rect -1028 5831 -964 5895
rect 1628 6412 1692 6476
rect -720 6334 -668 6386
rect -1957 5568 -1905 5578
rect -1957 5534 -1948 5568
rect -1948 5534 -1914 5568
rect -1914 5534 -1905 5568
rect -1957 5526 -1905 5534
rect -1765 5568 -1713 5578
rect -1765 5534 -1756 5568
rect -1756 5534 -1722 5568
rect -1722 5534 -1713 5568
rect -1765 5526 -1713 5534
rect -1572 5568 -1520 5579
rect -1572 5534 -1564 5568
rect -1564 5534 -1530 5568
rect -1530 5534 -1520 5568
rect -1572 5527 -1520 5534
rect -1380 5568 -1328 5579
rect -1380 5534 -1372 5568
rect -1372 5534 -1338 5568
rect -1338 5534 -1328 5568
rect -1380 5527 -1328 5534
rect -1188 5568 -1136 5579
rect -1188 5534 -1180 5568
rect -1180 5534 -1146 5568
rect -1146 5534 -1136 5568
rect -1188 5527 -1136 5534
rect -997 5568 -945 5579
rect -997 5534 -988 5568
rect -988 5534 -954 5568
rect -954 5534 -945 5568
rect -997 5527 -945 5534
rect -477 5829 -413 5893
rect -720 5527 -668 5579
rect -1957 4576 -1905 4586
rect -1957 4542 -1948 4576
rect -1948 4542 -1914 4576
rect -1914 4542 -1905 4576
rect -1957 4534 -1905 4542
rect -1765 4576 -1713 4586
rect -1765 4542 -1756 4576
rect -1756 4542 -1722 4576
rect -1722 4542 -1713 4576
rect -1765 4534 -1713 4542
rect -1573 4576 -1521 4586
rect -1573 4542 -1564 4576
rect -1564 4542 -1530 4576
rect -1530 4542 -1521 4576
rect -1573 4534 -1521 4542
rect -1381 4576 -1329 4586
rect -1381 4542 -1372 4576
rect -1372 4542 -1338 4576
rect -1338 4542 -1329 4576
rect -1381 4534 -1329 4542
rect -1190 4576 -1138 4586
rect -1190 4542 -1180 4576
rect -1180 4542 -1146 4576
rect -1146 4542 -1138 4576
rect -1190 4534 -1138 4542
rect -997 4576 -945 4586
rect -997 4542 -988 4576
rect -988 4542 -954 4576
rect -954 4542 -945 4576
rect -997 4534 -945 4542
rect -1024 4031 -960 4095
rect -720 4534 -668 4586
rect -1957 3768 -1905 3778
rect -1957 3734 -1948 3768
rect -1948 3734 -1914 3768
rect -1914 3734 -1905 3768
rect -1957 3726 -1905 3734
rect -1765 3768 -1713 3778
rect -1765 3734 -1756 3768
rect -1756 3734 -1722 3768
rect -1722 3734 -1713 3768
rect -1765 3726 -1713 3734
rect -1572 3768 -1520 3779
rect -1572 3734 -1564 3768
rect -1564 3734 -1530 3768
rect -1530 3734 -1520 3768
rect -1572 3727 -1520 3734
rect -1380 3768 -1328 3779
rect -1380 3734 -1372 3768
rect -1372 3734 -1338 3768
rect -1338 3734 -1328 3768
rect -1380 3727 -1328 3734
rect -1188 3768 -1136 3779
rect -1188 3734 -1180 3768
rect -1180 3734 -1146 3768
rect -1146 3734 -1136 3768
rect -1188 3727 -1136 3734
rect -997 3768 -945 3779
rect -997 3734 -988 3768
rect -988 3734 -954 3768
rect -954 3734 -945 3768
rect -997 3727 -945 3734
rect -434 4030 -370 4094
rect 8280 8134 8332 8186
rect 7043 7368 7095 7378
rect 7043 7334 7052 7368
rect 7052 7334 7086 7368
rect 7086 7334 7095 7368
rect 7043 7326 7095 7334
rect 7235 7368 7287 7378
rect 7235 7334 7244 7368
rect 7244 7334 7278 7368
rect 7278 7334 7287 7368
rect 7235 7326 7287 7334
rect 7428 7368 7480 7379
rect 7428 7334 7436 7368
rect 7436 7334 7470 7368
rect 7470 7334 7480 7368
rect 7428 7327 7480 7334
rect 7620 7368 7672 7379
rect 7620 7334 7628 7368
rect 7628 7334 7662 7368
rect 7662 7334 7672 7368
rect 7620 7327 7672 7334
rect 7812 7368 7864 7379
rect 7812 7334 7820 7368
rect 7820 7334 7854 7368
rect 7854 7334 7864 7368
rect 7812 7327 7864 7334
rect 8003 7368 8055 7379
rect 8003 7334 8012 7368
rect 8012 7334 8046 7368
rect 8046 7334 8055 7368
rect 8003 7327 8055 7334
rect 8280 7327 8332 7379
rect 7043 6376 7095 6386
rect 7043 6342 7052 6376
rect 7052 6342 7086 6376
rect 7086 6342 7095 6376
rect 7043 6334 7095 6342
rect 7235 6376 7287 6386
rect 7235 6342 7244 6376
rect 7244 6342 7278 6376
rect 7278 6342 7287 6376
rect 7235 6334 7287 6342
rect 7427 6376 7479 6386
rect 7427 6342 7436 6376
rect 7436 6342 7470 6376
rect 7470 6342 7479 6376
rect 7427 6334 7479 6342
rect 7619 6376 7671 6386
rect 7619 6342 7628 6376
rect 7628 6342 7662 6376
rect 7662 6342 7671 6376
rect 7619 6334 7671 6342
rect 7810 6376 7862 6386
rect 7810 6342 7820 6376
rect 7820 6342 7854 6376
rect 7854 6342 7862 6376
rect 7810 6334 7862 6342
rect 8003 6376 8055 6386
rect 8003 6342 8012 6376
rect 8012 6342 8046 6376
rect 8046 6342 8055 6376
rect 8003 6334 8055 6342
rect 6704 5831 6768 5895
rect 3157 5494 3221 5558
rect 8280 6334 8332 6386
rect 7043 5568 7095 5578
rect 7043 5534 7052 5568
rect 7052 5534 7086 5568
rect 7086 5534 7095 5568
rect 7043 5526 7095 5534
rect 7235 5568 7287 5578
rect 7235 5534 7244 5568
rect 7244 5534 7278 5568
rect 7278 5534 7287 5568
rect 7235 5526 7287 5534
rect 7428 5568 7480 5579
rect 7428 5534 7436 5568
rect 7436 5534 7470 5568
rect 7470 5534 7480 5568
rect 7428 5527 7480 5534
rect 7620 5568 7672 5579
rect 7620 5534 7628 5568
rect 7628 5534 7662 5568
rect 7662 5534 7672 5568
rect 7620 5527 7672 5534
rect 7812 5568 7864 5579
rect 7812 5534 7820 5568
rect 7820 5534 7854 5568
rect 7854 5534 7864 5568
rect 7812 5527 7864 5534
rect 8003 5568 8055 5579
rect 8003 5534 8012 5568
rect 8012 5534 8046 5568
rect 8046 5534 8055 5568
rect 8003 5527 8055 5534
rect 8280 5527 8332 5579
rect 3157 5020 3221 5084
rect 3768 4864 3832 4928
rect 6166 4868 6230 4932
rect 3106 4499 3170 4563
rect 5207 4326 5271 4390
rect 3308 4148 3372 4212
rect -720 3727 -668 3779
rect 333 3419 397 3483
rect 1631 3419 1695 3483
rect 333 3090 397 3154
rect -1957 2776 -1905 2786
rect -1957 2742 -1948 2776
rect -1948 2742 -1914 2776
rect -1914 2742 -1905 2776
rect -1957 2734 -1905 2742
rect -1765 2776 -1713 2786
rect -1765 2742 -1756 2776
rect -1756 2742 -1722 2776
rect -1722 2742 -1713 2776
rect -1765 2734 -1713 2742
rect -1573 2776 -1521 2786
rect -1573 2742 -1564 2776
rect -1564 2742 -1530 2776
rect -1530 2742 -1521 2776
rect -1573 2734 -1521 2742
rect -1381 2776 -1329 2786
rect -1381 2742 -1372 2776
rect -1372 2742 -1338 2776
rect -1338 2742 -1329 2776
rect -1381 2734 -1329 2742
rect -1190 2776 -1138 2786
rect -1190 2742 -1180 2776
rect -1180 2742 -1146 2776
rect -1146 2742 -1138 2776
rect -1190 2734 -1138 2742
rect -997 2776 -945 2786
rect -997 2742 -988 2776
rect -988 2742 -954 2776
rect -954 2742 -945 2776
rect -997 2734 -945 2742
rect -1027 2231 -963 2295
rect -720 2734 -668 2786
rect -1957 1968 -1905 1978
rect -1957 1934 -1948 1968
rect -1948 1934 -1914 1968
rect -1914 1934 -1905 1968
rect -1957 1926 -1905 1934
rect -1765 1968 -1713 1978
rect -1765 1934 -1756 1968
rect -1756 1934 -1722 1968
rect -1722 1934 -1713 1968
rect -1765 1926 -1713 1934
rect -1572 1968 -1520 1979
rect -1572 1934 -1564 1968
rect -1564 1934 -1530 1968
rect -1530 1934 -1520 1968
rect -1572 1927 -1520 1934
rect -1380 1968 -1328 1979
rect -1380 1934 -1372 1968
rect -1372 1934 -1338 1968
rect -1338 1934 -1328 1968
rect -1380 1927 -1328 1934
rect -1188 1968 -1136 1979
rect -1188 1934 -1180 1968
rect -1180 1934 -1146 1968
rect -1146 1934 -1136 1968
rect -1188 1927 -1136 1934
rect -997 1968 -945 1979
rect -997 1934 -988 1968
rect -988 1934 -954 1968
rect -954 1934 -945 1968
rect -997 1927 -945 1934
rect -434 2227 -370 2291
rect 7043 4576 7095 4586
rect 7043 4542 7052 4576
rect 7052 4542 7086 4576
rect 7086 4542 7095 4576
rect 7043 4534 7095 4542
rect 7235 4576 7287 4586
rect 7235 4542 7244 4576
rect 7244 4542 7278 4576
rect 7278 4542 7287 4576
rect 7235 4534 7287 4542
rect 7427 4576 7479 4586
rect 7427 4542 7436 4576
rect 7436 4542 7470 4576
rect 7470 4542 7479 4576
rect 7427 4534 7479 4542
rect 7619 4576 7671 4586
rect 7619 4542 7628 4576
rect 7628 4542 7662 4576
rect 7662 4542 7671 4576
rect 7619 4534 7671 4542
rect 7810 4576 7862 4586
rect 7810 4542 7820 4576
rect 7820 4542 7854 4576
rect 7854 4542 7862 4576
rect 7810 4534 7862 4542
rect 8003 4576 8055 4586
rect 8003 4542 8012 4576
rect 8012 4542 8046 4576
rect 8046 4542 8055 4576
rect 8003 4534 8055 4542
rect 6759 4031 6823 4095
rect 8280 4534 8332 4586
rect 4874 3578 4938 3642
rect 7043 3768 7095 3778
rect 7043 3734 7052 3768
rect 7052 3734 7086 3768
rect 7086 3734 7095 3768
rect 7043 3726 7095 3734
rect 7235 3768 7287 3778
rect 7235 3734 7244 3768
rect 7244 3734 7278 3768
rect 7278 3734 7287 3768
rect 7235 3726 7287 3734
rect 7428 3768 7480 3779
rect 7428 3734 7436 3768
rect 7436 3734 7470 3768
rect 7470 3734 7480 3768
rect 7428 3727 7480 3734
rect 7620 3768 7672 3779
rect 7620 3734 7628 3768
rect 7628 3734 7662 3768
rect 7662 3734 7672 3768
rect 7620 3727 7672 3734
rect 7812 3768 7864 3779
rect 7812 3734 7820 3768
rect 7820 3734 7854 3768
rect 7854 3734 7864 3768
rect 7812 3727 7864 3734
rect 8003 3768 8055 3779
rect 8003 3734 8012 3768
rect 8012 3734 8046 3768
rect 8046 3734 8055 3768
rect 8003 3727 8055 3734
rect 8280 3727 8332 3779
rect 7043 2776 7095 2786
rect 7043 2742 7052 2776
rect 7052 2742 7086 2776
rect 7086 2742 7095 2776
rect 7043 2734 7095 2742
rect 7235 2776 7287 2786
rect 7235 2742 7244 2776
rect 7244 2742 7278 2776
rect 7278 2742 7287 2776
rect 7235 2734 7287 2742
rect 7427 2776 7479 2786
rect 7427 2742 7436 2776
rect 7436 2742 7470 2776
rect 7470 2742 7479 2776
rect 7427 2734 7479 2742
rect 7619 2776 7671 2786
rect 7619 2742 7628 2776
rect 7628 2742 7662 2776
rect 7662 2742 7671 2776
rect 7619 2734 7671 2742
rect 7810 2776 7862 2786
rect 7810 2742 7820 2776
rect 7820 2742 7854 2776
rect 7854 2742 7862 2776
rect 7810 2734 7862 2742
rect 8003 2776 8055 2786
rect 8003 2742 8012 2776
rect 8012 2742 8046 2776
rect 8046 2742 8055 2776
rect 8003 2734 8055 2742
rect 6764 2233 6828 2297
rect 3308 2159 3372 2223
rect -720 1927 -668 1979
rect 8280 2734 8332 2786
rect 7043 1968 7095 1978
rect 7043 1934 7052 1968
rect 7052 1934 7086 1968
rect 7086 1934 7095 1968
rect 7043 1926 7095 1934
rect 7235 1968 7287 1978
rect 7235 1934 7244 1968
rect 7244 1934 7278 1968
rect 7278 1934 7287 1968
rect 7235 1926 7287 1934
rect 7428 1968 7480 1979
rect 7428 1934 7436 1968
rect 7436 1934 7470 1968
rect 7470 1934 7480 1968
rect 7428 1927 7480 1934
rect 7620 1968 7672 1979
rect 7620 1934 7628 1968
rect 7628 1934 7662 1968
rect 7662 1934 7672 1968
rect 7620 1927 7672 1934
rect 7812 1968 7864 1979
rect 7812 1934 7820 1968
rect 7820 1934 7854 1968
rect 7854 1934 7864 1968
rect 7812 1927 7864 1934
rect 8003 1968 8055 1979
rect 8003 1934 8012 1968
rect 8012 1934 8046 1968
rect 8046 1934 8055 1968
rect 8003 1927 8055 1934
rect 8280 1927 8332 1979
rect 2330 1576 2394 1640
rect -1957 976 -1905 986
rect -1957 942 -1948 976
rect -1948 942 -1914 976
rect -1914 942 -1905 976
rect -1957 934 -1905 942
rect -1765 976 -1713 986
rect -1765 942 -1756 976
rect -1756 942 -1722 976
rect -1722 942 -1713 976
rect -1765 934 -1713 942
rect -1573 976 -1521 986
rect -1573 942 -1564 976
rect -1564 942 -1530 976
rect -1530 942 -1521 976
rect -1573 934 -1521 942
rect -1381 976 -1329 986
rect -1381 942 -1372 976
rect -1372 942 -1338 976
rect -1338 942 -1329 976
rect -1381 934 -1329 942
rect -1190 976 -1138 986
rect -1190 942 -1180 976
rect -1180 942 -1146 976
rect -1146 942 -1138 976
rect -1190 934 -1138 942
rect -997 976 -945 986
rect -997 942 -988 976
rect -988 942 -954 976
rect -954 942 -945 976
rect -997 934 -945 942
rect -1020 433 -956 497
rect -720 934 -668 986
rect 3602 1462 3666 1526
rect 6152 1462 6216 1526
rect 170 1277 234 1341
rect 4326 1277 4390 1341
rect 7043 976 7095 986
rect 7043 942 7052 976
rect 7052 942 7086 976
rect 7086 942 7095 976
rect 7043 934 7095 942
rect 7235 976 7287 986
rect 7235 942 7244 976
rect 7244 942 7278 976
rect 7278 942 7287 976
rect 7235 934 7287 942
rect 7427 976 7479 986
rect 7427 942 7436 976
rect 7436 942 7470 976
rect 7470 942 7479 976
rect 7427 934 7479 942
rect 7619 976 7671 986
rect 7619 942 7628 976
rect 7628 942 7662 976
rect 7662 942 7671 976
rect 7619 934 7671 942
rect 7810 976 7862 986
rect 7810 942 7820 976
rect 7820 942 7854 976
rect 7854 942 7862 976
rect 7810 934 7862 942
rect 8003 976 8055 986
rect 8003 942 8012 976
rect 8012 942 8046 976
rect 8046 942 8055 976
rect 8003 934 8055 942
rect -1957 168 -1905 178
rect -1957 134 -1948 168
rect -1948 134 -1914 168
rect -1914 134 -1905 168
rect -1957 126 -1905 134
rect -1765 168 -1713 178
rect -1765 134 -1756 168
rect -1756 134 -1722 168
rect -1722 134 -1713 168
rect -1765 126 -1713 134
rect -1572 168 -1520 179
rect -1572 134 -1564 168
rect -1564 134 -1530 168
rect -1530 134 -1520 168
rect -1572 127 -1520 134
rect -1380 168 -1328 179
rect -1380 134 -1372 168
rect -1372 134 -1338 168
rect -1338 134 -1328 168
rect -1380 127 -1328 134
rect -1188 168 -1136 179
rect -1188 134 -1180 168
rect -1180 134 -1146 168
rect -1146 134 -1136 168
rect -1188 127 -1136 134
rect -997 168 -945 179
rect -997 134 -988 168
rect -988 134 -954 168
rect -954 134 -945 168
rect -997 127 -945 134
rect 6700 429 6764 493
rect -720 127 -668 179
rect 8280 934 8332 986
rect 7043 168 7095 178
rect 7043 134 7052 168
rect 7052 134 7086 168
rect 7086 134 7095 168
rect 7043 126 7095 134
rect 7235 168 7287 178
rect 7235 134 7244 168
rect 7244 134 7278 168
rect 7278 134 7287 168
rect 7235 126 7287 134
rect 7428 168 7480 179
rect 7428 134 7436 168
rect 7436 134 7470 168
rect 7470 134 7480 168
rect 7428 127 7480 134
rect 7620 168 7672 179
rect 7620 134 7628 168
rect 7628 134 7662 168
rect 7662 134 7672 168
rect 7620 127 7672 134
rect 7812 168 7864 179
rect 7812 134 7820 168
rect 7820 134 7854 168
rect 7854 134 7864 168
rect 7812 127 7864 134
rect 8003 168 8055 179
rect 8003 134 8012 168
rect 8012 134 8046 168
rect 8046 134 8055 168
rect 8003 127 8055 134
rect 8280 127 8332 179
rect -1957 -824 -1905 -814
rect -1957 -858 -1948 -824
rect -1948 -858 -1914 -824
rect -1914 -858 -1905 -824
rect -1957 -866 -1905 -858
rect -1765 -824 -1713 -814
rect -1765 -858 -1756 -824
rect -1756 -858 -1722 -824
rect -1722 -858 -1713 -824
rect -1765 -866 -1713 -858
rect -1573 -824 -1521 -814
rect -1573 -858 -1564 -824
rect -1564 -858 -1530 -824
rect -1530 -858 -1521 -824
rect -1573 -866 -1521 -858
rect -1381 -824 -1329 -814
rect -1381 -858 -1372 -824
rect -1372 -858 -1338 -824
rect -1338 -858 -1329 -824
rect -1381 -866 -1329 -858
rect -1190 -824 -1138 -814
rect -1190 -858 -1180 -824
rect -1180 -858 -1146 -824
rect -1146 -858 -1138 -824
rect -1190 -866 -1138 -858
rect -997 -824 -945 -814
rect -997 -858 -988 -824
rect -988 -858 -954 -824
rect -954 -858 -945 -824
rect -997 -866 -945 -858
rect -1019 -1368 -955 -1304
rect -720 -866 -668 -814
rect 7043 -824 7095 -814
rect 7043 -858 7052 -824
rect 7052 -858 7086 -824
rect 7086 -858 7095 -824
rect 7043 -866 7095 -858
rect 7235 -824 7287 -814
rect 7235 -858 7244 -824
rect 7244 -858 7278 -824
rect 7278 -858 7287 -824
rect 7235 -866 7287 -858
rect 7427 -824 7479 -814
rect 7427 -858 7436 -824
rect 7436 -858 7470 -824
rect 7470 -858 7479 -824
rect 7427 -866 7479 -858
rect 7619 -824 7671 -814
rect 7619 -858 7628 -824
rect 7628 -858 7662 -824
rect 7662 -858 7671 -824
rect 7619 -866 7671 -858
rect 7810 -824 7862 -814
rect 7810 -858 7820 -824
rect 7820 -858 7854 -824
rect 7854 -858 7862 -824
rect 7810 -866 7862 -858
rect 8003 -824 8055 -814
rect 8003 -858 8012 -824
rect 8012 -858 8046 -824
rect 8046 -858 8055 -824
rect 8003 -866 8055 -858
rect -1957 -1632 -1905 -1622
rect -1957 -1666 -1948 -1632
rect -1948 -1666 -1914 -1632
rect -1914 -1666 -1905 -1632
rect -1957 -1674 -1905 -1666
rect -1765 -1632 -1713 -1622
rect -1765 -1666 -1756 -1632
rect -1756 -1666 -1722 -1632
rect -1722 -1666 -1713 -1632
rect -1765 -1674 -1713 -1666
rect -1572 -1632 -1520 -1621
rect -1572 -1666 -1564 -1632
rect -1564 -1666 -1530 -1632
rect -1530 -1666 -1520 -1632
rect -1572 -1673 -1520 -1666
rect -1380 -1632 -1328 -1621
rect -1380 -1666 -1372 -1632
rect -1372 -1666 -1338 -1632
rect -1338 -1666 -1328 -1632
rect -1380 -1673 -1328 -1666
rect -1188 -1632 -1136 -1621
rect -1188 -1666 -1180 -1632
rect -1180 -1666 -1146 -1632
rect -1146 -1666 -1136 -1632
rect -1188 -1673 -1136 -1666
rect -997 -1632 -945 -1621
rect -997 -1666 -988 -1632
rect -988 -1666 -954 -1632
rect -954 -1666 -945 -1632
rect -997 -1673 -945 -1666
rect -502 -1365 -438 -1301
rect 6718 -1363 6782 -1299
rect -720 -1673 -668 -1621
rect 8280 -866 8332 -814
rect 7043 -1632 7095 -1622
rect 7043 -1666 7052 -1632
rect 7052 -1666 7086 -1632
rect 7086 -1666 7095 -1632
rect 7043 -1674 7095 -1666
rect 7235 -1632 7287 -1622
rect 7235 -1666 7244 -1632
rect 7244 -1666 7278 -1632
rect 7278 -1666 7287 -1632
rect 7235 -1674 7287 -1666
rect 7428 -1632 7480 -1621
rect 7428 -1666 7436 -1632
rect 7436 -1666 7470 -1632
rect 7470 -1666 7480 -1632
rect 7428 -1673 7480 -1666
rect 7620 -1632 7672 -1621
rect 7620 -1666 7628 -1632
rect 7628 -1666 7662 -1632
rect 7662 -1666 7672 -1632
rect 7620 -1673 7672 -1666
rect 7812 -1632 7864 -1621
rect 7812 -1666 7820 -1632
rect 7820 -1666 7854 -1632
rect 7854 -1666 7864 -1632
rect 7812 -1673 7864 -1666
rect 8003 -1632 8055 -1621
rect 8003 -1666 8012 -1632
rect 8012 -1666 8046 -1632
rect 8046 -1666 8055 -1632
rect 8003 -1673 8055 -1666
rect 8280 -1673 8332 -1621
<< metal2 >>
rect -2651 8198 -2587 8208
rect 8848 8198 8912 8208
rect -1957 8186 -1905 8196
rect -1765 8186 -1713 8196
rect -1573 8186 -1521 8196
rect -1381 8186 -1329 8196
rect -1190 8186 -1138 8196
rect -997 8186 -945 8196
rect -720 8186 -668 8196
rect 7043 8186 7095 8196
rect 7235 8186 7287 8196
rect 7427 8186 7479 8196
rect 7619 8186 7671 8196
rect 7810 8186 7862 8196
rect 8003 8186 8055 8196
rect 8280 8186 8332 8196
rect -2587 8134 -1957 8186
rect -1905 8134 -1765 8186
rect -1713 8134 -1573 8186
rect -1521 8134 -1381 8186
rect -1329 8134 -1190 8186
rect -1138 8134 -997 8186
rect -945 8134 -720 8186
rect 7036 8134 7043 8186
rect 7095 8134 7235 8186
rect 7287 8134 7427 8186
rect 7479 8134 7619 8186
rect 7671 8134 7810 8186
rect 7862 8134 8003 8186
rect 8055 8134 8280 8186
rect 8332 8134 8848 8186
rect -2651 8124 -2587 8134
rect -1957 8124 -1905 8134
rect -1765 8124 -1713 8134
rect -1573 8124 -1521 8134
rect -1381 8124 -1329 8134
rect -1190 8124 -1138 8134
rect -997 8124 -945 8134
rect -720 8124 -668 8134
rect 7043 8124 7095 8134
rect 7235 8124 7287 8134
rect 7427 8124 7479 8134
rect 7619 8124 7671 8134
rect 7810 8124 7862 8134
rect 8003 8124 8055 8134
rect 8280 8124 8332 8134
rect 8848 8124 8912 8134
rect -1022 7855 2060 7919
rect -1022 7695 -958 7855
rect -1022 7621 -958 7631
rect -2398 7390 -2334 7400
rect -1957 7379 -1905 7388
rect -1765 7379 -1713 7388
rect -1572 7379 -1520 7389
rect -1380 7379 -1328 7389
rect -1188 7379 -1136 7389
rect -997 7379 -945 7389
rect -720 7379 -668 7389
rect -1964 7378 -1572 7379
rect -2334 7326 -1957 7378
rect -1905 7327 -1765 7378
rect -2398 7316 -2334 7326
rect -1957 7316 -1905 7326
rect -1713 7327 -1572 7378
rect -1520 7327 -1380 7379
rect -1328 7327 -1188 7379
rect -1136 7327 -997 7379
rect -945 7327 -720 7379
rect -1765 7316 -1713 7326
rect -1572 7317 -1520 7327
rect -1380 7317 -1328 7327
rect -1188 7317 -1136 7327
rect -997 7317 -945 7327
rect -720 7317 -668 7327
rect 1996 6756 2060 7855
rect 6691 7697 6755 7707
rect 6691 7623 6755 7633
rect 8595 7391 8659 7401
rect 7043 7379 7095 7388
rect 7235 7379 7287 7388
rect 7428 7379 7480 7389
rect 7620 7379 7672 7389
rect 7812 7379 7864 7389
rect 8003 7379 8055 7389
rect 8280 7379 8332 7389
rect 7036 7378 7428 7379
rect 7036 7327 7043 7378
rect 7095 7327 7235 7378
rect 7043 7316 7095 7326
rect 7287 7327 7428 7378
rect 7480 7327 7620 7379
rect 7672 7327 7812 7379
rect 7864 7327 8003 7379
rect 8055 7327 8280 7379
rect 8332 7327 8595 7379
rect 7235 7316 7287 7326
rect 7428 7317 7480 7327
rect 7620 7317 7672 7327
rect 7812 7317 7864 7327
rect 8003 7317 8055 7327
rect 8280 7317 8332 7327
rect 8595 7317 8659 7327
rect 1996 6682 2060 6692
rect 1628 6476 1692 6486
rect -2651 6398 -2587 6408
rect 1628 6402 1692 6412
rect 8848 6398 8912 6408
rect -1957 6386 -1905 6396
rect -1765 6386 -1713 6396
rect -1573 6386 -1521 6396
rect -1381 6386 -1329 6396
rect -1190 6386 -1138 6396
rect -997 6386 -945 6396
rect -720 6386 -668 6396
rect 7043 6386 7095 6396
rect 7235 6386 7287 6396
rect 7427 6386 7479 6396
rect 7619 6386 7671 6396
rect 7810 6386 7862 6396
rect 8003 6386 8055 6396
rect 8280 6386 8332 6396
rect -2587 6334 -1957 6386
rect -1905 6334 -1765 6386
rect -1713 6334 -1573 6386
rect -1521 6334 -1381 6386
rect -1329 6334 -1190 6386
rect -1138 6334 -997 6386
rect -945 6334 -720 6386
rect 7036 6334 7043 6386
rect 7095 6334 7235 6386
rect 7287 6334 7427 6386
rect 7479 6334 7619 6386
rect 7671 6334 7810 6386
rect 7862 6334 8003 6386
rect 8055 6334 8280 6386
rect 8332 6334 8848 6386
rect -2651 6324 -2587 6334
rect -1957 6324 -1905 6334
rect -1765 6324 -1713 6334
rect -1573 6324 -1521 6334
rect -1381 6324 -1329 6334
rect -1190 6324 -1138 6334
rect -997 6324 -945 6334
rect -720 6324 -668 6334
rect 7043 6324 7095 6334
rect 7235 6324 7287 6334
rect 7427 6324 7479 6334
rect 7619 6324 7671 6334
rect 7810 6324 7862 6334
rect 8003 6324 8055 6334
rect 8280 6324 8332 6334
rect 8848 6324 8912 6334
rect -1028 5895 -964 5905
rect -1028 5726 -964 5831
rect -477 5893 -413 5903
rect -477 5819 -413 5829
rect 6704 5895 6768 5905
rect 6704 5821 6768 5831
rect 3410 5781 3474 5791
rect -1028 5662 -133 5726
rect -2398 5590 -2334 5600
rect -1957 5579 -1905 5588
rect -1765 5579 -1713 5588
rect -1572 5579 -1520 5589
rect -1380 5579 -1328 5589
rect -1188 5579 -1136 5589
rect -997 5579 -945 5589
rect -720 5579 -668 5589
rect -1964 5578 -1572 5579
rect -2334 5526 -1957 5578
rect -1905 5527 -1765 5578
rect -2398 5516 -2334 5526
rect -1957 5516 -1905 5526
rect -1713 5527 -1572 5578
rect -1520 5527 -1380 5579
rect -1328 5527 -1188 5579
rect -1136 5527 -997 5579
rect -945 5527 -720 5579
rect -1765 5516 -1713 5526
rect -1572 5517 -1520 5527
rect -1380 5517 -1328 5527
rect -1188 5517 -1136 5527
rect -997 5517 -945 5527
rect -720 5517 -668 5527
rect -197 5170 -133 5662
rect -197 5096 -133 5106
rect 1282 5612 1346 5622
rect -2651 4598 -2587 4608
rect -1957 4586 -1905 4596
rect -1765 4586 -1713 4596
rect -1573 4586 -1521 4596
rect -1381 4586 -1329 4596
rect -1190 4586 -1138 4596
rect -997 4586 -945 4596
rect -720 4586 -668 4596
rect -2587 4534 -1957 4586
rect -1905 4534 -1765 4586
rect -1713 4534 -1573 4586
rect -1521 4534 -1381 4586
rect -1329 4534 -1190 4586
rect -1138 4534 -997 4586
rect -945 4534 -720 4586
rect -2651 4524 -2587 4534
rect -1957 4524 -1905 4534
rect -1765 4524 -1713 4534
rect -1573 4524 -1521 4534
rect -1381 4524 -1329 4534
rect -1190 4524 -1138 4534
rect -997 4524 -945 4534
rect -720 4524 -668 4534
rect 1282 4219 1346 5548
rect 1630 5613 1694 5623
rect 1428 4219 1492 4229
rect -434 4155 1428 4219
rect -1024 4095 -960 4105
rect -1024 3923 -960 4031
rect -434 4094 -370 4155
rect 1428 4145 1492 4155
rect -434 4020 -370 4030
rect -1024 3859 -369 3923
rect -2398 3790 -2334 3800
rect -1957 3779 -1905 3788
rect -1765 3779 -1713 3788
rect -1572 3779 -1520 3789
rect -1380 3779 -1328 3789
rect -1188 3779 -1136 3789
rect -997 3779 -945 3789
rect -720 3779 -668 3789
rect -1964 3778 -1572 3779
rect -2334 3726 -1957 3778
rect -1905 3727 -1765 3778
rect -2398 3716 -2334 3726
rect -1957 3716 -1905 3726
rect -1713 3727 -1572 3778
rect -1520 3727 -1380 3779
rect -1328 3727 -1188 3779
rect -1136 3727 -997 3779
rect -945 3727 -720 3779
rect -1765 3716 -1713 3726
rect -1572 3717 -1520 3727
rect -1380 3717 -1328 3727
rect -1188 3717 -1136 3727
rect -997 3717 -945 3727
rect -720 3717 -668 3727
rect -433 3327 -369 3859
rect 1630 3843 1694 5549
rect 3157 5558 3221 5568
rect 3157 5484 3221 5494
rect 3410 5169 3474 5717
rect 8595 5591 8659 5601
rect 7043 5579 7095 5588
rect 7235 5579 7287 5588
rect 7428 5579 7480 5589
rect 7620 5579 7672 5589
rect 7812 5579 7864 5589
rect 8003 5579 8055 5589
rect 8280 5579 8332 5589
rect 7036 5578 7428 5579
rect 7036 5527 7043 5578
rect 7095 5527 7235 5578
rect 7043 5516 7095 5526
rect 7287 5527 7428 5578
rect 7480 5527 7620 5579
rect 7672 5527 7812 5579
rect 7864 5527 8003 5579
rect 8055 5527 8280 5579
rect 8332 5527 8595 5579
rect 7235 5516 7287 5526
rect 7428 5517 7480 5527
rect 7620 5517 7672 5527
rect 7812 5517 7864 5527
rect 8003 5517 8055 5527
rect 8280 5517 8332 5527
rect 8595 5517 8659 5527
rect 3410 5095 3474 5105
rect 4658 5106 4722 5116
rect 5418 5106 5482 5116
rect 3157 5084 3221 5094
rect 4722 5042 5418 5106
rect 4658 5032 4722 5042
rect 5418 5032 5482 5042
rect 3157 5010 3221 5020
rect 3768 4928 3832 4938
rect 3768 4854 3832 4864
rect 4084 4928 4148 4938
rect 5706 4928 5770 4938
rect 4148 4864 5706 4928
rect 4084 4854 4148 4864
rect 5706 4854 5770 4864
rect 6166 4932 6230 4942
rect 6166 4858 6230 4868
rect 8848 4598 8912 4608
rect 7043 4586 7095 4596
rect 7235 4586 7287 4596
rect 7427 4586 7479 4596
rect 7619 4586 7671 4596
rect 7810 4586 7862 4596
rect 8003 4586 8055 4596
rect 8280 4586 8332 4596
rect 3106 4563 3170 4573
rect 7036 4534 7043 4586
rect 7095 4534 7235 4586
rect 7287 4534 7427 4586
rect 7479 4534 7619 4586
rect 7671 4534 7810 4586
rect 7862 4534 8003 4586
rect 8055 4534 8280 4586
rect 8332 4534 8848 4586
rect 7043 4524 7095 4534
rect 7235 4524 7287 4534
rect 7427 4524 7479 4534
rect 7619 4524 7671 4534
rect 7810 4524 7862 4534
rect 8003 4524 8055 4534
rect 8280 4524 8332 4534
rect 8848 4524 8912 4534
rect 3106 4489 3170 4499
rect 5207 4390 5271 4400
rect 5207 4316 5271 4326
rect 3308 4212 3372 4222
rect 3308 4138 3372 4148
rect 6759 4095 6823 4105
rect 5952 4031 6759 4095
rect 4876 3980 4940 3990
rect 5206 3980 5270 3990
rect 4940 3916 5206 3980
rect 4876 3906 4940 3916
rect 5206 3906 5270 3916
rect 3306 3862 3370 3872
rect 1630 3779 1866 3843
rect 333 3483 397 3493
rect 333 3409 397 3419
rect 765 3483 829 3493
rect 1408 3483 1472 3493
rect 829 3419 1408 3483
rect 765 3409 829 3419
rect 1408 3409 1472 3419
rect 1631 3483 1695 3493
rect 1631 3409 1695 3419
rect 333 3327 397 3337
rect -433 3307 333 3327
rect -434 3263 333 3307
rect 397 3263 402 3327
rect -2651 2798 -2587 2808
rect -1957 2786 -1905 2796
rect -1765 2786 -1713 2796
rect -1573 2786 -1521 2796
rect -1381 2786 -1329 2796
rect -1190 2786 -1138 2796
rect -997 2786 -945 2796
rect -720 2786 -668 2796
rect -2587 2734 -1957 2786
rect -1905 2734 -1765 2786
rect -1713 2734 -1573 2786
rect -1521 2734 -1381 2786
rect -1329 2734 -1190 2786
rect -1138 2734 -997 2786
rect -945 2734 -720 2786
rect -2651 2724 -2587 2734
rect -1957 2724 -1905 2734
rect -1765 2724 -1713 2734
rect -1573 2724 -1521 2734
rect -1381 2724 -1329 2734
rect -1190 2724 -1138 2734
rect -997 2724 -945 2734
rect -720 2724 -668 2734
rect -434 2536 -370 3263
rect 333 3253 397 3263
rect 333 3154 397 3164
rect 333 3080 397 3090
rect 764 3153 828 3163
rect 1802 3153 1866 3779
rect 828 3089 1866 3153
rect 764 3079 828 3089
rect 3306 2623 3370 3798
rect 4874 3642 4938 3652
rect 4874 3568 4938 3578
rect 4510 3462 4574 3472
rect 5952 3462 6016 4031
rect 6759 4021 6823 4031
rect 8595 3791 8659 3801
rect 7043 3779 7095 3788
rect 7235 3779 7287 3788
rect 7428 3779 7480 3789
rect 7620 3779 7672 3789
rect 7812 3779 7864 3789
rect 8003 3779 8055 3789
rect 8280 3779 8332 3789
rect 7036 3778 7428 3779
rect 7036 3727 7043 3778
rect 7095 3727 7235 3778
rect 7043 3716 7095 3726
rect 7287 3727 7428 3778
rect 7480 3727 7620 3779
rect 7672 3727 7812 3779
rect 7864 3727 8003 3779
rect 8055 3727 8280 3779
rect 8332 3727 8595 3779
rect 7235 3716 7287 3726
rect 7428 3717 7480 3727
rect 7620 3717 7672 3727
rect 7812 3717 7864 3727
rect 8003 3717 8055 3727
rect 8280 3717 8332 3727
rect 8595 3717 8659 3727
rect 4574 3398 6016 3462
rect 4510 3388 4574 3398
rect 4508 3151 4572 3161
rect 4572 3087 6011 3151
rect 4508 3077 4572 3087
rect 3306 2549 3370 2559
rect -1027 2472 -370 2536
rect -1027 2295 -963 2472
rect -1027 2221 -963 2231
rect -434 2291 -370 2301
rect 5947 2297 6011 3087
rect 8848 2798 8912 2808
rect 7043 2786 7095 2796
rect 7235 2786 7287 2796
rect 7427 2786 7479 2796
rect 7619 2786 7671 2796
rect 7810 2786 7862 2796
rect 8003 2786 8055 2796
rect 8280 2786 8332 2796
rect 7036 2734 7043 2786
rect 7095 2734 7235 2786
rect 7287 2734 7427 2786
rect 7479 2734 7619 2786
rect 7671 2734 7810 2786
rect 7862 2734 8003 2786
rect 8055 2734 8280 2786
rect 8332 2734 8848 2786
rect 7043 2724 7095 2734
rect 7235 2724 7287 2734
rect 7427 2724 7479 2734
rect 7619 2724 7671 2734
rect 7810 2724 7862 2734
rect 8003 2724 8055 2734
rect 8280 2724 8332 2734
rect 8848 2724 8912 2734
rect 6764 2297 6828 2307
rect 5947 2233 6764 2297
rect -2398 1990 -2334 2000
rect -1957 1979 -1905 1988
rect -1765 1979 -1713 1988
rect -1572 1979 -1520 1989
rect -1380 1979 -1328 1989
rect -1188 1979 -1136 1989
rect -997 1979 -945 1989
rect -720 1979 -668 1989
rect -1964 1978 -1572 1979
rect -2334 1926 -1957 1978
rect -1905 1927 -1765 1978
rect -2398 1916 -2334 1926
rect -1957 1916 -1905 1926
rect -1713 1927 -1572 1978
rect -1520 1927 -1380 1979
rect -1328 1927 -1188 1979
rect -1136 1927 -997 1979
rect -945 1927 -720 1979
rect -1765 1916 -1713 1926
rect -1572 1917 -1520 1927
rect -1380 1917 -1328 1927
rect -1188 1917 -1136 1927
rect -997 1917 -945 1927
rect -720 1917 -668 1927
rect -434 1674 -370 2227
rect 3308 2223 3372 2233
rect 6764 2223 6828 2233
rect 3308 2149 3372 2159
rect 8595 1991 8659 2001
rect 7043 1979 7095 1988
rect 7235 1979 7287 1988
rect 7428 1979 7480 1989
rect 7620 1979 7672 1989
rect 7812 1979 7864 1989
rect 8003 1979 8055 1989
rect 8280 1979 8332 1989
rect 7036 1978 7428 1979
rect 7036 1927 7043 1978
rect 7095 1927 7235 1978
rect 7043 1916 7095 1926
rect 7287 1927 7428 1978
rect 7480 1927 7620 1979
rect 7672 1927 7812 1979
rect 7864 1927 8003 1979
rect 8055 1927 8280 1979
rect 8332 1927 8595 1979
rect 7235 1916 7287 1926
rect 7428 1917 7480 1927
rect 7620 1917 7672 1927
rect 7812 1917 7864 1927
rect 8003 1917 8055 1927
rect 8280 1917 8332 1927
rect 8595 1917 8659 1927
rect 4437 1704 4501 1714
rect 5426 1704 5490 1714
rect 540 1674 604 1684
rect 1830 1674 1894 1684
rect -434 1610 540 1674
rect 604 1610 1830 1674
rect 540 1600 604 1610
rect 1830 1600 1894 1610
rect 2330 1640 2394 1650
rect 4501 1640 5426 1704
rect 4437 1630 4501 1640
rect 5426 1630 5490 1640
rect 2330 1566 2394 1576
rect 3602 1526 3666 1536
rect 3602 1452 3666 1462
rect 3894 1522 3958 1532
rect 5736 1522 5800 1532
rect 3958 1458 5736 1522
rect 3894 1448 3958 1458
rect 5736 1448 5800 1458
rect 6152 1526 6216 1536
rect 6152 1452 6216 1462
rect 170 1341 234 1351
rect 170 1267 234 1277
rect 930 1341 994 1351
rect 3943 1341 4007 1351
rect 994 1277 3943 1341
rect 930 1267 994 1277
rect 3943 1267 4007 1277
rect 4326 1341 4390 1351
rect 4326 1267 4390 1277
rect -2651 998 -2587 1008
rect 8848 998 8912 1008
rect -1957 986 -1905 996
rect -1765 986 -1713 996
rect -1573 986 -1521 996
rect -1381 986 -1329 996
rect -1190 986 -1138 996
rect -997 986 -945 996
rect -720 986 -668 996
rect 7043 986 7095 996
rect 7235 986 7287 996
rect 7427 986 7479 996
rect 7619 986 7671 996
rect 7810 986 7862 996
rect 8003 986 8055 996
rect 8280 986 8332 996
rect -2587 934 -1957 986
rect -1905 934 -1765 986
rect -1713 934 -1573 986
rect -1521 934 -1381 986
rect -1329 934 -1190 986
rect -1138 934 -997 986
rect -945 934 -720 986
rect 7036 934 7043 986
rect 7095 934 7235 986
rect 7287 934 7427 986
rect 7479 934 7619 986
rect 7671 934 7810 986
rect 7862 934 8003 986
rect 8055 934 8280 986
rect 8332 934 8848 986
rect -2651 924 -2587 934
rect -1957 924 -1905 934
rect -1765 924 -1713 934
rect -1573 924 -1521 934
rect -1381 924 -1329 934
rect -1190 924 -1138 934
rect -997 924 -945 934
rect -720 924 -668 934
rect 7043 924 7095 934
rect 7235 924 7287 934
rect 7427 924 7479 934
rect 7619 924 7671 934
rect 7810 924 7862 934
rect 8003 924 8055 934
rect 8280 924 8332 934
rect 8848 924 8912 934
rect -1020 497 -956 507
rect -1020 348 -956 433
rect 6700 493 6764 503
rect 6700 419 6764 429
rect 1423 349 1487 359
rect -1020 285 1423 348
rect -1020 284 1487 285
rect 1423 275 1487 284
rect -2398 190 -2334 200
rect 8595 191 8659 201
rect -1957 179 -1905 188
rect -1765 179 -1713 188
rect -1572 179 -1520 189
rect -1380 179 -1328 189
rect -1188 179 -1136 189
rect -997 179 -945 189
rect -720 179 -668 189
rect 7043 179 7095 188
rect 7235 179 7287 188
rect 7428 179 7480 189
rect 7620 179 7672 189
rect 7812 179 7864 189
rect 8003 179 8055 189
rect 8280 179 8332 189
rect -1964 178 -1572 179
rect -2334 126 -1957 178
rect -1905 127 -1765 178
rect -2398 116 -2334 126
rect -1957 116 -1905 126
rect -1713 127 -1572 178
rect -1520 127 -1380 179
rect -1328 127 -1188 179
rect -1136 127 -997 179
rect -945 127 -720 179
rect 7036 178 7428 179
rect 7036 127 7043 178
rect -1765 116 -1713 126
rect -1572 117 -1520 127
rect -1380 117 -1328 127
rect -1188 117 -1136 127
rect -997 117 -945 127
rect -720 117 -668 127
rect 7095 127 7235 178
rect 7043 116 7095 126
rect 7287 127 7428 178
rect 7480 127 7620 179
rect 7672 127 7812 179
rect 7864 127 8003 179
rect 8055 127 8280 179
rect 8332 127 8595 179
rect 7235 116 7287 126
rect 7428 117 7480 127
rect 7620 117 7672 127
rect 7812 117 7864 127
rect 8003 117 8055 127
rect 8280 117 8332 127
rect 8595 117 8659 127
rect 160 -218 224 -208
rect -2651 -802 -2587 -792
rect -1957 -814 -1905 -804
rect -1765 -814 -1713 -804
rect -1573 -814 -1521 -804
rect -1381 -814 -1329 -804
rect -1190 -814 -1138 -804
rect -997 -814 -945 -804
rect -720 -814 -668 -804
rect -2587 -866 -1957 -814
rect -1905 -866 -1765 -814
rect -1713 -866 -1573 -814
rect -1521 -866 -1381 -814
rect -1329 -866 -1190 -814
rect -1138 -866 -997 -814
rect -945 -866 -720 -814
rect -2651 -876 -2587 -866
rect -1957 -876 -1905 -866
rect -1765 -876 -1713 -866
rect -1573 -876 -1521 -866
rect -1381 -876 -1329 -866
rect -1190 -876 -1138 -866
rect -997 -876 -945 -866
rect -720 -876 -668 -866
rect -364 -1074 -300 -1064
rect -1019 -1138 -364 -1074
rect -1019 -1304 -955 -1138
rect -364 -1148 -300 -1138
rect -1019 -1378 -955 -1368
rect -502 -1301 -438 -1291
rect 160 -1301 224 -282
rect 8848 -802 8912 -792
rect 7043 -814 7095 -804
rect 7235 -814 7287 -804
rect 7427 -814 7479 -804
rect 7619 -814 7671 -804
rect 7810 -814 7862 -804
rect 8003 -814 8055 -804
rect 8280 -814 8332 -804
rect 7036 -866 7043 -814
rect 7095 -866 7235 -814
rect 7287 -866 7427 -814
rect 7479 -866 7619 -814
rect 7671 -866 7810 -814
rect 7862 -866 8003 -814
rect 8055 -866 8280 -814
rect 8332 -866 8848 -814
rect 7043 -876 7095 -866
rect 7235 -876 7287 -866
rect 7427 -876 7479 -866
rect 7619 -876 7671 -866
rect 7810 -876 7862 -866
rect 8003 -876 8055 -866
rect 8280 -876 8332 -866
rect 8848 -876 8912 -866
rect -438 -1365 224 -1301
rect 6718 -1299 6782 -1289
rect -502 -1375 -438 -1365
rect 6718 -1373 6782 -1363
rect -2398 -1610 -2334 -1600
rect 8595 -1609 8659 -1599
rect -1957 -1621 -1905 -1612
rect -1765 -1621 -1713 -1612
rect -1572 -1621 -1520 -1611
rect -1380 -1621 -1328 -1611
rect -1188 -1621 -1136 -1611
rect -997 -1621 -945 -1611
rect -720 -1621 -668 -1611
rect 7043 -1621 7095 -1612
rect 7235 -1621 7287 -1612
rect 7428 -1621 7480 -1611
rect 7620 -1621 7672 -1611
rect 7812 -1621 7864 -1611
rect 8003 -1621 8055 -1611
rect 8280 -1621 8332 -1611
rect -1964 -1622 -1572 -1621
rect -2334 -1674 -1957 -1622
rect -1905 -1673 -1765 -1622
rect -2398 -1684 -2334 -1674
rect -1957 -1684 -1905 -1674
rect -1713 -1673 -1572 -1622
rect -1520 -1673 -1380 -1621
rect -1328 -1673 -1188 -1621
rect -1136 -1673 -997 -1621
rect -945 -1673 -720 -1621
rect 7036 -1622 7428 -1621
rect 7036 -1673 7043 -1622
rect -1765 -1684 -1713 -1674
rect -1572 -1683 -1520 -1673
rect -1380 -1683 -1328 -1673
rect -1188 -1683 -1136 -1673
rect -997 -1683 -945 -1673
rect -720 -1683 -668 -1673
rect 7095 -1673 7235 -1622
rect 7043 -1684 7095 -1674
rect 7287 -1673 7428 -1622
rect 7480 -1673 7620 -1621
rect 7672 -1673 7812 -1621
rect 7864 -1673 8003 -1621
rect 8055 -1673 8280 -1621
rect 8332 -1673 8595 -1621
rect 7235 -1684 7287 -1674
rect 7428 -1683 7480 -1673
rect 7620 -1683 7672 -1673
rect 7812 -1683 7864 -1673
rect 8003 -1683 8055 -1673
rect 8280 -1683 8332 -1673
rect 8595 -1683 8659 -1673
<< via2 >>
rect -2651 8134 -2587 8198
rect 8848 8134 8912 8198
rect -2398 7326 -2334 7390
rect 6691 7633 6755 7697
rect 8595 7327 8659 7391
rect 1996 6692 2060 6756
rect 1628 6412 1692 6476
rect -2651 6334 -2587 6398
rect 8848 6334 8912 6398
rect -477 5829 -413 5893
rect 6704 5831 6768 5895
rect -2398 5526 -2334 5590
rect 3410 5717 3474 5781
rect -197 5106 -133 5170
rect 1282 5548 1346 5612
rect -2651 4534 -2587 4598
rect 1630 5549 1694 5613
rect 1428 4155 1492 4219
rect -2398 3726 -2334 3790
rect 3157 5494 3221 5558
rect 8595 5527 8659 5591
rect 3410 5105 3474 5169
rect 3157 5020 3221 5084
rect 4658 5042 4722 5106
rect 5418 5042 5482 5106
rect 3768 4864 3832 4928
rect 4084 4864 4148 4928
rect 5706 4864 5770 4928
rect 6166 4868 6230 4932
rect 3106 4499 3170 4563
rect 8848 4534 8912 4598
rect 5207 4326 5271 4390
rect 3308 4148 3372 4212
rect 4876 3916 4940 3980
rect 5206 3916 5270 3980
rect 333 3419 397 3483
rect 765 3419 829 3483
rect 1408 3419 1472 3483
rect 1631 3419 1695 3483
rect 333 3263 397 3327
rect -2651 2734 -2587 2798
rect 333 3090 397 3154
rect 764 3089 828 3153
rect 3306 3798 3370 3862
rect 4874 3578 4938 3642
rect 8595 3727 8659 3791
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3306 2559 3370 2623
rect 8848 2734 8912 2798
rect -2398 1926 -2334 1990
rect 3308 2159 3372 2223
rect 8595 1927 8659 1991
rect 540 1610 604 1674
rect 1830 1610 1894 1674
rect 2330 1576 2394 1640
rect 4437 1640 4501 1704
rect 5426 1640 5490 1704
rect 3602 1462 3666 1526
rect 3894 1458 3958 1522
rect 5736 1458 5800 1522
rect 6152 1462 6216 1526
rect 170 1277 234 1341
rect 930 1277 994 1341
rect 3943 1277 4007 1341
rect 4326 1277 4390 1341
rect -2651 934 -2587 998
rect 8848 934 8912 998
rect 6700 429 6764 493
rect 1423 285 1487 349
rect -2398 126 -2334 190
rect 8595 127 8659 191
rect 160 -282 224 -218
rect -2651 -866 -2587 -802
rect -364 -1138 -300 -1074
rect 8848 -866 8912 -802
rect 6718 -1363 6782 -1299
rect -2398 -1674 -2334 -1610
rect 8595 -1673 8659 -1609
<< metal3 >>
rect -2651 8203 -2587 8208
rect -2661 8198 -2577 8203
rect -2661 8134 -2651 8198
rect -2587 8134 -2577 8198
rect -2661 8129 -2577 8134
rect -2651 6403 -2587 8129
rect -2398 7395 -2334 7400
rect -2408 7390 -2324 7395
rect -2408 7326 -2398 7390
rect -2334 7326 -2324 7390
rect -2408 7321 -2324 7326
rect -2661 6398 -2577 6403
rect -2661 6334 -2651 6398
rect -2587 6334 -2577 6398
rect -2661 6329 -2577 6334
rect -2651 4603 -2587 6329
rect -2398 5595 -2334 7321
rect -1800 7200 -642 8360
rect 0 7200 1158 8360
rect 1800 7200 2958 8360
rect 3600 7200 4758 8360
rect 5400 7200 6558 8360
rect 6681 7697 6765 7702
rect 6681 7633 6691 7697
rect 6755 7633 6765 7697
rect 6681 7628 6765 7633
rect 1975 6756 2080 6780
rect 6691 6779 6755 7628
rect 7200 7200 8358 8360
rect 8848 8203 8912 8208
rect 8838 8198 8922 8203
rect 8838 8134 8848 8198
rect 8912 8134 8922 8198
rect 8838 8129 8922 8134
rect 8595 7396 8659 7401
rect 8585 7391 8669 7396
rect 8585 7327 8595 7391
rect 8659 7327 8669 7391
rect 8585 7322 8669 7327
rect 1975 6692 1996 6756
rect 2060 6692 2080 6756
rect 1975 6669 2080 6692
rect 6191 6715 6755 6779
rect 6191 6560 6255 6715
rect -2408 5590 -2324 5595
rect -2408 5526 -2398 5590
rect -2334 5526 -2324 5590
rect -2408 5521 -2324 5526
rect -2661 4598 -2577 4603
rect -2661 4534 -2651 4598
rect -2587 4534 -2577 4598
rect -2661 4529 -2577 4534
rect -2651 4524 -2587 4529
rect -2398 3795 -2334 5521
rect -1800 5400 -642 6560
rect -497 5893 -391 5915
rect -497 5829 -477 5893
rect -413 5829 -391 5893
rect -497 5808 -391 5829
rect 0 5612 1158 6560
rect 1618 6476 1702 6481
rect 1800 6476 2958 6560
rect 1618 6412 1628 6476
rect 1692 6412 2958 6476
rect 1618 6407 1702 6412
rect 1272 5612 1356 5617
rect 0 5548 1282 5612
rect 1346 5548 1356 5612
rect 0 5400 1158 5548
rect 1272 5543 1356 5548
rect 1616 5613 1708 5646
rect 1616 5549 1630 5613
rect 1694 5549 1708 5613
rect 1616 5524 1708 5549
rect 1800 5400 2958 6412
rect 3600 6197 4758 6560
rect 3157 6133 4758 6197
rect 3157 5563 3221 6133
rect 3400 5781 3484 5810
rect 3400 5717 3410 5781
rect 3474 5717 3484 5781
rect 3400 5693 3484 5717
rect 3147 5558 3231 5563
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 3147 5489 3231 5494
rect 3600 5400 4758 6133
rect 5400 5400 6558 6560
rect 6686 5895 6784 5914
rect 6686 5831 6704 5895
rect 6768 5831 6784 5895
rect 6686 5814 6784 5831
rect 7200 5400 8358 6560
rect 8595 5596 8659 7322
rect 8848 6403 8912 8129
rect 8838 6398 8922 6403
rect 8838 6334 8848 6398
rect 8912 6334 8922 6398
rect 8838 6329 8922 6334
rect 8585 5591 8669 5596
rect 8585 5527 8595 5591
rect 8659 5527 8669 5591
rect 8585 5522 8669 5527
rect 544 5311 608 5400
rect 544 5247 5105 5311
rect -238 5170 -98 5201
rect -238 5106 -197 5170
rect -133 5106 -98 5170
rect -238 5072 -98 5106
rect 3379 5169 3508 5177
rect 3379 5105 3410 5169
rect 3474 5105 3508 5169
rect 3379 5097 3508 5105
rect 4648 5106 4732 5111
rect 3147 5084 3231 5089
rect 754 5020 3157 5084
rect 3221 5020 3231 5084
rect 4648 5042 4658 5106
rect 4722 5042 4732 5106
rect 4648 5037 4732 5042
rect 754 4760 818 5020
rect 3147 5015 3231 5020
rect 3758 4928 3842 4933
rect 1241 4864 3768 4928
rect 3832 4864 3842 4928
rect -2408 3790 -2324 3795
rect -2408 3726 -2398 3790
rect -2334 3726 -2324 3790
rect -2408 3721 -2324 3726
rect -1800 3600 -642 4760
rect 0 3600 1158 4760
rect 333 3488 397 3600
rect 323 3483 407 3488
rect 323 3419 333 3483
rect 397 3419 407 3483
rect 323 3414 407 3419
rect 743 3483 849 3501
rect 743 3419 765 3483
rect 829 3419 849 3483
rect 333 3332 397 3414
rect 743 3404 849 3419
rect 323 3327 407 3332
rect 323 3263 333 3327
rect 397 3263 407 3327
rect 323 3258 407 3263
rect 333 3159 397 3258
rect 323 3154 407 3159
rect 323 3090 333 3154
rect 397 3090 407 3154
rect 323 3085 407 3090
rect 745 3158 837 3183
rect 745 3153 838 3158
rect 745 3089 764 3153
rect 828 3089 838 3153
rect 333 2960 397 3085
rect 745 3084 838 3089
rect 745 3061 837 3084
rect -2651 2803 -2587 2808
rect -2661 2798 -2577 2803
rect -2661 2734 -2651 2798
rect -2587 2734 -2577 2798
rect -2661 2729 -2577 2734
rect -2651 1003 -2587 2729
rect -2398 1995 -2334 2000
rect -2408 1990 -2324 1995
rect -2408 1926 -2398 1990
rect -2334 1926 -2324 1990
rect -2408 1921 -2324 1926
rect -2661 998 -2577 1003
rect -2661 934 -2651 998
rect -2587 934 -2577 998
rect -2661 929 -2577 934
rect -2651 -797 -2587 929
rect -2398 195 -2334 1921
rect -1800 1800 -642 2960
rect 0 1800 1158 2960
rect 170 1346 234 1800
rect 530 1674 614 1679
rect 530 1610 540 1674
rect 604 1610 614 1674
rect 530 1605 614 1610
rect 160 1341 244 1346
rect 160 1277 170 1341
rect 234 1277 244 1341
rect 160 1272 244 1277
rect 540 1160 604 1605
rect 910 1341 1011 1357
rect 910 1277 930 1341
rect 994 1277 1011 1341
rect 910 1259 1011 1277
rect -2408 190 -2324 195
rect -2408 126 -2398 190
rect -2334 126 -2324 190
rect -2408 121 -2324 126
rect -2661 -802 -2577 -797
rect -2661 -866 -2651 -802
rect -2587 -866 -2577 -802
rect -2661 -871 -2577 -866
rect -2651 -876 -2587 -871
rect -2398 -1605 -2334 121
rect -1800 0 -642 1160
rect 0 354 1158 1160
rect 1241 354 1305 4864
rect 3758 4859 3842 4864
rect 4061 4928 4171 4944
rect 4061 4864 4084 4928
rect 4148 4864 4171 4928
rect 4061 4850 4171 4864
rect 4658 4760 4722 5037
rect 1418 4219 1502 4224
rect 1800 4219 2958 4760
rect 3081 4563 3190 4586
rect 3081 4499 3106 4563
rect 3170 4499 3190 4563
rect 3081 4479 3190 4499
rect 1418 4155 1428 4219
rect 1492 4155 2958 4219
rect 1418 4150 1502 4155
rect 1800 3600 2958 4155
rect 3298 4212 3382 4217
rect 3600 4212 4758 4760
rect 3298 4148 3308 4212
rect 3372 4148 4758 4212
rect 3298 4143 3382 4148
rect 3283 3862 3389 3885
rect 3283 3798 3306 3862
rect 3370 3798 3389 3862
rect 3283 3778 3389 3798
rect 3600 3600 4758 4148
rect 4862 3980 4953 4019
rect 4862 3916 4876 3980
rect 4940 3916 4953 3980
rect 4862 3879 4953 3916
rect 4864 3642 4948 3647
rect 1397 3483 1484 3517
rect 1397 3419 1408 3483
rect 1472 3419 1484 3483
rect 1397 3388 1484 3419
rect 1621 3483 1705 3488
rect 1621 3419 1631 3483
rect 1695 3419 1705 3483
rect 1621 3414 1705 3419
rect 2348 3432 2412 3600
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 4864 3573 4948 3578
rect 4479 3462 4604 3492
rect 0 290 1305 354
rect 1405 349 1503 380
rect 0 0 1158 290
rect 1405 285 1423 349
rect 1487 285 1503 349
rect 1631 365 1695 3414
rect 2348 3368 3912 3432
rect 4479 3398 4510 3462
rect 4574 3398 4604 3462
rect 4479 3371 4604 3398
rect 3848 2960 3912 3368
rect 4486 3151 4590 3171
rect 4486 3087 4508 3151
rect 4572 3087 4590 3151
rect 4486 3071 4590 3087
rect 1800 2223 2958 2960
rect 3284 2623 3390 2645
rect 3284 2559 3306 2623
rect 3370 2559 3390 2623
rect 3284 2538 3390 2559
rect 3298 2223 3382 2228
rect 1800 2159 3308 2223
rect 3372 2159 3382 2223
rect 1800 1800 2958 2159
rect 3298 2154 3382 2159
rect 3600 1800 4758 2960
rect 1830 1679 1894 1800
rect 4437 1709 4501 1800
rect 4427 1704 4511 1709
rect 1820 1674 1904 1679
rect 1820 1610 1830 1674
rect 1894 1610 1904 1674
rect 1820 1605 1904 1610
rect 2307 1640 2415 1666
rect 2307 1576 2330 1640
rect 2394 1576 2415 1640
rect 4427 1640 4437 1704
rect 4501 1640 4511 1704
rect 4427 1635 4511 1640
rect 2307 1553 2415 1576
rect 3592 1526 3676 1531
rect 3083 1462 3602 1526
rect 3666 1462 3676 1526
rect 1800 365 2958 1160
rect 1631 363 2958 365
rect 3083 363 3147 1462
rect 3592 1457 3676 1462
rect 3873 1522 3978 1546
rect 3873 1458 3894 1522
rect 3958 1458 3978 1522
rect 3873 1437 3978 1458
rect 3923 1341 4024 1360
rect 3923 1277 3943 1341
rect 4007 1277 4024 1341
rect 3923 1262 4024 1277
rect 4316 1341 4400 1346
rect 4316 1277 4326 1341
rect 4390 1277 4400 1341
rect 4316 1272 4400 1277
rect 4326 1160 4390 1272
rect 1631 301 3147 363
rect 1405 260 1503 285
rect 1800 299 3147 301
rect 3600 448 4758 1160
rect 4874 448 4938 3573
rect 5041 616 5105 5247
rect 5418 5111 5482 5400
rect 5408 5106 5492 5111
rect 5408 5042 5418 5106
rect 5482 5042 5492 5106
rect 5408 5037 5492 5042
rect 5683 4928 5793 4943
rect 6166 4937 6230 5400
rect 5683 4864 5706 4928
rect 5770 4864 5793 4928
rect 5683 4849 5793 4864
rect 6156 4932 6240 4937
rect 6156 4868 6166 4932
rect 6230 4868 6240 4932
rect 6156 4863 6240 4868
rect 5197 4390 5281 4395
rect 5400 4390 6558 4760
rect 5197 4326 5207 4390
rect 5271 4326 6558 4390
rect 5197 4321 5281 4326
rect 5193 3980 5284 4018
rect 5193 3916 5206 3980
rect 5270 3916 5284 3980
rect 5193 3878 5284 3916
rect 5400 3600 6558 4326
rect 7200 3600 8358 4760
rect 8595 3796 8659 5522
rect 8848 4603 8912 6329
rect 8838 4598 8922 4603
rect 8838 4534 8848 4598
rect 8912 4534 8922 4598
rect 8838 4529 8922 4534
rect 8585 3791 8669 3796
rect 8585 3727 8595 3791
rect 8659 3727 8669 3791
rect 8585 3722 8669 3727
rect 8595 3717 8659 3722
rect 5400 1800 6558 2960
rect 7200 1800 8358 2960
rect 8848 2803 8912 2808
rect 8838 2798 8922 2803
rect 8838 2734 8848 2798
rect 8912 2734 8922 2798
rect 8838 2729 8922 2734
rect 8595 1996 8659 2001
rect 8585 1991 8669 1996
rect 8585 1927 8595 1991
rect 8659 1927 8669 1991
rect 8585 1922 8669 1927
rect 5416 1704 5500 1709
rect 5416 1640 5426 1704
rect 5490 1640 5500 1704
rect 5416 1635 5500 1640
rect 5426 1160 5490 1635
rect 5715 1522 5820 1544
rect 6152 1531 6216 1800
rect 5715 1458 5736 1522
rect 5800 1458 5820 1522
rect 5715 1435 5820 1458
rect 6142 1526 6226 1531
rect 6142 1462 6152 1526
rect 6216 1462 6226 1526
rect 6142 1457 6226 1462
rect 5400 616 6558 1160
rect 5041 552 6558 616
rect 3600 384 4941 448
rect 1800 0 2958 299
rect 3600 0 4758 384
rect 5400 0 6558 552
rect 6683 493 6785 514
rect 6683 429 6700 493
rect 6764 429 6785 493
rect 6683 411 6785 429
rect 7200 0 8358 1160
rect 8595 196 8659 1922
rect 8848 1003 8912 2729
rect 8838 998 8922 1003
rect 8838 934 8848 998
rect 8912 934 8922 998
rect 8838 929 8922 934
rect 8585 191 8669 196
rect 8585 127 8595 191
rect 8659 127 8669 191
rect 8585 122 8669 127
rect 139 -218 245 -195
rect 139 -282 160 -218
rect 224 -282 245 -218
rect 139 -299 245 -282
rect 6179 -442 6243 0
rect 6179 -506 6782 -442
rect -2408 -1610 -2324 -1605
rect -2408 -1674 -2398 -1610
rect -2334 -1674 -2324 -1610
rect -2408 -1679 -2324 -1674
rect -2398 -1684 -2334 -1679
rect -1800 -1800 -642 -640
rect -378 -1074 -280 -1056
rect -378 -1138 -364 -1074
rect -300 -1138 -280 -1074
rect -378 -1159 -280 -1138
rect 0 -1800 1158 -640
rect 1800 -1800 2958 -640
rect 3600 -1800 4758 -640
rect 5400 -1800 6558 -640
rect 6718 -1294 6782 -506
rect 6708 -1299 6792 -1294
rect 6708 -1363 6718 -1299
rect 6782 -1363 6792 -1299
rect 6708 -1368 6792 -1363
rect 6718 -1372 6782 -1368
rect 7200 -1800 8358 -640
rect 8595 -1604 8659 122
rect 8848 -797 8912 929
rect 8838 -802 8922 -797
rect 8838 -866 8848 -802
rect 8912 -866 8922 -802
rect 8838 -871 8922 -866
rect 8585 -1609 8669 -1604
rect 8585 -1673 8595 -1609
rect 8659 -1673 8669 -1609
rect 8585 -1678 8669 -1673
rect 8595 -1683 8659 -1678
<< via3 >>
rect 1996 6692 2060 6756
rect -477 5829 -413 5893
rect 1630 5549 1694 5613
rect 3410 5717 3474 5781
rect 6704 5831 6768 5895
rect -197 5106 -133 5170
rect 3410 5105 3474 5169
rect 765 3419 829 3483
rect 764 3089 828 3153
rect 930 1277 994 1341
rect 4084 4864 4148 4928
rect 3106 4499 3170 4563
rect 3306 3798 3370 3862
rect 4876 3916 4940 3980
rect 1408 3419 1472 3483
rect 1423 285 1487 349
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3306 2559 3370 2623
rect 2330 1576 2394 1640
rect 3894 1458 3958 1522
rect 3943 1277 4007 1341
rect 5706 4864 5770 4928
rect 5206 3916 5270 3980
rect 5736 1458 5800 1522
rect 6700 429 6764 493
rect 160 -282 224 -218
rect -364 -1138 -300 -1074
<< mimcap >>
rect -1700 8220 -740 8260
rect -1700 7340 -1660 8220
rect -780 7340 -740 8220
rect -1700 7300 -740 7340
rect 100 8220 1060 8260
rect 100 7340 140 8220
rect 1020 7340 1060 8220
rect 100 7300 1060 7340
rect 1900 8220 2860 8260
rect 1900 7340 1940 8220
rect 2820 7340 2860 8220
rect 1900 7300 2860 7340
rect 3700 8220 4660 8260
rect 3700 7340 3740 8220
rect 4620 7340 4660 8220
rect 3700 7300 4660 7340
rect 5500 8220 6460 8260
rect 5500 7340 5540 8220
rect 6420 7340 6460 8220
rect 5500 7300 6460 7340
rect 7300 8220 8260 8260
rect 7300 7340 7340 8220
rect 8220 7340 8260 8220
rect 7300 7300 8260 7340
rect -1700 6420 -740 6460
rect -1700 5540 -1660 6420
rect -780 5540 -740 6420
rect -1700 5500 -740 5540
rect 100 6420 1060 6460
rect 100 5540 140 6420
rect 1020 5540 1060 6420
rect 100 5500 1060 5540
rect 1900 6420 2860 6460
rect 1900 5540 1940 6420
rect 2820 5540 2860 6420
rect 1900 5500 2860 5540
rect 3700 6420 4660 6460
rect 3700 5540 3740 6420
rect 4620 5540 4660 6420
rect 3700 5500 4660 5540
rect 5500 6420 6460 6460
rect 5500 5540 5540 6420
rect 6420 5540 6460 6420
rect 5500 5500 6460 5540
rect 7300 6420 8260 6460
rect 7300 5540 7340 6420
rect 8220 5540 8260 6420
rect 7300 5500 8260 5540
rect -1700 4620 -740 4660
rect -1700 3740 -1660 4620
rect -780 3740 -740 4620
rect -1700 3700 -740 3740
rect 100 4620 1060 4660
rect 100 3740 140 4620
rect 1020 3740 1060 4620
rect 100 3700 1060 3740
rect 1900 4620 2860 4660
rect 1900 3740 1940 4620
rect 2820 3740 2860 4620
rect 1900 3700 2860 3740
rect 3700 4620 4660 4660
rect 3700 3740 3740 4620
rect 4620 3740 4660 4620
rect 3700 3700 4660 3740
rect 5500 4620 6460 4660
rect 5500 3740 5540 4620
rect 6420 3740 6460 4620
rect 5500 3700 6460 3740
rect 7300 4620 8260 4660
rect 7300 3740 7340 4620
rect 8220 3740 8260 4620
rect 7300 3700 8260 3740
rect -1700 2820 -740 2860
rect -1700 1940 -1660 2820
rect -780 1940 -740 2820
rect -1700 1900 -740 1940
rect 100 2820 1060 2860
rect 100 1940 140 2820
rect 1020 1940 1060 2820
rect 100 1900 1060 1940
rect 1900 2820 2860 2860
rect 1900 1940 1940 2820
rect 2820 1940 2860 2820
rect 1900 1900 2860 1940
rect 3700 2820 4660 2860
rect 3700 1940 3740 2820
rect 4620 1940 4660 2820
rect 3700 1900 4660 1940
rect 5500 2820 6460 2860
rect 5500 1940 5540 2820
rect 6420 1940 6460 2820
rect 5500 1900 6460 1940
rect 7300 2820 8260 2860
rect 7300 1940 7340 2820
rect 8220 1940 8260 2820
rect 7300 1900 8260 1940
rect -1700 1020 -740 1060
rect -1700 140 -1660 1020
rect -780 140 -740 1020
rect -1700 100 -740 140
rect 100 1020 1060 1060
rect 100 140 140 1020
rect 1020 140 1060 1020
rect 100 100 1060 140
rect 1900 1020 2860 1060
rect 1900 140 1940 1020
rect 2820 140 2860 1020
rect 1900 100 2860 140
rect 3700 1020 4660 1060
rect 3700 140 3740 1020
rect 4620 140 4660 1020
rect 3700 100 4660 140
rect 5500 1020 6460 1060
rect 5500 140 5540 1020
rect 6420 140 6460 1020
rect 5500 100 6460 140
rect 7300 1020 8260 1060
rect 7300 140 7340 1020
rect 8220 140 8260 1020
rect 7300 100 8260 140
rect -1700 -780 -740 -740
rect -1700 -1660 -1660 -780
rect -780 -1660 -740 -780
rect -1700 -1700 -740 -1660
rect 100 -780 1060 -740
rect 100 -1660 140 -780
rect 1020 -1660 1060 -780
rect 100 -1700 1060 -1660
rect 1900 -780 2860 -740
rect 1900 -1660 1940 -780
rect 2820 -1660 2860 -780
rect 1900 -1700 2860 -1660
rect 3700 -780 4660 -740
rect 3700 -1660 3740 -780
rect 4620 -1660 4660 -780
rect 3700 -1700 4660 -1660
rect 5500 -780 6460 -740
rect 5500 -1660 5540 -780
rect 6420 -1660 6460 -780
rect 5500 -1700 6460 -1660
rect 7300 -780 8260 -740
rect 7300 -1660 7340 -780
rect 8220 -1660 8260 -780
rect 7300 -1700 8260 -1660
<< mimcapcontact >>
rect -1660 7340 -780 8220
rect 140 7340 1020 8220
rect 1940 7340 2820 8220
rect 3740 7340 4620 8220
rect 5540 7340 6420 8220
rect 7340 7340 8220 8220
rect -1660 5540 -780 6420
rect 140 5540 1020 6420
rect 1940 5540 2820 6420
rect 3740 5540 4620 6420
rect 5540 5540 6420 6420
rect 7340 5540 8220 6420
rect -1660 3740 -780 4620
rect 140 3740 1020 4620
rect 1940 3740 2820 4620
rect 3740 3740 4620 4620
rect 5540 3740 6420 4620
rect 7340 3740 8220 4620
rect -1660 1940 -780 2820
rect 140 1940 1020 2820
rect 1940 1940 2820 2820
rect 3740 1940 4620 2820
rect 5540 1940 6420 2820
rect 7340 1940 8220 2820
rect -1660 140 -780 1020
rect 140 140 1020 1020
rect 1940 140 2820 1020
rect 3740 140 4620 1020
rect 5540 140 6420 1020
rect 7340 140 8220 1020
rect -1660 -1660 -780 -780
rect 140 -1660 1020 -780
rect 1940 -1660 2820 -780
rect 3740 -1660 4620 -780
rect 5540 -1660 6420 -780
rect 7340 -1660 8220 -780
<< metal4 >>
rect 1995 6756 2061 6757
rect 1995 6692 1996 6756
rect 2060 6692 2061 6756
rect 1995 6691 2061 6692
rect 1996 6420 2060 6691
rect -478 5893 -412 5894
rect -478 5829 -477 5893
rect -413 5829 140 5893
rect -478 5828 -412 5829
rect 1629 5613 1695 5614
rect 1629 5549 1630 5613
rect 1694 5549 1940 5613
rect 1629 5548 1695 5549
rect 3409 5781 3475 5782
rect 3409 5717 3410 5781
rect 3474 5717 3740 5781
rect 3409 5716 3475 5717
rect 6703 5895 6769 5896
rect 6420 5831 6704 5895
rect 6768 5831 6769 5895
rect 6703 5830 6769 5831
rect 544 5311 608 5540
rect 544 5247 5105 5311
rect -198 5170 -132 5171
rect -198 5106 -197 5170
rect -133 5169 -132 5170
rect 3409 5169 3475 5170
rect -133 5106 3410 5169
rect -198 5105 3410 5106
rect 3474 5105 3475 5169
rect 320 4620 384 5105
rect 3409 5104 3475 5105
rect 4083 4928 4149 4929
rect 1242 4864 4084 4928
rect 4148 4864 4150 4928
rect 765 3484 829 3740
rect 764 3483 830 3484
rect 764 3419 765 3483
rect 829 3419 830 3483
rect 764 3418 830 3419
rect 763 3153 829 3154
rect 763 3089 764 3153
rect 828 3089 829 3153
rect 763 3088 829 3089
rect 764 2820 828 3088
rect -364 1985 140 2049
rect -364 -1073 -300 1985
rect 930 1342 994 1940
rect 929 1341 995 1342
rect 929 1277 930 1341
rect 994 1277 995 1341
rect 929 1276 995 1277
rect 1242 859 1306 4864
rect 4083 4863 4149 4864
rect 3105 4563 3171 4564
rect 2820 4499 3106 4563
rect 3170 4499 3171 4563
rect 3105 4498 3171 4499
rect 3305 3862 3371 3863
rect 3305 3798 3306 3862
rect 3370 3798 3740 3862
rect 3305 3797 3371 3798
rect 4875 3980 4941 3981
rect 4875 3916 4876 3980
rect 4940 3916 4941 3980
rect 4875 3915 4941 3916
rect 1407 3483 1473 3484
rect 1407 3419 1408 3483
rect 1472 3419 1473 3483
rect 1407 3418 1473 3419
rect 2348 3432 2412 3740
rect 4510 3463 4574 3740
rect 4509 3462 4575 3463
rect 1020 795 1306 859
rect 1408 813 1472 3418
rect 2348 3368 3912 3432
rect 4509 3398 4510 3462
rect 4574 3398 4575 3462
rect 4509 3397 4575 3398
rect 3848 2820 3912 3368
rect 4507 3151 4573 3152
rect 4507 3087 4508 3151
rect 4572 3087 4573 3151
rect 4507 3086 4573 3087
rect 4508 2820 4572 3086
rect 3305 2623 3371 2624
rect 2820 2559 3306 2623
rect 3370 2559 3371 2623
rect 3305 2558 3371 2559
rect 2330 1641 2394 1940
rect 2329 1640 2395 1641
rect 2329 1576 2330 1640
rect 2394 1576 2395 1640
rect 2329 1575 2395 1576
rect 3893 1522 3959 1523
rect 3083 1458 3894 1522
rect 3958 1458 3959 1522
rect 1408 749 1940 813
rect 1422 349 1488 350
rect 1420 285 1423 349
rect 1487 285 1940 349
rect 1422 284 1488 285
rect 3083 812 3147 1458
rect 3893 1457 3959 1458
rect 3943 1342 4007 1345
rect 3942 1341 4008 1342
rect 3942 1277 3943 1341
rect 4007 1277 4008 1341
rect 3942 1276 4008 1277
rect 3943 1020 4007 1276
rect 2820 748 3147 812
rect 4876 844 4940 3915
rect 4620 780 4940 844
rect 5041 616 5105 5247
rect 5706 4929 5770 5540
rect 5705 4928 5771 4929
rect 5705 4864 5706 4928
rect 5770 4864 5771 4928
rect 5705 4863 5771 4864
rect 5205 3980 5271 3981
rect 5205 3916 5206 3980
rect 5270 3916 5540 3980
rect 5205 3915 5271 3916
rect 5736 1523 5800 1940
rect 5735 1522 5801 1523
rect 5735 1458 5736 1522
rect 5800 1458 5801 1522
rect 5735 1457 5801 1458
rect 5041 552 5540 616
rect 6699 493 6765 494
rect 6420 429 6700 493
rect 6764 429 6766 493
rect 6699 428 6765 429
rect 160 -217 224 140
rect 159 -218 225 -217
rect 159 -282 160 -218
rect 224 -282 225 -218
rect 159 -283 225 -282
rect -365 -1074 -299 -1073
rect -365 -1138 -364 -1074
rect -300 -1138 -299 -1074
rect -365 -1139 -299 -1138
<< labels >>
flabel metal3 -2642 8019 -2642 8019 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal3 -2389 7236 -2389 7236 1 FreeSans 400 0 0 0 p2
port 7 n
flabel metal3 -2639 2626 -2639 2626 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal3 -2389 1840 -2389 1840 1 FreeSans 400 0 0 0 p1
port 9 n
flabel metal3 8645 -1537 8645 -1537 1 FreeSans 400 0 0 0 p1
port 9 n
flabel metal3 8898 -670 8898 -670 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal3 8648 7246 8648 7246 1 FreeSans 400 0 0 0 p2
port 7 n
flabel metal3 8904 8016 8904 8016 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal1 -3484 3369 -3484 3369 1 FreeSans 400 0 0 0 op
port 4 n
flabel metal1 -2872 3368 -2872 3368 1 FreeSans 400 0 0 0 on
port 1 n
flabel metal1 -2412 3371 -2412 3371 1 FreeSans 400 0 0 0 cmc
port 5 n
flabel metal1 8790 3295 8790 3295 1 FreeSans 400 0 0 0 cm
port 2 n
flabel metal1 9292 3298 9292 3298 1 FreeSans 400 0 0 0 bias_a
port 3 n
flabel metal1 -2046 8350 -2046 8350 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 7178 -2045 7178 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2043 6543 -2043 6543 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 5370 -2045 5370 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2043 4743 -2043 4743 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2047 3574 -2047 3574 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2047 2942 -2047 2942 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 1776 -2045 1776 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2043 1146 -2043 1146 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2047 -27 -2047 -27 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2045 -659 -2045 -659 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 -1822 -2045 -1822 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6957 -1822 6957 -1822 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6954 -659 6954 -659 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6957 -26 6957 -26 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6952 1141 6952 1141 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6952 1776 6952 1776 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6954 2944 6954 2944 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6954 3579 6954 3579 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6957 4740 6957 4740 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6954 5375 6954 5375 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6952 6547 6952 6547 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6954 7180 6954 7180 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6954 8345 6954 8345 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -646 -840 -646 -840 7 FreeSans 400 0 0 0 transmission_gate_11/en_b
flabel metal1 -645 -1336 -645 -1336 7 FreeSans 400 0 0 0 transmission_gate_11/in
flabel metal1 -645 -1647 -645 -1647 7 FreeSans 400 0 0 0 transmission_gate_11/en
flabel metal1 -2136 -1337 -2136 -1337 3 FreeSans 400 0 0 0 transmission_gate_11/out
flabel metal1 -2045 -691 -2045 -691 5 FreeSans 400 0 0 0 transmission_gate_11/VDD
flabel metal1 -2045 -1797 -2045 -1797 1 FreeSans 400 0 0 0 transmission_gate_11/VSS
flabel metal1 8354 -840 8354 -840 7 FreeSans 400 0 0 0 transmission_gate_2/en_b
flabel metal1 8355 -1336 8355 -1336 7 FreeSans 400 0 0 0 transmission_gate_2/in
flabel metal1 8355 -1647 8355 -1647 7 FreeSans 400 0 0 0 transmission_gate_2/en
flabel metal1 6864 -1337 6864 -1337 3 FreeSans 400 0 0 0 transmission_gate_2/out
flabel metal1 6955 -691 6955 -691 5 FreeSans 400 0 0 0 transmission_gate_2/VDD
flabel metal1 6955 -1797 6955 -1797 1 FreeSans 400 0 0 0 transmission_gate_2/VSS
flabel metal1 -646 960 -646 960 7 FreeSans 400 0 0 0 transmission_gate_10/en_b
flabel metal1 -645 464 -645 464 7 FreeSans 400 0 0 0 transmission_gate_10/in
flabel metal1 -645 153 -645 153 7 FreeSans 400 0 0 0 transmission_gate_10/en
flabel metal1 -2136 463 -2136 463 3 FreeSans 400 0 0 0 transmission_gate_10/out
flabel metal1 -2045 1109 -2045 1109 5 FreeSans 400 0 0 0 transmission_gate_10/VDD
flabel metal1 -2045 3 -2045 3 1 FreeSans 400 0 0 0 transmission_gate_10/VSS
flabel metal1 8354 960 8354 960 7 FreeSans 400 0 0 0 transmission_gate_0/en_b
flabel metal1 8355 464 8355 464 7 FreeSans 400 0 0 0 transmission_gate_0/in
flabel metal1 8355 153 8355 153 7 FreeSans 400 0 0 0 transmission_gate_0/en
flabel metal1 6864 463 6864 463 3 FreeSans 400 0 0 0 transmission_gate_0/out
flabel metal1 6955 1109 6955 1109 5 FreeSans 400 0 0 0 transmission_gate_0/VDD
flabel metal1 6955 3 6955 3 1 FreeSans 400 0 0 0 transmission_gate_0/VSS
flabel metal1 -646 2760 -646 2760 7 FreeSans 400 0 0 0 transmission_gate_9/en_b
flabel metal1 -645 2264 -645 2264 7 FreeSans 400 0 0 0 transmission_gate_9/in
flabel metal1 -645 1953 -645 1953 7 FreeSans 400 0 0 0 transmission_gate_9/en
flabel metal1 -2136 2263 -2136 2263 3 FreeSans 400 0 0 0 transmission_gate_9/out
flabel metal1 -2045 2909 -2045 2909 5 FreeSans 400 0 0 0 transmission_gate_9/VDD
flabel metal1 -2045 1803 -2045 1803 1 FreeSans 400 0 0 0 transmission_gate_9/VSS
flabel metal1 8354 2760 8354 2760 7 FreeSans 400 0 0 0 transmission_gate_1/en_b
flabel metal1 8355 2264 8355 2264 7 FreeSans 400 0 0 0 transmission_gate_1/in
flabel metal1 8355 1953 8355 1953 7 FreeSans 400 0 0 0 transmission_gate_1/en
flabel metal1 6864 2263 6864 2263 3 FreeSans 400 0 0 0 transmission_gate_1/out
flabel metal1 6955 2909 6955 2909 5 FreeSans 400 0 0 0 transmission_gate_1/VDD
flabel metal1 6955 1803 6955 1803 1 FreeSans 400 0 0 0 transmission_gate_1/VSS
flabel metal1 -646 4560 -646 4560 7 FreeSans 400 0 0 0 transmission_gate_8/en_b
flabel metal1 -645 4064 -645 4064 7 FreeSans 400 0 0 0 transmission_gate_8/in
flabel metal1 -645 3753 -645 3753 7 FreeSans 400 0 0 0 transmission_gate_8/en
flabel metal1 -2136 4063 -2136 4063 3 FreeSans 400 0 0 0 transmission_gate_8/out
flabel metal1 -2045 4709 -2045 4709 5 FreeSans 400 0 0 0 transmission_gate_8/VDD
flabel metal1 -2045 3603 -2045 3603 1 FreeSans 400 0 0 0 transmission_gate_8/VSS
flabel metal1 8354 4560 8354 4560 7 FreeSans 400 0 0 0 transmission_gate_3/en_b
flabel metal1 8355 4064 8355 4064 7 FreeSans 400 0 0 0 transmission_gate_3/in
flabel metal1 8355 3753 8355 3753 7 FreeSans 400 0 0 0 transmission_gate_3/en
flabel metal1 6864 4063 6864 4063 3 FreeSans 400 0 0 0 transmission_gate_3/out
flabel metal1 6955 4709 6955 4709 5 FreeSans 400 0 0 0 transmission_gate_3/VDD
flabel metal1 6955 3603 6955 3603 1 FreeSans 400 0 0 0 transmission_gate_3/VSS
flabel metal1 -646 6360 -646 6360 7 FreeSans 400 0 0 0 transmission_gate_7/en_b
flabel metal1 -645 5864 -645 5864 7 FreeSans 400 0 0 0 transmission_gate_7/in
flabel metal1 -645 5553 -645 5553 7 FreeSans 400 0 0 0 transmission_gate_7/en
flabel metal1 -2136 5863 -2136 5863 3 FreeSans 400 0 0 0 transmission_gate_7/out
flabel metal1 -2045 6509 -2045 6509 5 FreeSans 400 0 0 0 transmission_gate_7/VDD
flabel metal1 -2045 5403 -2045 5403 1 FreeSans 400 0 0 0 transmission_gate_7/VSS
flabel metal1 8354 6360 8354 6360 7 FreeSans 400 0 0 0 transmission_gate_4/en_b
flabel metal1 8355 5864 8355 5864 7 FreeSans 400 0 0 0 transmission_gate_4/in
flabel metal1 8355 5553 8355 5553 7 FreeSans 400 0 0 0 transmission_gate_4/en
flabel metal1 6864 5863 6864 5863 3 FreeSans 400 0 0 0 transmission_gate_4/out
flabel metal1 6955 6509 6955 6509 5 FreeSans 400 0 0 0 transmission_gate_4/VDD
flabel metal1 6955 5403 6955 5403 1 FreeSans 400 0 0 0 transmission_gate_4/VSS
flabel metal1 -646 8160 -646 8160 7 FreeSans 400 0 0 0 transmission_gate_6/en_b
flabel metal1 -645 7664 -645 7664 7 FreeSans 400 0 0 0 transmission_gate_6/in
flabel metal1 -645 7353 -645 7353 7 FreeSans 400 0 0 0 transmission_gate_6/en
flabel metal1 -2136 7663 -2136 7663 3 FreeSans 400 0 0 0 transmission_gate_6/out
flabel metal1 -2045 8309 -2045 8309 5 FreeSans 400 0 0 0 transmission_gate_6/VDD
flabel metal1 -2045 7203 -2045 7203 1 FreeSans 400 0 0 0 transmission_gate_6/VSS
flabel metal1 8354 8160 8354 8160 7 FreeSans 400 0 0 0 transmission_gate_5/en_b
flabel metal1 8355 7664 8355 7664 7 FreeSans 400 0 0 0 transmission_gate_5/in
flabel metal1 8355 7353 8355 7353 7 FreeSans 400 0 0 0 transmission_gate_5/en
flabel metal1 6864 7663 6864 7663 3 FreeSans 400 0 0 0 transmission_gate_5/out
flabel metal1 6955 8309 6955 8309 5 FreeSans 400 0 0 0 transmission_gate_5/VDD
flabel metal1 6955 7203 6955 7203 1 FreeSans 400 0 0 0 transmission_gate_5/VSS
<< end >>
