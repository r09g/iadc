magic
tech sky130A
timestamp 1654720150
<< error_p >>
rect -2062 86 -2033 89
rect -1852 86 -1823 89
rect -1642 86 -1613 89
rect -1432 86 -1403 89
rect -1222 86 -1193 89
rect -1012 86 -983 89
rect -802 86 -773 89
rect -592 86 -563 89
rect -382 86 -353 89
rect -172 86 -143 89
rect 38 86 67 89
rect 248 86 277 89
rect 458 86 487 89
rect 668 86 697 89
rect 878 86 907 89
rect 1088 86 1117 89
rect 1298 86 1327 89
rect 1508 86 1537 89
rect 1718 86 1747 89
rect 1928 86 1957 89
rect -2062 69 -2056 86
rect -1852 69 -1846 86
rect -1642 69 -1636 86
rect -1432 69 -1426 86
rect -1222 69 -1216 86
rect -1012 69 -1006 86
rect -802 69 -796 86
rect -592 69 -586 86
rect -382 69 -376 86
rect -172 69 -166 86
rect 38 69 44 86
rect 248 69 254 86
rect 458 69 464 86
rect 668 69 674 86
rect 878 69 884 86
rect 1088 69 1094 86
rect 1298 69 1304 86
rect 1508 69 1514 86
rect 1718 69 1724 86
rect 1928 69 1934 86
rect -2062 66 -2033 69
rect -1852 66 -1823 69
rect -1642 66 -1613 69
rect -1432 66 -1403 69
rect -1222 66 -1193 69
rect -1012 66 -983 69
rect -802 66 -773 69
rect -592 66 -563 69
rect -382 66 -353 69
rect -172 66 -143 69
rect 38 66 67 69
rect 248 66 277 69
rect 458 66 487 69
rect 668 66 697 69
rect 878 66 907 69
rect 1088 66 1117 69
rect 1298 66 1327 69
rect 1508 66 1537 69
rect 1718 66 1747 69
rect 1928 66 1957 69
rect -1957 -69 -1928 -66
rect -1747 -69 -1718 -66
rect -1537 -69 -1508 -66
rect -1327 -69 -1298 -66
rect -1117 -69 -1088 -66
rect -907 -69 -878 -66
rect -697 -69 -668 -66
rect -487 -69 -458 -66
rect -277 -69 -248 -66
rect -67 -69 -38 -66
rect 143 -69 172 -66
rect 353 -69 382 -66
rect 563 -69 592 -66
rect 773 -69 802 -66
rect 983 -69 1012 -66
rect 1193 -69 1222 -66
rect 1403 -69 1432 -66
rect 1613 -69 1642 -66
rect 1823 -69 1852 -66
rect 2033 -69 2062 -66
rect -1957 -86 -1951 -69
rect -1747 -86 -1741 -69
rect -1537 -86 -1531 -69
rect -1327 -86 -1321 -69
rect -1117 -86 -1111 -69
rect -907 -86 -901 -69
rect -697 -86 -691 -69
rect -487 -86 -481 -69
rect -277 -86 -271 -69
rect -67 -86 -61 -69
rect 143 -86 149 -69
rect 353 -86 359 -69
rect 563 -86 569 -69
rect 773 -86 779 -69
rect 983 -86 989 -69
rect 1193 -86 1199 -69
rect 1403 -86 1409 -69
rect 1613 -86 1619 -69
rect 1823 -86 1829 -69
rect 2033 -86 2039 -69
rect -1957 -89 -1928 -86
rect -1747 -89 -1718 -86
rect -1537 -89 -1508 -86
rect -1327 -89 -1298 -86
rect -1117 -89 -1088 -86
rect -907 -89 -878 -86
rect -697 -89 -668 -86
rect -487 -89 -458 -86
rect -277 -89 -248 -86
rect -67 -89 -38 -86
rect 143 -89 172 -86
rect 353 -89 382 -86
rect 563 -89 592 -86
rect 773 -89 802 -86
rect 983 -89 1012 -86
rect 1193 -89 1222 -86
rect 1403 -89 1432 -86
rect 1613 -89 1642 -86
rect 1823 -89 1852 -86
rect 2033 -89 2062 -86
<< nmos >>
rect -2160 -50 -2145 50
rect -2055 -50 -2040 50
rect -1950 -50 -1935 50
rect -1845 -50 -1830 50
rect -1740 -50 -1725 50
rect -1635 -50 -1620 50
rect -1530 -50 -1515 50
rect -1425 -50 -1410 50
rect -1320 -50 -1305 50
rect -1215 -50 -1200 50
rect -1110 -50 -1095 50
rect -1005 -50 -990 50
rect -900 -50 -885 50
rect -795 -50 -780 50
rect -690 -50 -675 50
rect -585 -50 -570 50
rect -480 -50 -465 50
rect -375 -50 -360 50
rect -270 -50 -255 50
rect -165 -50 -150 50
rect -60 -50 -45 50
rect 45 -50 60 50
rect 150 -50 165 50
rect 255 -50 270 50
rect 360 -50 375 50
rect 465 -50 480 50
rect 570 -50 585 50
rect 675 -50 690 50
rect 780 -50 795 50
rect 885 -50 900 50
rect 990 -50 1005 50
rect 1095 -50 1110 50
rect 1200 -50 1215 50
rect 1305 -50 1320 50
rect 1410 -50 1425 50
rect 1515 -50 1530 50
rect 1620 -50 1635 50
rect 1725 -50 1740 50
rect 1830 -50 1845 50
rect 1935 -50 1950 50
rect 2040 -50 2055 50
rect 2145 -50 2160 50
<< ndiff >>
rect -2191 44 -2160 50
rect -2191 -44 -2185 44
rect -2168 -44 -2160 44
rect -2191 -50 -2160 -44
rect -2145 44 -2114 50
rect -2145 -44 -2137 44
rect -2120 -44 -2114 44
rect -2145 -50 -2114 -44
rect -2086 44 -2055 50
rect -2086 -44 -2080 44
rect -2063 -44 -2055 44
rect -2086 -50 -2055 -44
rect -2040 44 -2009 50
rect -2040 -44 -2032 44
rect -2015 -44 -2009 44
rect -2040 -50 -2009 -44
rect -1981 44 -1950 50
rect -1981 -44 -1975 44
rect -1958 -44 -1950 44
rect -1981 -50 -1950 -44
rect -1935 44 -1904 50
rect -1935 -44 -1927 44
rect -1910 -44 -1904 44
rect -1935 -50 -1904 -44
rect -1876 44 -1845 50
rect -1876 -44 -1870 44
rect -1853 -44 -1845 44
rect -1876 -50 -1845 -44
rect -1830 44 -1799 50
rect -1830 -44 -1822 44
rect -1805 -44 -1799 44
rect -1830 -50 -1799 -44
rect -1771 44 -1740 50
rect -1771 -44 -1765 44
rect -1748 -44 -1740 44
rect -1771 -50 -1740 -44
rect -1725 44 -1694 50
rect -1725 -44 -1717 44
rect -1700 -44 -1694 44
rect -1725 -50 -1694 -44
rect -1666 44 -1635 50
rect -1666 -44 -1660 44
rect -1643 -44 -1635 44
rect -1666 -50 -1635 -44
rect -1620 44 -1589 50
rect -1620 -44 -1612 44
rect -1595 -44 -1589 44
rect -1620 -50 -1589 -44
rect -1561 44 -1530 50
rect -1561 -44 -1555 44
rect -1538 -44 -1530 44
rect -1561 -50 -1530 -44
rect -1515 44 -1484 50
rect -1515 -44 -1507 44
rect -1490 -44 -1484 44
rect -1515 -50 -1484 -44
rect -1456 44 -1425 50
rect -1456 -44 -1450 44
rect -1433 -44 -1425 44
rect -1456 -50 -1425 -44
rect -1410 44 -1379 50
rect -1410 -44 -1402 44
rect -1385 -44 -1379 44
rect -1410 -50 -1379 -44
rect -1351 44 -1320 50
rect -1351 -44 -1345 44
rect -1328 -44 -1320 44
rect -1351 -50 -1320 -44
rect -1305 44 -1274 50
rect -1305 -44 -1297 44
rect -1280 -44 -1274 44
rect -1305 -50 -1274 -44
rect -1246 44 -1215 50
rect -1246 -44 -1240 44
rect -1223 -44 -1215 44
rect -1246 -50 -1215 -44
rect -1200 44 -1169 50
rect -1200 -44 -1192 44
rect -1175 -44 -1169 44
rect -1200 -50 -1169 -44
rect -1141 44 -1110 50
rect -1141 -44 -1135 44
rect -1118 -44 -1110 44
rect -1141 -50 -1110 -44
rect -1095 44 -1064 50
rect -1095 -44 -1087 44
rect -1070 -44 -1064 44
rect -1095 -50 -1064 -44
rect -1036 44 -1005 50
rect -1036 -44 -1030 44
rect -1013 -44 -1005 44
rect -1036 -50 -1005 -44
rect -990 44 -959 50
rect -990 -44 -982 44
rect -965 -44 -959 44
rect -990 -50 -959 -44
rect -931 44 -900 50
rect -931 -44 -925 44
rect -908 -44 -900 44
rect -931 -50 -900 -44
rect -885 44 -854 50
rect -885 -44 -877 44
rect -860 -44 -854 44
rect -885 -50 -854 -44
rect -826 44 -795 50
rect -826 -44 -820 44
rect -803 -44 -795 44
rect -826 -50 -795 -44
rect -780 44 -749 50
rect -780 -44 -772 44
rect -755 -44 -749 44
rect -780 -50 -749 -44
rect -721 44 -690 50
rect -721 -44 -715 44
rect -698 -44 -690 44
rect -721 -50 -690 -44
rect -675 44 -644 50
rect -675 -44 -667 44
rect -650 -44 -644 44
rect -675 -50 -644 -44
rect -616 44 -585 50
rect -616 -44 -610 44
rect -593 -44 -585 44
rect -616 -50 -585 -44
rect -570 44 -539 50
rect -570 -44 -562 44
rect -545 -44 -539 44
rect -570 -50 -539 -44
rect -511 44 -480 50
rect -511 -44 -505 44
rect -488 -44 -480 44
rect -511 -50 -480 -44
rect -465 44 -434 50
rect -465 -44 -457 44
rect -440 -44 -434 44
rect -465 -50 -434 -44
rect -406 44 -375 50
rect -406 -44 -400 44
rect -383 -44 -375 44
rect -406 -50 -375 -44
rect -360 44 -329 50
rect -360 -44 -352 44
rect -335 -44 -329 44
rect -360 -50 -329 -44
rect -301 44 -270 50
rect -301 -44 -295 44
rect -278 -44 -270 44
rect -301 -50 -270 -44
rect -255 44 -224 50
rect -255 -44 -247 44
rect -230 -44 -224 44
rect -255 -50 -224 -44
rect -196 44 -165 50
rect -196 -44 -190 44
rect -173 -44 -165 44
rect -196 -50 -165 -44
rect -150 44 -119 50
rect -150 -44 -142 44
rect -125 -44 -119 44
rect -150 -50 -119 -44
rect -91 44 -60 50
rect -91 -44 -85 44
rect -68 -44 -60 44
rect -91 -50 -60 -44
rect -45 44 -14 50
rect -45 -44 -37 44
rect -20 -44 -14 44
rect -45 -50 -14 -44
rect 14 44 45 50
rect 14 -44 20 44
rect 37 -44 45 44
rect 14 -50 45 -44
rect 60 44 91 50
rect 60 -44 68 44
rect 85 -44 91 44
rect 60 -50 91 -44
rect 119 44 150 50
rect 119 -44 125 44
rect 142 -44 150 44
rect 119 -50 150 -44
rect 165 44 196 50
rect 165 -44 173 44
rect 190 -44 196 44
rect 165 -50 196 -44
rect 224 44 255 50
rect 224 -44 230 44
rect 247 -44 255 44
rect 224 -50 255 -44
rect 270 44 301 50
rect 270 -44 278 44
rect 295 -44 301 44
rect 270 -50 301 -44
rect 329 44 360 50
rect 329 -44 335 44
rect 352 -44 360 44
rect 329 -50 360 -44
rect 375 44 406 50
rect 375 -44 383 44
rect 400 -44 406 44
rect 375 -50 406 -44
rect 434 44 465 50
rect 434 -44 440 44
rect 457 -44 465 44
rect 434 -50 465 -44
rect 480 44 511 50
rect 480 -44 488 44
rect 505 -44 511 44
rect 480 -50 511 -44
rect 539 44 570 50
rect 539 -44 545 44
rect 562 -44 570 44
rect 539 -50 570 -44
rect 585 44 616 50
rect 585 -44 593 44
rect 610 -44 616 44
rect 585 -50 616 -44
rect 644 44 675 50
rect 644 -44 650 44
rect 667 -44 675 44
rect 644 -50 675 -44
rect 690 44 721 50
rect 690 -44 698 44
rect 715 -44 721 44
rect 690 -50 721 -44
rect 749 44 780 50
rect 749 -44 755 44
rect 772 -44 780 44
rect 749 -50 780 -44
rect 795 44 826 50
rect 795 -44 803 44
rect 820 -44 826 44
rect 795 -50 826 -44
rect 854 44 885 50
rect 854 -44 860 44
rect 877 -44 885 44
rect 854 -50 885 -44
rect 900 44 931 50
rect 900 -44 908 44
rect 925 -44 931 44
rect 900 -50 931 -44
rect 959 44 990 50
rect 959 -44 965 44
rect 982 -44 990 44
rect 959 -50 990 -44
rect 1005 44 1036 50
rect 1005 -44 1013 44
rect 1030 -44 1036 44
rect 1005 -50 1036 -44
rect 1064 44 1095 50
rect 1064 -44 1070 44
rect 1087 -44 1095 44
rect 1064 -50 1095 -44
rect 1110 44 1141 50
rect 1110 -44 1118 44
rect 1135 -44 1141 44
rect 1110 -50 1141 -44
rect 1169 44 1200 50
rect 1169 -44 1175 44
rect 1192 -44 1200 44
rect 1169 -50 1200 -44
rect 1215 44 1246 50
rect 1215 -44 1223 44
rect 1240 -44 1246 44
rect 1215 -50 1246 -44
rect 1274 44 1305 50
rect 1274 -44 1280 44
rect 1297 -44 1305 44
rect 1274 -50 1305 -44
rect 1320 44 1351 50
rect 1320 -44 1328 44
rect 1345 -44 1351 44
rect 1320 -50 1351 -44
rect 1379 44 1410 50
rect 1379 -44 1385 44
rect 1402 -44 1410 44
rect 1379 -50 1410 -44
rect 1425 44 1456 50
rect 1425 -44 1433 44
rect 1450 -44 1456 44
rect 1425 -50 1456 -44
rect 1484 44 1515 50
rect 1484 -44 1490 44
rect 1507 -44 1515 44
rect 1484 -50 1515 -44
rect 1530 44 1561 50
rect 1530 -44 1538 44
rect 1555 -44 1561 44
rect 1530 -50 1561 -44
rect 1589 44 1620 50
rect 1589 -44 1595 44
rect 1612 -44 1620 44
rect 1589 -50 1620 -44
rect 1635 44 1666 50
rect 1635 -44 1643 44
rect 1660 -44 1666 44
rect 1635 -50 1666 -44
rect 1694 44 1725 50
rect 1694 -44 1700 44
rect 1717 -44 1725 44
rect 1694 -50 1725 -44
rect 1740 44 1771 50
rect 1740 -44 1748 44
rect 1765 -44 1771 44
rect 1740 -50 1771 -44
rect 1799 44 1830 50
rect 1799 -44 1805 44
rect 1822 -44 1830 44
rect 1799 -50 1830 -44
rect 1845 44 1876 50
rect 1845 -44 1853 44
rect 1870 -44 1876 44
rect 1845 -50 1876 -44
rect 1904 44 1935 50
rect 1904 -44 1910 44
rect 1927 -44 1935 44
rect 1904 -50 1935 -44
rect 1950 44 1981 50
rect 1950 -44 1958 44
rect 1975 -44 1981 44
rect 1950 -50 1981 -44
rect 2009 44 2040 50
rect 2009 -44 2015 44
rect 2032 -44 2040 44
rect 2009 -50 2040 -44
rect 2055 44 2086 50
rect 2055 -44 2063 44
rect 2080 -44 2086 44
rect 2055 -50 2086 -44
rect 2114 44 2145 50
rect 2114 -44 2120 44
rect 2137 -44 2145 44
rect 2114 -50 2145 -44
rect 2160 44 2191 50
rect 2160 -44 2168 44
rect 2185 -44 2191 44
rect 2160 -50 2191 -44
<< ndiffc >>
rect -2185 -44 -2168 44
rect -2137 -44 -2120 44
rect -2080 -44 -2063 44
rect -2032 -44 -2015 44
rect -1975 -44 -1958 44
rect -1927 -44 -1910 44
rect -1870 -44 -1853 44
rect -1822 -44 -1805 44
rect -1765 -44 -1748 44
rect -1717 -44 -1700 44
rect -1660 -44 -1643 44
rect -1612 -44 -1595 44
rect -1555 -44 -1538 44
rect -1507 -44 -1490 44
rect -1450 -44 -1433 44
rect -1402 -44 -1385 44
rect -1345 -44 -1328 44
rect -1297 -44 -1280 44
rect -1240 -44 -1223 44
rect -1192 -44 -1175 44
rect -1135 -44 -1118 44
rect -1087 -44 -1070 44
rect -1030 -44 -1013 44
rect -982 -44 -965 44
rect -925 -44 -908 44
rect -877 -44 -860 44
rect -820 -44 -803 44
rect -772 -44 -755 44
rect -715 -44 -698 44
rect -667 -44 -650 44
rect -610 -44 -593 44
rect -562 -44 -545 44
rect -505 -44 -488 44
rect -457 -44 -440 44
rect -400 -44 -383 44
rect -352 -44 -335 44
rect -295 -44 -278 44
rect -247 -44 -230 44
rect -190 -44 -173 44
rect -142 -44 -125 44
rect -85 -44 -68 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 68 -44 85 44
rect 125 -44 142 44
rect 173 -44 190 44
rect 230 -44 247 44
rect 278 -44 295 44
rect 335 -44 352 44
rect 383 -44 400 44
rect 440 -44 457 44
rect 488 -44 505 44
rect 545 -44 562 44
rect 593 -44 610 44
rect 650 -44 667 44
rect 698 -44 715 44
rect 755 -44 772 44
rect 803 -44 820 44
rect 860 -44 877 44
rect 908 -44 925 44
rect 965 -44 982 44
rect 1013 -44 1030 44
rect 1070 -44 1087 44
rect 1118 -44 1135 44
rect 1175 -44 1192 44
rect 1223 -44 1240 44
rect 1280 -44 1297 44
rect 1328 -44 1345 44
rect 1385 -44 1402 44
rect 1433 -44 1450 44
rect 1490 -44 1507 44
rect 1538 -44 1555 44
rect 1595 -44 1612 44
rect 1643 -44 1660 44
rect 1700 -44 1717 44
rect 1748 -44 1765 44
rect 1805 -44 1822 44
rect 1853 -44 1870 44
rect 1910 -44 1927 44
rect 1958 -44 1975 44
rect 2015 -44 2032 44
rect 2063 -44 2080 44
rect 2120 -44 2137 44
rect 2168 -44 2185 44
<< poly >>
rect -2064 86 -2031 94
rect -2064 69 -2056 86
rect -2039 69 -2031 86
rect -2160 50 -2145 63
rect -2064 61 -2031 69
rect -1854 86 -1821 94
rect -1854 69 -1846 86
rect -1829 69 -1821 86
rect -2055 50 -2040 61
rect -1950 50 -1935 63
rect -1854 61 -1821 69
rect -1644 86 -1611 94
rect -1644 69 -1636 86
rect -1619 69 -1611 86
rect -1845 50 -1830 61
rect -1740 50 -1725 63
rect -1644 61 -1611 69
rect -1434 86 -1401 94
rect -1434 69 -1426 86
rect -1409 69 -1401 86
rect -1635 50 -1620 61
rect -1530 50 -1515 63
rect -1434 61 -1401 69
rect -1224 86 -1191 94
rect -1224 69 -1216 86
rect -1199 69 -1191 86
rect -1425 50 -1410 61
rect -1320 50 -1305 63
rect -1224 61 -1191 69
rect -1014 86 -981 94
rect -1014 69 -1006 86
rect -989 69 -981 86
rect -1215 50 -1200 61
rect -1110 50 -1095 63
rect -1014 61 -981 69
rect -804 86 -771 94
rect -804 69 -796 86
rect -779 69 -771 86
rect -1005 50 -990 61
rect -900 50 -885 63
rect -804 61 -771 69
rect -594 86 -561 94
rect -594 69 -586 86
rect -569 69 -561 86
rect -795 50 -780 61
rect -690 50 -675 63
rect -594 61 -561 69
rect -384 86 -351 94
rect -384 69 -376 86
rect -359 69 -351 86
rect -585 50 -570 61
rect -480 50 -465 63
rect -384 61 -351 69
rect -174 86 -141 94
rect -174 69 -166 86
rect -149 69 -141 86
rect -375 50 -360 61
rect -270 50 -255 63
rect -174 61 -141 69
rect 36 86 69 94
rect 36 69 44 86
rect 61 69 69 86
rect -165 50 -150 61
rect -60 50 -45 63
rect 36 61 69 69
rect 246 86 279 94
rect 246 69 254 86
rect 271 69 279 86
rect 45 50 60 61
rect 150 50 165 63
rect 246 61 279 69
rect 456 86 489 94
rect 456 69 464 86
rect 481 69 489 86
rect 255 50 270 61
rect 360 50 375 63
rect 456 61 489 69
rect 666 86 699 94
rect 666 69 674 86
rect 691 69 699 86
rect 465 50 480 61
rect 570 50 585 63
rect 666 61 699 69
rect 876 86 909 94
rect 876 69 884 86
rect 901 69 909 86
rect 675 50 690 61
rect 780 50 795 63
rect 876 61 909 69
rect 1086 86 1119 94
rect 1086 69 1094 86
rect 1111 69 1119 86
rect 885 50 900 61
rect 990 50 1005 63
rect 1086 61 1119 69
rect 1296 86 1329 94
rect 1296 69 1304 86
rect 1321 69 1329 86
rect 1095 50 1110 61
rect 1200 50 1215 63
rect 1296 61 1329 69
rect 1506 86 1539 94
rect 1506 69 1514 86
rect 1531 69 1539 86
rect 1305 50 1320 61
rect 1410 50 1425 63
rect 1506 61 1539 69
rect 1716 86 1749 94
rect 1716 69 1724 86
rect 1741 69 1749 86
rect 1515 50 1530 61
rect 1620 50 1635 63
rect 1716 61 1749 69
rect 1926 86 1959 94
rect 1926 69 1934 86
rect 1951 69 1959 86
rect 1725 50 1740 61
rect 1830 50 1845 63
rect 1926 61 1959 69
rect 2136 86 2169 94
rect 2136 69 2144 86
rect 2161 69 2169 86
rect 1935 50 1950 61
rect 2040 50 2055 63
rect 2136 61 2169 69
rect 2145 50 2160 61
rect -2160 -61 -2145 -50
rect -2169 -69 -2136 -61
rect -2055 -63 -2040 -50
rect -1950 -61 -1935 -50
rect -2169 -86 -2161 -69
rect -2144 -86 -2136 -69
rect -2169 -94 -2136 -86
rect -1959 -69 -1926 -61
rect -1845 -63 -1830 -50
rect -1740 -61 -1725 -50
rect -1959 -86 -1951 -69
rect -1934 -86 -1926 -69
rect -1959 -94 -1926 -86
rect -1749 -69 -1716 -61
rect -1635 -63 -1620 -50
rect -1530 -61 -1515 -50
rect -1749 -86 -1741 -69
rect -1724 -86 -1716 -69
rect -1749 -94 -1716 -86
rect -1539 -69 -1506 -61
rect -1425 -63 -1410 -50
rect -1320 -61 -1305 -50
rect -1539 -86 -1531 -69
rect -1514 -86 -1506 -69
rect -1539 -94 -1506 -86
rect -1329 -69 -1296 -61
rect -1215 -63 -1200 -50
rect -1110 -61 -1095 -50
rect -1329 -86 -1321 -69
rect -1304 -86 -1296 -69
rect -1329 -94 -1296 -86
rect -1119 -69 -1086 -61
rect -1005 -63 -990 -50
rect -900 -61 -885 -50
rect -1119 -86 -1111 -69
rect -1094 -86 -1086 -69
rect -1119 -94 -1086 -86
rect -909 -69 -876 -61
rect -795 -63 -780 -50
rect -690 -61 -675 -50
rect -909 -86 -901 -69
rect -884 -86 -876 -69
rect -909 -94 -876 -86
rect -699 -69 -666 -61
rect -585 -63 -570 -50
rect -480 -61 -465 -50
rect -699 -86 -691 -69
rect -674 -86 -666 -69
rect -699 -94 -666 -86
rect -489 -69 -456 -61
rect -375 -63 -360 -50
rect -270 -61 -255 -50
rect -489 -86 -481 -69
rect -464 -86 -456 -69
rect -489 -94 -456 -86
rect -279 -69 -246 -61
rect -165 -63 -150 -50
rect -60 -61 -45 -50
rect -279 -86 -271 -69
rect -254 -86 -246 -69
rect -279 -94 -246 -86
rect -69 -69 -36 -61
rect 45 -63 60 -50
rect 150 -61 165 -50
rect -69 -86 -61 -69
rect -44 -86 -36 -69
rect -69 -94 -36 -86
rect 141 -69 174 -61
rect 255 -63 270 -50
rect 360 -61 375 -50
rect 141 -86 149 -69
rect 166 -86 174 -69
rect 141 -94 174 -86
rect 351 -69 384 -61
rect 465 -63 480 -50
rect 570 -61 585 -50
rect 351 -86 359 -69
rect 376 -86 384 -69
rect 351 -94 384 -86
rect 561 -69 594 -61
rect 675 -63 690 -50
rect 780 -61 795 -50
rect 561 -86 569 -69
rect 586 -86 594 -69
rect 561 -94 594 -86
rect 771 -69 804 -61
rect 885 -63 900 -50
rect 990 -61 1005 -50
rect 771 -86 779 -69
rect 796 -86 804 -69
rect 771 -94 804 -86
rect 981 -69 1014 -61
rect 1095 -63 1110 -50
rect 1200 -61 1215 -50
rect 981 -86 989 -69
rect 1006 -86 1014 -69
rect 981 -94 1014 -86
rect 1191 -69 1224 -61
rect 1305 -63 1320 -50
rect 1410 -61 1425 -50
rect 1191 -86 1199 -69
rect 1216 -86 1224 -69
rect 1191 -94 1224 -86
rect 1401 -69 1434 -61
rect 1515 -63 1530 -50
rect 1620 -61 1635 -50
rect 1401 -86 1409 -69
rect 1426 -86 1434 -69
rect 1401 -94 1434 -86
rect 1611 -69 1644 -61
rect 1725 -63 1740 -50
rect 1830 -61 1845 -50
rect 1611 -86 1619 -69
rect 1636 -86 1644 -69
rect 1611 -94 1644 -86
rect 1821 -69 1854 -61
rect 1935 -63 1950 -50
rect 2040 -61 2055 -50
rect 1821 -86 1829 -69
rect 1846 -86 1854 -69
rect 1821 -94 1854 -86
rect 2031 -69 2064 -61
rect 2145 -63 2160 -50
rect 2031 -86 2039 -69
rect 2056 -86 2064 -69
rect 2031 -94 2064 -86
<< polycont >>
rect -2056 69 -2039 86
rect -1846 69 -1829 86
rect -1636 69 -1619 86
rect -1426 69 -1409 86
rect -1216 69 -1199 86
rect -1006 69 -989 86
rect -796 69 -779 86
rect -586 69 -569 86
rect -376 69 -359 86
rect -166 69 -149 86
rect 44 69 61 86
rect 254 69 271 86
rect 464 69 481 86
rect 674 69 691 86
rect 884 69 901 86
rect 1094 69 1111 86
rect 1304 69 1321 86
rect 1514 69 1531 86
rect 1724 69 1741 86
rect 1934 69 1951 86
rect 2144 69 2161 86
rect -2161 -86 -2144 -69
rect -1951 -86 -1934 -69
rect -1741 -86 -1724 -69
rect -1531 -86 -1514 -69
rect -1321 -86 -1304 -69
rect -1111 -86 -1094 -69
rect -901 -86 -884 -69
rect -691 -86 -674 -69
rect -481 -86 -464 -69
rect -271 -86 -254 -69
rect -61 -86 -44 -69
rect 149 -86 166 -69
rect 359 -86 376 -69
rect 569 -86 586 -69
rect 779 -86 796 -69
rect 989 -86 1006 -69
rect 1199 -86 1216 -69
rect 1409 -86 1426 -69
rect 1619 -86 1636 -69
rect 1829 -86 1846 -69
rect 2039 -86 2056 -69
<< locali >>
rect -2064 69 -2056 86
rect -2039 69 -2031 86
rect -1854 69 -1846 86
rect -1829 69 -1821 86
rect -1644 69 -1636 86
rect -1619 69 -1611 86
rect -1434 69 -1426 86
rect -1409 69 -1401 86
rect -1224 69 -1216 86
rect -1199 69 -1191 86
rect -1014 69 -1006 86
rect -989 69 -981 86
rect -804 69 -796 86
rect -779 69 -771 86
rect -594 69 -586 86
rect -569 69 -561 86
rect -384 69 -376 86
rect -359 69 -351 86
rect -174 69 -166 86
rect -149 69 -141 86
rect 36 69 44 86
rect 61 69 69 86
rect 246 69 254 86
rect 271 69 279 86
rect 456 69 464 86
rect 481 69 489 86
rect 666 69 674 86
rect 691 69 699 86
rect 876 69 884 86
rect 901 69 909 86
rect 1086 69 1094 86
rect 1111 69 1119 86
rect 1296 69 1304 86
rect 1321 69 1329 86
rect 1506 69 1514 86
rect 1531 69 1539 86
rect 1716 69 1724 86
rect 1741 69 1749 86
rect 1926 69 1934 86
rect 1951 69 1959 86
rect 2120 69 2144 86
rect 2161 69 2185 86
rect -2185 44 -2168 52
rect -2185 -69 -2168 -44
rect -2137 44 -2120 52
rect -2137 -69 -2120 -44
rect -2080 44 -2063 52
rect -2080 -52 -2063 -44
rect -2032 44 -2015 52
rect -2032 -52 -2015 -44
rect -1975 44 -1958 52
rect -1975 -52 -1958 -44
rect -1927 44 -1910 52
rect -1927 -52 -1910 -44
rect -1870 44 -1853 52
rect -1870 -52 -1853 -44
rect -1822 44 -1805 52
rect -1822 -52 -1805 -44
rect -1765 44 -1748 52
rect -1765 -52 -1748 -44
rect -1717 44 -1700 52
rect -1717 -52 -1700 -44
rect -1660 44 -1643 52
rect -1660 -52 -1643 -44
rect -1612 44 -1595 52
rect -1612 -52 -1595 -44
rect -1555 44 -1538 52
rect -1555 -52 -1538 -44
rect -1507 44 -1490 52
rect -1507 -52 -1490 -44
rect -1450 44 -1433 52
rect -1450 -52 -1433 -44
rect -1402 44 -1385 52
rect -1402 -52 -1385 -44
rect -1345 44 -1328 52
rect -1345 -52 -1328 -44
rect -1297 44 -1280 52
rect -1297 -52 -1280 -44
rect -1240 44 -1223 52
rect -1240 -52 -1223 -44
rect -1192 44 -1175 52
rect -1192 -52 -1175 -44
rect -1135 44 -1118 52
rect -1135 -52 -1118 -44
rect -1087 44 -1070 52
rect -1087 -52 -1070 -44
rect -1030 44 -1013 52
rect -1030 -52 -1013 -44
rect -982 44 -965 52
rect -982 -52 -965 -44
rect -925 44 -908 52
rect -925 -52 -908 -44
rect -877 44 -860 52
rect -877 -52 -860 -44
rect -820 44 -803 52
rect -820 -52 -803 -44
rect -772 44 -755 52
rect -772 -52 -755 -44
rect -715 44 -698 52
rect -715 -52 -698 -44
rect -667 44 -650 52
rect -667 -52 -650 -44
rect -610 44 -593 52
rect -610 -52 -593 -44
rect -562 44 -545 52
rect -562 -52 -545 -44
rect -505 44 -488 52
rect -505 -52 -488 -44
rect -457 44 -440 52
rect -457 -52 -440 -44
rect -400 44 -383 52
rect -400 -52 -383 -44
rect -352 44 -335 52
rect -352 -52 -335 -44
rect -295 44 -278 52
rect -295 -52 -278 -44
rect -247 44 -230 52
rect -247 -52 -230 -44
rect -190 44 -173 52
rect -190 -52 -173 -44
rect -142 44 -125 52
rect -142 -52 -125 -44
rect -85 44 -68 52
rect -85 -52 -68 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 68 44 85 52
rect 68 -52 85 -44
rect 125 44 142 52
rect 125 -52 142 -44
rect 173 44 190 52
rect 173 -52 190 -44
rect 230 44 247 52
rect 230 -52 247 -44
rect 278 44 295 52
rect 278 -52 295 -44
rect 335 44 352 52
rect 335 -52 352 -44
rect 383 44 400 52
rect 383 -52 400 -44
rect 440 44 457 52
rect 440 -52 457 -44
rect 488 44 505 52
rect 488 -52 505 -44
rect 545 44 562 52
rect 545 -52 562 -44
rect 593 44 610 52
rect 593 -52 610 -44
rect 650 44 667 52
rect 650 -52 667 -44
rect 698 44 715 52
rect 698 -52 715 -44
rect 755 44 772 52
rect 755 -52 772 -44
rect 803 44 820 52
rect 803 -52 820 -44
rect 860 44 877 52
rect 860 -52 877 -44
rect 908 44 925 52
rect 908 -52 925 -44
rect 965 44 982 52
rect 965 -52 982 -44
rect 1013 44 1030 52
rect 1013 -52 1030 -44
rect 1070 44 1087 52
rect 1070 -52 1087 -44
rect 1118 44 1135 52
rect 1118 -52 1135 -44
rect 1175 44 1192 52
rect 1175 -52 1192 -44
rect 1223 44 1240 52
rect 1223 -52 1240 -44
rect 1280 44 1297 52
rect 1280 -52 1297 -44
rect 1328 44 1345 52
rect 1328 -52 1345 -44
rect 1385 44 1402 52
rect 1385 -52 1402 -44
rect 1433 44 1450 52
rect 1433 -52 1450 -44
rect 1490 44 1507 52
rect 1490 -52 1507 -44
rect 1538 44 1555 52
rect 1538 -52 1555 -44
rect 1595 44 1612 52
rect 1595 -52 1612 -44
rect 1643 44 1660 52
rect 1643 -52 1660 -44
rect 1700 44 1717 52
rect 1700 -52 1717 -44
rect 1748 44 1765 52
rect 1748 -52 1765 -44
rect 1805 44 1822 52
rect 1805 -52 1822 -44
rect 1853 44 1870 52
rect 1853 -52 1870 -44
rect 1910 44 1927 52
rect 1910 -52 1927 -44
rect 1958 44 1975 52
rect 1958 -52 1975 -44
rect 2015 44 2032 52
rect 2015 -52 2032 -44
rect 2063 44 2080 52
rect 2063 -52 2080 -44
rect 2120 44 2137 69
rect 2120 -52 2137 -44
rect 2168 44 2185 69
rect 2168 -52 2185 -44
rect -2185 -86 -2161 -69
rect -2144 -86 -2120 -69
rect -1959 -86 -1951 -69
rect -1934 -86 -1926 -69
rect -1749 -86 -1741 -69
rect -1724 -86 -1716 -69
rect -1539 -86 -1531 -69
rect -1514 -86 -1506 -69
rect -1329 -86 -1321 -69
rect -1304 -86 -1296 -69
rect -1119 -86 -1111 -69
rect -1094 -86 -1086 -69
rect -909 -86 -901 -69
rect -884 -86 -876 -69
rect -699 -86 -691 -69
rect -674 -86 -666 -69
rect -489 -86 -481 -69
rect -464 -86 -456 -69
rect -279 -86 -271 -69
rect -254 -86 -246 -69
rect -69 -86 -61 -69
rect -44 -86 -36 -69
rect 141 -86 149 -69
rect 166 -86 174 -69
rect 351 -86 359 -69
rect 376 -86 384 -69
rect 561 -86 569 -69
rect 586 -86 594 -69
rect 771 -86 779 -69
rect 796 -86 804 -69
rect 981 -86 989 -69
rect 1006 -86 1014 -69
rect 1191 -86 1199 -69
rect 1216 -86 1224 -69
rect 1401 -86 1409 -69
rect 1426 -86 1434 -69
rect 1611 -86 1619 -69
rect 1636 -86 1644 -69
rect 1821 -86 1829 -69
rect 1846 -86 1854 -69
rect 2031 -86 2039 -69
rect 2056 -86 2064 -69
<< viali >>
rect -2056 69 -2039 86
rect -1846 69 -1829 86
rect -1636 69 -1619 86
rect -1426 69 -1409 86
rect -1216 69 -1199 86
rect -1006 69 -989 86
rect -796 69 -779 86
rect -586 69 -569 86
rect -376 69 -359 86
rect -166 69 -149 86
rect 44 69 61 86
rect 254 69 271 86
rect 464 69 481 86
rect 674 69 691 86
rect 884 69 901 86
rect 1094 69 1111 86
rect 1304 69 1321 86
rect 1514 69 1531 86
rect 1724 69 1741 86
rect 1934 69 1951 86
rect -2080 27 -2063 44
rect -2032 -44 -2015 -27
rect -1975 27 -1958 44
rect -1927 -44 -1910 -27
rect -1870 27 -1853 44
rect -1822 -44 -1805 -27
rect -1765 27 -1748 44
rect -1717 -44 -1700 -27
rect -1660 27 -1643 44
rect -1612 -44 -1595 -27
rect -1555 27 -1538 44
rect -1507 -44 -1490 -27
rect -1450 27 -1433 44
rect -1402 -44 -1385 -27
rect -1345 27 -1328 44
rect -1297 -44 -1280 -27
rect -1240 27 -1223 44
rect -1192 -44 -1175 -27
rect -1135 27 -1118 44
rect -1087 -44 -1070 -27
rect -1030 27 -1013 44
rect -982 -44 -965 -27
rect -925 27 -908 44
rect -877 -44 -860 -27
rect -820 27 -803 44
rect -772 -44 -755 -27
rect -715 27 -698 44
rect -667 -44 -650 -27
rect -610 27 -593 44
rect -562 -44 -545 -27
rect -505 27 -488 44
rect -457 -44 -440 -27
rect -400 27 -383 44
rect -352 -44 -335 -27
rect -295 27 -278 44
rect -247 -44 -230 -27
rect -190 27 -173 44
rect -142 -44 -125 -27
rect -85 27 -68 44
rect -37 -44 -20 -27
rect 20 27 37 44
rect 68 -44 85 -27
rect 125 27 142 44
rect 173 -44 190 -27
rect 230 27 247 44
rect 278 -44 295 -27
rect 335 27 352 44
rect 383 -44 400 -27
rect 440 27 457 44
rect 488 -44 505 -27
rect 545 27 562 44
rect 593 -44 610 -27
rect 650 27 667 44
rect 698 -44 715 -27
rect 755 27 772 44
rect 803 -44 820 -27
rect 860 27 877 44
rect 908 -44 925 -27
rect 965 27 982 44
rect 1013 -44 1030 -27
rect 1070 27 1087 44
rect 1118 -44 1135 -27
rect 1175 27 1192 44
rect 1223 -44 1240 -27
rect 1280 27 1297 44
rect 1328 -44 1345 -27
rect 1385 27 1402 44
rect 1433 -44 1450 -27
rect 1490 27 1507 44
rect 1538 -44 1555 -27
rect 1595 27 1612 44
rect 1643 -44 1660 -27
rect 1700 27 1717 44
rect 1748 -44 1765 -27
rect 1805 27 1822 44
rect 1853 -44 1870 -27
rect 1910 27 1927 44
rect 1958 -44 1975 -27
rect 2015 27 2032 44
rect 2063 -44 2080 -27
rect -1951 -86 -1934 -69
rect -1741 -86 -1724 -69
rect -1531 -86 -1514 -69
rect -1321 -86 -1304 -69
rect -1111 -86 -1094 -69
rect -901 -86 -884 -69
rect -691 -86 -674 -69
rect -481 -86 -464 -69
rect -271 -86 -254 -69
rect -61 -86 -44 -69
rect 149 -86 166 -69
rect 359 -86 376 -69
rect 569 -86 586 -69
rect 779 -86 796 -69
rect 989 -86 1006 -69
rect 1199 -86 1216 -69
rect 1409 -86 1426 -69
rect 1619 -86 1636 -69
rect 1829 -86 1846 -69
rect 2039 -86 2056 -69
<< metal1 >>
rect -2062 86 -2033 89
rect -2062 69 -2056 86
rect -2039 69 -2033 86
rect -2062 66 -2033 69
rect -1852 86 -1823 89
rect -1852 69 -1846 86
rect -1829 69 -1823 86
rect -1852 66 -1823 69
rect -1642 86 -1613 89
rect -1642 69 -1636 86
rect -1619 69 -1613 86
rect -1642 66 -1613 69
rect -1432 86 -1403 89
rect -1432 69 -1426 86
rect -1409 69 -1403 86
rect -1432 66 -1403 69
rect -1222 86 -1193 89
rect -1222 69 -1216 86
rect -1199 69 -1193 86
rect -1222 66 -1193 69
rect -1012 86 -983 89
rect -1012 69 -1006 86
rect -989 69 -983 86
rect -1012 66 -983 69
rect -802 86 -773 89
rect -802 69 -796 86
rect -779 69 -773 86
rect -802 66 -773 69
rect -592 86 -563 89
rect -592 69 -586 86
rect -569 69 -563 86
rect -592 66 -563 69
rect -382 86 -353 89
rect -382 69 -376 86
rect -359 69 -353 86
rect -382 66 -353 69
rect -172 86 -143 89
rect -172 69 -166 86
rect -149 69 -143 86
rect -172 66 -143 69
rect 38 86 67 89
rect 38 69 44 86
rect 61 69 67 86
rect 38 66 67 69
rect 248 86 277 89
rect 248 69 254 86
rect 271 69 277 86
rect 248 66 277 69
rect 458 86 487 89
rect 458 69 464 86
rect 481 69 487 86
rect 458 66 487 69
rect 668 86 697 89
rect 668 69 674 86
rect 691 69 697 86
rect 668 66 697 69
rect 878 86 907 89
rect 878 69 884 86
rect 901 69 907 86
rect 878 66 907 69
rect 1088 86 1117 89
rect 1088 69 1094 86
rect 1111 69 1117 86
rect 1088 66 1117 69
rect 1298 86 1327 89
rect 1298 69 1304 86
rect 1321 69 1327 86
rect 1298 66 1327 69
rect 1508 86 1537 89
rect 1508 69 1514 86
rect 1531 69 1537 86
rect 1508 66 1537 69
rect 1718 86 1747 89
rect 1718 69 1724 86
rect 1741 69 1747 86
rect 1718 66 1747 69
rect 1928 86 1957 89
rect 1928 69 1934 86
rect 1951 69 1957 86
rect 1928 66 1957 69
rect -2086 44 -2057 47
rect -1981 44 -1952 47
rect -1876 44 -1847 47
rect -1771 44 -1742 47
rect -1666 44 -1637 47
rect -1561 44 -1532 47
rect -1456 44 -1427 47
rect -1351 44 -1322 47
rect -1246 44 -1217 47
rect -1141 44 -1112 47
rect -1036 44 -1007 47
rect -931 44 -902 47
rect -826 44 -797 47
rect -721 44 -692 47
rect -616 44 -587 47
rect -511 44 -482 47
rect -406 44 -377 47
rect -301 44 -272 47
rect -196 44 -167 47
rect -91 44 -62 47
rect 14 44 43 47
rect 119 44 148 47
rect 224 44 253 47
rect 329 44 358 47
rect 434 44 463 47
rect 539 44 568 47
rect 644 44 673 47
rect 749 44 778 47
rect 854 44 883 47
rect 959 44 988 47
rect 1064 44 1093 47
rect 1169 44 1198 47
rect 1274 44 1303 47
rect 1379 44 1408 47
rect 1484 44 1513 47
rect 1589 44 1618 47
rect 1694 44 1723 47
rect 1799 44 1828 47
rect 1904 44 1933 47
rect 2009 44 2038 47
rect -2086 27 -2080 44
rect -2063 27 -1975 44
rect -1958 27 -1870 44
rect -1853 27 -1765 44
rect -1748 27 -1660 44
rect -1643 27 -1555 44
rect -1538 27 -1450 44
rect -1433 27 -1345 44
rect -1328 27 -1240 44
rect -1223 27 -1135 44
rect -1118 27 -1030 44
rect -1013 27 -925 44
rect -908 27 -820 44
rect -803 27 -715 44
rect -698 27 -610 44
rect -593 27 -505 44
rect -488 27 -400 44
rect -383 27 -295 44
rect -278 27 -190 44
rect -173 27 -85 44
rect -68 27 20 44
rect 37 27 125 44
rect 142 27 230 44
rect 247 27 335 44
rect 352 27 440 44
rect 457 27 545 44
rect 562 27 650 44
rect 667 27 755 44
rect 772 27 860 44
rect 877 27 965 44
rect 982 27 1070 44
rect 1087 27 1175 44
rect 1192 27 1280 44
rect 1297 27 1385 44
rect 1402 27 1490 44
rect 1507 27 1595 44
rect 1612 27 1700 44
rect 1717 27 1805 44
rect 1822 27 1910 44
rect 1927 27 2015 44
rect 2032 27 2086 44
rect -2086 24 -2057 27
rect -1981 24 -1952 27
rect -1876 24 -1847 27
rect -1771 24 -1742 27
rect -1666 24 -1637 27
rect -1561 24 -1532 27
rect -1456 24 -1427 27
rect -1351 24 -1322 27
rect -1246 24 -1217 27
rect -1141 24 -1112 27
rect -1036 24 -1007 27
rect -931 24 -902 27
rect -826 24 -797 27
rect -721 24 -692 27
rect -616 24 -587 27
rect -511 24 -482 27
rect -406 24 -377 27
rect -301 24 -272 27
rect -196 24 -167 27
rect -91 24 -62 27
rect 14 24 43 27
rect 119 24 148 27
rect 224 24 253 27
rect 329 24 358 27
rect 434 24 463 27
rect 539 24 568 27
rect 644 24 673 27
rect 749 24 778 27
rect 854 24 883 27
rect 959 24 988 27
rect 1064 24 1093 27
rect 1169 24 1198 27
rect 1274 24 1303 27
rect 1379 24 1408 27
rect 1484 24 1513 27
rect 1589 24 1618 27
rect 1694 24 1723 27
rect 1799 24 1828 27
rect 1904 24 1933 27
rect 2009 24 2038 27
rect -2038 -27 -2009 -24
rect -1933 -27 -1904 -24
rect -1828 -27 -1799 -24
rect -1723 -27 -1694 -24
rect -1618 -27 -1589 -24
rect -1513 -27 -1484 -24
rect -1408 -27 -1379 -24
rect -1303 -27 -1274 -24
rect -1198 -27 -1169 -24
rect -1093 -27 -1064 -24
rect -988 -27 -959 -24
rect -883 -27 -854 -24
rect -778 -27 -749 -24
rect -673 -27 -644 -24
rect -568 -27 -539 -24
rect -463 -27 -434 -24
rect -358 -27 -329 -24
rect -253 -27 -224 -24
rect -148 -27 -119 -24
rect -43 -27 -14 -24
rect 62 -27 91 -24
rect 167 -27 196 -24
rect 272 -27 301 -24
rect 377 -27 406 -24
rect 482 -27 511 -24
rect 587 -27 616 -24
rect 692 -27 721 -24
rect 797 -27 826 -24
rect 902 -27 931 -24
rect 1007 -27 1036 -24
rect 1112 -27 1141 -24
rect 1217 -27 1246 -24
rect 1322 -27 1351 -24
rect 1427 -27 1456 -24
rect 1532 -27 1561 -24
rect 1637 -27 1666 -24
rect 1742 -27 1771 -24
rect 1847 -27 1876 -24
rect 1952 -27 1981 -24
rect 2057 -27 2086 -24
rect -2086 -44 -2032 -27
rect -2015 -44 -1927 -27
rect -1910 -44 -1822 -27
rect -1805 -44 -1717 -27
rect -1700 -44 -1612 -27
rect -1595 -44 -1507 -27
rect -1490 -44 -1402 -27
rect -1385 -44 -1297 -27
rect -1280 -44 -1192 -27
rect -1175 -44 -1087 -27
rect -1070 -44 -982 -27
rect -965 -44 -877 -27
rect -860 -44 -772 -27
rect -755 -44 -667 -27
rect -650 -44 -562 -27
rect -545 -44 -457 -27
rect -440 -44 -352 -27
rect -335 -44 -247 -27
rect -230 -44 -142 -27
rect -125 -44 -37 -27
rect -20 -44 68 -27
rect 85 -44 173 -27
rect 190 -44 278 -27
rect 295 -44 383 -27
rect 400 -44 488 -27
rect 505 -44 593 -27
rect 610 -44 698 -27
rect 715 -44 803 -27
rect 820 -44 908 -27
rect 925 -44 1013 -27
rect 1030 -44 1118 -27
rect 1135 -44 1223 -27
rect 1240 -44 1328 -27
rect 1345 -44 1433 -27
rect 1450 -44 1538 -27
rect 1555 -44 1643 -27
rect 1660 -44 1748 -27
rect 1765 -44 1853 -27
rect 1870 -44 1958 -27
rect 1975 -44 2063 -27
rect 2080 -44 2086 -27
rect -2038 -47 -2009 -44
rect -1933 -47 -1904 -44
rect -1828 -47 -1799 -44
rect -1723 -47 -1694 -44
rect -1618 -47 -1589 -44
rect -1513 -47 -1484 -44
rect -1408 -47 -1379 -44
rect -1303 -47 -1274 -44
rect -1198 -47 -1169 -44
rect -1093 -47 -1064 -44
rect -988 -47 -959 -44
rect -883 -47 -854 -44
rect -778 -47 -749 -44
rect -673 -47 -644 -44
rect -568 -47 -539 -44
rect -463 -47 -434 -44
rect -358 -47 -329 -44
rect -253 -47 -224 -44
rect -148 -47 -119 -44
rect -43 -47 -14 -44
rect 62 -47 91 -44
rect 167 -47 196 -44
rect 272 -47 301 -44
rect 377 -47 406 -44
rect 482 -47 511 -44
rect 587 -47 616 -44
rect 692 -47 721 -44
rect 797 -47 826 -44
rect 902 -47 931 -44
rect 1007 -47 1036 -44
rect 1112 -47 1141 -44
rect 1217 -47 1246 -44
rect 1322 -47 1351 -44
rect 1427 -47 1456 -44
rect 1532 -47 1561 -44
rect 1637 -47 1666 -44
rect 1742 -47 1771 -44
rect 1847 -47 1876 -44
rect 1952 -47 1981 -44
rect 2057 -47 2086 -44
rect -1957 -69 -1928 -66
rect -1957 -86 -1951 -69
rect -1934 -86 -1928 -69
rect -1957 -89 -1928 -86
rect -1747 -69 -1718 -66
rect -1747 -86 -1741 -69
rect -1724 -86 -1718 -69
rect -1747 -89 -1718 -86
rect -1537 -69 -1508 -66
rect -1537 -86 -1531 -69
rect -1514 -86 -1508 -69
rect -1537 -89 -1508 -86
rect -1327 -69 -1298 -66
rect -1327 -86 -1321 -69
rect -1304 -86 -1298 -69
rect -1327 -89 -1298 -86
rect -1117 -69 -1088 -66
rect -1117 -86 -1111 -69
rect -1094 -86 -1088 -69
rect -1117 -89 -1088 -86
rect -907 -69 -878 -66
rect -907 -86 -901 -69
rect -884 -86 -878 -69
rect -907 -89 -878 -86
rect -697 -69 -668 -66
rect -697 -86 -691 -69
rect -674 -86 -668 -69
rect -697 -89 -668 -86
rect -487 -69 -458 -66
rect -487 -86 -481 -69
rect -464 -86 -458 -69
rect -487 -89 -458 -86
rect -277 -69 -248 -66
rect -277 -86 -271 -69
rect -254 -86 -248 -69
rect -277 -89 -248 -86
rect -67 -69 -38 -66
rect -67 -86 -61 -69
rect -44 -86 -38 -69
rect -67 -89 -38 -86
rect 143 -69 172 -66
rect 143 -86 149 -69
rect 166 -86 172 -69
rect 143 -89 172 -86
rect 353 -69 382 -66
rect 353 -86 359 -69
rect 376 -86 382 -69
rect 353 -89 382 -86
rect 563 -69 592 -66
rect 563 -86 569 -69
rect 586 -86 592 -69
rect 563 -89 592 -86
rect 773 -69 802 -66
rect 773 -86 779 -69
rect 796 -86 802 -69
rect 773 -89 802 -86
rect 983 -69 1012 -66
rect 983 -86 989 -69
rect 1006 -86 1012 -69
rect 983 -89 1012 -86
rect 1193 -69 1222 -66
rect 1193 -86 1199 -69
rect 1216 -86 1222 -69
rect 1193 -89 1222 -86
rect 1403 -69 1432 -66
rect 1403 -86 1409 -69
rect 1426 -86 1432 -69
rect 1403 -89 1432 -86
rect 1613 -69 1642 -66
rect 1613 -86 1619 -69
rect 1636 -86 1642 -69
rect 1613 -89 1642 -86
rect 1823 -69 1852 -66
rect 1823 -86 1829 -69
rect 1846 -86 1852 -69
rect 1823 -89 1852 -86
rect 2033 -69 2062 -66
rect 2033 -86 2039 -69
rect 2056 -86 2062 -69
rect 2033 -89 2062 -86
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 42 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
